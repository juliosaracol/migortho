module top (
            pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518, pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526, pi3527, pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535, pi3536, pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544, pi3545, pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553, pi3554, pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562, pi3563, pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571, pi3572, pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580, pi3581, pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589, pi3590, pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598, pi3599, pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607, pi3608, pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616, pi3617, pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625, pi3626, pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634, pi3635, pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643, pi3644, pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652, pi3653, pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661, pi3662, pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670, pi3671, pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679, pi3680, pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688, pi3689, pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697, pi3698, pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706, pi3707, pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715, pi3716, pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724, pi3725, pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733, pi3734, pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742, pi3743, pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751, pi3752, pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760, pi3761, pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769, pi3770, pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778, pi3779, pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787, pi3788, pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796, pi3797, pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805, pi3806, pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814, pi3815, pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823, pi3824, pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832, pi3833, pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841, pi3842, pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850, pi3851, pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859, pi3860, pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868, pi3869, pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877, pi3878, pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886, pi3887, pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895, pi3896, pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904, pi3905, pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913, pi3914, pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922, pi3923, pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931, pi3932, pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940, pi3941, pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949, pi3950, pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958, pi3959, pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967, pi3968, pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976, pi3977, pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985, pi3986, pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994, pi3995, pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003, pi4004, pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012, pi4013, pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021, pi4022, pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030, pi4031, pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039, pi4040, pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048, pi4049, pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057, pi4058, pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066, pi4067, pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075, pi4076, pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084, pi4085, pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093, pi4094, pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102, pi4103, pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111, pi4112, pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120, pi4121, pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129, pi4130, pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138, pi4139, pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147, pi4148, pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156, pi4157, pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165, pi4166, pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174, pi4175, pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183, pi4184, pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192, pi4193, pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201, pi4202, pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210, pi4211, pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219, pi4220, pi4221, pi4222, 
            po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535, po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544, po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553, po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562, po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571, po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580, po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589, po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598, po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607, po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616, po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625, po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634, po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643, po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652, po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661, po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670, po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679, po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688, po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697, po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706, po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715, po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724, po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733, po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742, po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751, po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760, po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769, po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778, po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787, po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796, po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805, po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814, po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823, po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832, po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841, po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850, po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859, po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868, po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877, po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886, po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895, po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904, po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913, po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922, po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931, po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940, po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949, po3950, po3951, po3952);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518, pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526, pi3527, pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535, pi3536, pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544, pi3545, pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553, pi3554, pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562, pi3563, pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571, pi3572, pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580, pi3581, pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589, pi3590, pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598, pi3599, pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607, pi3608, pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616, pi3617, pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625, pi3626, pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634, pi3635, pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643, pi3644, pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652, pi3653, pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661, pi3662, pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670, pi3671, pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679, pi3680, pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688, pi3689, pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697, pi3698, pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706, pi3707, pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715, pi3716, pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724, pi3725, pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733, pi3734, pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742, pi3743, pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751, pi3752, pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760, pi3761, pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769, pi3770, pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778, pi3779, pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787, pi3788, pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796, pi3797, pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805, pi3806, pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814, pi3815, pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823, pi3824, pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832, pi3833, pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841, pi3842, pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850, pi3851, pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859, pi3860, pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868, pi3869, pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877, pi3878, pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886, pi3887, pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895, pi3896, pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904, pi3905, pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913, pi3914, pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922, pi3923, pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931, pi3932, pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940, pi3941, pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949, pi3950, pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958, pi3959, pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967, pi3968, pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976, pi3977, pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985, pi3986, pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994, pi3995, pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003, pi4004, pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012, pi4013, pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021, pi4022, pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030, pi4031, pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039, pi4040, pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048, pi4049, pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057, pi4058, pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066, pi4067, pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075, pi4076, pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084, pi4085, pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093, pi4094, pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102, pi4103, pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111, pi4112, pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120, pi4121, pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129, pi4130, pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138, pi4139, pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147, pi4148, pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156, pi4157, pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165, pi4166, pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174, pi4175, pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183, pi4184, pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192, pi4193, pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201, pi4202, pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210, pi4211, pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219, pi4220, pi4221, pi4222;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535, po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544, po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553, po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562, po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571, po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580, po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589, po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598, po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607, po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616, po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625, po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634, po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643, po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652, po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661, po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670, po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679, po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688, po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697, po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706, po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715, po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724, po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733, po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742, po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751, po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760, po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769, po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778, po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787, po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796, po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805, po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814, po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823, po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832, po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841, po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850, po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859, po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868, po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877, po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886, po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895, po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904, po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913, po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922, po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931, po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940, po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949, po3950, po3951, po3952;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602, w18603, w18604, w18605, w18606, w18607, w18608, w18609, w18610, w18611, w18612, w18613, w18614, w18615, w18616, w18617, w18618, w18619, w18620, w18621, w18622, w18623, w18624, w18625, w18626, w18627, w18628, w18629, w18630, w18631, w18632, w18633, w18634, w18635, w18636, w18637, w18638, w18639, w18640, w18641, w18642, w18643, w18644, w18645, w18646, w18647, w18648, w18649, w18650, w18651, w18652, w18653, w18654, w18655, w18656, w18657, w18658, w18659, w18660, w18661, w18662, w18663, w18664, w18665, w18666, w18667, w18668, w18669, w18670, w18671, w18672, w18673, w18674, w18675, w18676, w18677, w18678, w18679, w18680, w18681, w18682, w18683, w18684, w18685, w18686, w18687, w18688, w18689, w18690, w18691, w18692, w18693, w18694, w18695, w18696, w18697, w18698, w18699, w18700, w18701, w18702, w18703, w18704, w18705, w18706, w18707, w18708, w18709, w18710, w18711, w18712, w18713, w18714, w18715, w18716, w18717, w18718, w18719, w18720, w18721, w18722, w18723, w18724, w18725, w18726, w18727, w18728, w18729, w18730, w18731, w18732, w18733, w18734, w18735, w18736, w18737, w18738, w18739, w18740, w18741, w18742, w18743, w18744, w18745, w18746, w18747, w18748, w18749, w18750, w18751, w18752, w18753, w18754, w18755, w18756, w18757, w18758, w18759, w18760, w18761, w18762, w18763, w18764, w18765, w18766, w18767, w18768, w18769, w18770, w18771, w18772, w18773, w18774, w18775, w18776, w18777, w18778, w18779, w18780, w18781, w18782, w18783, w18784, w18785, w18786, w18787, w18788, w18789, w18790, w18791, w18792, w18793, w18794, w18795, w18796, w18797, w18798, w18799, w18800, w18801, w18802, w18803, w18804, w18805, w18806, w18807, w18808, w18809, w18810, w18811, w18812, w18813, w18814, w18815, w18816, w18817, w18818, w18819, w18820, w18821, w18822, w18823, w18824, w18825, w18826, w18827, w18828, w18829, w18830, w18831, w18832, w18833, w18834, w18835, w18836, w18837, w18838, w18839, w18840, w18841, w18842, w18843, w18844, w18845, w18846, w18847, w18848, w18849, w18850, w18851, w18852, w18853, w18854, w18855, w18856, w18857, w18858, w18859, w18860, w18861, w18862, w18863, w18864, w18865, w18866, w18867, w18868, w18869, w18870, w18871, w18872, w18873, w18874, w18875, w18876, w18877, w18878, w18879, w18880, w18881, w18882, w18883, w18884, w18885, w18886, w18887, w18888, w18889, w18890, w18891, w18892, w18893, w18894, w18895, w18896, w18897, w18898, w18899, w18900, w18901, w18902, w18903, w18904, w18905, w18906, w18907, w18908, w18909, w18910, w18911, w18912, w18913, w18914, w18915, w18916, w18917, w18918, w18919, w18920, w18921, w18922, w18923, w18924, w18925, w18926, w18927, w18928, w18929, w18930, w18931, w18932, w18933, w18934, w18935, w18936, w18937, w18938, w18939, w18940, w18941, w18942, w18943, w18944, w18945, w18946, w18947, w18948, w18949, w18950, w18951, w18952, w18953, w18954, w18955, w18956, w18957, w18958, w18959, w18960, w18961, w18962, w18963, w18964, w18965, w18966, w18967, w18968, w18969, w18970, w18971, w18972, w18973, w18974, w18975, w18976, w18977, w18978, w18979, w18980, w18981, w18982, w18983, w18984, w18985, w18986, w18987, w18988, w18989, w18990, w18991, w18992, w18993, w18994, w18995, w18996, w18997, w18998, w18999, w19000, w19001, w19002, w19003, w19004, w19005, w19006, w19007, w19008, w19009, w19010, w19011, w19012, w19013, w19014, w19015, w19016, w19017, w19018, w19019, w19020, w19021, w19022, w19023, w19024, w19025, w19026, w19027, w19028, w19029, w19030, w19031, w19032, w19033, w19034, w19035, w19036, w19037, w19038, w19039, w19040, w19041, w19042, w19043, w19044, w19045, w19046, w19047, w19048, w19049, w19050, w19051, w19052, w19053, w19054, w19055, w19056, w19057, w19058, w19059, w19060, w19061, w19062, w19063, w19064, w19065, w19066, w19067, w19068, w19069, w19070, w19071, w19072, w19073, w19074, w19075, w19076, w19077, w19078, w19079, w19080, w19081, w19082, w19083, w19084, w19085, w19086, w19087, w19088, w19089, w19090, w19091, w19092, w19093, w19094, w19095, w19096, w19097, w19098, w19099, w19100, w19101, w19102, w19103, w19104, w19105, w19106, w19107, w19108, w19109, w19110, w19111, w19112, w19113, w19114, w19115, w19116, w19117, w19118, w19119, w19120, w19121, w19122, w19123, w19124, w19125, w19126, w19127, w19128, w19129, w19130, w19131, w19132, w19133, w19134, w19135, w19136, w19137, w19138, w19139, w19140, w19141, w19142, w19143, w19144, w19145, w19146, w19147, w19148, w19149, w19150, w19151, w19152, w19153, w19154, w19155, w19156, w19157, w19158, w19159, w19160, w19161, w19162, w19163, w19164, w19165, w19166, w19167, w19168, w19169, w19170, w19171, w19172, w19173, w19174, w19175, w19176, w19177, w19178, w19179, w19180, w19181, w19182, w19183, w19184, w19185, w19186, w19187, w19188, w19189, w19190, w19191, w19192, w19193, w19194, w19195, w19196, w19197, w19198, w19199, w19200, w19201, w19202, w19203, w19204, w19205, w19206, w19207, w19208, w19209, w19210, w19211, w19212, w19213, w19214, w19215, w19216, w19217, w19218, w19219, w19220, w19221, w19222, w19223, w19224, w19225, w19226, w19227, w19228, w19229, w19230, w19231, w19232, w19233, w19234, w19235, w19236, w19237, w19238, w19239, w19240, w19241, w19242, w19243, w19244, w19245, w19246, w19247, w19248, w19249, w19250, w19251, w19252, w19253, w19254, w19255, w19256, w19257, w19258, w19259, w19260, w19261, w19262, w19263, w19264, w19265, w19266, w19267, w19268, w19269, w19270, w19271, w19272, w19273, w19274, w19275, w19276, w19277, w19278, w19279, w19280, w19281, w19282, w19283, w19284, w19285, w19286, w19287, w19288, w19289, w19290, w19291, w19292, w19293, w19294, w19295, w19296, w19297, w19298, w19299, w19300, w19301, w19302, w19303, w19304, w19305, w19306, w19307, w19308, w19309, w19310, w19311, w19312, w19313, w19314, w19315, w19316, w19317, w19318, w19319, w19320, w19321, w19322, w19323, w19324, w19325, w19326, w19327, w19328, w19329, w19330, w19331, w19332, w19333, w19334, w19335, w19336, w19337, w19338, w19339, w19340, w19341, w19342, w19343, w19344, w19345, w19346, w19347, w19348, w19349, w19350, w19351, w19352, w19353, w19354, w19355, w19356, w19357, w19358, w19359, w19360, w19361, w19362, w19363, w19364, w19365, w19366, w19367, w19368, w19369, w19370, w19371, w19372, w19373, w19374, w19375, w19376, w19377, w19378, w19379, w19380, w19381, w19382, w19383, w19384, w19385, w19386, w19387, w19388, w19389, w19390, w19391, w19392, w19393, w19394, w19395, w19396, w19397, w19398, w19399, w19400, w19401, w19402, w19403, w19404, w19405, w19406, w19407, w19408, w19409, w19410, w19411, w19412, w19413, w19414, w19415, w19416, w19417, w19418, w19419, w19420, w19421, w19422, w19423, w19424, w19425, w19426, w19427, w19428, w19429, w19430, w19431, w19432, w19433, w19434, w19435, w19436, w19437, w19438, w19439, w19440, w19441, w19442, w19443, w19444, w19445, w19446, w19447, w19448, w19449, w19450, w19451, w19452, w19453, w19454, w19455, w19456, w19457, w19458, w19459, w19460, w19461, w19462, w19463, w19464, w19465, w19466, w19467, w19468, w19469, w19470, w19471, w19472, w19473, w19474, w19475, w19476, w19477, w19478, w19479, w19480, w19481, w19482, w19483, w19484, w19485, w19486, w19487, w19488, w19489, w19490, w19491, w19492, w19493, w19494, w19495, w19496, w19497, w19498, w19499, w19500, w19501, w19502, w19503, w19504, w19505, w19506, w19507, w19508, w19509, w19510, w19511, w19512, w19513, w19514, w19515, w19516, w19517, w19518, w19519, w19520, w19521, w19522, w19523, w19524, w19525, w19526, w19527, w19528, w19529, w19530, w19531, w19532, w19533, w19534, w19535, w19536, w19537, w19538, w19539, w19540, w19541, w19542, w19543, w19544, w19545, w19546, w19547, w19548, w19549, w19550, w19551, w19552, w19553, w19554, w19555, w19556, w19557, w19558, w19559, w19560, w19561, w19562, w19563, w19564, w19565, w19566, w19567, w19568, w19569, w19570, w19571, w19572, w19573, w19574, w19575, w19576, w19577, w19578, w19579, w19580, w19581, w19582, w19583, w19584, w19585, w19586, w19587, w19588, w19589, w19590, w19591, w19592, w19593, w19594, w19595, w19596, w19597, w19598, w19599, w19600, w19601, w19602, w19603, w19604, w19605, w19606, w19607, w19608, w19609, w19610, w19611, w19612, w19613, w19614, w19615, w19616, w19617, w19618, w19619, w19620, w19621, w19622, w19623, w19624, w19625, w19626, w19627, w19628, w19629, w19630, w19631, w19632, w19633, w19634, w19635, w19636, w19637, w19638, w19639, w19640, w19641, w19642, w19643, w19644, w19645, w19646, w19647, w19648, w19649, w19650, w19651, w19652, w19653, w19654, w19655, w19656, w19657, w19658, w19659, w19660, w19661, w19662, w19663, w19664, w19665, w19666, w19667, w19668, w19669, w19670, w19671, w19672, w19673, w19674, w19675, w19676, w19677, w19678, w19679, w19680, w19681, w19682, w19683, w19684, w19685, w19686, w19687, w19688, w19689, w19690, w19691, w19692, w19693, w19694, w19695, w19696, w19697, w19698, w19699, w19700, w19701, w19702, w19703, w19704, w19705, w19706, w19707, w19708, w19709, w19710, w19711, w19712, w19713, w19714, w19715, w19716, w19717, w19718, w19719, w19720, w19721, w19722, w19723, w19724, w19725, w19726, w19727, w19728, w19729, w19730, w19731, w19732, w19733, w19734, w19735, w19736, w19737, w19738, w19739, w19740, w19741, w19742, w19743, w19744, w19745, w19746, w19747, w19748, w19749, w19750, w19751, w19752, w19753, w19754, w19755, w19756, w19757, w19758, w19759, w19760, w19761, w19762, w19763, w19764, w19765, w19766, w19767, w19768, w19769, w19770, w19771, w19772, w19773, w19774, w19775, w19776, w19777, w19778, w19779, w19780, w19781, w19782, w19783, w19784, w19785, w19786, w19787, w19788, w19789, w19790, w19791, w19792, w19793, w19794, w19795, w19796, w19797, w19798, w19799, w19800, w19801, w19802, w19803, w19804, w19805, w19806, w19807, w19808, w19809, w19810, w19811, w19812, w19813, w19814, w19815, w19816, w19817, w19818, w19819, w19820, w19821, w19822, w19823, w19824, w19825, w19826, w19827, w19828, w19829, w19830, w19831, w19832, w19833, w19834, w19835, w19836, w19837, w19838, w19839, w19840, w19841, w19842, w19843, w19844, w19845, w19846, w19847, w19848, w19849, w19850, w19851, w19852, w19853, w19854, w19855, w19856, w19857, w19858, w19859, w19860, w19861, w19862, w19863, w19864, w19865, w19866, w19867, w19868, w19869, w19870, w19871, w19872, w19873, w19874, w19875, w19876, w19877, w19878, w19879, w19880, w19881, w19882, w19883, w19884, w19885, w19886, w19887, w19888, w19889, w19890, w19891, w19892, w19893, w19894, w19895, w19896, w19897, w19898, w19899, w19900, w19901, w19902, w19903, w19904, w19905, w19906, w19907, w19908, w19909, w19910, w19911, w19912, w19913, w19914, w19915, w19916, w19917, w19918, w19919, w19920, w19921, w19922, w19923, w19924, w19925, w19926, w19927, w19928, w19929, w19930, w19931, w19932, w19933, w19934, w19935, w19936, w19937, w19938, w19939, w19940, w19941, w19942, w19943, w19944, w19945, w19946, w19947, w19948, w19949, w19950, w19951, w19952, w19953, w19954, w19955, w19956, w19957, w19958, w19959, w19960, w19961, w19962, w19963, w19964, w19965, w19966, w19967, w19968, w19969, w19970, w19971, w19972, w19973, w19974, w19975, w19976, w19977, w19978, w19979, w19980, w19981, w19982, w19983, w19984, w19985, w19986, w19987, w19988, w19989, w19990, w19991, w19992, w19993, w19994, w19995, w19996, w19997, w19998, w19999, w20000, w20001, w20002, w20003, w20004, w20005, w20006, w20007, w20008, w20009, w20010, w20011, w20012, w20013, w20014, w20015, w20016, w20017, w20018, w20019, w20020, w20021, w20022, w20023, w20024, w20025, w20026, w20027, w20028, w20029, w20030, w20031, w20032, w20033, w20034, w20035, w20036, w20037, w20038, w20039, w20040, w20041, w20042, w20043, w20044, w20045, w20046, w20047, w20048, w20049, w20050, w20051, w20052, w20053, w20054, w20055, w20056, w20057, w20058, w20059, w20060, w20061, w20062, w20063, w20064, w20065, w20066, w20067, w20068, w20069, w20070, w20071, w20072, w20073, w20074, w20075, w20076, w20077, w20078, w20079, w20080, w20081, w20082, w20083, w20084, w20085, w20086, w20087, w20088, w20089, w20090, w20091, w20092, w20093, w20094, w20095, w20096, w20097, w20098, w20099, w20100, w20101, w20102, w20103, w20104, w20105, w20106, w20107, w20108, w20109, w20110, w20111, w20112, w20113, w20114, w20115, w20116, w20117, w20118, w20119, w20120, w20121, w20122, w20123, w20124, w20125, w20126, w20127, w20128, w20129, w20130, w20131, w20132, w20133, w20134, w20135, w20136, w20137, w20138, w20139, w20140, w20141, w20142, w20143, w20144, w20145, w20146, w20147, w20148, w20149, w20150, w20151, w20152, w20153, w20154, w20155, w20156, w20157, w20158, w20159, w20160, w20161, w20162, w20163, w20164, w20165, w20166, w20167, w20168, w20169, w20170, w20171, w20172, w20173, w20174, w20175, w20176, w20177, w20178, w20179, w20180, w20181, w20182, w20183, w20184, w20185, w20186, w20187, w20188, w20189, w20190, w20191, w20192, w20193, w20194, w20195, w20196, w20197, w20198, w20199, w20200, w20201, w20202, w20203, w20204, w20205, w20206, w20207, w20208, w20209, w20210, w20211, w20212, w20213, w20214, w20215, w20216, w20217, w20218, w20219, w20220, w20221, w20222, w20223, w20224, w20225, w20226, w20227, w20228, w20229, w20230, w20231, w20232, w20233, w20234, w20235, w20236, w20237, w20238, w20239, w20240, w20241, w20242, w20243, w20244, w20245, w20246, w20247, w20248, w20249, w20250, w20251, w20252, w20253, w20254, w20255, w20256, w20257, w20258, w20259, w20260, w20261, w20262, w20263, w20264, w20265, w20266, w20267, w20268, w20269, w20270, w20271, w20272, w20273, w20274, w20275, w20276, w20277, w20278, w20279, w20280, w20281, w20282, w20283, w20284, w20285, w20286, w20287, w20288, w20289, w20290, w20291, w20292, w20293, w20294, w20295, w20296, w20297, w20298, w20299, w20300, w20301, w20302, w20303, w20304, w20305, w20306, w20307, w20308, w20309, w20310, w20311, w20312, w20313, w20314, w20315, w20316, w20317, w20318, w20319, w20320, w20321, w20322, w20323, w20324, w20325, w20326, w20327, w20328, w20329, w20330, w20331, w20332, w20333, w20334, w20335, w20336, w20337, w20338, w20339, w20340, w20341, w20342, w20343, w20344, w20345, w20346, w20347, w20348, w20349, w20350, w20351, w20352, w20353, w20354, w20355, w20356, w20357, w20358, w20359, w20360, w20361, w20362, w20363, w20364, w20365, w20366, w20367, w20368, w20369, w20370, w20371, w20372, w20373, w20374, w20375, w20376, w20377, w20378, w20379, w20380, w20381, w20382, w20383, w20384, w20385, w20386, w20387, w20388, w20389, w20390, w20391, w20392, w20393, w20394, w20395, w20396, w20397, w20398, w20399, w20400, w20401, w20402, w20403, w20404, w20405, w20406, w20407, w20408, w20409, w20410, w20411, w20412, w20413, w20414, w20415, w20416, w20417, w20418, w20419, w20420, w20421, w20422, w20423, w20424, w20425, w20426, w20427, w20428, w20429, w20430, w20431, w20432, w20433, w20434, w20435, w20436, w20437, w20438, w20439, w20440, w20441, w20442, w20443, w20444, w20445, w20446, w20447, w20448, w20449, w20450, w20451, w20452, w20453, w20454, w20455, w20456, w20457, w20458, w20459, w20460, w20461, w20462, w20463, w20464, w20465, w20466, w20467, w20468, w20469, w20470, w20471, w20472, w20473, w20474, w20475, w20476, w20477, w20478, w20479, w20480, w20481, w20482, w20483, w20484, w20485, w20486, w20487, w20488, w20489, w20490, w20491, w20492, w20493, w20494, w20495, w20496, w20497, w20498, w20499, w20500, w20501, w20502, w20503, w20504, w20505, w20506, w20507, w20508, w20509, w20510, w20511, w20512, w20513, w20514, w20515, w20516, w20517, w20518, w20519, w20520, w20521, w20522, w20523, w20524, w20525, w20526, w20527, w20528, w20529, w20530, w20531, w20532, w20533, w20534, w20535, w20536, w20537, w20538, w20539, w20540, w20541, w20542, w20543, w20544, w20545, w20546, w20547, w20548, w20549, w20550, w20551, w20552, w20553, w20554, w20555, w20556, w20557, w20558, w20559, w20560, w20561, w20562, w20563, w20564, w20565, w20566, w20567, w20568, w20569, w20570, w20571, w20572, w20573, w20574, w20575, w20576, w20577, w20578, w20579, w20580, w20581, w20582, w20583, w20584, w20585, w20586, w20587, w20588, w20589, w20590, w20591, w20592, w20593, w20594, w20595, w20596, w20597, w20598, w20599, w20600, w20601, w20602, w20603, w20604, w20605, w20606, w20607, w20608, w20609, w20610, w20611, w20612, w20613, w20614, w20615, w20616, w20617, w20618, w20619, w20620, w20621, w20622, w20623, w20624, w20625, w20626, w20627, w20628, w20629, w20630, w20631, w20632, w20633, w20634, w20635, w20636, w20637, w20638, w20639, w20640, w20641, w20642, w20643, w20644, w20645, w20646, w20647, w20648, w20649, w20650, w20651, w20652, w20653, w20654, w20655, w20656, w20657, w20658, w20659, w20660, w20661, w20662, w20663, w20664, w20665, w20666, w20667, w20668, w20669, w20670, w20671, w20672, w20673, w20674, w20675, w20676, w20677, w20678, w20679, w20680, w20681, w20682, w20683, w20684, w20685, w20686, w20687, w20688, w20689, w20690, w20691, w20692, w20693, w20694, w20695, w20696, w20697, w20698, w20699, w20700, w20701, w20702, w20703, w20704, w20705, w20706, w20707, w20708, w20709, w20710, w20711, w20712, w20713, w20714, w20715, w20716, w20717, w20718, w20719, w20720, w20721, w20722, w20723, w20724, w20725, w20726, w20727, w20728, w20729, w20730, w20731, w20732, w20733, w20734, w20735, w20736, w20737, w20738, w20739, w20740, w20741, w20742, w20743, w20744, w20745, w20746, w20747, w20748, w20749, w20750, w20751, w20752, w20753, w20754, w20755, w20756, w20757, w20758, w20759, w20760, w20761, w20762, w20763, w20764, w20765, w20766, w20767, w20768, w20769, w20770, w20771, w20772, w20773, w20774, w20775, w20776, w20777, w20778, w20779, w20780, w20781, w20782, w20783, w20784, w20785, w20786, w20787, w20788, w20789, w20790, w20791, w20792, w20793, w20794, w20795, w20796, w20797, w20798, w20799, w20800, w20801, w20802, w20803, w20804, w20805, w20806, w20807, w20808, w20809, w20810, w20811, w20812, w20813, w20814, w20815, w20816, w20817, w20818, w20819, w20820, w20821, w20822, w20823, w20824, w20825, w20826, w20827, w20828, w20829, w20830, w20831, w20832, w20833, w20834, w20835, w20836, w20837, w20838, w20839, w20840, w20841, w20842, w20843, w20844, w20845, w20846, w20847, w20848, w20849, w20850, w20851, w20852, w20853, w20854, w20855, w20856, w20857, w20858, w20859, w20860, w20861, w20862, w20863, w20864, w20865, w20866, w20867, w20868, w20869, w20870, w20871, w20872, w20873, w20874, w20875, w20876, w20877, w20878, w20879, w20880, w20881, w20882, w20883, w20884, w20885, w20886, w20887, w20888, w20889, w20890, w20891, w20892, w20893, w20894, w20895, w20896, w20897, w20898, w20899, w20900, w20901, w20902, w20903, w20904, w20905, w20906, w20907, w20908, w20909, w20910, w20911, w20912, w20913, w20914, w20915, w20916, w20917, w20918, w20919, w20920, w20921, w20922, w20923, w20924, w20925, w20926, w20927, w20928, w20929, w20930, w20931, w20932, w20933, w20934, w20935, w20936, w20937, w20938, w20939, w20940, w20941, w20942, w20943, w20944, w20945, w20946, w20947, w20948, w20949, w20950, w20951, w20952, w20953, w20954, w20955, w20956, w20957, w20958, w20959, w20960, w20961, w20962, w20963, w20964, w20965, w20966, w20967, w20968, w20969, w20970, w20971, w20972, w20973, w20974, w20975, w20976, w20977, w20978, w20979, w20980, w20981, w20982, w20983, w20984, w20985, w20986, w20987, w20988, w20989, w20990, w20991, w20992, w20993, w20994, w20995, w20996, w20997, w20998, w20999, w21000, w21001, w21002, w21003, w21004, w21005, w21006, w21007, w21008, w21009, w21010, w21011, w21012, w21013, w21014, w21015, w21016, w21017, w21018, w21019, w21020, w21021, w21022, w21023, w21024, w21025, w21026, w21027, w21028, w21029, w21030, w21031, w21032, w21033, w21034, w21035, w21036, w21037, w21038, w21039, w21040, w21041, w21042, w21043, w21044, w21045, w21046, w21047, w21048, w21049, w21050, w21051, w21052, w21053, w21054, w21055, w21056, w21057, w21058, w21059, w21060, w21061, w21062, w21063, w21064, w21065, w21066, w21067, w21068, w21069, w21070, w21071, w21072, w21073, w21074, w21075, w21076, w21077, w21078, w21079, w21080, w21081, w21082, w21083, w21084, w21085, w21086, w21087, w21088, w21089, w21090, w21091, w21092, w21093, w21094, w21095, w21096, w21097, w21098, w21099, w21100, w21101, w21102, w21103, w21104, w21105, w21106, w21107, w21108, w21109, w21110, w21111, w21112, w21113, w21114, w21115, w21116, w21117, w21118, w21119, w21120, w21121, w21122, w21123, w21124, w21125, w21126, w21127, w21128, w21129, w21130, w21131, w21132, w21133, w21134, w21135, w21136, w21137, w21138, w21139, w21140, w21141, w21142, w21143, w21144, w21145, w21146, w21147, w21148, w21149, w21150, w21151, w21152, w21153, w21154, w21155, w21156, w21157, w21158, w21159, w21160, w21161, w21162, w21163, w21164, w21165, w21166, w21167, w21168, w21169, w21170, w21171, w21172, w21173, w21174, w21175, w21176, w21177, w21178, w21179, w21180, w21181, w21182, w21183, w21184, w21185, w21186, w21187, w21188, w21189, w21190, w21191, w21192, w21193, w21194, w21195, w21196, w21197, w21198, w21199, w21200, w21201, w21202, w21203, w21204, w21205, w21206, w21207, w21208, w21209, w21210, w21211, w21212, w21213, w21214, w21215, w21216, w21217, w21218, w21219, w21220, w21221, w21222, w21223, w21224, w21225, w21226, w21227, w21228, w21229, w21230, w21231, w21232, w21233, w21234, w21235, w21236, w21237, w21238, w21239, w21240, w21241, w21242, w21243, w21244, w21245, w21246, w21247, w21248, w21249, w21250, w21251, w21252, w21253, w21254, w21255, w21256, w21257, w21258, w21259, w21260, w21261, w21262, w21263, w21264, w21265, w21266, w21267, w21268, w21269, w21270, w21271, w21272, w21273, w21274, w21275, w21276, w21277, w21278, w21279, w21280, w21281, w21282, w21283, w21284, w21285, w21286, w21287, w21288, w21289, w21290, w21291, w21292, w21293, w21294, w21295, w21296, w21297, w21298, w21299, w21300, w21301, w21302, w21303, w21304, w21305, w21306, w21307, w21308, w21309, w21310, w21311, w21312, w21313, w21314, w21315, w21316, w21317, w21318, w21319, w21320, w21321, w21322, w21323, w21324, w21325, w21326, w21327, w21328, w21329, w21330, w21331, w21332, w21333, w21334, w21335, w21336, w21337, w21338, w21339, w21340, w21341, w21342, w21343, w21344, w21345, w21346, w21347, w21348, w21349, w21350, w21351, w21352, w21353, w21354, w21355, w21356, w21357, w21358, w21359, w21360, w21361, w21362, w21363, w21364, w21365, w21366, w21367, w21368, w21369, w21370, w21371, w21372, w21373, w21374, w21375, w21376, w21377, w21378, w21379, w21380, w21381, w21382, w21383, w21384, w21385, w21386, w21387, w21388, w21389, w21390, w21391, w21392, w21393, w21394, w21395, w21396, w21397, w21398, w21399, w21400, w21401, w21402, w21403, w21404, w21405, w21406, w21407, w21408, w21409, w21410, w21411, w21412, w21413, w21414, w21415, w21416, w21417, w21418, w21419, w21420, w21421, w21422, w21423, w21424, w21425, w21426, w21427, w21428, w21429, w21430, w21431, w21432, w21433, w21434, w21435, w21436, w21437, w21438, w21439, w21440, w21441, w21442, w21443, w21444, w21445, w21446, w21447, w21448, w21449, w21450, w21451, w21452, w21453, w21454, w21455, w21456, w21457, w21458, w21459, w21460, w21461, w21462, w21463, w21464, w21465, w21466, w21467, w21468, w21469, w21470, w21471, w21472, w21473, w21474, w21475, w21476, w21477, w21478, w21479, w21480, w21481, w21482, w21483, w21484, w21485, w21486, w21487, w21488, w21489, w21490, w21491, w21492, w21493, w21494, w21495, w21496, w21497, w21498, w21499, w21500, w21501, w21502, w21503, w21504, w21505, w21506, w21507, w21508, w21509, w21510, w21511, w21512, w21513, w21514, w21515, w21516, w21517, w21518, w21519, w21520, w21521, w21522, w21523, w21524, w21525, w21526, w21527, w21528, w21529, w21530, w21531, w21532, w21533, w21534, w21535, w21536, w21537, w21538, w21539, w21540, w21541, w21542, w21543, w21544, w21545, w21546, w21547, w21548, w21549, w21550, w21551, w21552, w21553, w21554, w21555, w21556, w21557, w21558, w21559, w21560, w21561, w21562, w21563, w21564, w21565, w21566, w21567, w21568, w21569, w21570, w21571, w21572, w21573, w21574, w21575, w21576, w21577, w21578, w21579, w21580, w21581, w21582, w21583, w21584, w21585, w21586, w21587, w21588, w21589, w21590, w21591, w21592, w21593, w21594, w21595, w21596, w21597, w21598, w21599, w21600, w21601, w21602, w21603, w21604, w21605, w21606, w21607, w21608, w21609, w21610, w21611, w21612, w21613, w21614, w21615, w21616, w21617, w21618, w21619, w21620, w21621, w21622, w21623, w21624, w21625, w21626, w21627, w21628, w21629, w21630, w21631, w21632, w21633, w21634, w21635, w21636, w21637, w21638, w21639, w21640, w21641, w21642, w21643, w21644, w21645, w21646, w21647, w21648, w21649, w21650, w21651, w21652, w21653, w21654, w21655, w21656, w21657, w21658, w21659, w21660, w21661, w21662, w21663, w21664, w21665, w21666, w21667, w21668, w21669, w21670, w21671, w21672, w21673, w21674, w21675, w21676, w21677, w21678, w21679, w21680, w21681, w21682, w21683, w21684, w21685, w21686, w21687, w21688, w21689, w21690, w21691, w21692, w21693, w21694, w21695, w21696, w21697, w21698, w21699, w21700, w21701, w21702, w21703, w21704, w21705, w21706, w21707, w21708, w21709, w21710, w21711, w21712, w21713, w21714, w21715, w21716, w21717, w21718, w21719, w21720, w21721, w21722, w21723, w21724, w21725, w21726, w21727, w21728, w21729, w21730, w21731, w21732, w21733, w21734, w21735, w21736, w21737, w21738, w21739, w21740, w21741, w21742, w21743, w21744, w21745, w21746, w21747, w21748, w21749, w21750, w21751, w21752, w21753, w21754, w21755, w21756, w21757, w21758, w21759, w21760, w21761, w21762, w21763, w21764, w21765, w21766, w21767, w21768, w21769, w21770, w21771, w21772, w21773, w21774, w21775, w21776, w21777, w21778, w21779, w21780, w21781, w21782, w21783, w21784, w21785, w21786, w21787, w21788, w21789, w21790, w21791, w21792, w21793, w21794, w21795, w21796, w21797, w21798, w21799, w21800, w21801, w21802, w21803, w21804, w21805, w21806, w21807, w21808, w21809, w21810, w21811, w21812, w21813, w21814, w21815, w21816, w21817, w21818, w21819, w21820, w21821, w21822, w21823, w21824, w21825, w21826, w21827, w21828, w21829, w21830, w21831, w21832, w21833, w21834, w21835, w21836, w21837, w21838, w21839, w21840, w21841, w21842, w21843, w21844, w21845, w21846, w21847, w21848, w21849, w21850, w21851, w21852, w21853, w21854, w21855, w21856, w21857, w21858, w21859, w21860, w21861, w21862, w21863, w21864, w21865, w21866, w21867, w21868, w21869, w21870, w21871, w21872, w21873, w21874, w21875, w21876, w21877, w21878, w21879, w21880, w21881, w21882, w21883, w21884, w21885, w21886, w21887, w21888, w21889, w21890, w21891, w21892, w21893, w21894, w21895, w21896, w21897, w21898, w21899, w21900, w21901, w21902, w21903, w21904, w21905, w21906, w21907, w21908, w21909, w21910, w21911, w21912, w21913, w21914, w21915, w21916, w21917, w21918, w21919, w21920, w21921, w21922, w21923, w21924, w21925, w21926, w21927, w21928, w21929, w21930, w21931, w21932, w21933, w21934, w21935, w21936, w21937, w21938, w21939, w21940, w21941, w21942, w21943, w21944, w21945, w21946, w21947, w21948, w21949, w21950, w21951, w21952, w21953, w21954, w21955, w21956, w21957, w21958, w21959, w21960, w21961, w21962, w21963, w21964, w21965, w21966, w21967, w21968, w21969, w21970, w21971, w21972, w21973, w21974, w21975, w21976, w21977, w21978, w21979, w21980, w21981, w21982, w21983, w21984, w21985, w21986, w21987, w21988, w21989, w21990, w21991, w21992, w21993, w21994, w21995, w21996, w21997, w21998, w21999, w22000, w22001, w22002, w22003, w22004, w22005, w22006, w22007, w22008, w22009, w22010, w22011, w22012, w22013, w22014, w22015, w22016, w22017, w22018, w22019, w22020, w22021, w22022, w22023, w22024, w22025, w22026, w22027, w22028, w22029, w22030, w22031, w22032, w22033, w22034, w22035, w22036, w22037, w22038, w22039, w22040, w22041, w22042, w22043, w22044, w22045, w22046, w22047, w22048, w22049, w22050, w22051, w22052, w22053, w22054, w22055, w22056, w22057, w22058, w22059, w22060, w22061, w22062, w22063, w22064, w22065, w22066, w22067, w22068, w22069, w22070, w22071, w22072, w22073, w22074, w22075, w22076, w22077, w22078, w22079, w22080, w22081, w22082, w22083, w22084, w22085, w22086, w22087, w22088, w22089, w22090, w22091, w22092, w22093, w22094, w22095, w22096, w22097, w22098, w22099, w22100, w22101, w22102, w22103, w22104, w22105, w22106, w22107, w22108, w22109, w22110, w22111, w22112, w22113, w22114, w22115, w22116, w22117, w22118, w22119, w22120, w22121, w22122, w22123, w22124, w22125, w22126, w22127, w22128, w22129, w22130, w22131, w22132, w22133, w22134, w22135, w22136, w22137, w22138, w22139, w22140, w22141, w22142, w22143, w22144, w22145, w22146, w22147, w22148, w22149, w22150, w22151, w22152, w22153, w22154, w22155, w22156, w22157, w22158, w22159, w22160, w22161, w22162, w22163, w22164, w22165, w22166, w22167, w22168, w22169, w22170, w22171, w22172, w22173, w22174, w22175, w22176, w22177, w22178, w22179, w22180, w22181, w22182, w22183, w22184, w22185, w22186, w22187, w22188, w22189, w22190, w22191, w22192, w22193, w22194, w22195, w22196, w22197, w22198, w22199, w22200, w22201, w22202, w22203, w22204, w22205, w22206, w22207, w22208, w22209, w22210, w22211, w22212, w22213, w22214, w22215, w22216, w22217, w22218, w22219, w22220, w22221, w22222, w22223, w22224, w22225, w22226, w22227, w22228, w22229, w22230, w22231, w22232, w22233, w22234, w22235, w22236, w22237, w22238, w22239, w22240, w22241, w22242, w22243, w22244, w22245, w22246, w22247, w22248, w22249, w22250, w22251, w22252, w22253, w22254, w22255, w22256, w22257, w22258, w22259, w22260, w22261, w22262, w22263, w22264, w22265, w22266, w22267, w22268, w22269, w22270, w22271, w22272, w22273, w22274, w22275, w22276, w22277, w22278, w22279, w22280, w22281, w22282, w22283, w22284, w22285, w22286, w22287, w22288, w22289, w22290, w22291, w22292, w22293, w22294, w22295, w22296, w22297, w22298, w22299, w22300, w22301, w22302, w22303, w22304, w22305, w22306, w22307, w22308, w22309, w22310, w22311, w22312, w22313, w22314, w22315, w22316, w22317, w22318, w22319, w22320, w22321, w22322, w22323, w22324, w22325, w22326, w22327, w22328, w22329, w22330, w22331, w22332, w22333, w22334, w22335, w22336, w22337, w22338, w22339, w22340, w22341, w22342, w22343, w22344, w22345, w22346, w22347, w22348, w22349, w22350, w22351, w22352, w22353, w22354, w22355, w22356, w22357, w22358, w22359, w22360, w22361, w22362, w22363, w22364, w22365, w22366, w22367, w22368, w22369, w22370, w22371, w22372, w22373, w22374, w22375, w22376, w22377, w22378, w22379, w22380, w22381, w22382, w22383, w22384, w22385, w22386, w22387, w22388, w22389, w22390, w22391, w22392, w22393, w22394, w22395, w22396, w22397, w22398, w22399, w22400, w22401, w22402, w22403, w22404, w22405, w22406, w22407, w22408, w22409, w22410, w22411, w22412, w22413, w22414, w22415, w22416, w22417, w22418, w22419, w22420, w22421, w22422, w22423, w22424, w22425, w22426, w22427, w22428, w22429, w22430, w22431, w22432, w22433, w22434, w22435, w22436, w22437, w22438, w22439, w22440, w22441, w22442, w22443, w22444, w22445, w22446, w22447, w22448, w22449, w22450, w22451, w22452, w22453, w22454, w22455, w22456, w22457, w22458, w22459, w22460, w22461, w22462, w22463, w22464, w22465, w22466, w22467, w22468, w22469, w22470, w22471, w22472, w22473, w22474, w22475, w22476, w22477, w22478, w22479, w22480, w22481, w22482, w22483, w22484, w22485, w22486, w22487, w22488, w22489, w22490, w22491, w22492, w22493, w22494, w22495, w22496, w22497, w22498, w22499, w22500, w22501, w22502, w22503, w22504, w22505, w22506, w22507, w22508, w22509, w22510, w22511, w22512, w22513, w22514, w22515, w22516, w22517, w22518, w22519, w22520, w22521, w22522, w22523, w22524, w22525, w22526, w22527, w22528, w22529, w22530, w22531, w22532, w22533, w22534, w22535, w22536, w22537, w22538, w22539, w22540, w22541, w22542, w22543, w22544, w22545, w22546, w22547, w22548, w22549, w22550, w22551, w22552, w22553, w22554, w22555, w22556, w22557, w22558, w22559, w22560, w22561, w22562, w22563, w22564, w22565, w22566, w22567, w22568, w22569, w22570, w22571, w22572, w22573, w22574, w22575, w22576, w22577, w22578, w22579, w22580, w22581, w22582, w22583, w22584, w22585, w22586, w22587, w22588, w22589, w22590, w22591, w22592, w22593, w22594, w22595, w22596, w22597, w22598, w22599, w22600, w22601, w22602, w22603, w22604, w22605, w22606, w22607, w22608, w22609, w22610, w22611, w22612, w22613, w22614, w22615, w22616, w22617, w22618, w22619, w22620, w22621, w22622, w22623, w22624, w22625, w22626, w22627, w22628, w22629, w22630, w22631, w22632, w22633, w22634, w22635, w22636, w22637, w22638, w22639, w22640, w22641, w22642, w22643, w22644, w22645, w22646, w22647, w22648, w22649, w22650, w22651, w22652, w22653, w22654, w22655, w22656, w22657, w22658, w22659, w22660, w22661, w22662, w22663, w22664, w22665, w22666, w22667, w22668, w22669, w22670, w22671, w22672, w22673, w22674, w22675, w22676, w22677, w22678, w22679, w22680, w22681, w22682, w22683, w22684, w22685, w22686, w22687, w22688, w22689, w22690, w22691, w22692, w22693, w22694, w22695, w22696, w22697, w22698, w22699, w22700, w22701, w22702, w22703, w22704, w22705, w22706, w22707, w22708, w22709, w22710, w22711, w22712, w22713, w22714, w22715, w22716, w22717, w22718, w22719, w22720, w22721, w22722, w22723, w22724, w22725, w22726, w22727, w22728, w22729, w22730, w22731, w22732, w22733, w22734, w22735, w22736, w22737, w22738, w22739, w22740, w22741, w22742, w22743, w22744, w22745, w22746, w22747, w22748, w22749, w22750, w22751, w22752, w22753, w22754, w22755, w22756, w22757, w22758, w22759, w22760, w22761, w22762, w22763, w22764, w22765, w22766, w22767, w22768, w22769, w22770, w22771, w22772, w22773, w22774, w22775, w22776, w22777, w22778, w22779, w22780, w22781, w22782, w22783, w22784, w22785, w22786, w22787, w22788, w22789, w22790, w22791, w22792, w22793, w22794, w22795, w22796, w22797, w22798, w22799, w22800, w22801, w22802, w22803, w22804, w22805, w22806, w22807, w22808, w22809, w22810, w22811, w22812, w22813, w22814, w22815, w22816, w22817, w22818, w22819, w22820, w22821, w22822, w22823, w22824, w22825, w22826, w22827, w22828, w22829, w22830, w22831, w22832, w22833, w22834, w22835, w22836, w22837, w22838, w22839, w22840, w22841, w22842, w22843, w22844, w22845, w22846, w22847, w22848, w22849, w22850, w22851, w22852, w22853, w22854, w22855, w22856, w22857, w22858, w22859, w22860, w22861, w22862, w22863, w22864, w22865, w22866, w22867, w22868, w22869, w22870, w22871, w22872, w22873, w22874, w22875, w22876, w22877, w22878, w22879, w22880, w22881, w22882, w22883, w22884, w22885, w22886, w22887, w22888, w22889, w22890, w22891, w22892, w22893, w22894, w22895, w22896, w22897, w22898, w22899, w22900, w22901, w22902, w22903, w22904, w22905, w22906, w22907, w22908, w22909, w22910, w22911, w22912, w22913, w22914, w22915, w22916, w22917, w22918, w22919, w22920, w22921, w22922, w22923, w22924, w22925, w22926, w22927, w22928, w22929, w22930, w22931, w22932, w22933, w22934, w22935, w22936, w22937, w22938, w22939, w22940, w22941, w22942, w22943, w22944, w22945, w22946, w22947, w22948, w22949, w22950, w22951, w22952, w22953, w22954, w22955, w22956, w22957, w22958, w22959, w22960, w22961, w22962, w22963, w22964, w22965, w22966, w22967, w22968, w22969, w22970, w22971, w22972, w22973, w22974, w22975, w22976, w22977, w22978, w22979, w22980, w22981, w22982, w22983, w22984, w22985, w22986, w22987, w22988, w22989, w22990, w22991, w22992, w22993, w22994, w22995, w22996, w22997, w22998, w22999, w23000, w23001, w23002, w23003, w23004, w23005, w23006, w23007, w23008, w23009, w23010, w23011, w23012, w23013, w23014, w23015, w23016, w23017, w23018, w23019, w23020, w23021, w23022, w23023, w23024, w23025, w23026, w23027, w23028, w23029, w23030, w23031, w23032, w23033, w23034, w23035, w23036, w23037, w23038, w23039, w23040, w23041, w23042, w23043, w23044, w23045, w23046, w23047, w23048, w23049, w23050, w23051, w23052, w23053, w23054, w23055, w23056, w23057, w23058, w23059, w23060, w23061, w23062, w23063, w23064, w23065, w23066, w23067, w23068, w23069, w23070, w23071, w23072, w23073, w23074, w23075, w23076, w23077, w23078, w23079, w23080, w23081, w23082, w23083, w23084, w23085, w23086, w23087, w23088, w23089, w23090, w23091, w23092, w23093, w23094, w23095, w23096, w23097, w23098, w23099, w23100, w23101, w23102, w23103, w23104, w23105, w23106, w23107, w23108, w23109, w23110, w23111, w23112, w23113, w23114, w23115, w23116, w23117, w23118, w23119, w23120, w23121, w23122, w23123, w23124, w23125, w23126, w23127, w23128, w23129, w23130, w23131, w23132, w23133, w23134, w23135, w23136, w23137, w23138, w23139, w23140, w23141, w23142, w23143, w23144, w23145, w23146, w23147, w23148, w23149, w23150, w23151, w23152, w23153, w23154, w23155, w23156, w23157, w23158, w23159, w23160, w23161, w23162, w23163, w23164, w23165, w23166, w23167, w23168, w23169, w23170, w23171, w23172, w23173, w23174, w23175, w23176, w23177, w23178, w23179, w23180, w23181, w23182, w23183, w23184, w23185, w23186, w23187, w23188, w23189, w23190, w23191, w23192, w23193, w23194, w23195, w23196, w23197, w23198, w23199, w23200, w23201, w23202, w23203, w23204, w23205, w23206, w23207, w23208, w23209, w23210, w23211, w23212, w23213, w23214, w23215, w23216, w23217, w23218, w23219, w23220, w23221, w23222, w23223, w23224, w23225, w23226, w23227, w23228, w23229, w23230, w23231, w23232, w23233, w23234, w23235, w23236, w23237, w23238, w23239, w23240, w23241, w23242, w23243, w23244, w23245, w23246, w23247, w23248, w23249, w23250, w23251, w23252, w23253, w23254, w23255, w23256, w23257, w23258, w23259, w23260, w23261, w23262, w23263, w23264, w23265, w23266, w23267, w23268, w23269, w23270, w23271, w23272, w23273, w23274, w23275, w23276, w23277, w23278, w23279, w23280, w23281, w23282, w23283, w23284, w23285, w23286, w23287, w23288, w23289, w23290, w23291, w23292, w23293, w23294, w23295, w23296, w23297, w23298, w23299, w23300, w23301, w23302, w23303, w23304, w23305, w23306, w23307, w23308, w23309, w23310, w23311, w23312, w23313, w23314, w23315, w23316, w23317, w23318, w23319, w23320, w23321, w23322, w23323, w23324, w23325, w23326, w23327, w23328, w23329, w23330, w23331, w23332, w23333, w23334, w23335, w23336, w23337, w23338, w23339, w23340, w23341, w23342, w23343, w23344, w23345, w23346, w23347, w23348, w23349, w23350, w23351, w23352, w23353, w23354, w23355, w23356, w23357, w23358, w23359, w23360, w23361, w23362, w23363, w23364, w23365, w23366, w23367, w23368, w23369, w23370, w23371, w23372, w23373, w23374, w23375, w23376, w23377, w23378, w23379, w23380, w23381, w23382, w23383, w23384, w23385, w23386, w23387, w23388, w23389, w23390, w23391, w23392, w23393, w23394, w23395, w23396, w23397, w23398, w23399, w23400, w23401, w23402, w23403, w23404, w23405, w23406, w23407, w23408, w23409, w23410, w23411, w23412, w23413, w23414, w23415, w23416, w23417, w23418, w23419, w23420, w23421, w23422, w23423, w23424, w23425, w23426, w23427, w23428, w23429, w23430, w23431, w23432, w23433, w23434, w23435, w23436, w23437, w23438, w23439, w23440, w23441, w23442, w23443, w23444, w23445, w23446, w23447, w23448, w23449, w23450, w23451, w23452, w23453, w23454, w23455, w23456, w23457, w23458, w23459, w23460, w23461, w23462, w23463, w23464, w23465, w23466, w23467, w23468, w23469, w23470, w23471, w23472, w23473, w23474, w23475, w23476, w23477, w23478, w23479, w23480, w23481, w23482, w23483, w23484, w23485, w23486, w23487, w23488, w23489, w23490, w23491, w23492, w23493, w23494, w23495, w23496, w23497, w23498, w23499, w23500, w23501, w23502, w23503, w23504, w23505, w23506, w23507, w23508, w23509, w23510, w23511, w23512, w23513, w23514, w23515, w23516, w23517, w23518, w23519, w23520, w23521, w23522, w23523, w23524, w23525, w23526, w23527, w23528, w23529, w23530, w23531, w23532, w23533, w23534, w23535, w23536, w23537, w23538, w23539, w23540, w23541, w23542, w23543, w23544, w23545, w23546, w23547, w23548, w23549, w23550, w23551, w23552, w23553, w23554, w23555, w23556, w23557, w23558, w23559, w23560, w23561, w23562, w23563, w23564, w23565, w23566, w23567, w23568, w23569, w23570, w23571, w23572, w23573, w23574, w23575, w23576, w23577, w23578, w23579, w23580, w23581, w23582, w23583, w23584, w23585, w23586, w23587, w23588, w23589, w23590, w23591, w23592, w23593, w23594, w23595, w23596, w23597, w23598, w23599, w23600, w23601, w23602, w23603, w23604, w23605, w23606, w23607, w23608, w23609, w23610, w23611, w23612, w23613, w23614, w23615, w23616, w23617, w23618, w23619, w23620, w23621, w23622, w23623, w23624, w23625, w23626, w23627, w23628, w23629, w23630, w23631, w23632, w23633, w23634, w23635, w23636, w23637, w23638, w23639, w23640, w23641, w23642, w23643, w23644, w23645, w23646, w23647, w23648, w23649, w23650, w23651, w23652, w23653, w23654, w23655, w23656, w23657, w23658, w23659, w23660, w23661, w23662, w23663, w23664, w23665, w23666, w23667, w23668, w23669, w23670, w23671, w23672, w23673, w23674, w23675, w23676, w23677, w23678, w23679, w23680, w23681, w23682, w23683, w23684, w23685, w23686, w23687, w23688, w23689, w23690, w23691, w23692, w23693, w23694, w23695, w23696, w23697, w23698, w23699, w23700, w23701, w23702, w23703, w23704, w23705, w23706, w23707, w23708, w23709, w23710, w23711, w23712, w23713, w23714, w23715, w23716, w23717, w23718, w23719, w23720, w23721, w23722, w23723, w23724, w23725, w23726, w23727, w23728, w23729, w23730, w23731, w23732, w23733, w23734, w23735, w23736, w23737, w23738, w23739, w23740, w23741, w23742, w23743, w23744, w23745, w23746, w23747, w23748, w23749, w23750, w23751, w23752, w23753, w23754, w23755, w23756, w23757, w23758, w23759, w23760, w23761, w23762, w23763, w23764, w23765, w23766, w23767, w23768, w23769, w23770, w23771, w23772, w23773, w23774, w23775, w23776, w23777, w23778, w23779, w23780, w23781, w23782, w23783, w23784, w23785, w23786, w23787, w23788, w23789, w23790, w23791, w23792, w23793, w23794, w23795, w23796, w23797, w23798, w23799, w23800, w23801, w23802, w23803, w23804, w23805, w23806, w23807, w23808, w23809, w23810, w23811, w23812, w23813, w23814, w23815, w23816, w23817, w23818, w23819, w23820, w23821, w23822, w23823, w23824, w23825, w23826, w23827, w23828, w23829, w23830, w23831, w23832, w23833, w23834, w23835, w23836, w23837, w23838, w23839, w23840, w23841, w23842, w23843, w23844, w23845, w23846, w23847, w23848, w23849, w23850, w23851, w23852, w23853, w23854, w23855, w23856, w23857, w23858, w23859, w23860, w23861, w23862, w23863, w23864, w23865, w23866, w23867, w23868, w23869, w23870, w23871, w23872, w23873, w23874, w23875, w23876, w23877, w23878, w23879, w23880, w23881, w23882, w23883, w23884, w23885, w23886, w23887, w23888, w23889, w23890, w23891, w23892, w23893, w23894, w23895, w23896, w23897, w23898, w23899, w23900, w23901, w23902, w23903, w23904, w23905, w23906, w23907, w23908, w23909, w23910, w23911, w23912, w23913, w23914, w23915, w23916, w23917, w23918, w23919, w23920, w23921, w23922, w23923, w23924, w23925, w23926, w23927, w23928, w23929, w23930, w23931, w23932, w23933, w23934, w23935, w23936, w23937, w23938, w23939, w23940, w23941, w23942, w23943, w23944, w23945, w23946, w23947, w23948, w23949, w23950, w23951, w23952, w23953, w23954, w23955, w23956, w23957, w23958, w23959, w23960, w23961, w23962, w23963, w23964, w23965, w23966, w23967, w23968, w23969, w23970, w23971, w23972, w23973, w23974, w23975, w23976, w23977, w23978, w23979, w23980, w23981, w23982, w23983, w23984, w23985, w23986, w23987, w23988, w23989, w23990, w23991, w23992, w23993, w23994, w23995, w23996, w23997, w23998, w23999, w24000, w24001, w24002, w24003, w24004, w24005, w24006, w24007, w24008, w24009, w24010, w24011, w24012, w24013, w24014, w24015, w24016, w24017, w24018, w24019, w24020, w24021, w24022, w24023, w24024, w24025, w24026, w24027, w24028, w24029, w24030, w24031, w24032, w24033, w24034, w24035, w24036, w24037, w24038, w24039, w24040, w24041, w24042, w24043, w24044, w24045, w24046, w24047, w24048, w24049, w24050, w24051, w24052, w24053, w24054, w24055, w24056, w24057, w24058, w24059, w24060, w24061, w24062, w24063, w24064, w24065, w24066, w24067, w24068, w24069, w24070, w24071, w24072, w24073, w24074, w24075, w24076, w24077, w24078, w24079, w24080, w24081, w24082, w24083, w24084, w24085, w24086, w24087, w24088, w24089, w24090, w24091, w24092, w24093, w24094, w24095, w24096, w24097, w24098, w24099, w24100, w24101, w24102, w24103, w24104, w24105, w24106, w24107, w24108, w24109, w24110, w24111, w24112, w24113, w24114, w24115, w24116, w24117, w24118, w24119, w24120, w24121, w24122, w24123, w24124, w24125, w24126, w24127, w24128, w24129, w24130, w24131, w24132, w24133, w24134, w24135, w24136, w24137, w24138, w24139, w24140, w24141, w24142, w24143, w24144, w24145, w24146, w24147, w24148, w24149, w24150, w24151, w24152, w24153, w24154, w24155, w24156, w24157, w24158, w24159, w24160, w24161, w24162, w24163, w24164, w24165, w24166, w24167, w24168, w24169, w24170, w24171, w24172, w24173, w24174, w24175, w24176, w24177, w24178, w24179, w24180, w24181, w24182, w24183, w24184, w24185, w24186, w24187, w24188, w24189, w24190, w24191, w24192, w24193, w24194, w24195, w24196, w24197, w24198, w24199, w24200, w24201, w24202, w24203, w24204, w24205, w24206, w24207, w24208, w24209, w24210, w24211, w24212, w24213, w24214, w24215, w24216, w24217, w24218, w24219, w24220, w24221, w24222, w24223, w24224, w24225, w24226, w24227, w24228, w24229, w24230, w24231, w24232, w24233, w24234, w24235, w24236, w24237, w24238, w24239, w24240, w24241, w24242, w24243, w24244, w24245, w24246, w24247, w24248, w24249, w24250, w24251, w24252, w24253, w24254, w24255, w24256, w24257, w24258, w24259, w24260, w24261, w24262, w24263, w24264, w24265, w24266, w24267, w24268, w24269, w24270, w24271, w24272, w24273, w24274, w24275, w24276, w24277, w24278, w24279, w24280, w24281, w24282, w24283, w24284, w24285, w24286, w24287, w24288, w24289, w24290, w24291, w24292, w24293, w24294, w24295, w24296, w24297, w24298, w24299, w24300, w24301, w24302, w24303, w24304, w24305, w24306, w24307, w24308, w24309, w24310, w24311, w24312, w24313, w24314, w24315, w24316, w24317, w24318, w24319, w24320, w24321, w24322, w24323, w24324, w24325, w24326, w24327, w24328, w24329, w24330, w24331, w24332, w24333, w24334, w24335, w24336, w24337, w24338, w24339, w24340, w24341, w24342, w24343, w24344, w24345, w24346, w24347, w24348, w24349, w24350, w24351, w24352, w24353, w24354, w24355, w24356, w24357, w24358, w24359, w24360, w24361, w24362, w24363, w24364, w24365, w24366, w24367, w24368, w24369, w24370, w24371, w24372, w24373, w24374, w24375, w24376, w24377, w24378, w24379, w24380, w24381, w24382, w24383, w24384, w24385, w24386, w24387, w24388, w24389, w24390, w24391, w24392, w24393, w24394, w24395, w24396, w24397, w24398, w24399, w24400, w24401, w24402, w24403, w24404, w24405, w24406, w24407, w24408, w24409, w24410, w24411, w24412, w24413, w24414, w24415, w24416, w24417, w24418, w24419, w24420, w24421, w24422, w24423, w24424, w24425, w24426, w24427, w24428, w24429, w24430, w24431, w24432, w24433, w24434, w24435, w24436, w24437, w24438, w24439, w24440, w24441, w24442, w24443, w24444, w24445, w24446, w24447, w24448, w24449, w24450, w24451, w24452, w24453, w24454, w24455, w24456, w24457, w24458, w24459, w24460, w24461, w24462, w24463, w24464, w24465, w24466, w24467, w24468, w24469, w24470, w24471, w24472, w24473, w24474, w24475, w24476, w24477, w24478, w24479, w24480, w24481, w24482, w24483, w24484, w24485, w24486, w24487, w24488, w24489, w24490, w24491, w24492, w24493, w24494, w24495, w24496, w24497, w24498, w24499, w24500, w24501, w24502, w24503, w24504, w24505, w24506, w24507, w24508, w24509, w24510, w24511, w24512, w24513, w24514, w24515, w24516, w24517, w24518, w24519, w24520, w24521, w24522, w24523, w24524, w24525, w24526, w24527, w24528, w24529, w24530, w24531, w24532, w24533, w24534, w24535, w24536, w24537, w24538, w24539, w24540, w24541, w24542, w24543, w24544, w24545, w24546, w24547, w24548, w24549, w24550, w24551, w24552, w24553, w24554, w24555, w24556, w24557, w24558, w24559, w24560, w24561, w24562, w24563, w24564, w24565, w24566, w24567, w24568, w24569, w24570, w24571, w24572, w24573, w24574, w24575, w24576, w24577, w24578, w24579, w24580, w24581, w24582, w24583, w24584, w24585, w24586, w24587, w24588, w24589, w24590, w24591, w24592, w24593, w24594, w24595, w24596, w24597, w24598, w24599, w24600, w24601, w24602, w24603, w24604, w24605, w24606, w24607, w24608, w24609, w24610, w24611, w24612, w24613, w24614, w24615, w24616, w24617, w24618, w24619, w24620, w24621, w24622, w24623, w24624, w24625, w24626, w24627, w24628, w24629, w24630, w24631, w24632, w24633, w24634, w24635, w24636, w24637, w24638, w24639, w24640, w24641, w24642, w24643, w24644, w24645, w24646, w24647, w24648, w24649, w24650, w24651, w24652, w24653, w24654, w24655, w24656, w24657, w24658, w24659, w24660, w24661, w24662, w24663, w24664, w24665, w24666, w24667, w24668, w24669, w24670, w24671, w24672, w24673, w24674, w24675, w24676, w24677, w24678, w24679, w24680, w24681, w24682, w24683, w24684, w24685, w24686, w24687, w24688, w24689, w24690, w24691, w24692, w24693, w24694, w24695, w24696, w24697, w24698, w24699, w24700, w24701, w24702, w24703, w24704, w24705, w24706, w24707, w24708, w24709, w24710, w24711, w24712, w24713, w24714, w24715, w24716, w24717, w24718, w24719, w24720, w24721, w24722, w24723, w24724, w24725, w24726, w24727, w24728, w24729, w24730, w24731, w24732, w24733, w24734, w24735, w24736, w24737, w24738, w24739, w24740, w24741, w24742, w24743, w24744, w24745, w24746, w24747, w24748, w24749, w24750, w24751, w24752, w24753, w24754, w24755, w24756, w24757, w24758, w24759, w24760, w24761, w24762, w24763, w24764, w24765, w24766, w24767, w24768, w24769, w24770, w24771, w24772, w24773, w24774, w24775, w24776, w24777, w24778, w24779, w24780, w24781, w24782, w24783, w24784, w24785, w24786, w24787, w24788, w24789, w24790, w24791, w24792, w24793, w24794, w24795, w24796, w24797, w24798, w24799, w24800, w24801, w24802, w24803, w24804, w24805, w24806, w24807, w24808, w24809, w24810, w24811, w24812, w24813, w24814, w24815, w24816, w24817, w24818, w24819, w24820, w24821, w24822, w24823, w24824, w24825, w24826, w24827, w24828, w24829, w24830, w24831, w24832, w24833, w24834, w24835, w24836, w24837, w24838, w24839, w24840, w24841, w24842, w24843, w24844, w24845, w24846, w24847, w24848, w24849, w24850, w24851, w24852, w24853, w24854, w24855, w24856, w24857, w24858, w24859, w24860, w24861, w24862, w24863, w24864, w24865, w24866, w24867, w24868, w24869, w24870, w24871, w24872, w24873, w24874, w24875, w24876, w24877, w24878, w24879, w24880, w24881, w24882, w24883, w24884, w24885, w24886, w24887, w24888, w24889, w24890, w24891, w24892, w24893, w24894, w24895, w24896, w24897, w24898, w24899, w24900, w24901, w24902, w24903, w24904, w24905, w24906, w24907, w24908, w24909, w24910, w24911, w24912, w24913, w24914, w24915, w24916, w24917, w24918, w24919, w24920, w24921, w24922, w24923, w24924, w24925, w24926, w24927, w24928, w24929, w24930, w24931, w24932, w24933, w24934, w24935, w24936, w24937, w24938, w24939, w24940, w24941, w24942, w24943, w24944, w24945, w24946, w24947, w24948, w24949, w24950, w24951, w24952, w24953, w24954, w24955, w24956, w24957, w24958, w24959, w24960, w24961, w24962, w24963, w24964, w24965, w24966, w24967, w24968, w24969, w24970, w24971, w24972, w24973, w24974, w24975, w24976, w24977, w24978, w24979, w24980, w24981, w24982, w24983, w24984, w24985, w24986, w24987, w24988, w24989, w24990, w24991, w24992, w24993, w24994, w24995, w24996, w24997, w24998, w24999, w25000, w25001, w25002, w25003, w25004, w25005, w25006, w25007, w25008, w25009, w25010, w25011, w25012, w25013, w25014, w25015, w25016, w25017, w25018, w25019, w25020, w25021, w25022, w25023, w25024, w25025, w25026, w25027, w25028, w25029, w25030, w25031, w25032, w25033, w25034, w25035, w25036, w25037, w25038, w25039, w25040, w25041, w25042, w25043, w25044, w25045, w25046, w25047, w25048, w25049, w25050, w25051, w25052, w25053, w25054, w25055, w25056, w25057, w25058, w25059, w25060, w25061, w25062, w25063, w25064, w25065, w25066, w25067, w25068, w25069, w25070, w25071, w25072, w25073, w25074, w25075, w25076, w25077, w25078, w25079, w25080, w25081, w25082, w25083, w25084, w25085, w25086, w25087, w25088, w25089, w25090, w25091, w25092, w25093, w25094, w25095, w25096, w25097, w25098, w25099, w25100, w25101, w25102, w25103, w25104, w25105, w25106, w25107, w25108, w25109, w25110, w25111, w25112, w25113, w25114, w25115, w25116, w25117, w25118, w25119, w25120, w25121, w25122, w25123, w25124, w25125, w25126, w25127, w25128, w25129, w25130, w25131, w25132, w25133, w25134, w25135, w25136, w25137, w25138, w25139, w25140, w25141, w25142, w25143, w25144, w25145, w25146, w25147, w25148, w25149, w25150, w25151, w25152, w25153, w25154, w25155, w25156, w25157, w25158, w25159, w25160, w25161, w25162, w25163, w25164, w25165, w25166, w25167, w25168, w25169, w25170, w25171, w25172, w25173, w25174, w25175, w25176, w25177, w25178, w25179, w25180, w25181, w25182, w25183, w25184, w25185, w25186, w25187, w25188, w25189, w25190, w25191, w25192, w25193, w25194, w25195, w25196, w25197, w25198, w25199, w25200, w25201, w25202, w25203, w25204, w25205, w25206, w25207, w25208, w25209, w25210, w25211, w25212, w25213, w25214, w25215, w25216, w25217, w25218, w25219, w25220, w25221, w25222, w25223, w25224, w25225, w25226, w25227, w25228, w25229, w25230, w25231, w25232, w25233, w25234, w25235, w25236, w25237, w25238, w25239, w25240, w25241, w25242, w25243, w25244, w25245, w25246, w25247, w25248, w25249, w25250, w25251, w25252, w25253, w25254, w25255, w25256, w25257, w25258, w25259, w25260, w25261, w25262, w25263, w25264, w25265, w25266, w25267, w25268, w25269, w25270, w25271, w25272, w25273, w25274, w25275, w25276, w25277, w25278, w25279, w25280, w25281, w25282, w25283, w25284, w25285, w25286, w25287, w25288, w25289, w25290, w25291, w25292, w25293, w25294, w25295, w25296, w25297, w25298, w25299, w25300, w25301, w25302, w25303, w25304, w25305, w25306, w25307, w25308, w25309, w25310, w25311, w25312, w25313, w25314, w25315, w25316, w25317, w25318, w25319, w25320, w25321, w25322, w25323, w25324, w25325, w25326, w25327, w25328, w25329, w25330, w25331, w25332, w25333, w25334, w25335, w25336, w25337, w25338, w25339, w25340, w25341, w25342, w25343, w25344, w25345, w25346, w25347, w25348, w25349, w25350, w25351, w25352, w25353, w25354, w25355, w25356, w25357, w25358, w25359, w25360, w25361, w25362, w25363, w25364, w25365, w25366, w25367, w25368, w25369, w25370, w25371, w25372, w25373, w25374, w25375, w25376, w25377, w25378, w25379, w25380, w25381, w25382, w25383, w25384, w25385, w25386, w25387, w25388, w25389, w25390, w25391, w25392, w25393, w25394, w25395, w25396, w25397, w25398, w25399, w25400, w25401, w25402, w25403, w25404, w25405, w25406, w25407, w25408, w25409, w25410, w25411, w25412, w25413, w25414, w25415, w25416, w25417, w25418, w25419, w25420, w25421, w25422, w25423, w25424, w25425, w25426, w25427, w25428, w25429, w25430, w25431, w25432, w25433, w25434, w25435, w25436, w25437, w25438, w25439, w25440, w25441, w25442, w25443, w25444, w25445, w25446, w25447, w25448, w25449, w25450, w25451, w25452, w25453, w25454, w25455, w25456, w25457, w25458, w25459, w25460, w25461, w25462, w25463, w25464, w25465, w25466, w25467, w25468, w25469, w25470, w25471, w25472, w25473, w25474, w25475, w25476, w25477, w25478, w25479, w25480, w25481, w25482, w25483, w25484, w25485, w25486, w25487, w25488, w25489, w25490, w25491, w25492, w25493, w25494, w25495, w25496, w25497, w25498, w25499, w25500, w25501, w25502, w25503, w25504, w25505, w25506, w25507, w25508, w25509, w25510, w25511, w25512, w25513, w25514, w25515, w25516, w25517, w25518, w25519, w25520, w25521, w25522, w25523, w25524, w25525, w25526, w25527, w25528, w25529, w25530, w25531, w25532, w25533, w25534, w25535, w25536, w25537, w25538, w25539, w25540, w25541, w25542, w25543, w25544, w25545, w25546, w25547, w25548, w25549, w25550, w25551, w25552, w25553, w25554, w25555, w25556, w25557, w25558, w25559, w25560, w25561, w25562, w25563, w25564, w25565, w25566, w25567, w25568, w25569, w25570, w25571, w25572, w25573, w25574, w25575, w25576, w25577, w25578, w25579, w25580, w25581, w25582, w25583, w25584, w25585, w25586, w25587, w25588, w25589, w25590, w25591, w25592, w25593, w25594, w25595, w25596, w25597, w25598, w25599, w25600, w25601, w25602, w25603, w25604, w25605, w25606, w25607, w25608, w25609, w25610, w25611, w25612, w25613, w25614, w25615, w25616, w25617, w25618, w25619, w25620, w25621, w25622, w25623, w25624, w25625, w25626, w25627, w25628, w25629, w25630, w25631, w25632, w25633, w25634, w25635, w25636, w25637, w25638, w25639, w25640, w25641, w25642, w25643, w25644, w25645, w25646, w25647, w25648, w25649, w25650, w25651, w25652, w25653, w25654, w25655, w25656, w25657, w25658, w25659, w25660, w25661, w25662, w25663, w25664, w25665, w25666, w25667, w25668, w25669, w25670, w25671, w25672, w25673, w25674, w25675, w25676, w25677, w25678, w25679, w25680, w25681, w25682, w25683, w25684, w25685, w25686, w25687, w25688, w25689, w25690, w25691, w25692, w25693, w25694, w25695, w25696, w25697, w25698, w25699, w25700, w25701, w25702, w25703, w25704, w25705, w25706, w25707, w25708, w25709, w25710, w25711, w25712, w25713, w25714, w25715, w25716, w25717, w25718, w25719, w25720, w25721, w25722, w25723, w25724, w25725, w25726, w25727, w25728, w25729, w25730, w25731, w25732, w25733, w25734, w25735, w25736, w25737, w25738, w25739, w25740, w25741, w25742, w25743, w25744, w25745, w25746, w25747, w25748, w25749, w25750, w25751, w25752, w25753, w25754, w25755, w25756, w25757, w25758, w25759, w25760, w25761, w25762, w25763, w25764, w25765, w25766, w25767, w25768, w25769, w25770, w25771, w25772, w25773, w25774, w25775, w25776, w25777, w25778, w25779, w25780, w25781, w25782, w25783, w25784, w25785, w25786, w25787, w25788, w25789, w25790, w25791, w25792, w25793, w25794, w25795, w25796, w25797, w25798, w25799, w25800, w25801, w25802, w25803, w25804, w25805, w25806, w25807, w25808, w25809, w25810, w25811, w25812, w25813, w25814, w25815, w25816, w25817, w25818, w25819, w25820, w25821, w25822, w25823, w25824, w25825, w25826, w25827, w25828, w25829, w25830, w25831, w25832, w25833, w25834, w25835, w25836, w25837, w25838, w25839, w25840, w25841, w25842, w25843, w25844, w25845, w25846, w25847, w25848, w25849, w25850, w25851, w25852, w25853, w25854, w25855, w25856, w25857, w25858, w25859, w25860, w25861, w25862, w25863, w25864, w25865, w25866, w25867, w25868, w25869, w25870, w25871, w25872, w25873, w25874, w25875, w25876, w25877, w25878, w25879, w25880, w25881, w25882, w25883, w25884, w25885, w25886, w25887, w25888, w25889, w25890, w25891, w25892, w25893, w25894, w25895, w25896, w25897, w25898, w25899, w25900, w25901, w25902, w25903, w25904, w25905, w25906, w25907, w25908, w25909, w25910, w25911, w25912, w25913, w25914, w25915, w25916, w25917, w25918, w25919, w25920, w25921, w25922, w25923, w25924, w25925, w25926, w25927, w25928, w25929, w25930, w25931, w25932, w25933, w25934, w25935, w25936, w25937, w25938, w25939, w25940, w25941, w25942, w25943, w25944, w25945, w25946, w25947, w25948, w25949, w25950, w25951, w25952, w25953, w25954, w25955, w25956, w25957, w25958, w25959, w25960, w25961, w25962, w25963, w25964, w25965, w25966, w25967, w25968, w25969, w25970, w25971, w25972, w25973, w25974, w25975, w25976, w25977, w25978, w25979, w25980, w25981, w25982, w25983, w25984, w25985, w25986, w25987, w25988, w25989, w25990, w25991, w25992, w25993, w25994, w25995, w25996, w25997, w25998, w25999, w26000, w26001, w26002, w26003, w26004, w26005, w26006, w26007, w26008, w26009, w26010, w26011, w26012, w26013, w26014, w26015, w26016, w26017, w26018, w26019, w26020, w26021, w26022, w26023, w26024, w26025, w26026, w26027, w26028, w26029, w26030, w26031, w26032, w26033, w26034, w26035, w26036, w26037, w26038, w26039, w26040, w26041, w26042, w26043, w26044, w26045, w26046, w26047, w26048, w26049, w26050, w26051, w26052, w26053, w26054, w26055, w26056, w26057, w26058, w26059, w26060, w26061, w26062, w26063, w26064, w26065, w26066, w26067, w26068, w26069, w26070, w26071, w26072, w26073, w26074, w26075, w26076, w26077, w26078, w26079, w26080, w26081, w26082, w26083, w26084, w26085, w26086, w26087, w26088, w26089, w26090, w26091, w26092, w26093, w26094, w26095, w26096, w26097, w26098, w26099, w26100, w26101, w26102, w26103, w26104, w26105, w26106, w26107, w26108, w26109, w26110, w26111, w26112, w26113, w26114, w26115, w26116, w26117, w26118, w26119, w26120, w26121, w26122, w26123, w26124, w26125, w26126, w26127, w26128, w26129, w26130, w26131, w26132, w26133, w26134, w26135, w26136, w26137, w26138, w26139, w26140, w26141, w26142, w26143, w26144, w26145, w26146, w26147, w26148, w26149, w26150, w26151, w26152, w26153, w26154, w26155, w26156, w26157, w26158, w26159, w26160, w26161, w26162, w26163, w26164, w26165, w26166, w26167, w26168, w26169, w26170, w26171, w26172, w26173, w26174, w26175, w26176, w26177, w26178, w26179, w26180, w26181, w26182, w26183, w26184, w26185, w26186, w26187, w26188, w26189, w26190, w26191, w26192, w26193, w26194, w26195, w26196, w26197, w26198, w26199, w26200, w26201, w26202, w26203, w26204, w26205, w26206, w26207, w26208, w26209, w26210, w26211, w26212, w26213, w26214, w26215, w26216, w26217, w26218, w26219, w26220, w26221, w26222, w26223, w26224, w26225, w26226, w26227, w26228, w26229, w26230, w26231, w26232, w26233, w26234, w26235, w26236, w26237, w26238, w26239, w26240, w26241, w26242, w26243, w26244, w26245, w26246, w26247, w26248, w26249, w26250, w26251, w26252, w26253, w26254, w26255, w26256, w26257, w26258, w26259, w26260, w26261, w26262, w26263, w26264, w26265, w26266, w26267, w26268, w26269, w26270, w26271, w26272, w26273, w26274, w26275, w26276, w26277, w26278, w26279, w26280, w26281, w26282, w26283, w26284, w26285, w26286, w26287, w26288, w26289, w26290, w26291, w26292, w26293, w26294, w26295, w26296, w26297, w26298, w26299, w26300, w26301, w26302, w26303, w26304, w26305, w26306, w26307, w26308, w26309, w26310, w26311, w26312, w26313, w26314, w26315, w26316, w26317, w26318, w26319, w26320, w26321, w26322, w26323, w26324, w26325, w26326, w26327, w26328, w26329, w26330, w26331, w26332, w26333, w26334, w26335, w26336, w26337, w26338, w26339, w26340, w26341, w26342, w26343, w26344, w26345, w26346, w26347, w26348, w26349, w26350, w26351, w26352, w26353, w26354, w26355, w26356, w26357, w26358, w26359, w26360, w26361, w26362, w26363, w26364, w26365, w26366, w26367, w26368, w26369, w26370, w26371, w26372, w26373, w26374, w26375, w26376, w26377, w26378, w26379, w26380, w26381, w26382, w26383, w26384, w26385, w26386, w26387, w26388, w26389, w26390, w26391, w26392, w26393, w26394, w26395, w26396, w26397, w26398, w26399, w26400, w26401, w26402, w26403, w26404, w26405, w26406, w26407, w26408, w26409, w26410, w26411, w26412, w26413, w26414, w26415, w26416, w26417, w26418, w26419, w26420, w26421, w26422, w26423, w26424, w26425, w26426, w26427, w26428, w26429, w26430, w26431, w26432, w26433, w26434, w26435, w26436, w26437, w26438, w26439, w26440, w26441, w26442, w26443, w26444, w26445, w26446, w26447, w26448, w26449, w26450, w26451, w26452, w26453, w26454, w26455, w26456, w26457, w26458, w26459, w26460, w26461, w26462, w26463, w26464, w26465, w26466, w26467, w26468, w26469, w26470, w26471, w26472, w26473, w26474, w26475, w26476, w26477, w26478, w26479, w26480, w26481, w26482, w26483, w26484, w26485, w26486, w26487, w26488, w26489, w26490, w26491, w26492, w26493, w26494, w26495, w26496, w26497, w26498, w26499, w26500, w26501, w26502, w26503, w26504, w26505, w26506, w26507, w26508, w26509, w26510, w26511, w26512, w26513, w26514, w26515, w26516, w26517, w26518, w26519, w26520, w26521, w26522, w26523, w26524, w26525, w26526, w26527, w26528, w26529, w26530, w26531, w26532, w26533, w26534, w26535, w26536, w26537, w26538, w26539, w26540, w26541, w26542, w26543, w26544, w26545, w26546, w26547, w26548, w26549, w26550, w26551, w26552, w26553, w26554, w26555, w26556, w26557, w26558, w26559, w26560, w26561, w26562, w26563, w26564, w26565, w26566, w26567, w26568, w26569, w26570, w26571, w26572, w26573, w26574, w26575, w26576, w26577, w26578, w26579, w26580, w26581, w26582, w26583, w26584, w26585, w26586, w26587, w26588, w26589, w26590, w26591, w26592, w26593, w26594, w26595, w26596, w26597, w26598, w26599, w26600, w26601, w26602, w26603, w26604, w26605, w26606, w26607, w26608, w26609, w26610, w26611, w26612, w26613, w26614, w26615, w26616, w26617, w26618, w26619, w26620, w26621, w26622, w26623, w26624, w26625, w26626, w26627, w26628, w26629, w26630, w26631, w26632, w26633, w26634, w26635, w26636, w26637, w26638, w26639, w26640, w26641, w26642, w26643, w26644, w26645, w26646, w26647, w26648, w26649, w26650, w26651, w26652, w26653, w26654, w26655, w26656, w26657, w26658, w26659, w26660, w26661, w26662, w26663, w26664, w26665, w26666, w26667, w26668, w26669, w26670, w26671, w26672, w26673, w26674, w26675, w26676, w26677, w26678, w26679, w26680, w26681, w26682, w26683, w26684, w26685, w26686, w26687, w26688, w26689, w26690, w26691, w26692, w26693, w26694, w26695, w26696, w26697, w26698, w26699, w26700, w26701, w26702, w26703, w26704, w26705, w26706, w26707, w26708, w26709, w26710, w26711, w26712, w26713, w26714, w26715, w26716, w26717, w26718, w26719, w26720, w26721, w26722, w26723, w26724, w26725, w26726, w26727, w26728, w26729, w26730, w26731, w26732, w26733, w26734, w26735, w26736, w26737, w26738, w26739, w26740, w26741, w26742, w26743, w26744, w26745, w26746, w26747, w26748, w26749, w26750, w26751, w26752, w26753, w26754, w26755, w26756, w26757, w26758, w26759, w26760, w26761, w26762, w26763, w26764, w26765, w26766, w26767, w26768, w26769, w26770, w26771, w26772, w26773, w26774, w26775, w26776, w26777, w26778, w26779, w26780, w26781, w26782, w26783, w26784, w26785, w26786, w26787, w26788, w26789, w26790, w26791, w26792, w26793, w26794, w26795, w26796, w26797, w26798, w26799, w26800, w26801, w26802, w26803, w26804, w26805, w26806, w26807, w26808, w26809, w26810, w26811, w26812, w26813, w26814, w26815, w26816, w26817, w26818, w26819, w26820, w26821, w26822, w26823, w26824, w26825, w26826, w26827, w26828, w26829, w26830, w26831, w26832, w26833, w26834, w26835, w26836, w26837, w26838, w26839, w26840, w26841, w26842, w26843, w26844, w26845, w26846, w26847, w26848, w26849, w26850, w26851, w26852, w26853, w26854, w26855, w26856, w26857, w26858, w26859, w26860, w26861, w26862, w26863, w26864, w26865, w26866, w26867, w26868, w26869, w26870, w26871, w26872, w26873, w26874, w26875, w26876, w26877, w26878, w26879, w26880, w26881, w26882, w26883, w26884, w26885, w26886, w26887, w26888, w26889, w26890, w26891, w26892, w26893, w26894, w26895, w26896, w26897, w26898, w26899, w26900, w26901, w26902, w26903, w26904, w26905, w26906, w26907, w26908, w26909, w26910, w26911, w26912, w26913, w26914, w26915, w26916, w26917, w26918, w26919, w26920, w26921, w26922, w26923, w26924, w26925, w26926, w26927, w26928, w26929, w26930, w26931, w26932, w26933, w26934, w26935, w26936, w26937, w26938, w26939, w26940, w26941, w26942, w26943, w26944, w26945, w26946, w26947, w26948, w26949, w26950, w26951, w26952, w26953, w26954, w26955, w26956, w26957, w26958, w26959, w26960, w26961, w26962, w26963, w26964, w26965, w26966, w26967, w26968, w26969, w26970, w26971, w26972, w26973, w26974, w26975, w26976, w26977, w26978, w26979, w26980, w26981, w26982, w26983, w26984, w26985, w26986, w26987, w26988, w26989, w26990, w26991, w26992, w26993, w26994, w26995, w26996, w26997, w26998, w26999, w27000, w27001, w27002, w27003, w27004, w27005, w27006, w27007, w27008, w27009, w27010, w27011, w27012, w27013, w27014, w27015, w27016, w27017, w27018, w27019, w27020, w27021, w27022, w27023, w27024, w27025, w27026, w27027, w27028, w27029, w27030, w27031, w27032, w27033, w27034, w27035, w27036, w27037, w27038, w27039, w27040, w27041, w27042, w27043, w27044, w27045, w27046, w27047, w27048, w27049, w27050, w27051, w27052, w27053, w27054, w27055, w27056, w27057, w27058, w27059, w27060, w27061, w27062, w27063, w27064, w27065, w27066, w27067, w27068, w27069, w27070, w27071, w27072, w27073, w27074, w27075, w27076, w27077, w27078, w27079, w27080, w27081, w27082, w27083, w27084, w27085, w27086, w27087, w27088, w27089, w27090, w27091, w27092, w27093, w27094, w27095, w27096, w27097, w27098, w27099, w27100, w27101, w27102, w27103, w27104, w27105, w27106, w27107, w27108, w27109, w27110, w27111, w27112, w27113, w27114, w27115, w27116, w27117, w27118, w27119, w27120, w27121, w27122, w27123, w27124, w27125, w27126, w27127, w27128, w27129, w27130, w27131, w27132, w27133, w27134, w27135, w27136, w27137, w27138, w27139, w27140, w27141, w27142, w27143, w27144, w27145, w27146, w27147, w27148, w27149, w27150, w27151, w27152, w27153, w27154, w27155, w27156, w27157, w27158, w27159, w27160, w27161, w27162, w27163, w27164, w27165, w27166, w27167, w27168, w27169, w27170, w27171, w27172, w27173, w27174, w27175, w27176, w27177, w27178, w27179, w27180, w27181, w27182, w27183, w27184, w27185, w27186, w27187, w27188, w27189, w27190, w27191, w27192, w27193, w27194, w27195, w27196, w27197, w27198, w27199, w27200, w27201, w27202, w27203, w27204, w27205, w27206, w27207, w27208, w27209, w27210, w27211, w27212, w27213, w27214, w27215, w27216, w27217, w27218, w27219, w27220, w27221, w27222, w27223, w27224, w27225, w27226, w27227, w27228, w27229, w27230, w27231, w27232, w27233, w27234, w27235, w27236, w27237, w27238, w27239, w27240, w27241, w27242, w27243, w27244, w27245, w27246, w27247, w27248, w27249, w27250, w27251, w27252, w27253, w27254, w27255, w27256, w27257, w27258, w27259, w27260, w27261, w27262, w27263, w27264, w27265, w27266, w27267, w27268, w27269, w27270, w27271, w27272, w27273, w27274, w27275, w27276, w27277, w27278, w27279, w27280, w27281, w27282, w27283, w27284, w27285, w27286, w27287, w27288, w27289, w27290, w27291, w27292, w27293, w27294, w27295, w27296, w27297, w27298, w27299, w27300, w27301, w27302, w27303, w27304, w27305, w27306, w27307, w27308, w27309, w27310, w27311, w27312, w27313, w27314, w27315, w27316, w27317, w27318, w27319, w27320, w27321, w27322, w27323, w27324, w27325, w27326, w27327, w27328, w27329, w27330, w27331, w27332, w27333, w27334, w27335, w27336, w27337, w27338, w27339, w27340, w27341, w27342, w27343, w27344, w27345, w27346, w27347, w27348, w27349, w27350, w27351, w27352, w27353, w27354, w27355, w27356, w27357, w27358, w27359, w27360, w27361, w27362, w27363, w27364, w27365, w27366, w27367, w27368, w27369, w27370, w27371, w27372, w27373, w27374, w27375, w27376, w27377, w27378, w27379, w27380, w27381, w27382, w27383, w27384, w27385, w27386, w27387, w27388, w27389, w27390, w27391, w27392, w27393, w27394, w27395, w27396, w27397, w27398, w27399, w27400, w27401, w27402, w27403, w27404, w27405, w27406, w27407, w27408, w27409, w27410, w27411, w27412, w27413, w27414, w27415, w27416, w27417, w27418, w27419, w27420, w27421, w27422, w27423, w27424, w27425, w27426, w27427, w27428, w27429, w27430, w27431, w27432, w27433, w27434, w27435, w27436, w27437, w27438, w27439, w27440, w27441, w27442, w27443, w27444, w27445, w27446, w27447, w27448, w27449, w27450, w27451, w27452, w27453, w27454, w27455, w27456, w27457, w27458, w27459, w27460, w27461, w27462, w27463, w27464, w27465, w27466, w27467, w27468, w27469, w27470, w27471, w27472, w27473, w27474, w27475, w27476, w27477, w27478, w27479, w27480, w27481, w27482, w27483, w27484, w27485, w27486, w27487, w27488, w27489, w27490, w27491, w27492, w27493, w27494, w27495, w27496, w27497, w27498, w27499, w27500, w27501, w27502, w27503, w27504, w27505, w27506, w27507, w27508, w27509, w27510, w27511, w27512, w27513, w27514, w27515, w27516, w27517, w27518, w27519, w27520, w27521, w27522, w27523, w27524, w27525, w27526, w27527, w27528, w27529, w27530, w27531, w27532, w27533, w27534, w27535, w27536, w27537, w27538, w27539, w27540, w27541, w27542, w27543, w27544, w27545, w27546, w27547, w27548, w27549, w27550, w27551, w27552, w27553, w27554, w27555, w27556, w27557, w27558, w27559, w27560, w27561, w27562, w27563, w27564, w27565, w27566, w27567, w27568, w27569, w27570, w27571, w27572, w27573, w27574, w27575, w27576, w27577, w27578, w27579, w27580, w27581, w27582, w27583, w27584, w27585, w27586, w27587, w27588, w27589, w27590, w27591, w27592, w27593, w27594, w27595, w27596, w27597, w27598, w27599, w27600, w27601, w27602, w27603, w27604, w27605, w27606, w27607, w27608, w27609, w27610, w27611, w27612, w27613, w27614, w27615, w27616, w27617, w27618, w27619, w27620, w27621, w27622, w27623, w27624, w27625, w27626, w27627, w27628, w27629, w27630, w27631, w27632, w27633, w27634, w27635, w27636, w27637, w27638, w27639, w27640, w27641, w27642, w27643, w27644, w27645, w27646, w27647, w27648, w27649, w27650, w27651, w27652, w27653, w27654, w27655, w27656, w27657, w27658, w27659, w27660, w27661, w27662, w27663, w27664, w27665, w27666, w27667, w27668, w27669, w27670, w27671, w27672, w27673, w27674, w27675, w27676, w27677, w27678, w27679, w27680, w27681, w27682, w27683, w27684, w27685, w27686, w27687, w27688, w27689, w27690, w27691, w27692, w27693, w27694, w27695, w27696, w27697, w27698, w27699, w27700, w27701, w27702, w27703, w27704, w27705, w27706, w27707, w27708, w27709, w27710, w27711, w27712, w27713, w27714, w27715, w27716, w27717, w27718, w27719, w27720, w27721, w27722, w27723, w27724, w27725, w27726, w27727, w27728, w27729, w27730, w27731, w27732, w27733, w27734, w27735, w27736, w27737, w27738, w27739, w27740, w27741, w27742, w27743, w27744, w27745, w27746, w27747, w27748, w27749, w27750, w27751, w27752, w27753, w27754, w27755, w27756, w27757, w27758, w27759, w27760, w27761, w27762, w27763, w27764, w27765, w27766, w27767, w27768, w27769, w27770, w27771, w27772, w27773, w27774, w27775, w27776, w27777, w27778, w27779, w27780, w27781, w27782, w27783, w27784, w27785, w27786, w27787, w27788, w27789, w27790, w27791, w27792, w27793, w27794, w27795, w27796, w27797, w27798, w27799, w27800, w27801, w27802, w27803, w27804, w27805, w27806, w27807, w27808, w27809, w27810, w27811, w27812, w27813, w27814, w27815, w27816, w27817, w27818, w27819, w27820, w27821, w27822, w27823, w27824, w27825, w27826, w27827, w27828, w27829, w27830, w27831, w27832, w27833, w27834, w27835, w27836, w27837, w27838, w27839, w27840, w27841, w27842, w27843, w27844, w27845, w27846, w27847, w27848, w27849, w27850, w27851, w27852, w27853, w27854, w27855, w27856, w27857, w27858, w27859, w27860, w27861, w27862, w27863, w27864, w27865, w27866, w27867, w27868, w27869, w27870, w27871, w27872, w27873, w27874, w27875, w27876, w27877, w27878, w27879, w27880, w27881, w27882, w27883, w27884, w27885, w27886, w27887, w27888, w27889, w27890, w27891, w27892, w27893, w27894, w27895, w27896, w27897, w27898, w27899, w27900, w27901, w27902, w27903, w27904, w27905, w27906, w27907, w27908, w27909, w27910, w27911, w27912, w27913, w27914, w27915, w27916, w27917, w27918, w27919, w27920, w27921, w27922, w27923, w27924, w27925, w27926, w27927, w27928, w27929, w27930, w27931, w27932, w27933, w27934, w27935, w27936, w27937, w27938, w27939, w27940, w27941, w27942, w27943, w27944, w27945, w27946, w27947, w27948, w27949, w27950, w27951, w27952, w27953, w27954, w27955, w27956, w27957, w27958, w27959, w27960, w27961, w27962, w27963, w27964, w27965, w27966, w27967, w27968, w27969, w27970, w27971, w27972, w27973, w27974, w27975, w27976, w27977, w27978, w27979, w27980, w27981, w27982, w27983, w27984, w27985, w27986, w27987, w27988, w27989, w27990, w27991, w27992, w27993, w27994, w27995, w27996, w27997, w27998, w27999, w28000, w28001, w28002, w28003, w28004, w28005, w28006, w28007, w28008, w28009, w28010, w28011, w28012, w28013, w28014, w28015, w28016, w28017, w28018, w28019, w28020, w28021, w28022, w28023, w28024, w28025, w28026, w28027, w28028, w28029, w28030, w28031, w28032, w28033, w28034, w28035, w28036, w28037, w28038, w28039, w28040, w28041, w28042, w28043, w28044, w28045, w28046, w28047, w28048, w28049, w28050, w28051, w28052, w28053, w28054, w28055, w28056, w28057, w28058, w28059, w28060, w28061, w28062, w28063, w28064, w28065, w28066, w28067, w28068, w28069, w28070, w28071, w28072, w28073, w28074, w28075, w28076, w28077, w28078, w28079, w28080, w28081, w28082, w28083, w28084, w28085, w28086, w28087, w28088, w28089, w28090, w28091, w28092, w28093, w28094, w28095, w28096, w28097, w28098, w28099, w28100, w28101, w28102, w28103, w28104, w28105, w28106, w28107, w28108, w28109, w28110, w28111, w28112, w28113, w28114, w28115, w28116, w28117, w28118, w28119, w28120, w28121, w28122, w28123, w28124, w28125, w28126, w28127, w28128, w28129, w28130, w28131, w28132, w28133, w28134, w28135, w28136, w28137, w28138, w28139, w28140, w28141, w28142, w28143, w28144, w28145, w28146, w28147, w28148, w28149, w28150, w28151, w28152, w28153, w28154, w28155, w28156, w28157, w28158, w28159, w28160, w28161, w28162, w28163, w28164, w28165, w28166, w28167, w28168, w28169, w28170, w28171, w28172, w28173, w28174, w28175, w28176, w28177, w28178, w28179, w28180, w28181, w28182, w28183, w28184, w28185, w28186, w28187, w28188, w28189, w28190, w28191, w28192, w28193, w28194, w28195, w28196, w28197, w28198, w28199, w28200, w28201, w28202, w28203, w28204, w28205, w28206, w28207, w28208, w28209, w28210, w28211, w28212, w28213, w28214, w28215, w28216, w28217, w28218, w28219, w28220, w28221, w28222, w28223, w28224, w28225, w28226, w28227, w28228, w28229, w28230, w28231, w28232, w28233, w28234, w28235, w28236, w28237, w28238, w28239, w28240, w28241, w28242, w28243, w28244, w28245, w28246, w28247, w28248, w28249, w28250, w28251, w28252, w28253, w28254, w28255, w28256, w28257, w28258, w28259, w28260, w28261, w28262, w28263, w28264, w28265, w28266, w28267, w28268, w28269, w28270, w28271, w28272, w28273, w28274, w28275, w28276, w28277, w28278, w28279, w28280, w28281, w28282, w28283, w28284, w28285, w28286, w28287, w28288, w28289, w28290, w28291, w28292, w28293, w28294, w28295, w28296, w28297, w28298, w28299, w28300, w28301, w28302, w28303, w28304, w28305, w28306, w28307, w28308, w28309, w28310, w28311, w28312, w28313, w28314, w28315, w28316, w28317, w28318, w28319, w28320, w28321, w28322, w28323, w28324, w28325, w28326, w28327, w28328, w28329, w28330, w28331, w28332, w28333, w28334, w28335, w28336, w28337, w28338, w28339, w28340, w28341, w28342, w28343, w28344, w28345, w28346, w28347, w28348, w28349, w28350, w28351, w28352, w28353, w28354, w28355, w28356, w28357, w28358, w28359, w28360, w28361, w28362, w28363, w28364, w28365, w28366, w28367, w28368, w28369, w28370, w28371, w28372, w28373, w28374, w28375, w28376, w28377, w28378, w28379, w28380, w28381, w28382, w28383, w28384, w28385, w28386, w28387, w28388, w28389, w28390, w28391, w28392, w28393, w28394, w28395, w28396, w28397, w28398, w28399, w28400, w28401, w28402, w28403, w28404, w28405, w28406, w28407, w28408, w28409, w28410, w28411, w28412, w28413, w28414, w28415, w28416, w28417, w28418, w28419, w28420, w28421, w28422, w28423, w28424, w28425, w28426, w28427, w28428, w28429, w28430, w28431, w28432, w28433, w28434, w28435, w28436, w28437, w28438, w28439, w28440, w28441, w28442, w28443, w28444, w28445, w28446, w28447, w28448, w28449, w28450, w28451, w28452, w28453, w28454, w28455, w28456, w28457, w28458, w28459, w28460, w28461, w28462, w28463, w28464, w28465, w28466, w28467, w28468, w28469, w28470, w28471, w28472, w28473, w28474, w28475, w28476, w28477, w28478, w28479, w28480, w28481, w28482, w28483, w28484, w28485, w28486, w28487, w28488, w28489, w28490, w28491, w28492, w28493, w28494, w28495, w28496, w28497, w28498, w28499, w28500, w28501, w28502, w28503, w28504, w28505, w28506, w28507, w28508, w28509, w28510, w28511, w28512, w28513, w28514, w28515, w28516, w28517, w28518, w28519, w28520, w28521, w28522, w28523, w28524, w28525, w28526, w28527, w28528, w28529, w28530, w28531, w28532, w28533, w28534, w28535, w28536, w28537, w28538, w28539, w28540, w28541, w28542, w28543, w28544, w28545, w28546, w28547, w28548, w28549, w28550, w28551, w28552, w28553, w28554, w28555, w28556, w28557, w28558, w28559, w28560, w28561, w28562, w28563, w28564, w28565, w28566, w28567, w28568, w28569, w28570, w28571, w28572, w28573, w28574, w28575, w28576, w28577, w28578, w28579, w28580, w28581, w28582, w28583, w28584, w28585, w28586, w28587, w28588, w28589, w28590, w28591, w28592, w28593, w28594, w28595, w28596, w28597, w28598, w28599, w28600, w28601, w28602, w28603, w28604, w28605, w28606, w28607, w28608, w28609, w28610, w28611, w28612, w28613, w28614, w28615, w28616, w28617, w28618, w28619, w28620, w28621, w28622, w28623, w28624, w28625, w28626, w28627, w28628, w28629, w28630, w28631, w28632, w28633, w28634, w28635, w28636, w28637, w28638, w28639, w28640, w28641, w28642, w28643, w28644, w28645, w28646, w28647, w28648, w28649, w28650, w28651, w28652, w28653, w28654, w28655, w28656, w28657, w28658, w28659, w28660, w28661, w28662, w28663, w28664, w28665, w28666, w28667, w28668, w28669, w28670, w28671, w28672, w28673, w28674, w28675, w28676, w28677, w28678, w28679, w28680, w28681, w28682, w28683, w28684, w28685, w28686, w28687, w28688, w28689, w28690, w28691, w28692, w28693, w28694, w28695, w28696, w28697, w28698, w28699, w28700, w28701, w28702, w28703, w28704, w28705, w28706, w28707, w28708, w28709, w28710, w28711, w28712, w28713, w28714, w28715, w28716, w28717, w28718, w28719, w28720, w28721, w28722, w28723, w28724, w28725, w28726, w28727, w28728, w28729, w28730, w28731, w28732, w28733, w28734, w28735, w28736, w28737, w28738, w28739, w28740, w28741, w28742, w28743, w28744, w28745, w28746, w28747, w28748, w28749, w28750, w28751, w28752, w28753, w28754, w28755, w28756, w28757, w28758, w28759, w28760, w28761, w28762, w28763, w28764, w28765, w28766, w28767, w28768, w28769, w28770, w28771, w28772, w28773, w28774, w28775, w28776, w28777, w28778, w28779, w28780, w28781, w28782, w28783, w28784, w28785, w28786, w28787, w28788, w28789, w28790, w28791, w28792, w28793, w28794, w28795, w28796, w28797, w28798, w28799, w28800, w28801, w28802, w28803, w28804, w28805, w28806, w28807, w28808, w28809, w28810, w28811, w28812, w28813, w28814, w28815, w28816, w28817, w28818, w28819, w28820, w28821, w28822, w28823, w28824, w28825, w28826, w28827, w28828, w28829, w28830, w28831, w28832, w28833, w28834, w28835, w28836, w28837, w28838, w28839, w28840, w28841, w28842, w28843, w28844, w28845, w28846, w28847, w28848, w28849, w28850, w28851, w28852, w28853, w28854, w28855, w28856, w28857, w28858, w28859, w28860, w28861, w28862, w28863, w28864, w28865, w28866, w28867, w28868, w28869, w28870, w28871, w28872, w28873, w28874, w28875, w28876, w28877, w28878, w28879, w28880, w28881, w28882, w28883, w28884, w28885, w28886, w28887, w28888, w28889, w28890, w28891, w28892, w28893, w28894, w28895, w28896, w28897, w28898, w28899, w28900, w28901, w28902, w28903, w28904, w28905, w28906, w28907, w28908, w28909, w28910, w28911, w28912, w28913, w28914, w28915, w28916, w28917, w28918, w28919, w28920, w28921, w28922, w28923, w28924, w28925, w28926, w28927, w28928, w28929, w28930, w28931, w28932, w28933, w28934, w28935, w28936, w28937, w28938, w28939, w28940, w28941, w28942, w28943, w28944, w28945, w28946, w28947, w28948, w28949, w28950, w28951, w28952, w28953, w28954, w28955, w28956, w28957, w28958, w28959, w28960, w28961, w28962, w28963, w28964, w28965, w28966, w28967, w28968, w28969, w28970, w28971, w28972, w28973, w28974, w28975, w28976, w28977, w28978, w28979, w28980, w28981, w28982, w28983, w28984, w28985, w28986, w28987, w28988, w28989, w28990, w28991, w28992, w28993, w28994, w28995, w28996, w28997, w28998, w28999, w29000, w29001, w29002, w29003, w29004, w29005, w29006, w29007, w29008, w29009, w29010, w29011, w29012, w29013, w29014, w29015, w29016, w29017, w29018, w29019, w29020, w29021, w29022, w29023, w29024, w29025, w29026, w29027, w29028, w29029, w29030, w29031, w29032, w29033, w29034, w29035, w29036, w29037, w29038, w29039, w29040, w29041, w29042, w29043, w29044, w29045, w29046, w29047, w29048, w29049, w29050, w29051, w29052, w29053, w29054, w29055, w29056, w29057, w29058, w29059, w29060, w29061, w29062, w29063, w29064, w29065, w29066, w29067, w29068, w29069, w29070, w29071, w29072, w29073, w29074, w29075, w29076, w29077, w29078, w29079, w29080, w29081, w29082, w29083, w29084, w29085, w29086, w29087, w29088, w29089, w29090, w29091, w29092, w29093, w29094, w29095, w29096, w29097, w29098, w29099, w29100, w29101, w29102, w29103, w29104, w29105, w29106, w29107, w29108, w29109, w29110, w29111, w29112, w29113, w29114, w29115, w29116, w29117, w29118, w29119, w29120, w29121, w29122, w29123, w29124, w29125, w29126, w29127, w29128, w29129, w29130, w29131, w29132, w29133, w29134, w29135, w29136, w29137, w29138, w29139, w29140, w29141, w29142, w29143, w29144, w29145, w29146, w29147, w29148, w29149, w29150, w29151, w29152, w29153, w29154, w29155, w29156, w29157, w29158, w29159, w29160, w29161, w29162, w29163, w29164, w29165, w29166, w29167, w29168, w29169, w29170, w29171, w29172, w29173, w29174, w29175, w29176, w29177, w29178, w29179, w29180, w29181, w29182, w29183, w29184, w29185, w29186, w29187, w29188, w29189, w29190, w29191, w29192, w29193, w29194, w29195, w29196, w29197, w29198, w29199, w29200, w29201, w29202, w29203, w29204, w29205, w29206, w29207, w29208, w29209, w29210, w29211, w29212, w29213, w29214, w29215, w29216, w29217, w29218, w29219, w29220, w29221, w29222, w29223, w29224, w29225, w29226, w29227, w29228, w29229, w29230, w29231, w29232, w29233, w29234, w29235, w29236, w29237, w29238, w29239, w29240, w29241, w29242, w29243, w29244, w29245, w29246, w29247, w29248, w29249, w29250, w29251, w29252, w29253, w29254, w29255, w29256, w29257, w29258, w29259, w29260, w29261, w29262, w29263, w29264, w29265, w29266, w29267, w29268, w29269, w29270, w29271, w29272, w29273, w29274, w29275, w29276, w29277, w29278, w29279, w29280, w29281, w29282, w29283, w29284, w29285, w29286, w29287, w29288, w29289, w29290, w29291, w29292, w29293, w29294, w29295, w29296, w29297, w29298, w29299, w29300, w29301, w29302, w29303, w29304, w29305, w29306, w29307, w29308, w29309, w29310, w29311, w29312, w29313, w29314, w29315, w29316, w29317, w29318, w29319, w29320, w29321, w29322, w29323, w29324, w29325, w29326, w29327, w29328, w29329, w29330, w29331, w29332, w29333, w29334, w29335, w29336, w29337, w29338, w29339, w29340, w29341, w29342, w29343, w29344, w29345, w29346, w29347, w29348, w29349, w29350, w29351, w29352, w29353, w29354, w29355, w29356, w29357, w29358, w29359, w29360, w29361, w29362, w29363, w29364, w29365, w29366, w29367, w29368, w29369, w29370, w29371, w29372, w29373, w29374, w29375, w29376, w29377, w29378, w29379, w29380, w29381, w29382, w29383, w29384, w29385, w29386, w29387, w29388, w29389, w29390, w29391, w29392, w29393, w29394, w29395, w29396, w29397, w29398, w29399, w29400, w29401, w29402, w29403, w29404, w29405, w29406, w29407, w29408, w29409, w29410, w29411, w29412, w29413, w29414, w29415, w29416, w29417, w29418, w29419, w29420, w29421, w29422, w29423, w29424, w29425, w29426, w29427, w29428, w29429, w29430, w29431, w29432, w29433, w29434, w29435, w29436, w29437, w29438, w29439, w29440, w29441, w29442, w29443, w29444, w29445, w29446, w29447, w29448, w29449, w29450, w29451, w29452, w29453, w29454, w29455, w29456, w29457, w29458, w29459, w29460, w29461, w29462, w29463, w29464, w29465, w29466, w29467, w29468, w29469, w29470, w29471, w29472, w29473, w29474, w29475, w29476, w29477, w29478, w29479, w29480, w29481, w29482, w29483, w29484, w29485, w29486, w29487, w29488, w29489, w29490, w29491, w29492, w29493, w29494, w29495, w29496, w29497, w29498, w29499, w29500, w29501, w29502, w29503, w29504, w29505, w29506, w29507, w29508, w29509, w29510, w29511, w29512, w29513, w29514, w29515, w29516, w29517, w29518, w29519, w29520, w29521, w29522, w29523, w29524, w29525, w29526, w29527, w29528, w29529, w29530, w29531, w29532, w29533, w29534, w29535, w29536, w29537, w29538, w29539, w29540, w29541, w29542, w29543, w29544, w29545, w29546, w29547, w29548, w29549, w29550, w29551, w29552, w29553, w29554, w29555, w29556, w29557, w29558, w29559, w29560, w29561, w29562, w29563, w29564, w29565, w29566, w29567, w29568, w29569, w29570, w29571, w29572, w29573, w29574, w29575, w29576, w29577, w29578, w29579, w29580, w29581, w29582, w29583, w29584, w29585, w29586, w29587, w29588, w29589, w29590, w29591, w29592, w29593, w29594, w29595, w29596, w29597, w29598, w29599, w29600, w29601, w29602, w29603, w29604, w29605, w29606, w29607, w29608, w29609, w29610, w29611, w29612, w29613, w29614, w29615, w29616, w29617, w29618, w29619, w29620, w29621, w29622, w29623, w29624, w29625, w29626, w29627, w29628, w29629, w29630, w29631, w29632, w29633, w29634, w29635, w29636, w29637, w29638, w29639, w29640, w29641, w29642, w29643, w29644, w29645, w29646, w29647, w29648, w29649, w29650, w29651, w29652, w29653, w29654, w29655, w29656, w29657, w29658, w29659, w29660, w29661, w29662, w29663, w29664, w29665, w29666, w29667, w29668, w29669, w29670, w29671, w29672, w29673, w29674, w29675, w29676, w29677, w29678, w29679, w29680, w29681, w29682, w29683, w29684, w29685, w29686, w29687, w29688, w29689, w29690, w29691, w29692, w29693, w29694, w29695, w29696, w29697, w29698, w29699, w29700, w29701, w29702, w29703, w29704, w29705, w29706, w29707, w29708, w29709, w29710, w29711, w29712, w29713, w29714, w29715, w29716, w29717, w29718, w29719, w29720, w29721, w29722, w29723, w29724, w29725, w29726, w29727, w29728, w29729, w29730, w29731, w29732, w29733, w29734, w29735, w29736, w29737, w29738, w29739, w29740, w29741, w29742, w29743, w29744, w29745, w29746, w29747, w29748, w29749, w29750, w29751, w29752, w29753, w29754, w29755, w29756, w29757, w29758, w29759, w29760, w29761, w29762, w29763, w29764, w29765, w29766, w29767, w29768, w29769, w29770, w29771, w29772, w29773, w29774, w29775, w29776, w29777, w29778, w29779, w29780, w29781, w29782, w29783, w29784, w29785, w29786, w29787, w29788, w29789, w29790, w29791, w29792, w29793, w29794, w29795, w29796, w29797, w29798, w29799, w29800, w29801, w29802, w29803, w29804, w29805, w29806, w29807, w29808, w29809, w29810, w29811, w29812, w29813, w29814, w29815, w29816, w29817, w29818, w29819, w29820, w29821, w29822, w29823, w29824, w29825, w29826, w29827, w29828, w29829, w29830, w29831, w29832, w29833, w29834, w29835, w29836, w29837, w29838, w29839, w29840, w29841, w29842, w29843, w29844, w29845, w29846, w29847, w29848, w29849, w29850, w29851, w29852, w29853, w29854, w29855, w29856, w29857, w29858, w29859, w29860, w29861, w29862, w29863, w29864, w29865, w29866, w29867, w29868, w29869, w29870, w29871, w29872, w29873, w29874, w29875, w29876, w29877, w29878, w29879, w29880, w29881, w29882, w29883, w29884, w29885, w29886, w29887, w29888, w29889, w29890, w29891, w29892, w29893, w29894, w29895, w29896, w29897, w29898, w29899, w29900, w29901, w29902, w29903, w29904, w29905, w29906, w29907, w29908, w29909, w29910, w29911, w29912, w29913, w29914, w29915, w29916, w29917, w29918, w29919, w29920, w29921, w29922, w29923, w29924, w29925, w29926, w29927, w29928, w29929, w29930, w29931, w29932, w29933, w29934, w29935, w29936, w29937, w29938, w29939, w29940, w29941, w29942, w29943, w29944, w29945, w29946, w29947, w29948, w29949, w29950, w29951, w29952, w29953, w29954, w29955, w29956, w29957, w29958, w29959, w29960, w29961, w29962, w29963, w29964, w29965, w29966, w29967, w29968, w29969, w29970, w29971, w29972, w29973, w29974, w29975, w29976, w29977, w29978, w29979, w29980, w29981, w29982, w29983, w29984, w29985, w29986, w29987, w29988, w29989, w29990, w29991, w29992, w29993, w29994, w29995, w29996, w29997, w29998, w29999, w30000, w30001, w30002, w30003, w30004, w30005, w30006, w30007, w30008, w30009, w30010, w30011, w30012, w30013, w30014, w30015, w30016, w30017, w30018, w30019, w30020, w30021, w30022, w30023, w30024, w30025, w30026, w30027, w30028, w30029, w30030, w30031, w30032, w30033, w30034, w30035, w30036, w30037, w30038, w30039, w30040, w30041, w30042, w30043, w30044, w30045, w30046, w30047, w30048, w30049, w30050, w30051, w30052, w30053, w30054, w30055, w30056, w30057, w30058, w30059, w30060, w30061, w30062, w30063, w30064, w30065, w30066, w30067, w30068, w30069, w30070, w30071, w30072, w30073, w30074, w30075, w30076, w30077, w30078, w30079, w30080, w30081, w30082, w30083, w30084, w30085, w30086, w30087, w30088, w30089, w30090, w30091, w30092, w30093, w30094, w30095, w30096, w30097, w30098, w30099, w30100, w30101, w30102, w30103, w30104, w30105, w30106, w30107, w30108, w30109, w30110, w30111, w30112, w30113, w30114, w30115, w30116, w30117, w30118, w30119, w30120, w30121, w30122, w30123, w30124, w30125, w30126, w30127, w30128, w30129, w30130, w30131, w30132, w30133, w30134, w30135, w30136, w30137, w30138, w30139, w30140, w30141, w30142, w30143, w30144, w30145, w30146, w30147, w30148, w30149, w30150, w30151, w30152, w30153, w30154, w30155, w30156, w30157, w30158, w30159, w30160, w30161, w30162, w30163, w30164, w30165, w30166, w30167, w30168, w30169, w30170, w30171, w30172, w30173, w30174, w30175, w30176, w30177, w30178, w30179, w30180, w30181, w30182, w30183, w30184, w30185, w30186, w30187, w30188, w30189, w30190, w30191, w30192, w30193, w30194, w30195, w30196, w30197, w30198, w30199, w30200, w30201, w30202, w30203, w30204, w30205, w30206, w30207, w30208, w30209, w30210, w30211, w30212, w30213, w30214, w30215, w30216, w30217, w30218, w30219, w30220, w30221, w30222, w30223, w30224, w30225, w30226, w30227, w30228, w30229, w30230, w30231, w30232, w30233, w30234, w30235, w30236, w30237, w30238, w30239, w30240, w30241, w30242, w30243, w30244, w30245, w30246, w30247, w30248, w30249, w30250, w30251, w30252, w30253, w30254, w30255, w30256, w30257, w30258, w30259, w30260, w30261, w30262, w30263, w30264, w30265, w30266, w30267, w30268, w30269, w30270, w30271, w30272, w30273, w30274, w30275, w30276, w30277, w30278, w30279, w30280, w30281, w30282, w30283, w30284, w30285, w30286, w30287, w30288, w30289, w30290, w30291, w30292, w30293, w30294, w30295, w30296, w30297, w30298, w30299, w30300, w30301, w30302, w30303, w30304, w30305, w30306, w30307, w30308, w30309, w30310, w30311, w30312, w30313, w30314, w30315, w30316, w30317, w30318, w30319, w30320, w30321, w30322, w30323, w30324, w30325, w30326, w30327, w30328, w30329, w30330, w30331, w30332, w30333, w30334, w30335, w30336, w30337, w30338, w30339, w30340, w30341, w30342, w30343, w30344, w30345, w30346, w30347, w30348, w30349, w30350, w30351, w30352, w30353, w30354, w30355, w30356, w30357, w30358, w30359, w30360, w30361, w30362, w30363, w30364, w30365, w30366, w30367, w30368, w30369, w30370, w30371, w30372, w30373, w30374, w30375, w30376, w30377, w30378, w30379, w30380, w30381, w30382, w30383, w30384, w30385, w30386, w30387, w30388, w30389, w30390, w30391, w30392, w30393, w30394, w30395, w30396, w30397, w30398, w30399, w30400, w30401, w30402, w30403, w30404, w30405, w30406, w30407, w30408, w30409, w30410, w30411, w30412, w30413, w30414, w30415, w30416, w30417, w30418, w30419, w30420, w30421, w30422, w30423, w30424, w30425, w30426, w30427, w30428, w30429, w30430, w30431, w30432, w30433, w30434, w30435, w30436, w30437, w30438, w30439, w30440, w30441, w30442, w30443, w30444, w30445, w30446, w30447, w30448, w30449, w30450, w30451, w30452, w30453, w30454, w30455, w30456, w30457, w30458, w30459, w30460, w30461, w30462, w30463, w30464, w30465, w30466, w30467, w30468, w30469, w30470, w30471, w30472, w30473, w30474, w30475, w30476, w30477, w30478, w30479, w30480, w30481, w30482, w30483, w30484, w30485, w30486, w30487, w30488, w30489, w30490, w30491, w30492, w30493, w30494, w30495, w30496, w30497, w30498, w30499, w30500, w30501, w30502, w30503, w30504, w30505, w30506, w30507, w30508, w30509, w30510, w30511, w30512, w30513, w30514, w30515, w30516, w30517, w30518, w30519, w30520, w30521, w30522, w30523, w30524, w30525, w30526, w30527, w30528, w30529, w30530, w30531, w30532, w30533, w30534, w30535, w30536, w30537, w30538, w30539, w30540, w30541, w30542, w30543, w30544, w30545, w30546, w30547, w30548, w30549, w30550, w30551, w30552, w30553, w30554, w30555, w30556, w30557, w30558, w30559, w30560, w30561, w30562, w30563, w30564, w30565, w30566, w30567, w30568, w30569, w30570, w30571, w30572, w30573, w30574, w30575, w30576, w30577, w30578, w30579, w30580, w30581, w30582, w30583, w30584, w30585, w30586, w30587, w30588, w30589, w30590, w30591, w30592, w30593, w30594, w30595, w30596, w30597, w30598, w30599, w30600, w30601, w30602, w30603, w30604, w30605, w30606, w30607, w30608, w30609, w30610, w30611, w30612, w30613, w30614, w30615, w30616, w30617, w30618, w30619, w30620, w30621, w30622, w30623, w30624, w30625, w30626, w30627, w30628, w30629, w30630, w30631, w30632, w30633, w30634, w30635, w30636, w30637, w30638, w30639, w30640, w30641, w30642, w30643, w30644, w30645, w30646, w30647, w30648, w30649, w30650, w30651, w30652, w30653, w30654, w30655, w30656, w30657, w30658, w30659, w30660, w30661, w30662, w30663, w30664, w30665, w30666, w30667, w30668, w30669, w30670, w30671, w30672, w30673, w30674, w30675, w30676, w30677, w30678, w30679, w30680, w30681, w30682, w30683, w30684, w30685, w30686, w30687, w30688, w30689, w30690, w30691, w30692, w30693, w30694, w30695, w30696, w30697, w30698, w30699, w30700, w30701, w30702, w30703, w30704, w30705, w30706, w30707, w30708, w30709, w30710, w30711, w30712, w30713, w30714, w30715, w30716, w30717, w30718, w30719, w30720, w30721, w30722, w30723, w30724, w30725, w30726, w30727, w30728, w30729, w30730, w30731, w30732, w30733, w30734, w30735, w30736, w30737, w30738, w30739, w30740, w30741, w30742, w30743, w30744, w30745, w30746, w30747, w30748, w30749, w30750, w30751, w30752, w30753, w30754, w30755, w30756, w30757, w30758, w30759, w30760, w30761, w30762, w30763, w30764, w30765, w30766, w30767, w30768, w30769, w30770, w30771, w30772, w30773, w30774, w30775, w30776, w30777, w30778, w30779, w30780, w30781, w30782, w30783, w30784, w30785, w30786, w30787, w30788, w30789, w30790, w30791, w30792, w30793, w30794, w30795, w30796, w30797, w30798, w30799, w30800, w30801, w30802, w30803, w30804, w30805, w30806, w30807, w30808, w30809, w30810, w30811, w30812, w30813, w30814, w30815, w30816, w30817, w30818, w30819, w30820, w30821, w30822, w30823, w30824, w30825, w30826, w30827, w30828, w30829, w30830, w30831, w30832, w30833, w30834, w30835, w30836, w30837, w30838, w30839, w30840, w30841, w30842, w30843, w30844, w30845, w30846, w30847, w30848, w30849, w30850, w30851, w30852, w30853, w30854, w30855, w30856, w30857, w30858, w30859, w30860, w30861, w30862, w30863, w30864, w30865, w30866, w30867, w30868, w30869, w30870, w30871, w30872, w30873, w30874, w30875, w30876, w30877, w30878, w30879, w30880, w30881, w30882, w30883, w30884, w30885, w30886, w30887, w30888, w30889, w30890, w30891, w30892, w30893, w30894, w30895, w30896, w30897, w30898, w30899, w30900, w30901, w30902, w30903, w30904, w30905, w30906, w30907, w30908, w30909, w30910, w30911, w30912, w30913, w30914, w30915, w30916, w30917, w30918, w30919, w30920, w30921, w30922, w30923, w30924, w30925, w30926, w30927, w30928, w30929, w30930, w30931, w30932, w30933, w30934, w30935, w30936, w30937, w30938, w30939, w30940, w30941, w30942, w30943, w30944, w30945, w30946, w30947, w30948, w30949, w30950, w30951, w30952, w30953, w30954, w30955, w30956, w30957, w30958, w30959, w30960, w30961, w30962, w30963, w30964, w30965, w30966, w30967, w30968, w30969, w30970, w30971, w30972, w30973, w30974, w30975, w30976, w30977, w30978, w30979, w30980, w30981, w30982, w30983, w30984, w30985, w30986, w30987, w30988, w30989, w30990, w30991, w30992, w30993, w30994, w30995, w30996, w30997, w30998, w30999, w31000, w31001, w31002, w31003, w31004, w31005, w31006, w31007, w31008, w31009, w31010, w31011, w31012, w31013, w31014, w31015, w31016, w31017, w31018, w31019, w31020, w31021, w31022, w31023, w31024, w31025, w31026, w31027, w31028, w31029, w31030, w31031, w31032, w31033, w31034, w31035, w31036, w31037, w31038, w31039, w31040, w31041, w31042, w31043, w31044, w31045, w31046, w31047, w31048, w31049, w31050, w31051, w31052, w31053, w31054, w31055, w31056, w31057, w31058, w31059, w31060, w31061, w31062, w31063, w31064, w31065, w31066, w31067, w31068, w31069, w31070, w31071, w31072, w31073, w31074, w31075, w31076, w31077, w31078, w31079, w31080, w31081, w31082, w31083, w31084, w31085, w31086, w31087, w31088, w31089, w31090, w31091, w31092, w31093, w31094, w31095, w31096, w31097, w31098, w31099, w31100, w31101, w31102, w31103, w31104, w31105, w31106, w31107, w31108, w31109, w31110, w31111, w31112, w31113, w31114, w31115, w31116, w31117, w31118, w31119, w31120, w31121, w31122, w31123, w31124, w31125, w31126, w31127, w31128, w31129, w31130, w31131, w31132, w31133, w31134, w31135, w31136, w31137, w31138, w31139, w31140, w31141, w31142, w31143, w31144, w31145, w31146, w31147, w31148, w31149, w31150, w31151, w31152, w31153, w31154, w31155, w31156, w31157, w31158, w31159, w31160, w31161, w31162, w31163, w31164, w31165, w31166, w31167, w31168, w31169, w31170, w31171, w31172, w31173, w31174, w31175, w31176, w31177, w31178, w31179, w31180, w31181, w31182, w31183, w31184, w31185, w31186, w31187, w31188, w31189, w31190, w31191, w31192, w31193, w31194, w31195, w31196, w31197, w31198, w31199, w31200, w31201, w31202, w31203, w31204, w31205, w31206, w31207, w31208, w31209, w31210, w31211, w31212, w31213, w31214, w31215, w31216, w31217, w31218, w31219, w31220, w31221, w31222, w31223, w31224, w31225, w31226, w31227, w31228, w31229, w31230, w31231, w31232, w31233, w31234, w31235, w31236, w31237, w31238, w31239, w31240, w31241, w31242, w31243, w31244, w31245, w31246, w31247, w31248, w31249, w31250, w31251, w31252, w31253, w31254, w31255, w31256, w31257, w31258, w31259, w31260, w31261, w31262, w31263, w31264, w31265, w31266, w31267, w31268, w31269, w31270, w31271, w31272, w31273, w31274, w31275, w31276, w31277, w31278, w31279, w31280, w31281, w31282, w31283, w31284, w31285, w31286, w31287, w31288, w31289, w31290, w31291, w31292, w31293, w31294, w31295, w31296, w31297, w31298, w31299, w31300, w31301, w31302, w31303, w31304, w31305, w31306, w31307, w31308, w31309, w31310, w31311, w31312, w31313, w31314, w31315, w31316, w31317, w31318, w31319, w31320, w31321, w31322, w31323, w31324, w31325, w31326, w31327, w31328, w31329, w31330, w31331, w31332, w31333, w31334, w31335, w31336, w31337, w31338, w31339, w31340, w31341, w31342, w31343, w31344, w31345, w31346, w31347, w31348, w31349, w31350, w31351, w31352, w31353, w31354, w31355, w31356, w31357, w31358, w31359, w31360, w31361, w31362, w31363, w31364, w31365, w31366, w31367, w31368, w31369, w31370, w31371, w31372, w31373, w31374, w31375, w31376, w31377, w31378, w31379, w31380, w31381, w31382, w31383, w31384, w31385, w31386, w31387, w31388, w31389, w31390, w31391, w31392, w31393, w31394, w31395, w31396, w31397, w31398, w31399, w31400, w31401, w31402, w31403, w31404, w31405, w31406, w31407, w31408, w31409, w31410, w31411, w31412, w31413, w31414, w31415, w31416, w31417, w31418, w31419, w31420, w31421, w31422, w31423, w31424, w31425, w31426, w31427, w31428, w31429, w31430, w31431, w31432, w31433, w31434, w31435, w31436, w31437, w31438, w31439, w31440, w31441, w31442, w31443, w31444, w31445, w31446, w31447, w31448, w31449, w31450, w31451, w31452, w31453, w31454, w31455, w31456, w31457, w31458, w31459, w31460, w31461, w31462, w31463, w31464, w31465, w31466, w31467, w31468, w31469, w31470, w31471, w31472, w31473, w31474, w31475, w31476, w31477, w31478, w31479, w31480, w31481, w31482, w31483, w31484, w31485, w31486, w31487, w31488, w31489, w31490, w31491, w31492, w31493, w31494, w31495, w31496, w31497, w31498, w31499, w31500, w31501, w31502, w31503, w31504, w31505, w31506, w31507, w31508, w31509, w31510, w31511, w31512, w31513, w31514, w31515, w31516, w31517, w31518, w31519, w31520, w31521, w31522, w31523, w31524, w31525, w31526, w31527, w31528, w31529, w31530, w31531, w31532, w31533, w31534, w31535, w31536, w31537, w31538, w31539, w31540, w31541, w31542, w31543, w31544, w31545, w31546, w31547, w31548, w31549, w31550, w31551, w31552, w31553, w31554, w31555, w31556, w31557, w31558, w31559, w31560, w31561, w31562, w31563, w31564, w31565, w31566, w31567, w31568, w31569, w31570, w31571, w31572, w31573, w31574, w31575, w31576, w31577, w31578, w31579, w31580, w31581, w31582, w31583, w31584, w31585, w31586, w31587, w31588, w31589, w31590, w31591, w31592, w31593, w31594, w31595, w31596, w31597, w31598, w31599, w31600, w31601, w31602, w31603, w31604, w31605, w31606, w31607, w31608, w31609, w31610, w31611, w31612, w31613, w31614, w31615, w31616, w31617, w31618, w31619, w31620, w31621, w31622, w31623, w31624, w31625, w31626, w31627, w31628, w31629, w31630, w31631, w31632, w31633, w31634, w31635, w31636, w31637, w31638, w31639, w31640, w31641, w31642, w31643, w31644, w31645, w31646, w31647, w31648, w31649, w31650, w31651, w31652, w31653, w31654, w31655, w31656, w31657, w31658, w31659, w31660, w31661, w31662, w31663, w31664, w31665, w31666, w31667, w31668, w31669, w31670, w31671, w31672, w31673, w31674, w31675, w31676, w31677, w31678, w31679, w31680, w31681, w31682, w31683, w31684, w31685, w31686, w31687, w31688, w31689, w31690, w31691, w31692, w31693, w31694, w31695, w31696, w31697, w31698, w31699, w31700, w31701, w31702, w31703, w31704, w31705, w31706, w31707, w31708, w31709, w31710, w31711, w31712, w31713, w31714, w31715, w31716, w31717, w31718, w31719, w31720, w31721, w31722, w31723, w31724, w31725, w31726, w31727, w31728, w31729, w31730, w31731, w31732, w31733, w31734, w31735, w31736, w31737, w31738, w31739, w31740, w31741, w31742, w31743, w31744, w31745, w31746, w31747, w31748, w31749, w31750, w31751, w31752, w31753, w31754, w31755, w31756, w31757, w31758, w31759, w31760, w31761, w31762, w31763, w31764, w31765, w31766, w31767, w31768, w31769, w31770, w31771, w31772, w31773, w31774, w31775, w31776, w31777, w31778, w31779, w31780, w31781, w31782, w31783, w31784, w31785, w31786, w31787, w31788, w31789, w31790, w31791, w31792, w31793, w31794, w31795, w31796, w31797, w31798, w31799, w31800, w31801, w31802, w31803, w31804, w31805, w31806, w31807, w31808, w31809, w31810, w31811, w31812, w31813, w31814, w31815, w31816, w31817, w31818, w31819, w31820, w31821, w31822, w31823, w31824, w31825, w31826, w31827, w31828, w31829, w31830, w31831, w31832, w31833, w31834, w31835, w31836, w31837, w31838, w31839, w31840, w31841, w31842, w31843, w31844, w31845, w31846, w31847, w31848, w31849, w31850, w31851, w31852, w31853, w31854, w31855, w31856, w31857, w31858, w31859, w31860, w31861, w31862, w31863, w31864, w31865, w31866, w31867, w31868, w31869, w31870, w31871, w31872, w31873, w31874, w31875, w31876, w31877, w31878, w31879, w31880, w31881, w31882, w31883, w31884, w31885, w31886, w31887, w31888, w31889, w31890, w31891, w31892, w31893, w31894, w31895, w31896, w31897, w31898, w31899, w31900, w31901, w31902, w31903, w31904, w31905, w31906, w31907, w31908, w31909, w31910, w31911, w31912, w31913, w31914, w31915, w31916, w31917, w31918, w31919, w31920, w31921, w31922, w31923, w31924, w31925, w31926, w31927, w31928, w31929, w31930, w31931, w31932, w31933, w31934, w31935, w31936, w31937, w31938, w31939, w31940, w31941, w31942, w31943, w31944, w31945, w31946, w31947, w31948, w31949, w31950, w31951, w31952, w31953, w31954, w31955, w31956, w31957, w31958, w31959, w31960, w31961, w31962, w31963, w31964, w31965, w31966, w31967, w31968, w31969, w31970, w31971, w31972, w31973, w31974, w31975, w31976, w31977, w31978, w31979, w31980, w31981, w31982, w31983, w31984, w31985, w31986, w31987, w31988, w31989, w31990, w31991, w31992, w31993, w31994, w31995, w31996, w31997, w31998, w31999, w32000, w32001, w32002, w32003, w32004, w32005, w32006, w32007, w32008, w32009, w32010, w32011, w32012, w32013, w32014, w32015, w32016, w32017, w32018, w32019, w32020, w32021, w32022, w32023, w32024, w32025, w32026, w32027, w32028, w32029, w32030, w32031, w32032, w32033, w32034, w32035, w32036, w32037, w32038, w32039, w32040, w32041, w32042, w32043, w32044, w32045, w32046, w32047, w32048, w32049, w32050, w32051, w32052, w32053, w32054, w32055, w32056, w32057, w32058, w32059, w32060, w32061, w32062, w32063, w32064, w32065, w32066, w32067, w32068, w32069, w32070, w32071, w32072, w32073, w32074, w32075, w32076, w32077, w32078, w32079, w32080, w32081, w32082, w32083, w32084, w32085, w32086, w32087, w32088, w32089, w32090, w32091, w32092, w32093, w32094, w32095, w32096, w32097, w32098, w32099, w32100, w32101, w32102, w32103, w32104, w32105, w32106, w32107, w32108, w32109, w32110, w32111, w32112, w32113, w32114, w32115, w32116, w32117, w32118, w32119, w32120, w32121, w32122, w32123, w32124, w32125, w32126, w32127, w32128, w32129, w32130, w32131, w32132, w32133, w32134, w32135, w32136, w32137, w32138, w32139, w32140, w32141, w32142, w32143, w32144, w32145, w32146, w32147, w32148, w32149, w32150, w32151, w32152, w32153, w32154, w32155, w32156, w32157, w32158, w32159, w32160, w32161, w32162, w32163, w32164, w32165, w32166, w32167, w32168, w32169, w32170, w32171, w32172, w32173, w32174, w32175, w32176, w32177, w32178, w32179, w32180, w32181, w32182, w32183, w32184, w32185, w32186, w32187, w32188, w32189, w32190, w32191, w32192, w32193, w32194, w32195, w32196, w32197, w32198, w32199, w32200, w32201, w32202, w32203, w32204, w32205, w32206, w32207, w32208, w32209, w32210, w32211, w32212, w32213, w32214, w32215, w32216, w32217, w32218, w32219, w32220, w32221, w32222, w32223, w32224, w32225, w32226, w32227, w32228, w32229, w32230, w32231, w32232, w32233, w32234, w32235, w32236, w32237, w32238, w32239, w32240, w32241, w32242, w32243, w32244, w32245, w32246, w32247, w32248, w32249, w32250, w32251, w32252, w32253, w32254, w32255, w32256, w32257, w32258, w32259, w32260, w32261, w32262, w32263, w32264, w32265, w32266, w32267, w32268, w32269, w32270, w32271, w32272, w32273, w32274, w32275, w32276, w32277, w32278, w32279, w32280, w32281, w32282, w32283, w32284, w32285, w32286, w32287, w32288, w32289, w32290, w32291, w32292, w32293, w32294, w32295, w32296, w32297, w32298, w32299, w32300, w32301, w32302, w32303, w32304, w32305, w32306, w32307, w32308, w32309, w32310, w32311, w32312, w32313, w32314, w32315, w32316, w32317, w32318, w32319, w32320, w32321, w32322, w32323, w32324, w32325, w32326, w32327, w32328, w32329, w32330, w32331, w32332, w32333, w32334, w32335, w32336, w32337, w32338, w32339, w32340, w32341, w32342, w32343, w32344, w32345, w32346, w32347, w32348, w32349, w32350, w32351, w32352, w32353, w32354, w32355, w32356, w32357, w32358, w32359, w32360, w32361, w32362, w32363, w32364, w32365, w32366, w32367, w32368, w32369, w32370, w32371, w32372, w32373, w32374, w32375, w32376, w32377, w32378, w32379, w32380, w32381, w32382, w32383, w32384, w32385, w32386, w32387, w32388, w32389, w32390, w32391, w32392, w32393, w32394, w32395, w32396, w32397, w32398, w32399, w32400, w32401, w32402, w32403, w32404, w32405, w32406, w32407, w32408, w32409, w32410, w32411, w32412, w32413, w32414, w32415, w32416, w32417, w32418, w32419, w32420, w32421, w32422, w32423, w32424, w32425, w32426, w32427, w32428, w32429, w32430, w32431, w32432, w32433, w32434, w32435, w32436, w32437, w32438, w32439, w32440, w32441, w32442, w32443, w32444, w32445, w32446, w32447, w32448, w32449, w32450, w32451, w32452, w32453, w32454, w32455, w32456, w32457, w32458, w32459, w32460, w32461, w32462, w32463, w32464, w32465, w32466, w32467, w32468, w32469, w32470, w32471, w32472, w32473, w32474, w32475, w32476, w32477, w32478, w32479, w32480, w32481, w32482, w32483, w32484, w32485, w32486, w32487, w32488, w32489, w32490, w32491, w32492, w32493, w32494, w32495, w32496, w32497, w32498, w32499, w32500, w32501, w32502, w32503, w32504, w32505, w32506, w32507, w32508, w32509, w32510, w32511, w32512, w32513, w32514, w32515, w32516, w32517, w32518, w32519, w32520, w32521, w32522, w32523, w32524, w32525, w32526, w32527, w32528, w32529, w32530, w32531, w32532, w32533, w32534, w32535, w32536, w32537, w32538, w32539, w32540, w32541, w32542, w32543, w32544, w32545, w32546, w32547, w32548, w32549, w32550, w32551, w32552, w32553, w32554, w32555, w32556, w32557, w32558, w32559, w32560, w32561, w32562, w32563, w32564, w32565, w32566, w32567, w32568, w32569, w32570, w32571, w32572, w32573, w32574, w32575, w32576, w32577, w32578, w32579, w32580, w32581, w32582, w32583, w32584, w32585, w32586, w32587, w32588, w32589, w32590, w32591, w32592, w32593, w32594, w32595, w32596, w32597, w32598, w32599, w32600, w32601, w32602, w32603, w32604, w32605, w32606, w32607, w32608, w32609, w32610, w32611, w32612, w32613, w32614, w32615, w32616, w32617, w32618, w32619, w32620, w32621, w32622, w32623, w32624, w32625, w32626, w32627, w32628, w32629, w32630, w32631, w32632, w32633, w32634, w32635, w32636, w32637, w32638, w32639, w32640, w32641, w32642, w32643, w32644, w32645, w32646, w32647, w32648, w32649, w32650, w32651, w32652, w32653, w32654, w32655, w32656, w32657, w32658, w32659, w32660, w32661, w32662, w32663, w32664, w32665, w32666, w32667, w32668, w32669, w32670, w32671, w32672, w32673, w32674, w32675, w32676, w32677, w32678, w32679, w32680, w32681, w32682, w32683, w32684, w32685, w32686, w32687, w32688, w32689, w32690, w32691, w32692, w32693, w32694, w32695, w32696, w32697, w32698, w32699, w32700, w32701, w32702, w32703, w32704, w32705, w32706, w32707, w32708, w32709, w32710, w32711, w32712, w32713, w32714, w32715, w32716, w32717, w32718, w32719, w32720, w32721, w32722, w32723, w32724, w32725, w32726, w32727, w32728, w32729, w32730, w32731, w32732, w32733, w32734, w32735, w32736, w32737, w32738, w32739, w32740, w32741, w32742, w32743, w32744, w32745, w32746, w32747, w32748, w32749, w32750, w32751, w32752, w32753, w32754, w32755, w32756, w32757, w32758, w32759, w32760, w32761, w32762, w32763, w32764, w32765, w32766, w32767, w32768, w32769, w32770, w32771, w32772, w32773, w32774, w32775, w32776, w32777, w32778, w32779, w32780, w32781, w32782, w32783, w32784, w32785, w32786, w32787, w32788, w32789, w32790, w32791, w32792, w32793, w32794, w32795, w32796, w32797, w32798, w32799, w32800, w32801, w32802, w32803, w32804, w32805, w32806, w32807, w32808, w32809, w32810, w32811, w32812, w32813, w32814, w32815, w32816, w32817, w32818, w32819, w32820, w32821, w32822, w32823, w32824, w32825, w32826, w32827, w32828, w32829, w32830, w32831, w32832, w32833, w32834, w32835, w32836, w32837, w32838, w32839, w32840, w32841, w32842, w32843, w32844, w32845, w32846, w32847, w32848, w32849, w32850, w32851, w32852, w32853, w32854, w32855, w32856, w32857, w32858, w32859, w32860, w32861, w32862, w32863, w32864, w32865, w32866, w32867, w32868, w32869, w32870, w32871, w32872, w32873, w32874, w32875, w32876, w32877, w32878, w32879, w32880, w32881, w32882, w32883, w32884, w32885, w32886, w32887, w32888, w32889, w32890, w32891, w32892, w32893, w32894, w32895, w32896, w32897, w32898, w32899, w32900, w32901, w32902, w32903, w32904, w32905, w32906, w32907, w32908, w32909, w32910, w32911, w32912, w32913, w32914, w32915, w32916, w32917, w32918, w32919, w32920, w32921, w32922, w32923, w32924, w32925, w32926, w32927, w32928, w32929, w32930, w32931, w32932, w32933, w32934, w32935, w32936, w32937, w32938, w32939, w32940, w32941, w32942, w32943, w32944, w32945, w32946, w32947, w32948, w32949, w32950, w32951, w32952, w32953, w32954, w32955, w32956, w32957, w32958, w32959, w32960, w32961, w32962, w32963, w32964, w32965, w32966, w32967, w32968, w32969, w32970, w32971, w32972, w32973, w32974, w32975, w32976, w32977, w32978, w32979, w32980, w32981, w32982, w32983, w32984, w32985, w32986, w32987, w32988, w32989, w32990, w32991, w32992, w32993, w32994, w32995, w32996, w32997, w32998, w32999, w33000, w33001, w33002, w33003, w33004, w33005, w33006, w33007, w33008, w33009, w33010, w33011, w33012, w33013, w33014, w33015, w33016, w33017, w33018, w33019, w33020, w33021, w33022, w33023, w33024, w33025, w33026, w33027, w33028, w33029, w33030, w33031, w33032, w33033, w33034, w33035, w33036, w33037, w33038, w33039, w33040, w33041, w33042, w33043, w33044, w33045, w33046, w33047, w33048, w33049, w33050, w33051, w33052, w33053, w33054, w33055, w33056, w33057, w33058, w33059, w33060, w33061, w33062, w33063, w33064, w33065, w33066, w33067, w33068, w33069, w33070, w33071, w33072, w33073, w33074, w33075, w33076, w33077, w33078, w33079, w33080, w33081, w33082, w33083, w33084, w33085, w33086, w33087, w33088, w33089, w33090, w33091, w33092, w33093, w33094, w33095, w33096, w33097, w33098, w33099, w33100, w33101, w33102, w33103, w33104, w33105, w33106, w33107, w33108, w33109, w33110, w33111, w33112, w33113, w33114, w33115, w33116, w33117, w33118, w33119, w33120, w33121, w33122, w33123, w33124, w33125, w33126, w33127, w33128, w33129, w33130, w33131, w33132, w33133, w33134, w33135, w33136, w33137, w33138, w33139, w33140, w33141, w33142, w33143, w33144, w33145, w33146, w33147, w33148, w33149, w33150, w33151, w33152, w33153, w33154, w33155, w33156, w33157, w33158, w33159, w33160, w33161, w33162, w33163, w33164, w33165, w33166, w33167, w33168, w33169, w33170, w33171, w33172, w33173, w33174, w33175, w33176, w33177, w33178, w33179, w33180, w33181, w33182, w33183, w33184, w33185, w33186, w33187, w33188, w33189, w33190, w33191, w33192, w33193, w33194, w33195, w33196, w33197, w33198, w33199, w33200, w33201, w33202, w33203, w33204, w33205, w33206, w33207, w33208, w33209, w33210, w33211, w33212, w33213, w33214, w33215, w33216, w33217, w33218, w33219, w33220, w33221, w33222, w33223, w33224, w33225, w33226, w33227, w33228, w33229, w33230, w33231, w33232, w33233, w33234, w33235, w33236, w33237, w33238, w33239, w33240, w33241, w33242, w33243, w33244, w33245, w33246, w33247, w33248, w33249, w33250, w33251, w33252, w33253, w33254, w33255, w33256, w33257, w33258, w33259, w33260, w33261, w33262, w33263, w33264, w33265, w33266, w33267, w33268, w33269, w33270, w33271, w33272, w33273, w33274, w33275, w33276, w33277, w33278, w33279, w33280, w33281, w33282, w33283, w33284, w33285, w33286, w33287, w33288, w33289, w33290, w33291, w33292, w33293, w33294, w33295, w33296, w33297, w33298, w33299, w33300, w33301, w33302, w33303, w33304, w33305, w33306, w33307, w33308, w33309, w33310, w33311, w33312, w33313, w33314, w33315, w33316, w33317, w33318, w33319, w33320, w33321, w33322, w33323, w33324, w33325, w33326, w33327, w33328, w33329, w33330, w33331, w33332, w33333, w33334, w33335, w33336, w33337, w33338, w33339, w33340, w33341, w33342, w33343, w33344, w33345, w33346, w33347, w33348, w33349, w33350, w33351, w33352, w33353, w33354, w33355, w33356, w33357, w33358, w33359, w33360, w33361, w33362, w33363, w33364, w33365, w33366, w33367, w33368, w33369, w33370, w33371, w33372, w33373, w33374, w33375, w33376, w33377, w33378, w33379, w33380, w33381, w33382, w33383, w33384, w33385, w33386, w33387, w33388, w33389, w33390, w33391, w33392, w33393, w33394, w33395, w33396, w33397, w33398, w33399, w33400, w33401, w33402, w33403, w33404, w33405, w33406, w33407, w33408, w33409, w33410, w33411, w33412, w33413, w33414, w33415, w33416, w33417, w33418, w33419, w33420, w33421, w33422, w33423, w33424, w33425, w33426, w33427, w33428, w33429, w33430, w33431, w33432, w33433, w33434, w33435, w33436, w33437, w33438, w33439, w33440, w33441, w33442, w33443, w33444, w33445, w33446, w33447, w33448, w33449, w33450, w33451, w33452, w33453, w33454, w33455, w33456, w33457, w33458, w33459, w33460, w33461, w33462, w33463, w33464, w33465, w33466, w33467, w33468, w33469, w33470, w33471, w33472, w33473, w33474, w33475, w33476, w33477, w33478, w33479, w33480, w33481, w33482, w33483, w33484, w33485, w33486, w33487, w33488, w33489, w33490, w33491, w33492, w33493, w33494, w33495, w33496, w33497, w33498, w33499, w33500, w33501, w33502, w33503, w33504, w33505, w33506, w33507, w33508, w33509, w33510, w33511, w33512, w33513, w33514, w33515, w33516, w33517, w33518, w33519, w33520, w33521, w33522, w33523, w33524, w33525, w33526, w33527, w33528, w33529, w33530, w33531, w33532, w33533, w33534, w33535, w33536, w33537, w33538, w33539, w33540, w33541, w33542, w33543, w33544, w33545, w33546, w33547, w33548, w33549, w33550, w33551, w33552, w33553, w33554, w33555, w33556, w33557, w33558, w33559, w33560, w33561, w33562, w33563, w33564, w33565, w33566, w33567, w33568, w33569, w33570, w33571, w33572, w33573, w33574, w33575, w33576, w33577, w33578, w33579, w33580, w33581, w33582, w33583, w33584, w33585, w33586, w33587, w33588, w33589, w33590, w33591, w33592, w33593, w33594, w33595, w33596, w33597, w33598, w33599, w33600, w33601, w33602, w33603, w33604, w33605, w33606, w33607, w33608, w33609, w33610, w33611, w33612, w33613, w33614, w33615, w33616, w33617, w33618, w33619, w33620, w33621, w33622, w33623, w33624, w33625, w33626, w33627, w33628, w33629, w33630, w33631, w33632, w33633, w33634, w33635, w33636, w33637, w33638, w33639, w33640, w33641, w33642, w33643, w33644, w33645, w33646, w33647, w33648, w33649, w33650, w33651, w33652, w33653, w33654, w33655, w33656, w33657, w33658, w33659, w33660, w33661, w33662, w33663, w33664, w33665, w33666, w33667, w33668, w33669, w33670, w33671, w33672, w33673, w33674, w33675, w33676, w33677, w33678, w33679, w33680, w33681, w33682, w33683, w33684, w33685, w33686, w33687, w33688, w33689, w33690, w33691, w33692, w33693, w33694, w33695, w33696, w33697, w33698, w33699, w33700, w33701, w33702, w33703, w33704, w33705, w33706, w33707, w33708, w33709, w33710, w33711, w33712, w33713, w33714, w33715, w33716, w33717, w33718, w33719, w33720, w33721, w33722, w33723, w33724, w33725, w33726, w33727, w33728, w33729, w33730, w33731, w33732, w33733, w33734, w33735, w33736, w33737, w33738, w33739, w33740, w33741, w33742, w33743, w33744, w33745, w33746, w33747, w33748, w33749, w33750, w33751, w33752, w33753, w33754, w33755, w33756, w33757, w33758, w33759, w33760, w33761, w33762, w33763, w33764, w33765, w33766, w33767, w33768, w33769, w33770, w33771, w33772, w33773, w33774, w33775, w33776, w33777, w33778, w33779, w33780, w33781, w33782, w33783, w33784, w33785, w33786, w33787, w33788, w33789, w33790, w33791, w33792, w33793, w33794, w33795, w33796, w33797, w33798, w33799, w33800, w33801, w33802, w33803, w33804, w33805, w33806, w33807, w33808, w33809, w33810, w33811, w33812, w33813, w33814, w33815, w33816, w33817, w33818, w33819, w33820, w33821, w33822, w33823, w33824, w33825, w33826, w33827, w33828, w33829, w33830, w33831, w33832, w33833, w33834, w33835, w33836, w33837, w33838, w33839, w33840, w33841, w33842, w33843, w33844, w33845, w33846, w33847, w33848, w33849, w33850, w33851, w33852, w33853, w33854, w33855, w33856, w33857, w33858, w33859, w33860, w33861, w33862, w33863, w33864, w33865, w33866, w33867, w33868, w33869, w33870, w33871, w33872, w33873, w33874, w33875, w33876, w33877, w33878, w33879, w33880, w33881, w33882, w33883, w33884, w33885, w33886, w33887, w33888, w33889, w33890, w33891, w33892, w33893, w33894, w33895, w33896, w33897, w33898, w33899, w33900, w33901, w33902, w33903, w33904, w33905, w33906, w33907, w33908, w33909, w33910, w33911, w33912, w33913, w33914, w33915, w33916, w33917, w33918, w33919, w33920, w33921, w33922, w33923, w33924, w33925, w33926, w33927, w33928, w33929, w33930, w33931, w33932, w33933, w33934, w33935, w33936, w33937, w33938, w33939, w33940, w33941, w33942, w33943, w33944, w33945, w33946, w33947, w33948, w33949, w33950, w33951, w33952, w33953, w33954, w33955, w33956, w33957, w33958, w33959, w33960, w33961, w33962, w33963, w33964, w33965, w33966, w33967, w33968, w33969, w33970, w33971, w33972, w33973, w33974, w33975, w33976, w33977, w33978, w33979, w33980, w33981, w33982, w33983, w33984, w33985, w33986, w33987, w33988, w33989, w33990, w33991, w33992, w33993, w33994, w33995, w33996, w33997, w33998, w33999, w34000, w34001, w34002, w34003, w34004, w34005, w34006, w34007, w34008, w34009, w34010, w34011, w34012, w34013, w34014, w34015, w34016, w34017, w34018, w34019, w34020, w34021, w34022, w34023, w34024, w34025, w34026, w34027, w34028, w34029, w34030, w34031, w34032, w34033, w34034, w34035, w34036, w34037, w34038, w34039, w34040, w34041, w34042, w34043, w34044, w34045, w34046, w34047, w34048, w34049, w34050, w34051, w34052, w34053, w34054, w34055, w34056, w34057, w34058, w34059, w34060, w34061, w34062, w34063, w34064, w34065, w34066, w34067, w34068, w34069, w34070, w34071, w34072, w34073, w34074, w34075, w34076, w34077, w34078, w34079, w34080, w34081, w34082, w34083, w34084, w34085, w34086, w34087, w34088, w34089, w34090, w34091, w34092, w34093, w34094, w34095, w34096, w34097, w34098, w34099, w34100, w34101, w34102, w34103, w34104, w34105, w34106, w34107, w34108, w34109, w34110, w34111, w34112, w34113, w34114, w34115, w34116, w34117, w34118, w34119, w34120, w34121, w34122, w34123, w34124, w34125, w34126, w34127, w34128, w34129, w34130, w34131, w34132, w34133, w34134, w34135, w34136, w34137, w34138, w34139, w34140, w34141, w34142, w34143, w34144, w34145, w34146, w34147, w34148, w34149, w34150, w34151, w34152, w34153, w34154, w34155, w34156, w34157, w34158, w34159, w34160, w34161, w34162, w34163, w34164, w34165, w34166, w34167, w34168, w34169, w34170, w34171, w34172, w34173, w34174, w34175, w34176, w34177, w34178, w34179, w34180, w34181, w34182, w34183, w34184, w34185, w34186, w34187, w34188, w34189, w34190, w34191, w34192, w34193, w34194, w34195, w34196, w34197, w34198, w34199, w34200, w34201, w34202, w34203, w34204, w34205, w34206, w34207, w34208, w34209, w34210, w34211, w34212, w34213, w34214, w34215, w34216, w34217, w34218, w34219, w34220, w34221, w34222, w34223, w34224, w34225, w34226, w34227, w34228, w34229, w34230, w34231, w34232, w34233, w34234, w34235, w34236, w34237, w34238, w34239, w34240, w34241, w34242, w34243, w34244, w34245, w34246, w34247, w34248, w34249, w34250, w34251, w34252, w34253, w34254, w34255, w34256, w34257, w34258, w34259, w34260, w34261, w34262, w34263, w34264, w34265, w34266, w34267, w34268, w34269, w34270, w34271, w34272, w34273, w34274, w34275, w34276, w34277, w34278, w34279, w34280, w34281, w34282, w34283, w34284, w34285, w34286, w34287, w34288, w34289, w34290, w34291, w34292, w34293, w34294, w34295, w34296, w34297, w34298, w34299, w34300, w34301, w34302, w34303, w34304, w34305, w34306, w34307, w34308, w34309, w34310, w34311, w34312, w34313, w34314, w34315, w34316, w34317, w34318, w34319, w34320, w34321, w34322, w34323, w34324, w34325, w34326, w34327, w34328, w34329, w34330, w34331, w34332, w34333, w34334, w34335, w34336, w34337, w34338, w34339, w34340, w34341, w34342, w34343, w34344, w34345, w34346, w34347, w34348, w34349, w34350, w34351, w34352, w34353, w34354, w34355, w34356, w34357, w34358, w34359, w34360, w34361, w34362, w34363, w34364, w34365, w34366, w34367, w34368, w34369, w34370, w34371, w34372, w34373, w34374, w34375, w34376, w34377, w34378, w34379, w34380, w34381, w34382, w34383, w34384, w34385, w34386, w34387, w34388, w34389, w34390, w34391, w34392, w34393, w34394, w34395, w34396, w34397, w34398, w34399, w34400, w34401, w34402, w34403, w34404, w34405, w34406, w34407, w34408, w34409, w34410, w34411, w34412, w34413, w34414, w34415, w34416, w34417, w34418, w34419, w34420, w34421, w34422, w34423, w34424, w34425, w34426, w34427, w34428, w34429, w34430, w34431, w34432, w34433, w34434, w34435, w34436, w34437, w34438, w34439, w34440, w34441, w34442, w34443, w34444, w34445, w34446, w34447, w34448, w34449, w34450, w34451, w34452, w34453, w34454, w34455, w34456, w34457, w34458, w34459, w34460, w34461, w34462, w34463, w34464, w34465, w34466, w34467, w34468, w34469, w34470, w34471, w34472, w34473, w34474, w34475, w34476, w34477, w34478, w34479, w34480, w34481, w34482, w34483, w34484, w34485, w34486, w34487, w34488, w34489, w34490, w34491, w34492, w34493, w34494, w34495, w34496, w34497, w34498, w34499, w34500, w34501, w34502, w34503, w34504, w34505, w34506, w34507, w34508, w34509, w34510, w34511, w34512, w34513, w34514, w34515, w34516, w34517, w34518, w34519, w34520, w34521, w34522, w34523, w34524, w34525, w34526, w34527, w34528, w34529, w34530, w34531, w34532, w34533, w34534, w34535, w34536, w34537, w34538, w34539, w34540, w34541, w34542, w34543, w34544, w34545, w34546, w34547, w34548, w34549, w34550, w34551, w34552, w34553, w34554, w34555, w34556, w34557, w34558, w34559, w34560, w34561, w34562, w34563, w34564, w34565, w34566, w34567, w34568, w34569, w34570, w34571, w34572, w34573, w34574, w34575, w34576, w34577, w34578, w34579, w34580, w34581, w34582, w34583, w34584, w34585, w34586, w34587, w34588, w34589, w34590, w34591, w34592, w34593, w34594, w34595, w34596, w34597, w34598, w34599, w34600, w34601, w34602, w34603, w34604, w34605, w34606, w34607, w34608, w34609, w34610, w34611, w34612, w34613, w34614, w34615, w34616, w34617, w34618, w34619, w34620, w34621, w34622, w34623, w34624, w34625, w34626, w34627, w34628, w34629, w34630, w34631, w34632, w34633, w34634, w34635, w34636, w34637, w34638, w34639, w34640, w34641, w34642, w34643, w34644, w34645, w34646, w34647, w34648, w34649, w34650, w34651, w34652, w34653, w34654, w34655, w34656, w34657, w34658, w34659, w34660, w34661, w34662, w34663, w34664, w34665, w34666, w34667, w34668, w34669, w34670, w34671, w34672, w34673, w34674, w34675, w34676, w34677, w34678, w34679, w34680, w34681, w34682, w34683, w34684, w34685, w34686, w34687, w34688, w34689, w34690, w34691, w34692, w34693, w34694, w34695, w34696, w34697, w34698, w34699, w34700, w34701, w34702, w34703, w34704, w34705, w34706, w34707, w34708, w34709, w34710, w34711, w34712, w34713, w34714, w34715, w34716, w34717, w34718, w34719, w34720, w34721, w34722, w34723, w34724, w34725, w34726, w34727, w34728, w34729, w34730, w34731, w34732, w34733, w34734, w34735, w34736, w34737, w34738, w34739, w34740, w34741, w34742, w34743, w34744, w34745, w34746, w34747, w34748, w34749, w34750, w34751, w34752, w34753, w34754, w34755, w34756, w34757, w34758, w34759, w34760, w34761, w34762, w34763, w34764, w34765, w34766, w34767, w34768, w34769, w34770, w34771, w34772, w34773, w34774, w34775, w34776, w34777, w34778, w34779, w34780, w34781, w34782, w34783, w34784, w34785, w34786, w34787, w34788, w34789, w34790, w34791, w34792, w34793, w34794, w34795, w34796, w34797, w34798, w34799, w34800, w34801, w34802, w34803, w34804, w34805, w34806, w34807, w34808, w34809, w34810, w34811, w34812, w34813, w34814, w34815, w34816, w34817, w34818, w34819, w34820, w34821, w34822, w34823, w34824, w34825, w34826, w34827, w34828, w34829, w34830, w34831, w34832, w34833, w34834, w34835, w34836, w34837, w34838, w34839, w34840, w34841, w34842, w34843, w34844, w34845, w34846, w34847, w34848, w34849, w34850, w34851, w34852, w34853, w34854, w34855, w34856, w34857, w34858, w34859, w34860, w34861, w34862, w34863, w34864, w34865, w34866, w34867, w34868, w34869, w34870, w34871, w34872, w34873, w34874, w34875, w34876, w34877, w34878, w34879, w34880, w34881, w34882, w34883, w34884, w34885, w34886, w34887, w34888, w34889, w34890, w34891, w34892, w34893, w34894, w34895, w34896, w34897, w34898, w34899, w34900, w34901, w34902, w34903, w34904, w34905, w34906, w34907, w34908, w34909, w34910, w34911, w34912, w34913, w34914, w34915, w34916, w34917, w34918, w34919, w34920, w34921, w34922, w34923, w34924, w34925, w34926, w34927, w34928, w34929, w34930, w34931, w34932, w34933, w34934, w34935, w34936, w34937, w34938, w34939, w34940, w34941, w34942, w34943, w34944, w34945, w34946, w34947, w34948, w34949, w34950, w34951, w34952, w34953, w34954, w34955, w34956, w34957, w34958, w34959, w34960, w34961, w34962, w34963, w34964, w34965, w34966, w34967, w34968, w34969, w34970, w34971, w34972, w34973, w34974, w34975, w34976, w34977, w34978, w34979, w34980, w34981, w34982, w34983, w34984, w34985, w34986, w34987, w34988, w34989, w34990, w34991, w34992, w34993, w34994, w34995, w34996, w34997, w34998, w34999, w35000, w35001, w35002, w35003, w35004, w35005, w35006, w35007, w35008, w35009, w35010, w35011, w35012, w35013, w35014, w35015, w35016, w35017, w35018, w35019, w35020, w35021, w35022, w35023, w35024, w35025, w35026, w35027, w35028, w35029, w35030, w35031, w35032, w35033, w35034, w35035, w35036, w35037, w35038, w35039, w35040, w35041, w35042, w35043, w35044, w35045, w35046, w35047, w35048, w35049, w35050, w35051, w35052, w35053, w35054, w35055, w35056, w35057, w35058, w35059, w35060, w35061, w35062, w35063, w35064, w35065, w35066, w35067, w35068, w35069, w35070, w35071, w35072, w35073, w35074, w35075, w35076, w35077, w35078, w35079, w35080, w35081, w35082, w35083, w35084, w35085, w35086, w35087, w35088, w35089, w35090, w35091, w35092, w35093, w35094, w35095, w35096, w35097, w35098, w35099, w35100, w35101, w35102, w35103, w35104, w35105, w35106, w35107, w35108, w35109, w35110, w35111, w35112, w35113, w35114, w35115, w35116, w35117, w35118, w35119, w35120, w35121, w35122, w35123, w35124, w35125, w35126, w35127, w35128, w35129, w35130, w35131, w35132, w35133, w35134, w35135, w35136, w35137, w35138, w35139, w35140, w35141, w35142, w35143, w35144, w35145, w35146, w35147, w35148, w35149, w35150, w35151, w35152, w35153, w35154, w35155, w35156, w35157, w35158, w35159, w35160, w35161, w35162, w35163, w35164, w35165, w35166, w35167, w35168, w35169, w35170, w35171, w35172, w35173, w35174, w35175, w35176, w35177, w35178, w35179, w35180, w35181, w35182, w35183, w35184, w35185, w35186, w35187, w35188, w35189, w35190, w35191, w35192, w35193, w35194, w35195, w35196, w35197, w35198, w35199, w35200, w35201, w35202, w35203, w35204, w35205, w35206, w35207, w35208, w35209, w35210, w35211, w35212, w35213, w35214, w35215, w35216, w35217, w35218, w35219, w35220, w35221, w35222, w35223, w35224, w35225, w35226, w35227, w35228, w35229, w35230, w35231, w35232, w35233, w35234, w35235, w35236, w35237, w35238, w35239, w35240, w35241, w35242, w35243, w35244, w35245, w35246, w35247, w35248, w35249, w35250, w35251, w35252, w35253, w35254, w35255, w35256, w35257, w35258, w35259, w35260, w35261, w35262, w35263, w35264, w35265, w35266, w35267, w35268, w35269, w35270, w35271, w35272, w35273, w35274, w35275, w35276, w35277, w35278, w35279, w35280, w35281, w35282, w35283, w35284, w35285, w35286, w35287, w35288, w35289, w35290, w35291, w35292, w35293, w35294, w35295, w35296, w35297, w35298, w35299, w35300, w35301, w35302, w35303, w35304, w35305, w35306, w35307, w35308, w35309, w35310, w35311, w35312, w35313, w35314, w35315, w35316, w35317, w35318, w35319, w35320, w35321, w35322, w35323, w35324, w35325, w35326, w35327, w35328, w35329, w35330, w35331, w35332, w35333, w35334, w35335, w35336, w35337, w35338, w35339, w35340, w35341, w35342, w35343, w35344, w35345, w35346, w35347, w35348, w35349, w35350, w35351, w35352, w35353, w35354, w35355, w35356, w35357, w35358, w35359, w35360, w35361, w35362, w35363, w35364, w35365, w35366, w35367, w35368, w35369, w35370, w35371, w35372, w35373, w35374, w35375, w35376, w35377, w35378, w35379, w35380, w35381, w35382, w35383, w35384, w35385, w35386, w35387, w35388, w35389, w35390, w35391, w35392, w35393, w35394, w35395, w35396, w35397, w35398, w35399, w35400, w35401, w35402, w35403, w35404, w35405, w35406, w35407, w35408, w35409, w35410, w35411, w35412, w35413, w35414, w35415, w35416, w35417, w35418, w35419, w35420, w35421, w35422, w35423, w35424, w35425, w35426, w35427, w35428, w35429, w35430, w35431, w35432, w35433, w35434, w35435, w35436, w35437, w35438, w35439, w35440, w35441, w35442, w35443, w35444, w35445, w35446, w35447, w35448, w35449, w35450, w35451, w35452, w35453, w35454, w35455, w35456, w35457, w35458, w35459, w35460, w35461, w35462, w35463, w35464, w35465, w35466, w35467, w35468, w35469, w35470, w35471, w35472, w35473, w35474, w35475, w35476, w35477, w35478, w35479, w35480, w35481, w35482, w35483, w35484, w35485, w35486, w35487, w35488, w35489, w35490, w35491, w35492, w35493, w35494, w35495, w35496, w35497, w35498, w35499, w35500, w35501, w35502, w35503, w35504, w35505, w35506, w35507, w35508, w35509, w35510, w35511, w35512, w35513, w35514, w35515, w35516, w35517, w35518, w35519, w35520, w35521, w35522, w35523, w35524, w35525, w35526, w35527, w35528, w35529, w35530, w35531, w35532, w35533, w35534, w35535, w35536, w35537, w35538, w35539, w35540, w35541, w35542, w35543, w35544, w35545, w35546, w35547, w35548, w35549, w35550, w35551, w35552, w35553, w35554, w35555, w35556, w35557, w35558, w35559, w35560, w35561, w35562, w35563, w35564, w35565, w35566, w35567, w35568, w35569, w35570, w35571, w35572, w35573, w35574, w35575, w35576, w35577, w35578, w35579, w35580, w35581, w35582, w35583, w35584, w35585, w35586, w35587, w35588, w35589, w35590, w35591, w35592, w35593, w35594, w35595, w35596, w35597, w35598, w35599, w35600, w35601, w35602, w35603, w35604, w35605, w35606, w35607, w35608, w35609, w35610, w35611, w35612, w35613, w35614, w35615, w35616, w35617, w35618, w35619, w35620, w35621, w35622, w35623, w35624, w35625, w35626, w35627, w35628, w35629, w35630, w35631, w35632, w35633, w35634, w35635, w35636, w35637, w35638, w35639, w35640, w35641, w35642, w35643, w35644, w35645, w35646, w35647, w35648, w35649, w35650, w35651, w35652, w35653, w35654, w35655, w35656, w35657, w35658, w35659, w35660, w35661, w35662, w35663, w35664, w35665, w35666, w35667, w35668, w35669, w35670, w35671, w35672, w35673, w35674, w35675, w35676, w35677, w35678, w35679, w35680, w35681, w35682, w35683, w35684, w35685, w35686, w35687, w35688, w35689, w35690, w35691, w35692, w35693, w35694, w35695, w35696, w35697, w35698, w35699, w35700, w35701, w35702, w35703, w35704, w35705, w35706, w35707, w35708, w35709, w35710, w35711, w35712, w35713, w35714, w35715, w35716, w35717, w35718, w35719, w35720, w35721, w35722, w35723, w35724, w35725, w35726, w35727, w35728, w35729, w35730, w35731, w35732, w35733, w35734, w35735, w35736, w35737, w35738, w35739, w35740, w35741, w35742, w35743, w35744, w35745, w35746, w35747, w35748, w35749, w35750, w35751, w35752, w35753, w35754, w35755, w35756, w35757, w35758, w35759, w35760, w35761, w35762, w35763, w35764, w35765, w35766, w35767, w35768, w35769, w35770, w35771, w35772, w35773, w35774, w35775, w35776, w35777, w35778, w35779, w35780, w35781, w35782, w35783, w35784, w35785, w35786, w35787, w35788, w35789, w35790, w35791, w35792, w35793, w35794, w35795, w35796, w35797, w35798, w35799, w35800, w35801, w35802, w35803, w35804, w35805, w35806, w35807, w35808, w35809, w35810, w35811, w35812, w35813, w35814, w35815, w35816, w35817, w35818, w35819, w35820, w35821, w35822, w35823, w35824, w35825, w35826, w35827, w35828, w35829, w35830, w35831, w35832, w35833, w35834, w35835, w35836, w35837, w35838, w35839, w35840, w35841, w35842, w35843, w35844, w35845, w35846, w35847, w35848, w35849, w35850, w35851, w35852, w35853, w35854, w35855, w35856, w35857, w35858, w35859, w35860, w35861, w35862, w35863, w35864, w35865, w35866, w35867, w35868, w35869, w35870, w35871, w35872, w35873, w35874, w35875, w35876, w35877, w35878, w35879, w35880, w35881, w35882, w35883, w35884, w35885, w35886, w35887, w35888, w35889, w35890, w35891, w35892, w35893, w35894, w35895, w35896, w35897, w35898, w35899, w35900, w35901, w35902, w35903, w35904, w35905, w35906, w35907, w35908, w35909, w35910, w35911, w35912, w35913, w35914, w35915, w35916, w35917, w35918, w35919, w35920, w35921, w35922, w35923, w35924, w35925, w35926, w35927, w35928, w35929, w35930, w35931, w35932, w35933, w35934, w35935, w35936, w35937, w35938, w35939, w35940, w35941, w35942, w35943, w35944, w35945, w35946, w35947, w35948, w35949, w35950, w35951, w35952, w35953, w35954, w35955, w35956, w35957, w35958, w35959, w35960, w35961, w35962, w35963, w35964, w35965, w35966, w35967, w35968, w35969, w35970, w35971, w35972, w35973, w35974, w35975, w35976, w35977, w35978, w35979, w35980, w35981, w35982, w35983, w35984, w35985, w35986, w35987, w35988, w35989, w35990, w35991, w35992, w35993, w35994, w35995, w35996, w35997, w35998, w35999, w36000, w36001, w36002, w36003, w36004, w36005, w36006, w36007, w36008, w36009, w36010, w36011, w36012, w36013, w36014, w36015, w36016, w36017, w36018, w36019, w36020, w36021, w36022, w36023, w36024, w36025, w36026, w36027, w36028, w36029, w36030, w36031, w36032, w36033, w36034, w36035, w36036, w36037, w36038, w36039, w36040, w36041, w36042, w36043, w36044, w36045, w36046, w36047, w36048, w36049, w36050, w36051, w36052, w36053, w36054, w36055, w36056, w36057, w36058, w36059, w36060, w36061, w36062, w36063, w36064, w36065, w36066, w36067, w36068, w36069, w36070, w36071, w36072, w36073, w36074, w36075, w36076, w36077, w36078, w36079, w36080, w36081, w36082, w36083, w36084, w36085, w36086, w36087, w36088, w36089, w36090, w36091, w36092, w36093, w36094, w36095, w36096, w36097, w36098, w36099, w36100, w36101, w36102, w36103, w36104, w36105, w36106, w36107, w36108, w36109, w36110, w36111, w36112, w36113, w36114, w36115, w36116, w36117, w36118, w36119, w36120, w36121, w36122, w36123, w36124, w36125, w36126, w36127, w36128, w36129, w36130, w36131, w36132, w36133, w36134, w36135, w36136, w36137, w36138, w36139, w36140, w36141, w36142, w36143, w36144, w36145, w36146, w36147, w36148, w36149, w36150, w36151, w36152, w36153, w36154, w36155, w36156, w36157, w36158, w36159, w36160, w36161, w36162, w36163, w36164, w36165, w36166, w36167, w36168, w36169, w36170, w36171, w36172, w36173, w36174, w36175, w36176, w36177, w36178, w36179, w36180, w36181, w36182, w36183, w36184, w36185, w36186, w36187, w36188, w36189, w36190, w36191, w36192, w36193, w36194, w36195, w36196, w36197, w36198, w36199, w36200, w36201, w36202, w36203, w36204, w36205, w36206, w36207, w36208, w36209, w36210, w36211, w36212, w36213, w36214, w36215, w36216, w36217, w36218, w36219, w36220, w36221, w36222, w36223, w36224, w36225, w36226, w36227, w36228, w36229, w36230, w36231, w36232, w36233, w36234, w36235, w36236, w36237, w36238, w36239, w36240, w36241, w36242, w36243, w36244, w36245, w36246, w36247, w36248, w36249, w36250, w36251, w36252, w36253, w36254, w36255, w36256, w36257, w36258, w36259, w36260, w36261, w36262, w36263, w36264, w36265, w36266, w36267, w36268, w36269, w36270, w36271, w36272, w36273, w36274, w36275, w36276, w36277, w36278, w36279, w36280, w36281, w36282, w36283, w36284, w36285, w36286, w36287, w36288, w36289, w36290, w36291, w36292, w36293, w36294, w36295, w36296, w36297, w36298, w36299, w36300, w36301, w36302, w36303, w36304, w36305, w36306, w36307, w36308, w36309, w36310, w36311, w36312, w36313, w36314, w36315, w36316, w36317, w36318, w36319, w36320, w36321, w36322, w36323, w36324, w36325, w36326, w36327, w36328, w36329, w36330, w36331, w36332, w36333, w36334, w36335, w36336, w36337, w36338, w36339, w36340, w36341, w36342, w36343, w36344, w36345, w36346, w36347, w36348, w36349, w36350, w36351, w36352, w36353, w36354, w36355, w36356, w36357, w36358, w36359, w36360, w36361, w36362, w36363, w36364, w36365, w36366, w36367, w36368, w36369, w36370, w36371, w36372, w36373, w36374, w36375, w36376, w36377, w36378, w36379, w36380, w36381, w36382, w36383, w36384, w36385, w36386, w36387, w36388, w36389, w36390, w36391, w36392, w36393, w36394, w36395, w36396, w36397, w36398, w36399, w36400, w36401, w36402, w36403, w36404, w36405, w36406, w36407, w36408, w36409, w36410, w36411, w36412, w36413, w36414, w36415, w36416, w36417, w36418, w36419, w36420, w36421, w36422, w36423, w36424, w36425, w36426, w36427, w36428, w36429, w36430, w36431, w36432, w36433, w36434, w36435, w36436, w36437, w36438, w36439, w36440, w36441, w36442, w36443, w36444, w36445, w36446, w36447, w36448, w36449, w36450, w36451, w36452, w36453, w36454, w36455, w36456, w36457, w36458, w36459, w36460, w36461, w36462, w36463, w36464, w36465, w36466, w36467, w36468, w36469, w36470, w36471, w36472, w36473, w36474, w36475, w36476, w36477, w36478, w36479, w36480, w36481, w36482, w36483, w36484, w36485, w36486, w36487, w36488, w36489, w36490, w36491, w36492, w36493, w36494, w36495, w36496, w36497, w36498, w36499, w36500, w36501, w36502, w36503, w36504, w36505, w36506, w36507, w36508, w36509, w36510, w36511, w36512, w36513, w36514, w36515, w36516, w36517, w36518, w36519, w36520, w36521, w36522, w36523, w36524, w36525, w36526, w36527, w36528, w36529, w36530, w36531, w36532, w36533, w36534, w36535, w36536, w36537, w36538, w36539, w36540, w36541, w36542, w36543, w36544, w36545, w36546, w36547, w36548, w36549, w36550, w36551, w36552, w36553, w36554, w36555, w36556, w36557, w36558, w36559, w36560, w36561, w36562, w36563, w36564, w36565, w36566, w36567, w36568, w36569, w36570, w36571, w36572, w36573, w36574, w36575, w36576, w36577, w36578, w36579, w36580, w36581, w36582, w36583, w36584, w36585, w36586, w36587, w36588, w36589, w36590, w36591, w36592, w36593, w36594, w36595, w36596, w36597, w36598, w36599, w36600, w36601, w36602, w36603, w36604, w36605, w36606, w36607, w36608, w36609, w36610, w36611, w36612, w36613, w36614, w36615, w36616, w36617, w36618, w36619, w36620, w36621, w36622, w36623, w36624, w36625, w36626, w36627, w36628, w36629, w36630, w36631, w36632, w36633, w36634, w36635, w36636, w36637, w36638, w36639, w36640, w36641, w36642, w36643, w36644, w36645, w36646, w36647, w36648, w36649, w36650, w36651, w36652, w36653, w36654, w36655, w36656, w36657, w36658, w36659, w36660, w36661, w36662, w36663, w36664, w36665, w36666, w36667, w36668, w36669, w36670, w36671, w36672, w36673, w36674, w36675, w36676, w36677, w36678, w36679, w36680, w36681, w36682, w36683, w36684, w36685, w36686, w36687, w36688, w36689, w36690, w36691, w36692, w36693, w36694, w36695, w36696, w36697, w36698, w36699, w36700, w36701, w36702, w36703, w36704, w36705, w36706, w36707, w36708, w36709, w36710, w36711, w36712, w36713, w36714, w36715, w36716, w36717, w36718, w36719, w36720, w36721, w36722, w36723, w36724, w36725, w36726, w36727, w36728, w36729, w36730, w36731, w36732, w36733, w36734, w36735, w36736, w36737, w36738, w36739, w36740, w36741, w36742, w36743, w36744, w36745, w36746, w36747, w36748, w36749, w36750, w36751, w36752, w36753, w36754, w36755, w36756, w36757, w36758, w36759, w36760, w36761, w36762, w36763, w36764, w36765, w36766, w36767, w36768, w36769, w36770, w36771, w36772, w36773, w36774, w36775, w36776, w36777, w36778, w36779, w36780, w36781, w36782, w36783, w36784, w36785, w36786, w36787, w36788, w36789, w36790, w36791, w36792, w36793, w36794, w36795, w36796, w36797, w36798, w36799, w36800, w36801, w36802, w36803, w36804, w36805, w36806, w36807, w36808, w36809, w36810, w36811, w36812, w36813, w36814, w36815, w36816, w36817, w36818, w36819, w36820, w36821, w36822, w36823, w36824, w36825, w36826, w36827, w36828, w36829, w36830, w36831, w36832, w36833, w36834, w36835, w36836, w36837, w36838, w36839, w36840, w36841, w36842, w36843, w36844, w36845, w36846, w36847, w36848, w36849, w36850, w36851, w36852, w36853, w36854, w36855, w36856, w36857, w36858, w36859, w36860, w36861, w36862, w36863, w36864, w36865, w36866, w36867, w36868, w36869, w36870, w36871, w36872, w36873, w36874, w36875, w36876, w36877, w36878, w36879, w36880, w36881, w36882, w36883, w36884, w36885, w36886, w36887, w36888, w36889, w36890, w36891, w36892, w36893, w36894, w36895, w36896, w36897, w36898, w36899, w36900, w36901, w36902, w36903, w36904, w36905, w36906, w36907, w36908, w36909, w36910, w36911, w36912, w36913, w36914, w36915, w36916, w36917, w36918, w36919, w36920, w36921, w36922, w36923, w36924, w36925, w36926, w36927, w36928, w36929, w36930, w36931, w36932, w36933, w36934, w36935, w36936, w36937, w36938, w36939, w36940, w36941, w36942, w36943, w36944, w36945, w36946, w36947, w36948, w36949, w36950, w36951, w36952, w36953, w36954, w36955, w36956, w36957, w36958, w36959, w36960, w36961, w36962, w36963, w36964, w36965, w36966, w36967, w36968, w36969, w36970, w36971, w36972, w36973, w36974, w36975, w36976, w36977, w36978, w36979, w36980, w36981, w36982, w36983, w36984, w36985, w36986, w36987, w36988, w36989, w36990, w36991, w36992, w36993, w36994, w36995, w36996, w36997, w36998, w36999, w37000, w37001, w37002, w37003, w37004, w37005, w37006, w37007, w37008, w37009, w37010, w37011, w37012, w37013, w37014, w37015, w37016, w37017, w37018, w37019, w37020, w37021, w37022, w37023, w37024, w37025, w37026, w37027, w37028, w37029, w37030, w37031, w37032, w37033, w37034, w37035, w37036, w37037, w37038, w37039, w37040, w37041, w37042, w37043, w37044, w37045, w37046, w37047, w37048, w37049, w37050, w37051, w37052, w37053, w37054, w37055, w37056, w37057, w37058, w37059, w37060, w37061, w37062, w37063, w37064, w37065, w37066, w37067, w37068, w37069, w37070, w37071, w37072, w37073, w37074, w37075, w37076, w37077, w37078, w37079, w37080, w37081, w37082, w37083, w37084, w37085, w37086, w37087, w37088, w37089, w37090, w37091, w37092, w37093, w37094, w37095, w37096, w37097, w37098, w37099, w37100, w37101, w37102, w37103, w37104, w37105, w37106, w37107, w37108, w37109, w37110, w37111, w37112, w37113, w37114, w37115, w37116, w37117, w37118, w37119, w37120, w37121, w37122, w37123, w37124, w37125, w37126, w37127, w37128, w37129, w37130, w37131, w37132, w37133, w37134, w37135, w37136, w37137, w37138, w37139, w37140, w37141, w37142, w37143, w37144, w37145, w37146, w37147, w37148, w37149, w37150, w37151, w37152, w37153, w37154, w37155, w37156, w37157, w37158, w37159, w37160, w37161, w37162, w37163, w37164, w37165, w37166, w37167, w37168, w37169, w37170, w37171, w37172, w37173, w37174, w37175, w37176, w37177, w37178, w37179, w37180, w37181, w37182, w37183, w37184, w37185, w37186, w37187, w37188, w37189, w37190, w37191, w37192, w37193, w37194, w37195, w37196, w37197, w37198, w37199, w37200, w37201, w37202, w37203, w37204, w37205, w37206, w37207, w37208, w37209, w37210, w37211, w37212, w37213, w37214, w37215, w37216, w37217, w37218, w37219, w37220, w37221, w37222, w37223, w37224, w37225, w37226, w37227, w37228, w37229, w37230, w37231, w37232, w37233, w37234, w37235, w37236, w37237, w37238, w37239, w37240, w37241, w37242, w37243, w37244, w37245, w37246, w37247, w37248, w37249, w37250, w37251, w37252, w37253, w37254, w37255, w37256, w37257, w37258, w37259, w37260, w37261, w37262, w37263, w37264, w37265, w37266, w37267, w37268, w37269, w37270, w37271, w37272, w37273, w37274, w37275, w37276, w37277, w37278, w37279, w37280, w37281, w37282, w37283, w37284, w37285, w37286, w37287, w37288, w37289, w37290, w37291, w37292, w37293, w37294, w37295, w37296, w37297, w37298, w37299, w37300, w37301, w37302, w37303, w37304, w37305, w37306, w37307, w37308, w37309, w37310, w37311, w37312, w37313, w37314, w37315, w37316, w37317, w37318, w37319, w37320, w37321, w37322, w37323, w37324, w37325, w37326, w37327, w37328, w37329, w37330, w37331, w37332, w37333, w37334, w37335, w37336, w37337, w37338, w37339, w37340, w37341, w37342, w37343, w37344, w37345, w37346, w37347, w37348, w37349, w37350, w37351, w37352, w37353, w37354, w37355, w37356, w37357, w37358, w37359, w37360, w37361, w37362, w37363, w37364, w37365, w37366, w37367, w37368, w37369, w37370, w37371, w37372, w37373, w37374, w37375, w37376, w37377, w37378, w37379, w37380, w37381, w37382, w37383, w37384, w37385, w37386, w37387, w37388, w37389, w37390, w37391, w37392, w37393, w37394, w37395, w37396, w37397, w37398, w37399, w37400, w37401, w37402, w37403, w37404, w37405, w37406, w37407, w37408, w37409, w37410, w37411, w37412, w37413, w37414, w37415, w37416, w37417, w37418, w37419, w37420, w37421, w37422, w37423, w37424, w37425, w37426, w37427, w37428, w37429, w37430, w37431, w37432, w37433, w37434, w37435, w37436, w37437, w37438, w37439, w37440, w37441, w37442, w37443, w37444, w37445, w37446, w37447, w37448, w37449, w37450, w37451, w37452, w37453, w37454, w37455, w37456, w37457, w37458, w37459, w37460, w37461, w37462, w37463, w37464, w37465, w37466, w37467, w37468, w37469, w37470, w37471, w37472, w37473, w37474, w37475, w37476, w37477, w37478, w37479, w37480, w37481, w37482, w37483, w37484, w37485, w37486, w37487, w37488, w37489, w37490, w37491, w37492, w37493, w37494, w37495, w37496, w37497, w37498, w37499, w37500, w37501, w37502, w37503, w37504, w37505, w37506, w37507, w37508, w37509, w37510, w37511, w37512, w37513, w37514, w37515, w37516, w37517, w37518, w37519, w37520, w37521, w37522, w37523, w37524, w37525, w37526, w37527, w37528, w37529, w37530, w37531, w37532, w37533, w37534, w37535, w37536, w37537, w37538, w37539, w37540, w37541, w37542, w37543, w37544, w37545, w37546, w37547, w37548, w37549, w37550, w37551, w37552, w37553, w37554, w37555, w37556, w37557, w37558, w37559, w37560, w37561, w37562, w37563, w37564, w37565, w37566, w37567, w37568, w37569, w37570, w37571, w37572, w37573, w37574, w37575, w37576, w37577, w37578, w37579, w37580, w37581, w37582, w37583, w37584, w37585, w37586, w37587, w37588, w37589, w37590, w37591, w37592, w37593, w37594, w37595, w37596, w37597, w37598, w37599, w37600, w37601, w37602, w37603, w37604, w37605, w37606, w37607, w37608, w37609, w37610, w37611, w37612, w37613, w37614, w37615, w37616, w37617, w37618, w37619, w37620, w37621, w37622, w37623, w37624, w37625, w37626, w37627, w37628, w37629, w37630, w37631, w37632, w37633, w37634, w37635, w37636, w37637, w37638, w37639, w37640, w37641, w37642, w37643, w37644, w37645, w37646, w37647, w37648, w37649, w37650, w37651, w37652, w37653, w37654, w37655, w37656, w37657, w37658, w37659, w37660, w37661, w37662, w37663, w37664, w37665, w37666, w37667, w37668, w37669, w37670, w37671, w37672, w37673, w37674, w37675, w37676, w37677, w37678, w37679, w37680, w37681, w37682, w37683, w37684, w37685, w37686, w37687, w37688, w37689, w37690, w37691, w37692, w37693, w37694, w37695, w37696, w37697, w37698, w37699, w37700, w37701, w37702, w37703, w37704, w37705, w37706, w37707, w37708, w37709, w37710, w37711, w37712, w37713, w37714, w37715, w37716, w37717, w37718, w37719, w37720, w37721, w37722, w37723, w37724, w37725, w37726, w37727, w37728, w37729, w37730, w37731, w37732, w37733, w37734, w37735, w37736, w37737, w37738, w37739, w37740, w37741, w37742, w37743, w37744, w37745, w37746, w37747, w37748, w37749, w37750, w37751, w37752, w37753, w37754, w37755, w37756, w37757, w37758, w37759, w37760, w37761, w37762, w37763, w37764, w37765, w37766, w37767, w37768, w37769, w37770, w37771, w37772, w37773, w37774, w37775, w37776, w37777, w37778, w37779, w37780, w37781, w37782, w37783, w37784, w37785, w37786, w37787, w37788, w37789, w37790, w37791, w37792, w37793, w37794, w37795, w37796, w37797, w37798, w37799, w37800, w37801, w37802, w37803, w37804, w37805, w37806, w37807, w37808, w37809, w37810, w37811, w37812, w37813, w37814, w37815, w37816, w37817, w37818, w37819, w37820, w37821, w37822, w37823, w37824, w37825, w37826, w37827, w37828, w37829, w37830, w37831, w37832, w37833, w37834, w37835, w37836, w37837, w37838, w37839, w37840, w37841, w37842, w37843, w37844, w37845, w37846, w37847, w37848, w37849, w37850, w37851, w37852, w37853, w37854, w37855, w37856, w37857, w37858, w37859, w37860, w37861, w37862, w37863, w37864, w37865, w37866, w37867, w37868, w37869, w37870, w37871, w37872, w37873, w37874, w37875, w37876, w37877, w37878, w37879, w37880, w37881, w37882, w37883, w37884, w37885, w37886, w37887, w37888, w37889, w37890, w37891, w37892, w37893, w37894, w37895, w37896, w37897, w37898, w37899, w37900, w37901, w37902, w37903, w37904, w37905, w37906, w37907, w37908, w37909, w37910, w37911, w37912, w37913, w37914, w37915, w37916, w37917, w37918, w37919, w37920, w37921, w37922, w37923, w37924, w37925, w37926, w37927, w37928, w37929, w37930, w37931, w37932, w37933, w37934, w37935, w37936, w37937, w37938, w37939, w37940, w37941, w37942, w37943, w37944, w37945, w37946, w37947, w37948, w37949, w37950, w37951, w37952, w37953, w37954, w37955, w37956, w37957, w37958, w37959, w37960, w37961, w37962, w37963, w37964, w37965, w37966, w37967, w37968, w37969, w37970, w37971, w37972, w37973, w37974, w37975, w37976, w37977, w37978, w37979, w37980, w37981, w37982, w37983, w37984, w37985, w37986, w37987, w37988, w37989, w37990, w37991, w37992, w37993, w37994, w37995, w37996, w37997, w37998, w37999, w38000, w38001, w38002, w38003, w38004, w38005, w38006, w38007, w38008, w38009, w38010, w38011, w38012, w38013, w38014, w38015, w38016, w38017, w38018, w38019, w38020, w38021, w38022, w38023, w38024, w38025, w38026, w38027, w38028, w38029, w38030, w38031, w38032, w38033, w38034, w38035, w38036, w38037, w38038, w38039, w38040, w38041, w38042, w38043, w38044, w38045, w38046, w38047, w38048, w38049, w38050, w38051, w38052, w38053, w38054, w38055, w38056, w38057, w38058, w38059, w38060, w38061, w38062, w38063, w38064, w38065, w38066, w38067, w38068, w38069, w38070, w38071, w38072, w38073, w38074, w38075, w38076, w38077, w38078, w38079, w38080, w38081, w38082, w38083, w38084, w38085, w38086, w38087, w38088, w38089, w38090, w38091, w38092, w38093, w38094, w38095, w38096, w38097, w38098, w38099, w38100, w38101, w38102, w38103, w38104, w38105, w38106, w38107, w38108, w38109, w38110, w38111, w38112, w38113, w38114, w38115, w38116, w38117, w38118, w38119, w38120, w38121, w38122, w38123, w38124, w38125, w38126, w38127, w38128, w38129, w38130, w38131, w38132, w38133, w38134, w38135, w38136, w38137, w38138, w38139, w38140, w38141, w38142, w38143, w38144, w38145, w38146, w38147, w38148, w38149, w38150, w38151, w38152, w38153, w38154, w38155, w38156, w38157, w38158, w38159, w38160, w38161, w38162, w38163, w38164, w38165, w38166, w38167, w38168, w38169, w38170, w38171, w38172, w38173, w38174, w38175, w38176, w38177, w38178, w38179, w38180, w38181, w38182, w38183, w38184, w38185, w38186, w38187, w38188, w38189, w38190, w38191, w38192, w38193, w38194, w38195, w38196, w38197, w38198, w38199, w38200, w38201, w38202, w38203, w38204, w38205, w38206, w38207, w38208, w38209, w38210, w38211, w38212, w38213, w38214, w38215, w38216, w38217, w38218, w38219, w38220, w38221, w38222, w38223, w38224, w38225, w38226, w38227, w38228, w38229, w38230, w38231, w38232, w38233, w38234, w38235, w38236, w38237, w38238, w38239, w38240, w38241, w38242, w38243, w38244, w38245, w38246, w38247, w38248, w38249, w38250, w38251, w38252, w38253, w38254, w38255, w38256, w38257, w38258, w38259, w38260, w38261, w38262, w38263, w38264, w38265, w38266, w38267, w38268, w38269, w38270, w38271, w38272, w38273, w38274, w38275, w38276, w38277, w38278, w38279, w38280, w38281, w38282, w38283, w38284, w38285, w38286, w38287, w38288, w38289, w38290, w38291, w38292, w38293, w38294, w38295, w38296, w38297, w38298, w38299, w38300, w38301, w38302, w38303, w38304, w38305, w38306, w38307, w38308, w38309, w38310, w38311, w38312, w38313, w38314, w38315, w38316, w38317, w38318, w38319, w38320, w38321, w38322, w38323, w38324, w38325, w38326, w38327, w38328, w38329, w38330, w38331, w38332, w38333, w38334, w38335, w38336, w38337, w38338, w38339, w38340, w38341, w38342, w38343, w38344, w38345, w38346, w38347, w38348, w38349, w38350, w38351, w38352, w38353, w38354, w38355, w38356, w38357, w38358, w38359, w38360, w38361, w38362, w38363, w38364, w38365, w38366, w38367, w38368, w38369, w38370, w38371, w38372, w38373, w38374, w38375, w38376, w38377, w38378, w38379, w38380, w38381, w38382, w38383, w38384, w38385, w38386, w38387, w38388, w38389, w38390, w38391, w38392, w38393, w38394, w38395, w38396, w38397, w38398, w38399, w38400, w38401, w38402, w38403, w38404, w38405, w38406, w38407, w38408, w38409, w38410, w38411, w38412, w38413, w38414, w38415, w38416, w38417, w38418, w38419, w38420, w38421, w38422, w38423, w38424, w38425, w38426, w38427, w38428, w38429, w38430, w38431, w38432, w38433, w38434, w38435, w38436, w38437, w38438, w38439, w38440, w38441, w38442, w38443, w38444, w38445, w38446, w38447, w38448, w38449, w38450, w38451, w38452, w38453, w38454, w38455, w38456, w38457, w38458, w38459, w38460, w38461, w38462, w38463, w38464, w38465, w38466, w38467, w38468, w38469, w38470, w38471, w38472, w38473, w38474, w38475, w38476, w38477, w38478, w38479, w38480, w38481, w38482, w38483, w38484, w38485, w38486, w38487, w38488, w38489, w38490, w38491, w38492, w38493, w38494, w38495, w38496, w38497, w38498, w38499, w38500, w38501, w38502, w38503, w38504, w38505, w38506, w38507, w38508, w38509, w38510, w38511, w38512, w38513, w38514, w38515, w38516, w38517, w38518, w38519, w38520, w38521, w38522, w38523, w38524, w38525, w38526, w38527, w38528, w38529, w38530, w38531, w38532, w38533, w38534, w38535, w38536, w38537, w38538, w38539, w38540, w38541, w38542, w38543, w38544, w38545, w38546, w38547, w38548, w38549, w38550, w38551, w38552, w38553, w38554, w38555, w38556, w38557, w38558, w38559, w38560, w38561, w38562, w38563, w38564, w38565, w38566, w38567, w38568, w38569, w38570, w38571, w38572, w38573, w38574, w38575, w38576, w38577, w38578, w38579, w38580, w38581, w38582, w38583, w38584, w38585, w38586, w38587, w38588, w38589, w38590, w38591, w38592, w38593, w38594, w38595, w38596, w38597, w38598, w38599, w38600, w38601, w38602, w38603, w38604, w38605, w38606, w38607, w38608, w38609, w38610, w38611, w38612, w38613, w38614, w38615, w38616, w38617, w38618, w38619, w38620, w38621, w38622, w38623, w38624, w38625, w38626, w38627, w38628, w38629, w38630, w38631, w38632, w38633, w38634, w38635, w38636, w38637, w38638, w38639, w38640, w38641, w38642, w38643, w38644, w38645, w38646, w38647, w38648, w38649, w38650, w38651, w38652, w38653, w38654, w38655, w38656, w38657, w38658, w38659, w38660, w38661, w38662, w38663, w38664, w38665, w38666, w38667, w38668, w38669, w38670, w38671, w38672, w38673, w38674, w38675, w38676, w38677, w38678, w38679, w38680, w38681, w38682, w38683, w38684, w38685, w38686, w38687, w38688, w38689, w38690, w38691, w38692, w38693, w38694, w38695, w38696, w38697, w38698, w38699, w38700, w38701, w38702, w38703, w38704, w38705, w38706, w38707, w38708, w38709, w38710, w38711, w38712, w38713, w38714, w38715, w38716, w38717, w38718, w38719, w38720, w38721, w38722, w38723, w38724, w38725, w38726, w38727, w38728, w38729, w38730, w38731, w38732, w38733, w38734, w38735, w38736, w38737, w38738, w38739, w38740, w38741, w38742, w38743, w38744, w38745, w38746, w38747, w38748, w38749, w38750, w38751, w38752, w38753, w38754, w38755, w38756, w38757, w38758, w38759, w38760, w38761, w38762, w38763, w38764, w38765, w38766, w38767, w38768, w38769, w38770, w38771, w38772, w38773, w38774, w38775, w38776, w38777, w38778, w38779, w38780, w38781, w38782, w38783, w38784, w38785, w38786, w38787, w38788, w38789, w38790, w38791, w38792, w38793, w38794, w38795, w38796, w38797, w38798, w38799, w38800, w38801, w38802, w38803, w38804, w38805, w38806, w38807, w38808, w38809, w38810, w38811, w38812, w38813, w38814, w38815, w38816, w38817, w38818, w38819, w38820, w38821, w38822, w38823, w38824, w38825, w38826, w38827, w38828, w38829, w38830, w38831, w38832, w38833, w38834, w38835, w38836, w38837, w38838, w38839, w38840, w38841, w38842, w38843, w38844, w38845, w38846, w38847, w38848, w38849, w38850, w38851, w38852, w38853, w38854, w38855, w38856, w38857, w38858, w38859, w38860, w38861, w38862, w38863, w38864, w38865, w38866, w38867, w38868, w38869, w38870, w38871, w38872, w38873, w38874, w38875, w38876, w38877, w38878, w38879, w38880, w38881, w38882, w38883, w38884, w38885, w38886, w38887, w38888, w38889, w38890, w38891, w38892, w38893, w38894, w38895, w38896, w38897, w38898, w38899, w38900, w38901, w38902, w38903, w38904, w38905, w38906, w38907, w38908, w38909, w38910, w38911, w38912, w38913, w38914, w38915, w38916, w38917, w38918, w38919, w38920, w38921, w38922, w38923, w38924, w38925, w38926, w38927, w38928, w38929, w38930, w38931, w38932, w38933, w38934, w38935, w38936, w38937, w38938, w38939, w38940, w38941, w38942, w38943, w38944, w38945, w38946, w38947, w38948, w38949, w38950, w38951, w38952, w38953, w38954, w38955, w38956, w38957, w38958, w38959, w38960, w38961, w38962, w38963, w38964, w38965, w38966, w38967, w38968, w38969, w38970, w38971, w38972, w38973, w38974, w38975, w38976, w38977, w38978, w38979, w38980, w38981, w38982, w38983, w38984, w38985, w38986, w38987, w38988, w38989, w38990, w38991, w38992, w38993, w38994, w38995, w38996, w38997, w38998, w38999, w39000, w39001, w39002, w39003, w39004, w39005, w39006, w39007, w39008, w39009, w39010, w39011, w39012, w39013, w39014, w39015, w39016, w39017, w39018, w39019, w39020, w39021, w39022, w39023, w39024, w39025, w39026, w39027, w39028, w39029, w39030, w39031, w39032, w39033, w39034, w39035, w39036, w39037, w39038, w39039, w39040, w39041, w39042, w39043, w39044, w39045, w39046, w39047, w39048, w39049, w39050, w39051, w39052, w39053, w39054, w39055, w39056, w39057, w39058, w39059, w39060, w39061, w39062, w39063, w39064, w39065, w39066, w39067, w39068, w39069, w39070, w39071, w39072, w39073, w39074, w39075, w39076, w39077, w39078, w39079, w39080, w39081, w39082, w39083, w39084, w39085, w39086, w39087, w39088, w39089, w39090, w39091, w39092, w39093, w39094, w39095, w39096, w39097, w39098, w39099, w39100, w39101, w39102, w39103, w39104, w39105, w39106, w39107, w39108, w39109, w39110, w39111, w39112, w39113, w39114, w39115, w39116, w39117, w39118, w39119, w39120, w39121, w39122, w39123, w39124, w39125, w39126, w39127, w39128, w39129, w39130, w39131, w39132, w39133, w39134, w39135, w39136, w39137, w39138, w39139, w39140, w39141, w39142, w39143, w39144, w39145, w39146, w39147, w39148, w39149, w39150, w39151, w39152, w39153, w39154, w39155, w39156, w39157, w39158, w39159, w39160, w39161, w39162, w39163, w39164, w39165, w39166, w39167, w39168, w39169, w39170, w39171, w39172, w39173, w39174, w39175, w39176, w39177, w39178, w39179, w39180, w39181, w39182, w39183, w39184, w39185, w39186, w39187, w39188, w39189, w39190, w39191, w39192, w39193, w39194, w39195, w39196, w39197, w39198, w39199, w39200, w39201, w39202, w39203, w39204, w39205, w39206, w39207, w39208, w39209, w39210, w39211, w39212, w39213, w39214, w39215, w39216, w39217, w39218, w39219, w39220, w39221, w39222, w39223, w39224, w39225, w39226, w39227, w39228, w39229, w39230, w39231, w39232, w39233, w39234, w39235, w39236, w39237, w39238, w39239, w39240, w39241, w39242, w39243, w39244, w39245, w39246, w39247, w39248, w39249, w39250, w39251, w39252, w39253, w39254, w39255, w39256, w39257, w39258, w39259, w39260, w39261, w39262, w39263, w39264, w39265, w39266, w39267, w39268, w39269, w39270, w39271, w39272, w39273, w39274, w39275, w39276, w39277, w39278, w39279, w39280, w39281, w39282, w39283, w39284, w39285, w39286, w39287, w39288, w39289, w39290, w39291, w39292, w39293, w39294, w39295, w39296, w39297, w39298, w39299, w39300, w39301, w39302, w39303, w39304, w39305, w39306, w39307, w39308, w39309, w39310, w39311, w39312, w39313, w39314, w39315, w39316, w39317, w39318, w39319, w39320, w39321, w39322, w39323, w39324, w39325, w39326, w39327, w39328, w39329, w39330, w39331, w39332, w39333, w39334, w39335, w39336, w39337, w39338, w39339, w39340, w39341, w39342, w39343, w39344, w39345, w39346, w39347, w39348, w39349, w39350, w39351, w39352, w39353, w39354, w39355, w39356, w39357, w39358, w39359, w39360, w39361, w39362, w39363, w39364, w39365, w39366, w39367, w39368, w39369, w39370, w39371, w39372, w39373, w39374, w39375, w39376, w39377, w39378, w39379, w39380, w39381, w39382, w39383, w39384, w39385, w39386, w39387, w39388, w39389, w39390, w39391, w39392, w39393, w39394, w39395, w39396, w39397, w39398, w39399, w39400, w39401, w39402, w39403, w39404, w39405, w39406, w39407, w39408, w39409, w39410, w39411, w39412, w39413, w39414, w39415, w39416, w39417, w39418, w39419, w39420, w39421, w39422, w39423, w39424, w39425, w39426, w39427, w39428, w39429, w39430, w39431, w39432, w39433, w39434, w39435, w39436, w39437, w39438, w39439, w39440, w39441, w39442, w39443, w39444, w39445, w39446, w39447, w39448, w39449, w39450, w39451, w39452, w39453, w39454, w39455, w39456, w39457, w39458, w39459, w39460, w39461, w39462, w39463, w39464, w39465, w39466, w39467, w39468, w39469, w39470, w39471, w39472, w39473, w39474, w39475, w39476, w39477, w39478, w39479, w39480, w39481, w39482, w39483, w39484, w39485, w39486, w39487, w39488, w39489, w39490, w39491, w39492, w39493, w39494, w39495, w39496, w39497, w39498, w39499, w39500, w39501, w39502, w39503, w39504, w39505, w39506, w39507, w39508, w39509, w39510, w39511, w39512, w39513, w39514, w39515, w39516, w39517, w39518, w39519, w39520, w39521, w39522, w39523, w39524, w39525, w39526, w39527, w39528, w39529, w39530, w39531, w39532, w39533, w39534, w39535, w39536, w39537, w39538, w39539, w39540, w39541, w39542, w39543, w39544, w39545, w39546, w39547, w39548, w39549, w39550, w39551, w39552, w39553, w39554, w39555, w39556, w39557, w39558, w39559, w39560, w39561, w39562, w39563, w39564, w39565, w39566, w39567, w39568, w39569, w39570, w39571, w39572, w39573, w39574, w39575, w39576, w39577, w39578, w39579, w39580, w39581, w39582, w39583, w39584, w39585, w39586, w39587, w39588, w39589, w39590, w39591, w39592, w39593, w39594, w39595, w39596, w39597, w39598, w39599, w39600, w39601, w39602, w39603, w39604, w39605, w39606, w39607, w39608, w39609, w39610, w39611, w39612, w39613, w39614, w39615, w39616, w39617, w39618, w39619, w39620, w39621, w39622, w39623, w39624, w39625, w39626, w39627, w39628, w39629, w39630, w39631, w39632, w39633, w39634, w39635, w39636, w39637, w39638, w39639, w39640, w39641, w39642, w39643, w39644, w39645, w39646, w39647, w39648, w39649, w39650, w39651, w39652, w39653, w39654, w39655, w39656, w39657, w39658, w39659, w39660, w39661, w39662, w39663, w39664, w39665, w39666, w39667, w39668, w39669, w39670, w39671, w39672, w39673, w39674, w39675, w39676, w39677, w39678, w39679, w39680, w39681, w39682, w39683, w39684, w39685, w39686, w39687, w39688, w39689, w39690, w39691, w39692, w39693, w39694, w39695, w39696, w39697, w39698, w39699, w39700, w39701, w39702, w39703, w39704, w39705, w39706, w39707, w39708, w39709, w39710, w39711, w39712, w39713, w39714, w39715, w39716, w39717, w39718, w39719, w39720, w39721, w39722, w39723, w39724, w39725, w39726, w39727, w39728, w39729, w39730, w39731, w39732, w39733, w39734, w39735, w39736, w39737, w39738, w39739, w39740, w39741, w39742, w39743, w39744, w39745, w39746, w39747, w39748, w39749, w39750, w39751, w39752, w39753, w39754, w39755, w39756, w39757, w39758, w39759, w39760, w39761, w39762, w39763, w39764, w39765, w39766, w39767, w39768, w39769, w39770, w39771, w39772, w39773, w39774, w39775, w39776, w39777, w39778, w39779, w39780, w39781, w39782, w39783, w39784, w39785, w39786, w39787, w39788, w39789, w39790, w39791, w39792, w39793, w39794, w39795, w39796, w39797, w39798, w39799, w39800, w39801, w39802, w39803, w39804, w39805, w39806, w39807, w39808, w39809, w39810, w39811, w39812, w39813, w39814, w39815, w39816, w39817, w39818, w39819, w39820, w39821, w39822, w39823, w39824, w39825, w39826, w39827, w39828, w39829, w39830, w39831, w39832, w39833, w39834, w39835, w39836, w39837, w39838, w39839, w39840, w39841, w39842, w39843, w39844, w39845, w39846, w39847, w39848, w39849, w39850, w39851, w39852, w39853, w39854, w39855, w39856, w39857, w39858, w39859, w39860, w39861, w39862, w39863, w39864, w39865, w39866, w39867, w39868, w39869, w39870, w39871, w39872, w39873, w39874, w39875, w39876, w39877, w39878, w39879, w39880, w39881, w39882, w39883, w39884, w39885, w39886, w39887, w39888, w39889, w39890, w39891, w39892, w39893, w39894, w39895, w39896, w39897, w39898, w39899, w39900, w39901, w39902, w39903, w39904, w39905, w39906, w39907, w39908, w39909, w39910, w39911, w39912, w39913, w39914, w39915, w39916, w39917, w39918, w39919, w39920, w39921, w39922, w39923, w39924, w39925, w39926, w39927, w39928, w39929, w39930, w39931, w39932, w39933, w39934, w39935, w39936, w39937, w39938, w39939, w39940, w39941, w39942, w39943, w39944, w39945, w39946, w39947, w39948, w39949, w39950, w39951, w39952, w39953, w39954, w39955, w39956, w39957, w39958, w39959, w39960, w39961, w39962, w39963, w39964, w39965, w39966, w39967, w39968, w39969, w39970, w39971, w39972, w39973, w39974, w39975, w39976, w39977, w39978, w39979, w39980, w39981, w39982, w39983, w39984, w39985, w39986, w39987, w39988, w39989, w39990, w39991, w39992, w39993, w39994, w39995, w39996, w39997, w39998, w39999, w40000, w40001, w40002, w40003, w40004, w40005, w40006, w40007, w40008, w40009, w40010, w40011, w40012, w40013, w40014, w40015, w40016, w40017, w40018, w40019, w40020, w40021, w40022, w40023, w40024, w40025, w40026, w40027, w40028, w40029, w40030, w40031, w40032, w40033, w40034, w40035, w40036, w40037, w40038, w40039, w40040, w40041, w40042, w40043, w40044, w40045, w40046, w40047, w40048, w40049, w40050, w40051, w40052, w40053, w40054, w40055, w40056, w40057, w40058, w40059, w40060, w40061, w40062, w40063, w40064, w40065, w40066, w40067, w40068, w40069, w40070, w40071, w40072, w40073, w40074, w40075, w40076, w40077, w40078, w40079, w40080, w40081, w40082, w40083, w40084, w40085, w40086, w40087, w40088, w40089, w40090, w40091, w40092, w40093, w40094, w40095, w40096, w40097, w40098, w40099, w40100, w40101, w40102, w40103, w40104, w40105, w40106, w40107, w40108, w40109, w40110, w40111, w40112, w40113, w40114, w40115, w40116, w40117, w40118, w40119, w40120, w40121, w40122, w40123, w40124, w40125, w40126, w40127, w40128, w40129, w40130, w40131, w40132, w40133, w40134, w40135, w40136, w40137, w40138, w40139, w40140, w40141, w40142, w40143, w40144, w40145, w40146, w40147, w40148, w40149, w40150, w40151, w40152, w40153, w40154, w40155, w40156, w40157, w40158, w40159, w40160, w40161, w40162, w40163, w40164, w40165, w40166, w40167, w40168, w40169, w40170, w40171, w40172, w40173, w40174, w40175, w40176, w40177, w40178, w40179, w40180, w40181, w40182, w40183, w40184, w40185, w40186, w40187, w40188, w40189, w40190, w40191, w40192, w40193, w40194, w40195, w40196, w40197, w40198, w40199, w40200, w40201, w40202, w40203, w40204, w40205, w40206, w40207, w40208, w40209, w40210, w40211;
assign w0 = pi3649 & pi3650;
assign w1 = pi3415 & w0;
assign w2 = pi0939 & w0;
assign w3 = pi2604 & w0;
assign w4 = ~pi3653 & pi3655;
assign w5 = ~pi3654 & ~pi3655;
assign w6 = ~w4 & ~w5;
assign w7 = ~w3 & w6;
assign w8 = w0 & w35533;
assign w9 = (~w8 & ~w7) | (~w8 & w35534) | (~w7 & w35534);
assign w10 = ~w1 & w9;
assign w11 = ~pi1835 & pi2386;
assign w12 = pi3294 & ~pi3324;
assign w13 = pi3322 & pi3323;
assign w14 = w12 & ~w13;
assign w15 = ~pi1776 & pi2825;
assign w16 = pi1776 & ~pi2825;
assign w17 = pi2114 & ~w16;
assign w18 = ~w15 & w17;
assign w19 = ~pi1462 & ~pi2785;
assign w20 = ~pi1928 & w19;
assign w21 = ~pi1462 & pi2785;
assign w22 = ~pi1780 & w21;
assign w23 = pi1462 & ~pi1772;
assign w24 = ~w22 & ~w23;
assign w25 = (pi2825 & ~w24) | (pi2825 & w35535) | (~w24 & w35535);
assign w26 = ~pi1785 & ~pi2799;
assign w27 = pi1785 & pi2799;
assign w28 = pi1462 & ~w27;
assign w29 = (~pi2114 & ~w28) | (~pi2114 & w35536) | (~w28 & w35536);
assign w30 = ~w25 & w29;
assign w31 = pi1945 & ~pi2785;
assign w32 = pi1779 & pi2785;
assign w33 = ~w31 & ~w32;
assign w34 = pi2799 & ~w33;
assign w35 = (~pi1462 & ~w33) | (~pi1462 & w35537) | (~w33 & w35537);
assign w36 = ~w34 & w35;
assign w37 = w24 & w35538;
assign w38 = ~w36 & ~w37;
assign w39 = w30 & w38;
assign w40 = ~w18 & ~w39;
assign w41 = pi1462 & ~pi1773;
assign w42 = ~pi1786 & w21;
assign w43 = (~pi2114 & w42) | (~pi2114 & w35539) | (w42 & w35539);
assign w44 = ~pi2114 & w19;
assign w45 = w19 & w35540;
assign w46 = ~pi1777 & pi2114;
assign w47 = ~w45 & ~w46;
assign w48 = ~w43 & w47;
assign w49 = ~pi2798 & w48;
assign w50 = ~pi1778 & w21;
assign w51 = pi1462 & ~pi1784;
assign w52 = (~pi2114 & w50) | (~pi2114 & w35541) | (w50 & w35541);
assign w53 = ~pi1774 & pi2114;
assign w54 = (~w53 & ~w44) | (~w53 & w35542) | (~w44 & w35542);
assign w55 = ~w52 & w54;
assign w56 = ~pi2600 & w55;
assign w57 = pi2798 & ~w48;
assign w58 = ~w56 & ~w57;
assign w59 = ~w49 & w58;
assign w60 = ~pi1941 & pi2114;
assign w61 = pi1943 & w21;
assign w62 = pi1462 & pi1939;
assign w63 = ~pi2114 & ~w62;
assign w64 = ~w61 & w63;
assign w65 = ~w64 & w35543;
assign w66 = ~pi1940 & pi2114;
assign w67 = pi1942 & w21;
assign w68 = pi1462 & pi1938;
assign w69 = ~pi2114 & ~w68;
assign w70 = ~w67 & w69;
assign w71 = (pi2113 & w70) | (pi2113 & w35544) | (w70 & w35544);
assign w72 = (pi2082 & w64) | (pi2082 & w35545) | (w64 & w35545);
assign w73 = ~w71 & ~w72;
assign w74 = ~w65 & w73;
assign w75 = pi2600 & ~w55;
assign w76 = ~w70 & w35546;
assign w77 = pi1775 & pi2799;
assign w78 = ~pi1775 & ~pi2799;
assign w79 = pi2114 & ~w78;
assign w80 = ~w77 & w79;
assign w81 = ~w76 & ~w80;
assign w82 = ~w75 & w81;
assign w83 = w74 & w82;
assign w84 = w59 & w83;
assign w85 = ~w40 & w84;
assign w86 = w84 & w35547;
assign w87 = pi1860 & w12;
assign w88 = ~pi3294 & pi3324;
assign w89 = ~pi3419 & w88;
assign w90 = ~w87 & ~w89;
assign w91 = w13 & ~w90;
assign w92 = pi0783 & ~pi3631;
assign w93 = ~pi3682 & w92;
assign w94 = pi3631 & pi3682;
assign w95 = ~w93 & ~w94;
assign w96 = ~pi3322 & ~pi3323;
assign w97 = ~pi3294 & ~pi3324;
assign w98 = ~pi2114 & ~pi2813;
assign w99 = w97 & w98;
assign w100 = w96 & w99;
assign w101 = w99 & w35548;
assign w102 = ~w95 & w101;
assign w103 = pi3324 & pi3682;
assign w104 = ~pi3322 & ~w103;
assign w105 = pi3322 & pi3324;
assign w106 = ~pi3294 & ~w105;
assign w107 = ~w104 & w106;
assign w108 = ~w102 & ~w107;
assign w109 = ~w91 & w108;
assign w110 = pi3322 & ~pi3323;
assign w111 = ~w12 & ~w88;
assign w112 = w110 & ~w111;
assign w113 = w108 & w35549;
assign w114 = ~w86 & w113;
assign w115 = ~pi3294 & w110;
assign w116 = w12 & w96;
assign w117 = ~pi1035 & pi2978;
assign w118 = pi3344 & w117;
assign w119 = w116 & w118;
assign w120 = ~w115 & ~w119;
assign w121 = w84 & w35550;
assign w122 = (w14 & ~w84) | (w14 & w35551) | (~w84 & w35551);
assign w123 = pi2504 & ~pi2759;
assign w124 = ~pi2505 & pi3281;
assign w125 = ~w123 & ~w124;
assign w126 = ~pi2049 & pi2503;
assign w127 = ~pi2522 & pi3199;
assign w128 = ~w126 & ~w127;
assign w129 = w125 & w128;
assign w130 = pi2049 & ~pi2503;
assign w131 = pi3099 & ~w130;
assign w132 = ~pi2505 & pi3343;
assign w133 = pi3281 & pi3343;
assign w134 = ~w132 & ~w133;
assign w135 = pi2522 & ~pi3199;
assign w136 = ~pi2504 & pi2759;
assign w137 = ~w135 & ~w136;
assign w138 = ~w134 & w137;
assign w139 = w131 & w138;
assign w140 = w129 & w139;
assign w141 = ~pi2522 & pi3281;
assign w142 = pi2522 & ~pi3281;
assign w143 = ~w141 & ~w142;
assign w144 = pi2505 & ~pi3343;
assign w145 = w143 & ~w144;
assign w146 = ~pi2503 & pi2759;
assign w147 = pi2503 & ~pi2759;
assign w148 = ~w146 & ~w147;
assign w149 = ~pi2504 & pi3199;
assign w150 = pi2504 & ~pi3199;
assign w151 = ~w149 & ~w150;
assign w152 = pi2049 & ~pi3099;
assign w153 = ~w132 & w152;
assign w154 = w151 & w153;
assign w155 = w148 & w154;
assign w156 = w145 & w155;
assign w157 = (pi3322 & ~w155) | (pi3322 & w35552) | (~w155 & w35552);
assign w158 = ~w140 & w157;
assign w159 = ~pi2813 & ~pi3322;
assign w160 = pi3631 & w159;
assign w161 = ~w44 & w160;
assign w162 = (~w161 & w158) | (~w161 & w35553) | (w158 & w35553);
assign w163 = w97 & ~w162;
assign w164 = ~w122 & ~w163;
assign w165 = ~w121 & w164;
assign w166 = w19 & ~w93;
assign w167 = ~pi3631 & ~w19;
assign w168 = w100 & ~w167;
assign w169 = ~w166 & w168;
assign w170 = pi3294 & ~pi3323;
assign w171 = pi3324 & ~w170;
assign w172 = ~pi3323 & ~pi3324;
assign w173 = pi3294 & pi3322;
assign w174 = ~w172 & ~w173;
assign w175 = ~w171 & w174;
assign w176 = ~w91 & ~w175;
assign w177 = ~w169 & w176;
assign w178 = ~w165 & w35554;
assign w179 = ~pi3322 & pi3323;
assign w180 = ~w111 & w179;
assign w181 = (pi1462 & w178) | (pi1462 & w35555) | (w178 & w35555);
assign w182 = (pi2785 & w178) | (pi2785 & w35556) | (w178 & w35556);
assign w183 = ~w181 & ~w182;
assign w184 = ~w165 & w35557;
assign w185 = w96 & ~w111;
assign w186 = ~w184 & ~w185;
assign w187 = ~pi3305 & pi3390;
assign w188 = pi3324 & ~w187;
assign w189 = (pi3626 & w188) | (pi3626 & w35558) | (w188 & w35558);
assign w190 = w186 & w189;
assign w191 = w183 & w190;
assign w192 = ~pi3452 & ~w191;
assign w193 = (w178 & w35559) | (w178 & w35560) | (w35559 & w35560);
assign w194 = (w178 & w35561) | (w178 & w35562) | (w35561 & w35562);
assign w195 = (pi1783 & w184) | (pi1783 & w35563) | (w184 & w35563);
assign w196 = ~w194 & ~w195;
assign w197 = ~w193 & w196;
assign w198 = pi1601 & ~pi3626;
assign w199 = pi3622 & pi3626;
assign w200 = ~w198 & ~w199;
assign w201 = ~pi3452 & pi3620;
assign w202 = pi3626 & ~w201;
assign w203 = pi3099 & ~pi3626;
assign w204 = ~w201 & ~w203;
assign w205 = pi0799 & ~pi3592;
assign w206 = ~pi0793 & ~pi3595;
assign w207 = pi0793 & pi3593;
assign w208 = pi0957 & ~w207;
assign w209 = ~w206 & w208;
assign w210 = ~pi0793 & ~pi3609;
assign w211 = pi0793 & ~pi3605;
assign w212 = ~pi0957 & ~w211;
assign w213 = (pi1009 & ~w212) | (pi1009 & w35564) | (~w212 & w35564);
assign w214 = ~w209 & w213;
assign w215 = pi0793 & ~pi3613;
assign w216 = ~pi0793 & ~pi3618;
assign w217 = ~pi0957 & ~w216;
assign w218 = ~w215 & w217;
assign w219 = ~pi0793 & ~pi3601;
assign w220 = pi0793 & ~pi3598;
assign w221 = pi0957 & ~w220;
assign w222 = (~pi1009 & ~w221) | (~pi1009 & w35565) | (~w221 & w35565);
assign w223 = ~w218 & w222;
assign w224 = ~w214 & ~w223;
assign w225 = ~pi0795 & ~w224;
assign w226 = ~pi0793 & ~pi3607;
assign w227 = pi0793 & ~pi3603;
assign w228 = ~pi0957 & ~w227;
assign w229 = ~w226 & w228;
assign w230 = ~pi0793 & ~pi3594;
assign w231 = pi0793 & pi3592;
assign w232 = pi0957 & ~w231;
assign w233 = ~w230 & w232;
assign w234 = ~w229 & ~w233;
assign w235 = pi1009 & ~w234;
assign w236 = pi0793 & ~pi3611;
assign w237 = ~pi0793 & ~pi3615;
assign w238 = ~pi0957 & ~w237;
assign w239 = ~w236 & w238;
assign w240 = ~pi0793 & ~pi3599;
assign w241 = pi0793 & ~pi3596;
assign w242 = pi0957 & ~w241;
assign w243 = ~w240 & w242;
assign w244 = ~w239 & ~w243;
assign w245 = (pi0795 & w244) | (pi0795 & w35566) | (w244 & w35566);
assign w246 = ~w235 & w245;
assign w247 = ~pi0799 & ~w246;
assign w248 = (~w205 & ~w247) | (~w205 & w35567) | (~w247 & w35567);
assign w249 = ~pi0958 & ~w248;
assign w250 = pi0893 & ~pi3461;
assign w251 = ~pi0885 & pi3604;
assign w252 = pi0885 & pi3471;
assign w253 = pi0741 & ~w252;
assign w254 = ~w251 & w253;
assign w255 = ~pi0885 & pi3606;
assign w256 = pi0885 & ~pi3597;
assign w257 = ~pi0741 & ~w256;
assign w258 = (pi0884 & ~w257) | (pi0884 & w35568) | (~w257 & w35568);
assign w259 = ~w254 & w258;
assign w260 = pi0885 & pi3614;
assign w261 = ~pi0885 & pi3623;
assign w262 = ~pi0741 & ~w261;
assign w263 = ~w260 & w262;
assign w264 = ~pi0885 & pi3619;
assign w265 = pi0885 & pi3612;
assign w266 = pi0741 & ~w265;
assign w267 = (~pi0884 & ~w266) | (~pi0884 & w35569) | (~w266 & w35569);
assign w268 = ~w263 & w267;
assign w269 = ~w259 & ~w268;
assign w270 = ~pi0739 & ~w269;
assign w271 = ~pi0885 & pi3602;
assign w272 = pi0885 & pi3473;
assign w273 = ~pi0741 & ~w272;
assign w274 = ~w271 & w273;
assign w275 = ~pi0885 & pi3600;
assign w276 = pi0885 & pi3461;
assign w277 = pi0741 & ~w276;
assign w278 = ~w275 & w277;
assign w279 = ~w274 & ~w278;
assign w280 = pi0884 & ~w279;
assign w281 = ~pi0885 & pi3617;
assign w282 = pi0885 & pi3610;
assign w283 = ~pi0741 & ~w282;
assign w284 = ~w281 & w283;
assign w285 = ~pi0885 & pi3616;
assign w286 = pi0885 & pi3608;
assign w287 = pi0741 & ~w286;
assign w288 = ~w285 & w287;
assign w289 = ~w284 & ~w288;
assign w290 = (pi0739 & w289) | (pi0739 & w35570) | (w289 & w35570);
assign w291 = ~w280 & w290;
assign w292 = ~pi0893 & ~w291;
assign w293 = (~w250 & ~w292) | (~w250 & w35571) | (~w292 & w35571);
assign w294 = ~pi0886 & w293;
assign w295 = ~pi0960 & pi1746;
assign w296 = pi0960 & ~pi1746;
assign w297 = ~w295 & ~w296;
assign w298 = ~pi0888 & pi1739;
assign w299 = pi0888 & ~pi1739;
assign w300 = ~w298 & ~w299;
assign w301 = ~pi0954 & pi1002;
assign w302 = pi0796 & pi0962;
assign w303 = pi0954 & ~pi1002;
assign w304 = ~w302 & ~w303;
assign w305 = ~w301 & w304;
assign w306 = ~pi0956 & pi1002;
assign w307 = pi0956 & ~pi1002;
assign w308 = ~w302 & ~w307;
assign w309 = ~w306 & w308;
assign w310 = ~pi0881 & pi1001;
assign w311 = pi0890 & pi0947;
assign w312 = pi0881 & ~pi1001;
assign w313 = ~w311 & ~w312;
assign w314 = ~w310 & w313;
assign w315 = ~pi0880 & pi1001;
assign w316 = pi0880 & ~pi1001;
assign w317 = ~w311 & ~w316;
assign w318 = ~w315 & w317;
assign w319 = ~pi2515 & ~pi3645;
assign w320 = ~pi3632 & ~pi3677;
assign w321 = ~pi0565 & pi3547;
assign w322 = pi2813 & pi3643;
assign w323 = ~w321 & ~w322;
assign w324 = ~pi3452 & pi3548;
assign w325 = ~pi3215 & pi3505;
assign w326 = ~pi3528 & ~w325;
assign w327 = ~pi0404 & ~pi0684;
assign w328 = ~pi3190 & ~pi3515;
assign w329 = w327 & w328;
assign w330 = ~pi3148 & w329;
assign w331 = (~w324 & ~w330) | (~w324 & w35572) | (~w330 & w35572);
assign w332 = ~pi3522 & ~pi3523;
assign w333 = ~pi0565 & w40088;
assign w334 = pi2813 & pi3526;
assign w335 = ~pi3416 & ~pi3583;
assign w336 = ~pi1046 & pi3416;
assign w337 = ~pi2800 & w336;
assign w338 = ~w335 & ~w337;
assign w339 = ~w337 & w35574;
assign w340 = ~w334 & ~w339;
assign w341 = ~w333 & w340;
assign w342 = ~w333 & w35575;
assign w343 = ~pi3551 & w342;
assign w344 = pi3585 & pi3631;
assign w345 = ~pi3416 & ~pi3515;
assign w346 = ~w344 & w345;
assign w347 = ~pi0784 & ~pi1449;
assign w348 = w323 & w347;
assign w349 = w346 & w348;
assign w350 = ~w333 & w35576;
assign w351 = ~pi1642 & ~pi3376;
assign w352 = ~pi3304 & w351;
assign w353 = w351 & w35577;
assign w354 = pi3641 & ~w353;
assign w355 = pi1860 & pi3641;
assign w356 = ~pi2601 & ~w355;
assign w357 = ~w354 & w356;
assign w358 = ~w350 & ~w357;
assign w359 = ~w343 & ~w358;
assign w360 = ~pi0692 & pi3216;
assign w361 = ~pi3426 & w360;
assign w362 = w359 & ~w361;
assign w363 = (w354 & ~w342) | (w354 & w35579) | (~w342 & w35579);
assign w364 = (~w363 & ~w359) | (~w363 & w35580) | (~w359 & w35580);
assign w365 = ~pi3395 & ~pi3424;
assign w366 = ~pi3427 & ~pi3429;
assign w367 = w365 & w366;
assign w368 = w367 & w35582;
assign w369 = (~pi3426 & w368) | (~pi3426 & w35583) | (w368 & w35583);
assign w370 = ~pi3551 & w341;
assign w371 = (w369 & ~w341) | (w369 & w35584) | (~w341 & w35584);
assign w372 = ~pi3436 & pi3451;
assign w373 = ~w367 & w35585;
assign w374 = pi0403 & ~pi0417;
assign w375 = pi0416 & w374;
assign w376 = pi0419 & pi0420;
assign w377 = ~pi0416 & ~pi0417;
assign w378 = ~pi0403 & ~pi0418;
assign w379 = w377 & w378;
assign w380 = ~pi0421 & w379;
assign w381 = w379 & w35586;
assign w382 = w379 & w35587;
assign w383 = (~pi0412 & w382) | (~pi0412 & w35588) | (w382 & w35588);
assign w384 = pi0411 & w383;
assign w385 = pi0414 & ~pi0415;
assign w386 = ~w382 & w35589;
assign w387 = (~w373 & w384) | (~w373 & w35590) | (w384 & w35590);
assign w388 = ~w371 & w387;
assign w389 = w367 & w35591;
assign w390 = (~pi0994 & ~w389) | (~pi0994 & w35592) | (~w389 & w35592);
assign w391 = ~pi3426 & ~w390;
assign w392 = (w391 & ~w341) | (w391 & w35593) | (~w341 & w35593);
assign w393 = pi3436 & pi3451;
assign w394 = ~w367 & w35594;
assign w395 = (~pi0411 & w382) | (~pi0411 & w35595) | (w382 & w35595);
assign w396 = pi0412 & w395;
assign w397 = ~pi0414 & pi0415;
assign w398 = ~w382 & w35596;
assign w399 = ~w396 & ~w398;
assign w400 = (~w394 & w396) | (~w394 & w35597) | (w396 & w35597);
assign w401 = ~w392 & w400;
assign w402 = ~w388 & ~w401;
assign w403 = w367 & w35598;
assign w404 = (~pi3426 & w403) | (~pi3426 & w35599) | (w403 & w35599);
assign w405 = ~w370 & w404;
assign w406 = ~w367 & w35600;
assign w407 = ~w382 & w35601;
assign w408 = ~w395 & ~w407;
assign w409 = w399 & ~w408;
assign w410 = w399 & w35602;
assign w411 = ~w405 & w410;
assign w412 = w367 & w35603;
assign w413 = (~pi3426 & w412) | (~pi3426 & w35604) | (w412 & w35604);
assign w414 = ~w370 & w413;
assign w415 = ~w382 & w35605;
assign w416 = ~w383 & ~w415;
assign w417 = ~w367 & w35606;
assign w418 = w408 & ~w417;
assign w419 = w416 & w418;
assign w420 = ~w414 & w419;
assign w421 = ~w411 & ~w420;
assign w422 = w402 & w421;
assign w423 = (w362 & ~w421) | (w362 & w35607) | (~w421 & w35607);
assign w424 = ~w364 & ~w423;
assign w425 = ~pi0634 & ~pi0638;
assign w426 = ~pi0639 & w425;
assign w427 = ~pi0640 & ~pi0641;
assign w428 = w426 & w427;
assign w429 = ~pi0637 & ~pi0736;
assign w430 = ~pi0636 & w429;
assign w431 = ~pi0658 & ~pi0735;
assign w432 = w430 & w431;
assign w433 = w430 & w35608;
assign w434 = w428 & w433;
assign w435 = ~pi0613 & ~pi0614;
assign w436 = w434 & w435;
assign w437 = w434 & w35609;
assign w438 = ~pi0613 & ~pi0753;
assign w439 = ~pi0614 & w438;
assign w440 = ~w430 & ~w431;
assign w441 = w439 & ~w440;
assign w442 = ~w433 & ~w441;
assign w443 = w425 & w35610;
assign w444 = (~pi0641 & w425) | (~pi0641 & w35611) | (w425 & w35611);
assign w445 = ~w443 & ~w444;
assign w446 = pi0658 & pi0735;
assign w447 = ~pi0612 & ~w446;
assign w448 = ~w432 & ~w447;
assign w449 = pi0636 & ~w429;
assign w450 = pi0753 & ~w435;
assign w451 = pi0637 & pi0736;
assign w452 = pi0613 & pi0614;
assign w453 = ~w451 & ~w452;
assign w454 = ~w450 & w453;
assign w455 = ~w449 & w454;
assign w456 = ~w448 & w455;
assign w457 = ~w445 & w456;
assign w458 = w433 & w439;
assign w459 = pi0634 & pi0638;
assign w460 = w433 & w35612;
assign w461 = w425 & w35611;
assign w462 = ~w460 & ~w461;
assign w463 = w457 & w35613;
assign w464 = w433 & w35614;
assign w465 = pi0640 & ~w464;
assign w466 = w463 & ~w465;
assign w467 = (pi0753 & ~w463) | (pi0753 & w35615) | (~w463 & w35615);
assign w468 = (w463 & w35616) | (w463 & w35617) | (w35616 & w35617);
assign w469 = pi0666 & ~w468;
assign w470 = (w463 & w35619) | (w463 & w35620) | (w35619 & w35620);
assign w471 = pi0534 & pi0643;
assign w472 = ~w470 & w471;
assign w473 = (~pi0534 & w470) | (~pi0534 & w35621) | (w470 & w35621);
assign w474 = w434 & w466;
assign w475 = w466 & w35622;
assign w476 = (~w439 & ~w463) | (~w439 & w35623) | (~w463 & w35623);
assign w477 = (pi0756 & w475) | (pi0756 & w35624) | (w475 & w35624);
assign w478 = ~pi0535 & ~w477;
assign w479 = w457 & w35625;
assign w480 = w430 & w479;
assign w481 = w479 & w35626;
assign w482 = w479 & w35627;
assign w483 = w438 & w35628;
assign w484 = ~pi0612 & w483;
assign w485 = (~w484 & ~w463) | (~w484 & w35629) | (~w463 & w35629);
assign w486 = ~w482 & ~w485;
assign w487 = (~pi0533 & w486) | (~pi0533 & w35630) | (w486 & w35630);
assign w488 = (~w483 & ~w463) | (~w483 & w35631) | (~w463 & w35631);
assign w489 = (pi0757 & w474) | (pi0757 & w35632) | (w474 & w35632);
assign w490 = ~pi0536 & ~w489;
assign w491 = ~w487 & ~w490;
assign w492 = pi0535 & w477;
assign w493 = ~w478 & ~w492;
assign w494 = pi0536 & pi0757;
assign w495 = (w494 & w474) | (w494 & w35633) | (w474 & w35633);
assign w496 = w493 & ~w495;
assign w497 = ~w491 & w496;
assign w498 = (~w478 & ~w496) | (~w478 & w35634) | (~w496 & w35634);
assign w499 = ~w473 & w498;
assign w500 = ~w469 & w40089;
assign w501 = pi0569 & pi0667;
assign w502 = (w501 & ~w463) | (w501 & w599) | (~w463 & w599);
assign w503 = ~pi0510 & ~w502;
assign w504 = pi0510 & w502;
assign w505 = (pi0665 & ~w463) | (pi0665 & w35637) | (~w463 & w35637);
assign w506 = ~w504 & ~w505;
assign w507 = ~w503 & ~w506;
assign w508 = ~pi0509 & ~w507;
assign w509 = (pi0509 & w502) | (pi0509 & w35638) | (w502 & w35638);
assign w510 = ~w506 & w509;
assign w511 = ~pi0639 & w427;
assign w512 = w463 & w35639;
assign w513 = (pi0664 & w463) | (pi0664 & w35640) | (w463 & w35640);
assign w514 = ~w512 & w513;
assign w515 = ~w510 & ~w514;
assign w516 = ~w508 & ~w515;
assign w517 = ~pi0508 & ~w516;
assign w518 = w433 & w35641;
assign w519 = ~w479 & w518;
assign w520 = (pi0634 & ~w463) | (pi0634 & w35642) | (~w463 & w35642);
assign w521 = w519 & ~w520;
assign w522 = pi0663 & ~w521;
assign w523 = (w522 & w516) | (w522 & w35643) | (w516 & w35643);
assign w524 = w463 & w35644;
assign w525 = ~w519 & ~w524;
assign w526 = pi0662 & w525;
assign w527 = w525 & w35645;
assign w528 = pi0508 & w516;
assign w529 = (~w527 & ~w516) | (~w527 & w35646) | (~w516 & w35646);
assign w530 = ~w523 & w529;
assign w531 = w483 & w35647;
assign w532 = w483 & w35648;
assign w533 = (~w532 & ~w463) | (~w532 & w35649) | (~w463 & w35649);
assign w534 = ~pi0736 & w479;
assign w535 = w479 & w429;
assign w536 = ~w533 & ~w535;
assign w537 = (pi0637 & ~w463) | (pi0637 & w35650) | (~w463 & w35650);
assign w538 = (pi0642 & ~w536) | (pi0642 & w681) | (~w536 & w681);
assign w539 = ~pi0505 & ~w538;
assign w540 = (~w458 & ~w463) | (~w458 & w35651) | (~w463 & w35651);
assign w541 = ~w534 & ~w540;
assign w542 = ~w541 & w35652;
assign w543 = (~pi0506 & w541) | (~pi0506 & w35653) | (w541 & w35653);
assign w544 = ~w542 & ~w543;
assign w545 = (~pi0507 & ~w525) | (~pi0507 & w35654) | (~w525 & w35654);
assign w546 = w544 & ~w545;
assign w547 = ~w539 & w546;
assign w548 = ~w541 & w35655;
assign w549 = ~w538 & ~w548;
assign w550 = (w549 & w530) | (w549 & w35656) | (w530 & w35656);
assign w551 = ~pi0505 & ~w542;
assign w552 = ~w480 & ~w533;
assign w553 = (~pi0567 & w552) | (~pi0567 & w35657) | (w552 & w35657);
assign w554 = (~w531 & ~w463) | (~w531 & w35658) | (~w463 & w35658);
assign w555 = ~w481 & ~w554;
assign w556 = (~pi0566 & w555) | (~pi0566 & w6550) | (w555 & w6550);
assign w557 = ~w553 & ~w556;
assign w558 = ~w551 & w557;
assign w559 = w546 & w557;
assign w560 = (~w558 & w530) | (~w558 & w35659) | (w530 & w35659);
assign w561 = ~w550 & ~w560;
assign w562 = (~w473 & w477) | (~w473 & w35660) | (w477 & w35660);
assign w563 = (w562 & ~w493) | (w562 & w35661) | (~w493 & w35661);
assign w564 = ~w486 & w35662;
assign w565 = ~w487 & ~w564;
assign w566 = ~w555 & w35663;
assign w567 = ~w552 & w35664;
assign w568 = ~w566 & ~w567;
assign w569 = ~w556 & ~w568;
assign w570 = w565 & ~w569;
assign w571 = ~w569 & w35665;
assign w572 = ~w563 & w571;
assign w573 = ~w469 & w572;
assign w574 = (~w500 & w561) | (~w500 & w35666) | (w561 & w35666);
assign w575 = pi0568 & w574;
assign w576 = ~pi0568 & pi0634;
assign w577 = pi0568 & ~pi0634;
assign w578 = ~w576 & ~w577;
assign w579 = ~pi0508 & ~w578;
assign w580 = pi0508 & w578;
assign w581 = ~w579 & w40090;
assign w582 = ~w527 & ~w545;
assign w583 = ~pi0568 & pi0638;
assign w584 = pi0568 & ~pi0638;
assign w585 = ~w583 & ~w584;
assign w586 = ~w582 & w585;
assign w587 = w582 & ~w585;
assign w588 = ~w586 & ~w587;
assign w589 = w581 & ~w588;
assign w590 = ~w581 & w588;
assign w591 = ~w589 & ~w590;
assign w592 = ~pi0568 & pi0640;
assign w593 = pi0568 & ~pi0640;
assign w594 = ~w592 & ~w593;
assign w595 = ~pi0510 & ~w594;
assign w596 = pi0510 & w594;
assign w597 = ~w595 & ~w596;
assign w598 = ~w505 & w597;
assign w599 = ~pi0641 & w501;
assign w600 = w501 & w35668;
assign w601 = pi0665 & ~w597;
assign w602 = (w601 & ~w463) | (w601 & w35669) | (~w463 & w35669);
assign w603 = ~w600 & ~w602;
assign w604 = ~w598 & w603;
assign w605 = pi0568 & ~pi0641;
assign w606 = ~pi0569 & w605;
assign w607 = ~pi0569 & pi0641;
assign w608 = ~w605 & ~w607;
assign w609 = ~w501 & ~w608;
assign w610 = (w609 & w463) | (w609 & w35671) | (w463 & w35671);
assign w611 = ~w604 & ~w610;
assign w612 = (~w595 & w505) | (~w595 & w35672) | (w505 & w35672);
assign w613 = ~w611 & ~w612;
assign w614 = ~w579 & ~w580;
assign w615 = (w614 & w521) | (w614 & w35673) | (w521 & w35673);
assign w616 = ~w521 & w35674;
assign w617 = ~w615 & ~w616;
assign w618 = ~w613 & ~w617;
assign w619 = ~pi0568 & pi0639;
assign w620 = pi0568 & ~pi0639;
assign w621 = ~w619 & ~w620;
assign w622 = ~pi0509 & ~w621;
assign w623 = pi0509 & w621;
assign w624 = (~w622 & w514) | (~w622 & w35675) | (w514 & w35675);
assign w625 = ~w618 & ~w624;
assign w626 = w514 & w623;
assign w627 = (w626 & w611) | (w626 & w35676) | (w611 & w35676);
assign w628 = ~w604 & w35677;
assign w629 = ~w514 & w622;
assign w630 = ~w617 & ~w629;
assign w631 = ~w628 & ~w630;
assign w632 = ~w627 & w631;
assign w633 = ~w625 & ~w632;
assign w634 = w591 & w633;
assign w635 = ~pi0568 & pi0736;
assign w636 = pi0568 & ~pi0736;
assign w637 = ~w635 & ~w636;
assign w638 = ~w544 & w637;
assign w639 = w544 & ~w637;
assign w640 = ~w638 & ~w639;
assign w641 = (w525 & w35678) | (w525 & w35679) | (w35678 & w35679);
assign w642 = ~w527 & ~w641;
assign w643 = w640 & w642;
assign w644 = ~w640 & ~w642;
assign w645 = ~w643 & ~w644;
assign w646 = ~w589 & w645;
assign w647 = ~w634 & w646;
assign w648 = ~pi0568 & pi0658;
assign w649 = pi0568 & ~pi0658;
assign w650 = ~w648 & ~w649;
assign w651 = (~w650 & w555) | (~w650 & w35680) | (w555 & w35680);
assign w652 = ~w556 & ~w651;
assign w653 = ~pi0568 & pi0612;
assign w654 = pi0568 & ~pi0612;
assign w655 = ~w653 & ~w654;
assign w656 = w565 & w655;
assign w657 = ~w565 & ~w655;
assign w658 = ~w656 & ~w657;
assign w659 = ~w652 & ~w658;
assign w660 = ~w556 & ~w566;
assign w661 = w650 & ~w660;
assign w662 = ~w650 & w660;
assign w663 = ~w661 & ~w662;
assign w664 = ~w552 & w35681;
assign w665 = ~pi0567 & pi0568;
assign w666 = pi0567 & ~pi0568;
assign w667 = ~w665 & ~w666;
assign w668 = (w463 & w35683) | (w463 & w35684) | (w35683 & w35684);
assign w669 = w667 & ~w668;
assign w670 = ~w667 & w668;
assign w671 = ~w669 & ~w670;
assign w672 = ~w664 & w671;
assign w673 = ~w552 & w35685;
assign w674 = ~w672 & ~w673;
assign w675 = (~w553 & w672) | (~w553 & w35686) | (w672 & w35686);
assign w676 = ~w567 & ~w675;
assign w677 = w663 & w676;
assign w678 = ~w659 & ~w677;
assign w679 = w637 & ~w543;
assign w680 = ~w542 & ~w679;
assign w681 = pi0642 & w537;
assign w682 = ~w681 & w40091;
assign w683 = ~pi0505 & pi0568;
assign w684 = pi0505 & ~pi0568;
assign w685 = ~w683 & ~w684;
assign w686 = w682 & w685;
assign w687 = ~w682 & ~w685;
assign w688 = ~w686 & ~w687;
assign w689 = w680 & ~w688;
assign w690 = pi0568 & pi0642;
assign w691 = (w690 & ~w463) | (w690 & w35688) | (~w463 & w35688);
assign w692 = (~w691 & w536) | (~w691 & w35689) | (w536 & w35689);
assign w693 = ~pi0505 & w692;
assign w694 = ~pi0568 & pi0637;
assign w695 = pi0568 & ~pi0637;
assign w696 = ~w694 & ~w695;
assign w697 = (w696 & w692) | (w696 & w35690) | (w692 & w35690);
assign w698 = ~w693 & w697;
assign w699 = pi0505 & w538;
assign w700 = (~w699 & w672) | (~w699 & w35691) | (w672 & w35691);
assign w701 = ~w698 & w700;
assign w702 = ~w643 & w35692;
assign w703 = w678 & w702;
assign w704 = ~w647 & w703;
assign w705 = (~w696 & w541) | (~w696 & w35693) | (w541 & w35693);
assign w706 = ~w679 & w705;
assign w707 = ~w539 & ~w706;
assign w708 = (~w637 & w541) | (~w637 & w35694) | (w541 & w35694);
assign w709 = w696 & ~w543;
assign w710 = ~w708 & w709;
assign w711 = ~w699 & ~w710;
assign w712 = ~w707 & w711;
assign w713 = w699 & w710;
assign w714 = ~w674 & ~w713;
assign w715 = ~w712 & ~w714;
assign w716 = ~w663 & ~w676;
assign w717 = ~w715 & ~w716;
assign w718 = w678 & ~w717;
assign w719 = w652 & w658;
assign w720 = ~w490 & ~w495;
assign w721 = ~pi0568 & pi0735;
assign w722 = pi0568 & ~pi0735;
assign w723 = ~w721 & ~w722;
assign w724 = (w723 & w490) | (w723 & w35695) | (w490 & w35695);
assign w725 = ~w490 & w746;
assign w726 = ~w724 & ~w725;
assign w727 = (~w655 & w486) | (~w655 & w35696) | (w486 & w35696);
assign w728 = ~w487 & ~w727;
assign w729 = w726 & ~w728;
assign w730 = ~w726 & w728;
assign w731 = ~w729 & ~w730;
assign w732 = ~w719 & w731;
assign w733 = pi0568 & ~pi0614;
assign w734 = ~pi0568 & pi0614;
assign w735 = ~w733 & ~w734;
assign w736 = (~w735 & ~w477) | (~w735 & w35697) | (~w477 & w35697);
assign w737 = ~w478 & ~w736;
assign w738 = ~pi0568 & pi0613;
assign w739 = pi0568 & ~pi0613;
assign w740 = ~w738 & ~w739;
assign w741 = ~w472 & ~w473;
assign w742 = w740 & w741;
assign w743 = ~w740 & ~w741;
assign w744 = ~w742 & ~w743;
assign w745 = w737 & w744;
assign w746 = ~w495 & ~w723;
assign w747 = ~pi0535 & w735;
assign w748 = pi0535 & ~w735;
assign w749 = ~w747 & ~w748;
assign w750 = w477 & w749;
assign w751 = ~w477 & ~w749;
assign w752 = ~w750 & ~w751;
assign w753 = ~w490 & ~w752;
assign w754 = ~w752 & w35698;
assign w755 = ~w745 & ~w754;
assign w756 = w434 & w35699;
assign w757 = ~w756 & w40092;
assign w758 = ~w473 & w740;
assign w759 = w466 & w35701;
assign w760 = (~pi0568 & ~w463) | (~pi0568 & w35702) | (~w463 & w35702);
assign w761 = ~w467 & ~w760;
assign w762 = ~w759 & w761;
assign w763 = w471 & ~w762;
assign w764 = (w757 & w763) | (w757 & w35703) | (w763 & w35703);
assign w765 = (~pi0568 & ~w434) | (~pi0568 & w35704) | (~w434 & w35704);
assign w766 = ~w764 & w765;
assign w767 = w755 & w766;
assign w768 = w732 & w767;
assign w769 = ~w718 & w768;
assign w770 = ~w704 & w769;
assign w771 = ~w763 & w35705;
assign w772 = ~w495 & w752;
assign w773 = ~w753 & ~w772;
assign w774 = ~pi0614 & pi0735;
assign w775 = pi0614 & ~pi0735;
assign w776 = ~w774 & ~w775;
assign w777 = ~w490 & w35706;
assign w778 = w493 & w777;
assign w779 = ~w490 & w35707;
assign w780 = ~w493 & w779;
assign w781 = ~w778 & ~w780;
assign w782 = ~w773 & w781;
assign w783 = ~w737 & ~w744;
assign w784 = ~w729 & ~w783;
assign w785 = ~w782 & w784;
assign w786 = ~w755 & ~w783;
assign w787 = ~w785 & ~w786;
assign w788 = (~w771 & w785) | (~w771 & w35708) | (w785 & w35708);
assign w789 = w766 & ~w788;
assign w790 = ~w770 & ~w789;
assign w791 = w731 & w35709;
assign w792 = ~w718 & w791;
assign w793 = ~w704 & w792;
assign w794 = w434 & w35710;
assign w795 = w788 & w794;
assign w796 = ~w793 & w795;
assign w797 = w790 & ~w796;
assign w798 = ~w575 & w797;
assign w799 = w496 & w570;
assign w800 = ~w561 & w799;
assign w801 = pi0643 & w470;
assign w802 = ~w741 & ~w801;
assign w803 = w802 & w40093;
assign w804 = ~w471 & w499;
assign w805 = ~w800 & w804;
assign w806 = ~w803 & ~w805;
assign w807 = (w806 & ~w797) | (w806 & w35712) | (~w797 & w35712);
assign w808 = (~w754 & w782) | (~w754 & w35713) | (w782 & w35713);
assign w809 = w731 & w35714;
assign w810 = ~w718 & w809;
assign w811 = (~w808 & w704) | (~w808 & w35715) | (w704 & w35715);
assign w812 = ~w745 & ~w783;
assign w813 = ~w801 & w812;
assign w814 = w811 & w813;
assign w815 = ~w801 & ~w812;
assign w816 = ~w811 & w815;
assign w817 = ~w814 & ~w816;
assign w818 = w798 & w817;
assign w819 = ~w807 & ~w818;
assign w820 = ~w818 & w35716;
assign w821 = pi2598 & pi3641;
assign w822 = w352 & w821;
assign w823 = w352 & w35717;
assign w824 = pi1642 & ~pi3376;
assign w825 = pi3641 & w824;
assign w826 = w824 & w35718;
assign w827 = pi3304 & pi3641;
assign w828 = w351 & w827;
assign w829 = pi1727 & w828;
assign w830 = pi3376 & pi3641;
assign w831 = pi1436 & w830;
assign w832 = ~w829 & w35719;
assign w833 = ~w823 & w832;
assign w834 = w352 & w35720;
assign w835 = w824 & w35721;
assign w836 = pi1737 & w828;
assign w837 = pi1446 & w830;
assign w838 = ~w836 & w35722;
assign w839 = ~w834 & w838;
assign w840 = w833 & ~w839;
assign w841 = ~w369 & ~w373;
assign w842 = ~pi3551 & ~w373;
assign w843 = ~w333 & w35723;
assign w844 = ~w841 & ~w843;
assign w845 = w840 & ~w844;
assign w846 = ~w404 & ~w406;
assign w847 = ~pi3551 & ~w406;
assign w848 = ~w333 & w35724;
assign w849 = ~w846 & ~w848;
assign w850 = w833 & w839;
assign w851 = ~w849 & w850;
assign w852 = ~w845 & ~w851;
assign w853 = (~w394 & w390) | (~w394 & w35725) | (w390 & w35725);
assign w854 = ~pi3551 & ~w394;
assign w855 = ~w333 & w35726;
assign w856 = ~w853 & ~w855;
assign w857 = ~w833 & w839;
assign w858 = ~w856 & w857;
assign w859 = w352 & w35727;
assign w860 = w824 & w35728;
assign w861 = pi1736 & w828;
assign w862 = pi1445 & w830;
assign w863 = ~w861 & w35729;
assign w864 = ~w859 & w863;
assign w865 = ~w833 & ~w839;
assign w866 = (~w864 & ~w865) | (~w864 & w35730) | (~w865 & w35730);
assign w867 = w413 & ~w864;
assign w868 = ~w370 & w867;
assign w869 = ~w866 & ~w868;
assign w870 = ~w858 & ~w869;
assign w871 = (w363 & ~w870) | (w363 & w35731) | (~w870 & w35731);
assign w872 = ~w362 & w871;
assign w873 = (~w364 & ~w871) | (~w364 & w35732) | (~w871 & w35732);
assign w874 = ~pi2382 & w367;
assign w875 = ~w423 & w874;
assign w876 = w873 & ~w875;
assign w877 = ~w414 & w35733;
assign w878 = ~w405 & w35734;
assign w879 = ~w877 & ~w878;
assign w880 = ~w371 & w35735;
assign w881 = ~w392 & w35736;
assign w882 = ~w880 & ~w881;
assign w883 = w879 & w882;
assign w884 = ~w424 & w883;
assign w885 = w876 & ~w884;
assign w886 = w342 & w35737;
assign w887 = ~w344 & w886;
assign w888 = ~pi2601 & w355;
assign w889 = w353 & w888;
assign w890 = ~pi0779 & ~pi3680;
assign w891 = pi0752 & ~w890;
assign w892 = pi0783 & pi3585;
assign w893 = ~pi2986 & ~pi2990;
assign w894 = w892 & w893;
assign w895 = ~pi1861 & w894;
assign w896 = w894 & w35738;
assign w897 = w894 & w35739;
assign w898 = w891 & w897;
assign w899 = w889 & w898;
assign w900 = (w899 & ~w886) | (w899 & w35740) | (~w886 & w35740);
assign w901 = ~pi1840 & pi1861;
assign w902 = w894 & w901;
assign w903 = w891 & w902;
assign w904 = ~pi3099 & w889;
assign w905 = ~w900 & ~w40129;
assign w906 = ~pi3481 & ~pi3546;
assign w907 = (w906 & w331) | (w906 & w35742) | (w331 & w35742);
assign w908 = pi0565 & ~w907;
assign w909 = ~pi3589 & w347;
assign w910 = w347 & w35743;
assign w911 = ~pi3505 & ~pi3545;
assign w912 = (~pi3362 & ~w329) | (~pi3362 & w35744) | (~w329 & w35744);
assign w913 = (pi3148 & ~w912) | (pi3148 & w35745) | (~w912 & w35745);
assign w914 = pi3452 & pi3526;
assign w915 = ~w913 & ~w914;
assign w916 = ~pi2813 & pi3362;
assign w917 = pi0565 & pi3526;
assign w918 = w909 & w917;
assign w919 = (~w916 & ~w909) | (~w916 & w35746) | (~w909 & w35746);
assign w920 = ~pi3505 & ~pi3548;
assign w921 = w329 & w35747;
assign w922 = ~pi3452 & pi3526;
assign w923 = (pi0541 & w921) | (pi0541 & w35748) | (w921 & w35748);
assign w924 = pi3215 & w921;
assign w925 = ~pi3412 & ~pi3515;
assign w926 = (~pi3548 & ~w925) | (~pi3548 & w35749) | (~w925 & w35749);
assign w927 = ~w924 & w926;
assign w928 = ~w923 & w927;
assign w929 = w927 & w35750;
assign w930 = w915 & w929;
assign w931 = ~pi3236 & pi3523;
assign w932 = ~pi3522 & ~w931;
assign w933 = w930 & w35751;
assign w934 = w359 & w361;
assign w935 = w933 & ~w934;
assign w936 = (pi2529 & w934) | (pi2529 & w35752) | (w934 & w35752);
assign w937 = (~pi1422 & ~w342) | (~pi1422 & w35753) | (~w342 & w35753);
assign w938 = (pi2601 & w353) | (pi2601 & w35754) | (w353 & w35754);
assign w939 = (w353 & w35755) | (w353 & w35756) | (w35755 & w35756);
assign w940 = pi3412 & pi3481;
assign w941 = ~pi3515 & w940;
assign w942 = w940 & w35759;
assign w943 = (w342 & w35760) | (w342 & w35761) | (w35760 & w35761);
assign w944 = ~w936 & w35762;
assign w945 = ~pi0779 & ~w905;
assign w946 = w364 & ~w945;
assign w947 = ~w944 & w946;
assign w948 = w873 & w875;
assign w949 = ~pi3364 & ~pi3385;
assign w950 = ~pi3359 & ~pi3399;
assign w951 = ~pi3387 & ~pi3388;
assign w952 = w950 & w951;
assign w953 = w949 & w952;
assign w954 = ~pi3365 & ~pi3386;
assign w955 = pi3363 & w954;
assign w956 = w953 & w955;
assign w957 = ~pi3363 & w954;
assign w958 = w949 & w957;
assign w959 = pi3359 & ~pi3399;
assign w960 = w951 & w959;
assign w961 = w958 & w960;
assign w962 = ~w956 & ~w961;
assign w963 = w952 & w957;
assign w964 = ~pi3364 & pi3385;
assign w965 = w963 & w964;
assign w966 = pi3364 & ~pi3385;
assign w967 = w963 & w966;
assign w968 = ~w965 & ~w967;
assign w969 = w962 & w968;
assign w970 = w957 & w35763;
assign w971 = ~pi3387 & pi3388;
assign w972 = w970 & w971;
assign w973 = w952 & w35764;
assign w974 = ~pi3365 & pi3386;
assign w975 = w973 & w974;
assign w976 = ~w972 & ~w975;
assign w977 = pi3387 & ~pi3388;
assign w978 = w970 & w977;
assign w979 = pi3365 & ~pi3386;
assign w980 = w973 & w979;
assign w981 = ~w978 & ~w980;
assign w982 = w976 & w981;
assign w983 = w969 & w982;
assign w984 = pi3871 & w983;
assign w985 = w973 & w35765;
assign w986 = w973 & w35766;
assign w987 = w970 & w35767;
assign w988 = ~w986 & ~w987;
assign w989 = ~w985 & w988;
assign w990 = w963 & w35768;
assign w991 = w953 & w35769;
assign w992 = w958 & w35770;
assign w993 = ~w991 & ~w992;
assign w994 = ~w990 & w993;
assign w995 = w970 & w35771;
assign w996 = w963 & w35772;
assign w997 = w952 & w958;
assign w998 = ~w996 & ~w997;
assign w999 = ~w995 & w998;
assign w1000 = w994 & w999;
assign w1001 = w989 & w1000;
assign w1002 = ~w984 & w1001;
assign w1003 = w940 & w35773;
assign w1004 = pi1044 & ~pi1256;
assign w1005 = ~pi1044 & ~pi1158;
assign w1006 = pi1014 & ~w1005;
assign w1007 = ~w1004 & w1006;
assign w1008 = ~pi1014 & pi1044;
assign w1009 = pi1284 & w1008;
assign w1010 = ~pi1014 & ~pi1044;
assign w1011 = pi1186 & w1010;
assign w1012 = ~w1009 & ~w1011;
assign w1013 = ~w1007 & w1012;
assign w1014 = ~pi1043 & pi1044;
assign w1015 = w1014 & w35774;
assign w1016 = (~w1015 & w1013) | (~w1015 & w35775) | (w1013 & w35775);
assign w1017 = ~pi0976 & ~w1016;
assign w1018 = pi1044 & pi1298;
assign w1019 = ~pi1044 & pi1200;
assign w1020 = ~w1018 & ~w1019;
assign w1021 = ~pi1043 & w1020;
assign w1022 = pi1043 & pi1044;
assign w1023 = ~pi1242 & w1022;
assign w1024 = pi0976 & pi1014;
assign w1025 = pi1043 & ~pi1044;
assign w1026 = ~pi1144 & w1025;
assign w1027 = w1024 & ~w1026;
assign w1028 = ~w1023 & w1027;
assign w1029 = ~w1021 & w1028;
assign w1030 = pi0976 & ~pi1014;
assign w1031 = pi1172 & w1025;
assign w1032 = pi1270 & w1022;
assign w1033 = pi1116 & w1014;
assign w1034 = ~w1032 & ~w1033;
assign w1035 = (w1030 & ~w1034) | (w1030 & w35776) | (~w1034 & w35776);
assign w1036 = ~pi0976 & ~pi1014;
assign w1037 = w1014 & w1036;
assign w1038 = pi1130 & w1037;
assign w1039 = ~pi1043 & ~pi1044;
assign w1040 = w1036 & w1039;
assign w1041 = pi1326 & w1040;
assign w1042 = ~w1038 & ~w1041;
assign w1043 = w1030 & w1039;
assign w1044 = pi1228 & w1043;
assign w1045 = ~pi0976 & pi1014;
assign w1046 = w1039 & w1045;
assign w1047 = pi1214 & w1046;
assign w1048 = ~w1044 & ~w1047;
assign w1049 = w1042 & w1048;
assign w1050 = ~w1035 & w1049;
assign w1051 = ~w1029 & w1050;
assign w1052 = ~w1017 & w1051;
assign w1053 = (pi1331 & ~w1051) | (pi1331 & w35777) | (~w1051 & w35777);
assign w1054 = ~pi3233 & ~pi3329;
assign w1055 = pi3512 & ~w1054;
assign w1056 = pi0381 & pi1057;
assign w1057 = pi0593 & pi1359;
assign w1058 = ~w1056 & ~w1057;
assign w1059 = ~w1055 & w1058;
assign w1060 = (pi0650 & w1053) | (pi0650 & w35778) | (w1053 & w35778);
assign w1061 = pi1339 & pi2253;
assign w1062 = pi1346 & pi2671;
assign w1063 = ~w1061 & ~w1062;
assign w1064 = pi1337 & pi2225;
assign w1065 = pi1352 & pi2446;
assign w1066 = ~w1064 & ~w1065;
assign w1067 = w1063 & w1066;
assign w1068 = pi1353 & pi1984;
assign w1069 = pi1351 & pi2269;
assign w1070 = ~w1068 & ~w1069;
assign w1071 = pi1600 & pi2211;
assign w1072 = pi1345 & pi2657;
assign w1073 = ~w1071 & ~w1072;
assign w1074 = w1070 & w1073;
assign w1075 = pi1347 & pi2685;
assign w1076 = pi1338 & pi2239;
assign w1077 = ~w1075 & ~w1076;
assign w1078 = pi1350 & pi2436;
assign w1079 = pi1348 & pi2695;
assign w1080 = ~w1078 & ~w1079;
assign w1081 = w1077 & w1080;
assign w1082 = w1074 & w1081;
assign w1083 = (pi0722 & ~w1082) | (pi0722 & w35779) | (~w1082 & w35779);
assign w1084 = pi1340 & pi2288;
assign w1085 = pi1349 & pi2735;
assign w1086 = ~w1084 & ~w1085;
assign w1087 = pi1354 & pi2533;
assign w1088 = pi1343 & pi2324;
assign w1089 = ~w1087 & ~w1088;
assign w1090 = w1086 & w1089;
assign w1091 = pi1341 & pi2122;
assign w1092 = pi1056 & pi2543;
assign w1093 = ~w1091 & ~w1092;
assign w1094 = pi1357 & pi2467;
assign w1095 = pi1055 & pi2725;
assign w1096 = ~w1094 & ~w1095;
assign w1097 = w1093 & w1096;
assign w1098 = pi1356 & pi2755;
assign w1099 = pi1342 & pi2310;
assign w1100 = ~w1098 & ~w1099;
assign w1101 = pi1355 & pi2525;
assign w1102 = pi1054 & pi2717;
assign w1103 = ~w1101 & ~w1102;
assign w1104 = w1100 & w1103;
assign w1105 = w1097 & w1104;
assign w1106 = (pi0539 & ~w1105) | (pi0539 & w35780) | (~w1105 & w35780);
assign w1107 = pi0189 & pi1336;
assign w1108 = pi1332 & pi2579;
assign w1109 = ~w1107 & ~w1108;
assign w1110 = pi1333 & pi1744;
assign w1111 = pi1335 & pi2594;
assign w1112 = ~w1110 & ~w1111;
assign w1113 = w1109 & w1112;
assign w1114 = pi0762 & ~w1113;
assign w1115 = ~w1106 & ~w1114;
assign w1116 = ~w1083 & w1115;
assign w1117 = pi0979 & pi2189;
assign w1118 = ~pi0979 & pi2949;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = pi0837 & ~w1119;
assign w1121 = pi0979 & pi2173;
assign w1122 = ~pi0979 & pi2803;
assign w1123 = ~w1121 & ~w1122;
assign w1124 = pi0836 & ~w1123;
assign w1125 = ~w1120 & ~w1124;
assign w1126 = pi0979 & pi2155;
assign w1127 = ~pi0979 & pi2927;
assign w1128 = ~w1126 & ~w1127;
assign w1129 = pi0767 & ~w1128;
assign w1130 = pi0979 & pi1965;
assign w1131 = ~pi0979 & pi2430;
assign w1132 = ~w1130 & ~w1131;
assign w1133 = pi0768 & ~w1132;
assign w1134 = pi0179 & ~pi0979;
assign w1135 = pi0164 & pi0979;
assign w1136 = ~w1134 & ~w1135;
assign w1137 = pi0838 & ~w1136;
assign w1138 = ~w1133 & ~w1137;
assign w1139 = ~w1129 & w1138;
assign w1140 = (pi0576 & ~w1139) | (pi0576 & w35781) | (~w1139 & w35781);
assign w1141 = pi0053 & ~pi0979;
assign w1142 = pi0051 & pi0979;
assign w1143 = ~w1141 & ~w1142;
assign w1144 = pi0719 & ~w1143;
assign w1145 = pi0241 & ~pi0979;
assign w1146 = pi0240 & pi0979;
assign w1147 = ~w1145 & ~w1146;
assign w1148 = pi0721 & ~w1147;
assign w1149 = pi0979 & pi2608;
assign w1150 = ~pi0979 & pi2614;
assign w1151 = ~w1149 & ~w1150;
assign w1152 = pi0763 & ~w1151;
assign w1153 = ~w1148 & ~w1152;
assign w1154 = ~w1144 & w1153;
assign w1155 = pi0979 & pi2621;
assign w1156 = ~pi0979 & pi2627;
assign w1157 = ~w1155 & ~w1156;
assign w1158 = pi0764 & ~w1157;
assign w1159 = pi0120 & ~pi0979;
assign w1160 = pi0117 & pi0979;
assign w1161 = ~w1159 & ~w1160;
assign w1162 = pi0720 & ~w1161;
assign w1163 = ~w1158 & ~w1162;
assign w1164 = pi0979 & pi3174;
assign w1165 = ~pi0979 & pi2641;
assign w1166 = ~w1164 & ~w1165;
assign w1167 = pi0765 & ~w1166;
assign w1168 = pi0979 & pi3143;
assign w1169 = ~pi0979 & pi2895;
assign w1170 = ~w1168 & ~w1169;
assign w1171 = pi0766 & ~w1170;
assign w1172 = ~w1167 & ~w1171;
assign w1173 = w1163 & w1172;
assign w1174 = w1154 & w1173;
assign w1175 = pi0524 & ~w1174;
assign w1176 = pi0203 & ~pi0979;
assign w1177 = pi0199 & pi0979;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = pi1599 & ~w1178;
assign w1180 = pi0486 & ~pi0979;
assign w1181 = pi0483 & pi0979;
assign w1182 = ~w1180 & ~w1181;
assign w1183 = pi0718 & ~w1182;
assign w1184 = ~w1179 & ~w1183;
assign w1185 = pi0184 & ~pi0979;
assign w1186 = pi0183 & pi0979;
assign w1187 = ~w1185 & ~w1186;
assign w1188 = pi0716 & ~w1187;
assign w1189 = pi0272 & ~pi0979;
assign w1190 = pi0271 & pi0979;
assign w1191 = ~w1189 & ~w1190;
assign w1192 = pi0761 & ~w1191;
assign w1193 = pi0979 & pi2136;
assign w1194 = ~pi0979 & pi2853;
assign w1195 = ~w1193 & ~w1194;
assign w1196 = pi0717 & ~w1195;
assign w1197 = ~w1192 & ~w1196;
assign w1198 = ~w1188 & w1197;
assign w1199 = (pi0538 & ~w1198) | (pi0538 & w35782) | (~w1198 & w35782);
assign w1200 = ~w1175 & w35783;
assign w1201 = w1116 & w1200;
assign w1202 = ~w1060 & w1201;
assign w1203 = ~w941 & ~w1202;
assign w1204 = ~pi1034 & ~pi1039;
assign w1205 = pi2112 & w1204;
assign w1206 = pi1036 & pi1037;
assign w1207 = pi1038 & w1206;
assign w1208 = pi1013 & pi1028;
assign w1209 = pi1029 & pi1030;
assign w1210 = pi1031 & pi1035;
assign w1211 = w1209 & w1210;
assign w1212 = w1208 & w1211;
assign w1213 = w1207 & w1212;
assign w1214 = pi1012 & ~pi1033;
assign w1215 = ~pi1032 & w1214;
assign w1216 = w1212 & w35784;
assign w1217 = w1205 & w1216;
assign w1218 = w1216 & w35785;
assign w1219 = ~pi1012 & ~pi1032;
assign w1220 = pi2112 & w1219;
assign w1221 = w1212 & w35786;
assign w1222 = pi1034 & ~pi1039;
assign w1223 = ~pi1033 & w1222;
assign w1224 = w1221 & w35787;
assign w1225 = ~pi1034 & pi1039;
assign w1226 = pi2112 & w1225;
assign w1227 = w1216 & w1226;
assign w1228 = w1216 & w35788;
assign w1229 = ~w1224 & ~w1228;
assign w1230 = ~w1218 & w1229;
assign w1231 = ~pi1012 & pi1032;
assign w1232 = ~pi1033 & w1231;
assign w1233 = pi2112 & w1222;
assign w1234 = w1232 & w1233;
assign w1235 = pi0972 & w1234;
assign w1236 = pi1034 & pi1039;
assign w1237 = pi2112 & w1236;
assign w1238 = w1232 & w1237;
assign w1239 = pi2053 & w1238;
assign w1240 = ~w1235 & ~w1239;
assign w1241 = pi1033 & w1231;
assign w1242 = w1233 & w1241;
assign w1243 = pi0303 & w1242;
assign w1244 = pi1032 & w1214;
assign w1245 = w1233 & w1244;
assign w1246 = pi0961 & w1245;
assign w1247 = ~w1243 & ~w1246;
assign w1248 = w1240 & w1247;
assign w1249 = w1215 & w1237;
assign w1250 = pi1750 & w1249;
assign w1251 = w1205 & w1244;
assign w1252 = pi0889 & w1251;
assign w1253 = ~w1250 & ~w1252;
assign w1254 = w1205 & w1232;
assign w1255 = pi0897 & w1254;
assign w1256 = pi1012 & pi1033;
assign w1257 = pi1032 & w1256;
assign w1258 = w1233 & w1257;
assign w1259 = pi1783 & w1258;
assign w1260 = ~w1255 & ~w1259;
assign w1261 = w1253 & w1260;
assign w1262 = w1248 & w1261;
assign w1263 = w1215 & w1233;
assign w1264 = pi1762 & w1263;
assign w1265 = ~pi1033 & w1219;
assign w1266 = w1237 & w1265;
assign w1267 = pi1019 & w1266;
assign w1268 = w1205 & w1257;
assign w1269 = pi1837 & w1268;
assign w1270 = ~w1267 & ~w1269;
assign w1271 = ~w1264 & w1270;
assign w1272 = w1237 & w1257;
assign w1273 = pi2111 & w1272;
assign w1274 = pi1033 & w1219;
assign w1275 = w1205 & w1274;
assign w1276 = pi2102 & w1275;
assign w1277 = ~w1273 & ~w1276;
assign w1278 = w1226 & w1232;
assign w1279 = pi1874 & w1278;
assign w1280 = w1226 & w1244;
assign w1281 = pi1909 & w1280;
assign w1282 = ~w1279 & ~w1281;
assign w1283 = w1277 & w1282;
assign w1284 = w1271 & w1283;
assign w1285 = w1262 & w1284;
assign w1286 = ~pi1033 & w1225;
assign w1287 = w1221 & w35789;
assign w1288 = w1237 & w1244;
assign w1289 = pi0796 & w1288;
assign w1290 = w1288 & w35790;
assign w1291 = w1205 & w1241;
assign w1292 = pi0890 & w1291;
assign w1293 = w1291 & w35791;
assign w1294 = w1237 & w1241;
assign w1295 = pi1880 & w1294;
assign w1296 = w1205 & w1265;
assign w1297 = pi0819 & w1296;
assign w1298 = ~w1295 & ~w1297;
assign w1299 = w1298 & w35792;
assign w1300 = ~w1287 & w1299;
assign w1301 = w1285 & w35793;
assign w1302 = pi1934 & ~w1301;
assign w1303 = ~w1203 & ~w1302;
assign w1304 = ~w1203 & w35794;
assign w1305 = pi1787 & pi2833;
assign w1306 = w958 & w35795;
assign w1307 = (w1306 & w1304) | (w1306 & w35796) | (w1304 & w35796);
assign w1308 = ~w1002 & ~w1307;
assign w1309 = ~w849 & w35797;
assign w1310 = pi1984 & w1309;
assign w1311 = w865 & w35798;
assign w1312 = ~w414 & w35799;
assign w1313 = ~w1310 & ~w1312;
assign w1314 = ~w844 & w35800;
assign w1315 = pi2269 & w1314;
assign w1316 = ~w856 & w35801;
assign w1317 = pi2446 & w1316;
assign w1318 = ~w1315 & ~w1317;
assign w1319 = w1313 & w1318;
assign w1320 = w872 & ~w1319;
assign w1321 = (~w1320 & ~w1308) | (~w1320 & w35802) | (~w1308 & w35802);
assign w1322 = ~w947 & w1321;
assign w1323 = (w1322 & w820) | (w1322 & w35803) | (w820 & w35803);
assign w1324 = (w938 & ~w886) | (w938 & w35804) | (~w886 & w35804);
assign w1325 = pi1459 & w1324;
assign w1326 = ~pi2409 & ~w889;
assign w1327 = ~pi2500 & w889;
assign w1328 = ~w1326 & ~w1327;
assign w1329 = (w886 & w35805) | (w886 & w35806) | (w35805 & w35806);
assign w1330 = ~w1325 & ~w1329;
assign w1331 = (w1330 & ~w1323) | (w1330 & w35807) | (~w1323 & w35807);
assign w1332 = pi1460 & w1324;
assign w1333 = ~pi2473 & ~w889;
assign w1334 = ~pi2501 & w889;
assign w1335 = ~w1333 & ~w1334;
assign w1336 = (w886 & w35808) | (w886 & w35809) | (w35808 & w35809);
assign w1337 = ~w1332 & ~w1336;
assign w1338 = w1337 & w1331;
assign w1339 = ~pi1450 & w1324;
assign w1340 = pi2404 & ~w889;
assign w1341 = pi2493 & w889;
assign w1342 = ~w1340 & ~w1341;
assign w1343 = (w886 & w35810) | (w886 & w35811) | (w35810 & w35811);
assign w1344 = ~w1339 & ~w1343;
assign w1345 = pi1451 & w1324;
assign w1346 = ~pi2405 & ~w889;
assign w1347 = ~pi2494 & w889;
assign w1348 = ~w1346 & ~w1347;
assign w1349 = (w886 & w35812) | (w886 & w35813) | (w35812 & w35813);
assign w1350 = ~w1345 & ~w1349;
assign w1351 = ~w1344 & w1350;
assign w1352 = (~w787 & w704) | (~w787 & w35814) | (w704 & w35814);
assign w1353 = ~w764 & ~w771;
assign w1354 = ~w1352 & w1353;
assign w1355 = w1352 & ~w1353;
assign w1356 = ~w1354 & ~w1355;
assign w1357 = w798 & ~w1356;
assign w1358 = (w498 & w35815) | (w498 & w35816) | (w35815 & w35816);
assign w1359 = (w1358 & w561) | (w1358 & w35817) | (w561 & w35817);
assign w1360 = w574 & ~w1359;
assign w1361 = pi0666 & w468;
assign w1362 = pi0568 & pi0666;
assign w1363 = (w498 & w35818) | (w498 & w35819) | (w35818 & w35819);
assign w1364 = ~w1361 & ~w1363;
assign w1365 = w572 & ~w1361;
assign w1366 = ~w561 & w1365;
assign w1367 = ~w1364 & ~w1366;
assign w1368 = (~w1367 & w797) | (~w1367 & w35820) | (w797 & w35820);
assign w1369 = ~w1357 & w1368;
assign w1370 = ~w1357 & w35821;
assign w1371 = ~w371 & w35822;
assign w1372 = ~w414 & w35823;
assign w1373 = ~w1371 & ~w1372;
assign w1374 = ~w405 & w35824;
assign w1375 = ~w392 & w35825;
assign w1376 = ~w1374 & ~w1375;
assign w1377 = w1373 & w1376;
assign w1378 = ~w424 & w1377;
assign w1379 = w876 & ~w1378;
assign w1380 = w940 & w35826;
assign w1381 = pi1043 & w1024;
assign w1382 = w1024 & w1025;
assign w1383 = pi1143 & w1382;
assign w1384 = pi1227 & w1043;
assign w1385 = w1025 & w1036;
assign w1386 = pi1185 & w1385;
assign w1387 = ~w1384 & ~w1386;
assign w1388 = w1025 & w1045;
assign w1389 = pi1157 & w1388;
assign w1390 = w1022 & w1030;
assign w1391 = pi1269 & w1390;
assign w1392 = ~w1389 & ~w1391;
assign w1393 = w1387 & w1392;
assign w1394 = ~w1383 & w1393;
assign w1395 = pi1325 & w1039;
assign w1396 = pi1283 & w1022;
assign w1397 = pi1129 & w1014;
assign w1398 = ~w1396 & ~w1397;
assign w1399 = (w1036 & ~w1398) | (w1036 & w35827) | (~w1398 & w35827);
assign w1400 = w1039 & w35828;
assign w1401 = ~w1024 & ~w1400;
assign w1402 = pi1297 & w1014;
assign w1403 = pi1241 & w1022;
assign w1404 = pi0976 & ~pi1199;
assign w1405 = w1039 & ~w1404;
assign w1406 = ~w1403 & ~w1405;
assign w1407 = ~w1402 & w1406;
assign w1408 = ~w1401 & ~w1407;
assign w1409 = w1014 & w1030;
assign w1410 = pi1115 & w1409;
assign w1411 = w1025 & w1030;
assign w1412 = pi1171 & w1411;
assign w1413 = ~w1410 & ~w1412;
assign w1414 = w1022 & w1045;
assign w1415 = pi1255 & w1414;
assign w1416 = w1014 & w1045;
assign w1417 = pi1311 & w1416;
assign w1418 = ~w1415 & ~w1417;
assign w1419 = w1413 & w1418;
assign w1420 = ~w1408 & w1419;
assign w1421 = ~w1399 & w1420;
assign w1422 = w1394 & w1421;
assign w1423 = (pi1331 & ~w1421) | (pi1331 & w35829) | (~w1421 & w35829);
assign w1424 = pi3519 & ~w1054;
assign w1425 = pi0378 & pi1057;
assign w1426 = pi0573 & pi1359;
assign w1427 = ~w1425 & ~w1426;
assign w1428 = ~w1424 & w1427;
assign w1429 = (pi0650 & w1423) | (pi0650 & w35830) | (w1423 & w35830);
assign w1430 = pi0979 & pi2172;
assign w1431 = ~pi0979 & pi2936;
assign w1432 = ~w1430 & ~w1431;
assign w1433 = pi0836 & ~w1432;
assign w1434 = pi0979 & pi2154;
assign w1435 = ~pi0979 & pi2926;
assign w1436 = ~w1434 & ~w1435;
assign w1437 = pi0767 & ~w1436;
assign w1438 = ~w1433 & ~w1437;
assign w1439 = pi0979 & pi2188;
assign w1440 = ~pi0979 & pi2948;
assign w1441 = ~w1439 & ~w1440;
assign w1442 = pi0837 & ~w1441;
assign w1443 = pi0979 & pi1964;
assign w1444 = ~pi0979 & pi2429;
assign w1445 = ~w1443 & ~w1444;
assign w1446 = pi0768 & ~w1445;
assign w1447 = pi0178 & ~pi0979;
assign w1448 = pi0163 & pi0979;
assign w1449 = ~w1447 & ~w1448;
assign w1450 = pi0838 & ~w1449;
assign w1451 = ~w1446 & ~w1450;
assign w1452 = ~w1442 & w1451;
assign w1453 = w1438 & w1452;
assign w1454 = (pi0576 & ~w1452) | (pi0576 & w35831) | (~w1452 & w35831);
assign w1455 = pi1352 & pi2445;
assign w1456 = pi1347 & pi2684;
assign w1457 = ~w1455 & ~w1456;
assign w1458 = pi1353 & pi1983;
assign w1459 = pi1351 & pi2268;
assign w1460 = ~w1458 & ~w1459;
assign w1461 = w1457 & w1460;
assign w1462 = pi1346 & pi2670;
assign w1463 = pi1348 & pi2694;
assign w1464 = ~w1462 & ~w1463;
assign w1465 = pi1350 & pi2435;
assign w1466 = pi1345 & pi2656;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = w1464 & w1467;
assign w1469 = w1461 & w1468;
assign w1470 = pi0722 & ~w1469;
assign w1471 = pi1337 & pi2224;
assign w1472 = pi1338 & pi2238;
assign w1473 = ~w1471 & ~w1472;
assign w1474 = pi1600 & pi2210;
assign w1475 = pi1339 & pi2252;
assign w1476 = ~w1474 & ~w1475;
assign w1477 = w1473 & w1476;
assign w1478 = pi0722 & ~w1477;
assign w1479 = pi1341 & pi2300;
assign w1480 = pi1342 & pi2309;
assign w1481 = ~w1479 & ~w1480;
assign w1482 = pi1343 & pi2323;
assign w1483 = pi1340 & pi2287;
assign w1484 = ~w1482 & ~w1483;
assign w1485 = w1481 & w1484;
assign w1486 = pi0539 & ~w1485;
assign w1487 = ~w1478 & ~w1486;
assign w1488 = pi1357 & pi2410;
assign w1489 = pi1355 & pi2458;
assign w1490 = ~w1488 & ~w1489;
assign w1491 = pi1056 & pi2744;
assign w1492 = pi1356 & pi2530;
assign w1493 = ~w1491 & ~w1492;
assign w1494 = w1490 & w1493;
assign w1495 = pi1054 & pi2716;
assign w1496 = pi1349 & pi2561;
assign w1497 = ~w1495 & ~w1496;
assign w1498 = pi1354 & pi2748;
assign w1499 = pi1055 & pi2774;
assign w1500 = ~w1498 & ~w1499;
assign w1501 = w1497 & w1500;
assign w1502 = w1494 & w1501;
assign w1503 = pi0539 & ~w1502;
assign w1504 = w1487 & ~w1503;
assign w1505 = ~w1470 & w1504;
assign w1506 = ~w1454 & w1505;
assign w1507 = pi0118 & ~pi0979;
assign w1508 = pi0116 & pi0979;
assign w1509 = ~w1507 & ~w1508;
assign w1510 = pi0720 & ~w1509;
assign w1511 = pi0979 & pi2607;
assign w1512 = ~pi0979 & pi2613;
assign w1513 = ~w1511 & ~w1512;
assign w1514 = pi0763 & ~w1513;
assign w1515 = pi0229 & ~pi0979;
assign w1516 = pi0228 & pi0979;
assign w1517 = ~w1515 & ~w1516;
assign w1518 = pi0721 & ~w1517;
assign w1519 = ~w1514 & ~w1518;
assign w1520 = ~w1510 & w1519;
assign w1521 = pi0979 & pi3119;
assign w1522 = ~pi0979 & pi2969;
assign w1523 = ~w1521 & ~w1522;
assign w1524 = pi0766 & ~w1523;
assign w1525 = ~w1144 & ~w1524;
assign w1526 = pi0979 & pi2620;
assign w1527 = ~pi0979 & pi2626;
assign w1528 = ~w1526 & ~w1527;
assign w1529 = pi0764 & ~w1528;
assign w1530 = pi0979 & pi3173;
assign w1531 = ~pi0979 & pi2640;
assign w1532 = ~w1530 & ~w1531;
assign w1533 = pi0765 & ~w1532;
assign w1534 = ~w1529 & ~w1533;
assign w1535 = w1525 & w1534;
assign w1536 = w1520 & w1535;
assign w1537 = pi0524 & ~w1536;
assign w1538 = pi0265 & ~pi0979;
assign w1539 = pi0261 & pi0979;
assign w1540 = ~w1538 & ~w1539;
assign w1541 = pi0716 & ~w1540;
assign w1542 = pi0979 & pi2135;
assign w1543 = ~pi0979 & pi2852;
assign w1544 = ~w1542 & ~w1543;
assign w1545 = pi0717 & ~w1544;
assign w1546 = pi0310 & ~pi0979;
assign w1547 = pi0308 & pi0979;
assign w1548 = ~w1546 & ~w1547;
assign w1549 = pi0761 & ~w1548;
assign w1550 = ~w1545 & ~w1549;
assign w1551 = ~w1541 & w1550;
assign w1552 = (pi0538 & ~w1551) | (pi0538 & w35782) | (~w1551 & w35782);
assign w1553 = ~w1537 & ~w1552;
assign w1554 = w1506 & w1553;
assign w1555 = ~w1429 & w1554;
assign w1556 = ~w941 & ~w1555;
assign w1557 = w1221 & w35832;
assign w1558 = w1221 & w35833;
assign w1559 = w1216 & w35834;
assign w1560 = ~w1558 & ~w1559;
assign w1561 = ~w1557 & w1560;
assign w1562 = pi0960 & w1245;
assign w1563 = pi1905 & w1238;
assign w1564 = pi0888 & w1251;
assign w1565 = ~w1563 & ~w1564;
assign w1566 = ~w1562 & w1565;
assign w1567 = pi0796 & ~pi1845;
assign w1568 = ~pi0796 & ~pi0962;
assign w1569 = ~w1567 & ~w1568;
assign w1570 = w1288 & w1569;
assign w1571 = pi1930 & w1272;
assign w1572 = ~w1570 & ~w1571;
assign w1573 = pi0981 & w1234;
assign w1574 = ~pi0890 & ~pi0947;
assign w1575 = pi0890 & ~pi1843;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = w1291 & w1576;
assign w1578 = ~w1573 & ~w1577;
assign w1579 = w1572 & w1578;
assign w1580 = pi2100 & w1280;
assign w1581 = pi1836 & w1268;
assign w1582 = ~w1580 & ~w1581;
assign w1583 = pi1782 & w1258;
assign w1584 = pi1879 & w1294;
assign w1585 = ~w1583 & ~w1584;
assign w1586 = w1582 & w1585;
assign w1587 = w1579 & w1586;
assign w1588 = w1566 & w1587;
assign w1589 = w1216 & w35835;
assign w1590 = pi1761 & w1263;
assign w1591 = pi0870 & w1254;
assign w1592 = ~w1590 & ~w1591;
assign w1593 = pi0909 & w1296;
assign w1594 = pi0277 & w1242;
assign w1595 = ~w1593 & ~w1594;
assign w1596 = w1592 & w1595;
assign w1597 = pi1890 & w1278;
assign w1598 = pi1749 & w1249;
assign w1599 = ~w1597 & ~w1598;
assign w1600 = pi2101 & w1275;
assign w1601 = pi0974 & w1266;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = w1599 & w1602;
assign w1604 = w1596 & w1603;
assign w1605 = ~w1589 & w1604;
assign w1606 = w1588 & w1605;
assign w1607 = pi0762 & ~w941;
assign w1608 = pi1333 & pi1743;
assign w1609 = pi1335 & pi2593;
assign w1610 = ~w1608 & ~w1609;
assign w1611 = pi0606 & pi1336;
assign w1612 = pi1332 & pi2578;
assign w1613 = ~w1611 & ~w1612;
assign w1614 = w1610 & w1613;
assign w1615 = w1607 & ~w1614;
assign w1616 = (w1606 & w35837) | (w1606 & w35838) | (w35837 & w35838);
assign w1617 = ~w1556 & w1616;
assign w1618 = ~w1556 & w35839;
assign w1619 = pi1787 & pi2817;
assign w1620 = w958 & w35840;
assign w1621 = pi3872 & w983;
assign w1622 = w973 & w35842;
assign w1623 = w973 & w35843;
assign w1624 = w970 & w35844;
assign w1625 = ~w1623 & ~w1624;
assign w1626 = ~w1622 & w1625;
assign w1627 = w958 & w35845;
assign w1628 = w963 & w35846;
assign w1629 = w953 & w35847;
assign w1630 = ~w1628 & ~w1629;
assign w1631 = ~w1627 & w1630;
assign w1632 = w970 & w35848;
assign w1633 = w963 & w35849;
assign w1634 = ~w997 & ~w1633;
assign w1635 = ~w1632 & w1634;
assign w1636 = w1631 & w1635;
assign w1637 = w1626 & w1636;
assign w1638 = ~w1621 & w1637;
assign w1639 = ~w1638 & w40095;
assign w1640 = w948 & w1639;
assign w1641 = (pi2647 & w934) | (pi2647 & w35852) | (w934 & w35852);
assign w1642 = (w353 & w35853) | (w353 & w35854) | (w35853 & w35854);
assign w1643 = w940 & w35857;
assign w1644 = (w342 & w35858) | (w342 & w35859) | (w35858 & w35859);
assign w1645 = ~w1641 & w35860;
assign w1646 = w364 & ~w1645;
assign w1647 = pi1983 & w1309;
assign w1648 = ~w414 & w35861;
assign w1649 = ~w1647 & ~w1648;
assign w1650 = pi2445 & w1316;
assign w1651 = pi2268 & w1314;
assign w1652 = ~w1650 & ~w1651;
assign w1653 = w1649 & w1652;
assign w1654 = w872 & ~w1653;
assign w1655 = ~w1646 & ~w1654;
assign w1656 = ~w1640 & w1655;
assign w1657 = (w1656 & w1370) | (w1656 & w35862) | (w1370 & w35862);
assign w1658 = pi1142 & w1382;
assign w1659 = w1014 & w1024;
assign w1660 = pi1296 & w1659;
assign w1661 = w1022 & w1024;
assign w1662 = pi1240 & w1661;
assign w1663 = ~w1660 & ~w1662;
assign w1664 = pi1184 & w1385;
assign w1665 = pi1226 & w1043;
assign w1666 = ~w1664 & ~w1665;
assign w1667 = w1663 & w1666;
assign w1668 = ~w1658 & w1667;
assign w1669 = w1039 & w35863;
assign w1670 = pi1014 & ~pi1310;
assign w1671 = ~pi1014 & ~pi1128;
assign w1672 = w1014 & ~w1671;
assign w1673 = ~w1670 & w1672;
assign w1674 = (~pi0976 & w1673) | (~pi0976 & w35864) | (w1673 & w35864);
assign w1675 = pi1170 & w1411;
assign w1676 = pi1156 & w1388;
assign w1677 = ~w1675 & ~w1676;
assign w1678 = w1022 & w1036;
assign w1679 = pi1282 & w1678;
assign w1680 = pi1114 & w1409;
assign w1681 = ~w1679 & ~w1680;
assign w1682 = w1677 & w1681;
assign w1683 = pi1254 & w1414;
assign w1684 = pi1268 & w1390;
assign w1685 = ~w1683 & ~w1684;
assign w1686 = pi1324 & w1040;
assign w1687 = w1024 & w1039;
assign w1688 = pi1198 & w1687;
assign w1689 = ~w1686 & ~w1688;
assign w1690 = w1685 & w1689;
assign w1691 = w1682 & w1690;
assign w1692 = ~w1674 & w1691;
assign w1693 = w1668 & w1692;
assign w1694 = w1692 & w35865;
assign w1695 = pi1150 & w1025;
assign w1696 = pi1248 & w1022;
assign w1697 = ~w1695 & ~w1696;
assign w1698 = pi1014 & ~w1697;
assign w1699 = w1014 & w35866;
assign w1700 = pi1043 & ~pi1178;
assign w1701 = ~pi1043 & ~pi1318;
assign w1702 = w1010 & ~w1701;
assign w1703 = ~w1700 & w1702;
assign w1704 = w1039 & w35867;
assign w1705 = ~w1703 & w35868;
assign w1706 = ~w1698 & w1705;
assign w1707 = ~pi0976 & ~w1706;
assign w1708 = pi1043 & ~pi1234;
assign w1709 = ~pi1043 & ~pi1290;
assign w1710 = pi1014 & pi1044;
assign w1711 = ~w1709 & w1710;
assign w1712 = ~w1708 & w1711;
assign w1713 = ~pi1014 & pi1043;
assign w1714 = pi1044 & pi1262;
assign w1715 = ~pi1044 & pi1164;
assign w1716 = ~w1714 & ~w1715;
assign w1717 = w1713 & ~w1716;
assign w1718 = w1039 & w35869;
assign w1719 = ~w1717 & ~w1718;
assign w1720 = (pi0976 & ~w1719) | (pi0976 & w35870) | (~w1719 & w35870);
assign w1721 = pi1136 & w1382;
assign w1722 = pi1108 & w1409;
assign w1723 = pi1220 & w1043;
assign w1724 = ~w1722 & ~w1723;
assign w1725 = pi1276 & w1678;
assign w1726 = pi1122 & w1037;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = w1724 & w1727;
assign w1729 = ~w1721 & w1728;
assign w1730 = ~w1720 & w1729;
assign w1731 = ~w1707 & w1730;
assign w1732 = w1730 & w35871;
assign w1733 = ~w1694 & ~w1732;
assign w1734 = w1039 & w35872;
assign w1735 = pi1043 & ~pi1259;
assign w1736 = ~pi1043 & ~pi1315;
assign w1737 = w1710 & ~w1736;
assign w1738 = ~w1735 & w1737;
assign w1739 = pi1044 & ~pi1287;
assign w1740 = ~pi1044 & ~pi1189;
assign w1741 = w1713 & ~w1740;
assign w1742 = ~w1739 & w1741;
assign w1743 = ~w1738 & ~w1742;
assign w1744 = (~pi0976 & ~w1743) | (~pi0976 & w35873) | (~w1743 & w35873);
assign w1745 = pi1245 & w1661;
assign w1746 = pi1161 & w1388;
assign w1747 = pi1133 & w1037;
assign w1748 = ~w1746 & ~w1747;
assign w1749 = ~w1745 & w1748;
assign w1750 = pi1329 & w1040;
assign w1751 = pi1273 & w1390;
assign w1752 = ~w1750 & ~w1751;
assign w1753 = pi1119 & w1409;
assign w1754 = ~pi1043 & w1024;
assign w1755 = pi1044 & pi1301;
assign w1756 = ~pi1044 & pi1203;
assign w1757 = ~w1755 & ~w1756;
assign w1758 = w1754 & ~w1757;
assign w1759 = ~w1753 & ~w1758;
assign w1760 = w1752 & w1759;
assign w1761 = pi1147 & w1382;
assign w1762 = ~pi1044 & w1030;
assign w1763 = ~pi1044 & pi1175;
assign w1764 = pi1043 & ~w1763;
assign w1765 = ~pi1231 & w1039;
assign w1766 = ~w1764 & ~w1765;
assign w1767 = w1762 & w1766;
assign w1768 = ~w1761 & ~w1767;
assign w1769 = w1760 & w1768;
assign w1770 = w1769 & w35874;
assign w1771 = ~pi2516 & ~w1770;
assign w1772 = (~pi2477 & ~w1730) | (~pi2477 & w35875) | (~w1730 & w35875);
assign w1773 = ~w1771 & ~w1772;
assign w1774 = w1733 & w1773;
assign w1775 = (~pi1014 & ~w1022) | (~pi1014 & w35876) | (~w1022 & w35876);
assign w1776 = pi1305 & w1014;
assign w1777 = pi1207 & w1039;
assign w1778 = ~w1776 & ~w1777;
assign w1779 = pi1014 & ~pi1249;
assign w1780 = w1022 & ~w1779;
assign w1781 = pi1151 & w1025;
assign w1782 = ~w1780 & ~w1781;
assign w1783 = w1778 & w1782;
assign w1784 = ~w1783 & w35877;
assign w1785 = pi1044 & pi1291;
assign w1786 = ~pi1044 & pi1193;
assign w1787 = ~w1785 & ~w1786;
assign w1788 = ~pi1043 & w1787;
assign w1789 = ~pi1235 & w1022;
assign w1790 = ~pi1137 & w1025;
assign w1791 = w1024 & ~w1790;
assign w1792 = ~w1789 & w1791;
assign w1793 = ~w1788 & w1792;
assign w1794 = pi1109 & w1014;
assign w1795 = pi1165 & w1025;
assign w1796 = ~w1794 & ~w1795;
assign w1797 = pi1221 & w1039;
assign w1798 = pi1263 & w1022;
assign w1799 = ~w1797 & ~w1798;
assign w1800 = w1796 & w1799;
assign w1801 = w1030 & ~w1800;
assign w1802 = pi1319 & w1040;
assign w1803 = pi1123 & w1037;
assign w1804 = pi1179 & w1385;
assign w1805 = ~w1803 & ~w1804;
assign w1806 = ~w1802 & w1805;
assign w1807 = ~w1801 & w1806;
assign w1808 = w1807 & w35878;
assign w1809 = ~pi2478 & w1808;
assign w1810 = pi2478 & ~w1808;
assign w1811 = ~w1809 & ~w1810;
assign w1812 = pi1188 & w1385;
assign w1813 = pi1118 & w1409;
assign w1814 = ~w1812 & ~w1813;
assign w1815 = pi1328 & w1040;
assign w1816 = pi1044 & pi1300;
assign w1817 = ~pi1044 & pi1202;
assign w1818 = ~w1816 & ~w1817;
assign w1819 = w1754 & ~w1818;
assign w1820 = ~w1815 & ~w1819;
assign w1821 = w1814 & w1820;
assign w1822 = pi1146 & w1382;
assign w1823 = pi1043 & pi1174;
assign w1824 = ~pi1043 & pi1230;
assign w1825 = ~w1823 & ~w1824;
assign w1826 = w1762 & ~w1825;
assign w1827 = pi1244 & w1661;
assign w1828 = ~w1826 & ~w1827;
assign w1829 = ~w1822 & w1828;
assign w1830 = w1821 & w1829;
assign w1831 = pi1314 & w1014;
assign w1832 = pi1216 & w1039;
assign w1833 = ~w1831 & ~w1832;
assign w1834 = pi1258 & w1022;
assign w1835 = pi1160 & w1025;
assign w1836 = ~w1834 & ~w1835;
assign w1837 = w1833 & w1836;
assign w1838 = w1045 & ~w1837;
assign w1839 = pi1272 & w1390;
assign w1840 = pi1286 & w1678;
assign w1841 = pi1132 & w1037;
assign w1842 = ~w1840 & ~w1841;
assign w1843 = ~w1839 & w1842;
assign w1844 = ~w1838 & w1843;
assign w1845 = w1830 & w1844;
assign w1846 = pi2517 & w1845;
assign w1847 = pi1117 & w1409;
assign w1848 = pi1257 & w1414;
assign w1849 = ~w1847 & ~w1848;
assign w1850 = pi1201 & w1687;
assign w1851 = pi1299 & w1659;
assign w1852 = ~w1850 & ~w1851;
assign w1853 = pi1044 & pi1243;
assign w1854 = ~pi1044 & pi1145;
assign w1855 = ~w1853 & ~w1854;
assign w1856 = w1381 & ~w1855;
assign w1857 = pi1043 & pi1173;
assign w1858 = ~pi1043 & pi1229;
assign w1859 = ~w1857 & ~w1858;
assign w1860 = w1762 & ~w1859;
assign w1861 = ~w1856 & ~w1860;
assign w1862 = w1852 & w1861;
assign w1863 = w1849 & w1862;
assign w1864 = pi1285 & w1678;
assign w1865 = pi1271 & w1390;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = pi1131 & w1037;
assign w1868 = pi1215 & w1046;
assign w1869 = ~w1867 & ~w1868;
assign w1870 = w1866 & w1869;
assign w1871 = pi1327 & w1040;
assign w1872 = pi1187 & w1385;
assign w1873 = ~w1871 & ~w1872;
assign w1874 = pi1313 & w1416;
assign w1875 = pi1159 & w1388;
assign w1876 = ~w1874 & ~w1875;
assign w1877 = w1873 & w1876;
assign w1878 = w1870 & w1877;
assign w1879 = w1863 & w1878;
assign w1880 = ~pi2518 & w1879;
assign w1881 = pi2518 & ~w1879;
assign w1882 = ~w1880 & ~w1881;
assign w1883 = ~w1846 & ~w1882;
assign w1884 = ~w1811 & w1883;
assign w1885 = w1774 & w1884;
assign w1886 = (~pi2483 & ~w1692) | (~pi2483 & w35879) | (~w1692 & w35879);
assign w1887 = pi1209 & w1046;
assign w1888 = pi1251 & w1414;
assign w1889 = ~w1887 & ~w1888;
assign w1890 = pi1237 & w1661;
assign w1891 = pi1279 & w1678;
assign w1892 = ~w1890 & ~w1891;
assign w1893 = pi1125 & w1037;
assign w1894 = pi1181 & w1385;
assign w1895 = ~w1893 & ~w1894;
assign w1896 = w1892 & w1895;
assign w1897 = w1889 & w1896;
assign w1898 = pi1153 & w1388;
assign w1899 = pi0976 & ~pi1139;
assign w1900 = (~w1899 & w1898) | (~w1899 & w35880) | (w1898 & w35880);
assign w1901 = pi1111 & w1014;
assign w1902 = pi1167 & w1025;
assign w1903 = ~w1901 & ~w1902;
assign w1904 = pi1265 & w1022;
assign w1905 = pi1223 & w1039;
assign w1906 = ~w1904 & ~w1905;
assign w1907 = w1903 & w1906;
assign w1908 = w1030 & ~w1907;
assign w1909 = pi1307 & w1416;
assign w1910 = pi1195 & w1687;
assign w1911 = ~w1909 & ~w1910;
assign w1912 = pi1293 & w1659;
assign w1913 = pi1321 & w1040;
assign w1914 = ~w1912 & ~w1913;
assign w1915 = w1911 & w1914;
assign w1916 = ~w1908 & w1915;
assign w1917 = ~w1900 & w1916;
assign w1918 = w1897 & w1917;
assign w1919 = w1917 & w35881;
assign w1920 = ~w1886 & ~w1919;
assign w1921 = pi2516 & w1770;
assign w1922 = (~pi2480 & ~w1917) | (~pi2480 & w35882) | (~w1917 & w35882);
assign w1923 = ~w1921 & ~w1922;
assign w1924 = w1920 & w1923;
assign w1925 = pi1127 & w1008;
assign w1926 = pi1323 & w1010;
assign w1927 = ~w1925 & ~w1926;
assign w1928 = ~pi1043 & ~w1927;
assign w1929 = pi1253 & w1710;
assign w1930 = pi1183 & w1010;
assign w1931 = ~w1929 & ~w1930;
assign w1932 = pi1043 & ~w1931;
assign w1933 = w1014 & w35883;
assign w1934 = w1039 & w35884;
assign w1935 = ~w1933 & ~w1934;
assign w1936 = ~w1932 & w1935;
assign w1937 = (~pi0976 & ~w1936) | (~pi0976 & w35885) | (~w1936 & w35885);
assign w1938 = pi1281 & w1678;
assign w1939 = pi1197 & w1687;
assign w1940 = pi1155 & w1388;
assign w1941 = ~w1939 & ~w1940;
assign w1942 = ~w1938 & w1941;
assign w1943 = pi1239 & w1661;
assign w1944 = pi1295 & w1659;
assign w1945 = ~w1943 & ~w1944;
assign w1946 = pi1225 & w1043;
assign w1947 = pi1267 & w1390;
assign w1948 = ~w1946 & ~w1947;
assign w1949 = w1945 & w1948;
assign w1950 = pi1141 & w1382;
assign w1951 = pi1169 & w1411;
assign w1952 = pi1113 & w1409;
assign w1953 = ~w1951 & ~w1952;
assign w1954 = ~w1950 & w1953;
assign w1955 = w1949 & w1954;
assign w1956 = w1942 & w1955;
assign w1957 = ~w1937 & w1956;
assign w1958 = (~pi2482 & ~w1956) | (~pi2482 & w35886) | (~w1956 & w35886);
assign w1959 = w1956 & w35887;
assign w1960 = ~w1958 & ~w1959;
assign w1961 = (~pi2485 & ~w1051) | (~pi2485 & w35888) | (~w1051 & w35888);
assign w1962 = w1051 & w35889;
assign w1963 = ~w1961 & ~w1962;
assign w1964 = w1960 & w1963;
assign w1965 = w1924 & w1964;
assign w1966 = w1885 & w1965;
assign w1967 = w1421 & w35890;
assign w1968 = ~pi2517 & ~w1845;
assign w1969 = (~pi2484 & ~w1421) | (~pi2484 & w35891) | (~w1421 & w35891);
assign w1970 = ~w1968 & ~w1969;
assign w1971 = ~w1967 & w1970;
assign w1972 = w1970 & w35892;
assign w1973 = w1885 & w35893;
assign w1974 = ~pi2016 & pi2516;
assign w1975 = pi2012 & ~pi2480;
assign w1976 = pi2375 & ~pi2484;
assign w1977 = ~w1975 & ~w1976;
assign w1978 = ~w1974 & w1977;
assign w1979 = ~pi2378 & pi2517;
assign w1980 = pi2014 & ~pi2482;
assign w1981 = ~w1979 & ~w1980;
assign w1982 = ~pi2375 & pi2484;
assign w1983 = ~pi2014 & pi2482;
assign w1984 = ~w1982 & ~w1983;
assign w1985 = w1981 & w1984;
assign w1986 = ~pi2012 & pi2480;
assign w1987 = pi2763 & ~w1986;
assign w1988 = pi2378 & ~pi2517;
assign w1989 = pi2016 & ~pi2516;
assign w1990 = ~w1988 & ~w1989;
assign w1991 = w1987 & w1990;
assign w1992 = w1985 & w1991;
assign w1993 = w1978 & w1992;
assign w1994 = pi1140 & w1382;
assign w1995 = pi1238 & w1661;
assign w1996 = pi1308 & w1416;
assign w1997 = ~w1995 & ~w1996;
assign w1998 = pi1126 & w1037;
assign w1999 = pi1280 & w1678;
assign w2000 = ~w1998 & ~w1999;
assign w2001 = w1997 & w2000;
assign w2002 = ~w1994 & w2001;
assign w2003 = pi1252 & w1022;
assign w2004 = pi1210 & w1039;
assign w2005 = pi1154 & w1025;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = (w1045 & ~w2006) | (w1045 & w35894) | (~w2006 & w35894);
assign w2008 = pi1112 & w1014;
assign w2009 = pi1266 & w1022;
assign w2010 = ~w2008 & ~w2009;
assign w2011 = pi1168 & w1025;
assign w2012 = pi1224 & w1039;
assign w2013 = ~w2011 & ~w2012;
assign w2014 = w2010 & w2013;
assign w2015 = w1030 & ~w2014;
assign w2016 = pi1294 & w1659;
assign w2017 = pi1322 & w1040;
assign w2018 = ~w2016 & ~w2017;
assign w2019 = pi1196 & w1687;
assign w2020 = pi1182 & w1385;
assign w2021 = ~w2019 & ~w2020;
assign w2022 = w2018 & w2021;
assign w2023 = ~w2015 & w2022;
assign w2024 = ~w2007 & w2023;
assign w2025 = w2002 & w2024;
assign w2026 = (~pi2481 & ~w2024) | (~pi2481 & w35895) | (~w2024 & w35895);
assign w2027 = pi1148 & w1025;
assign w2028 = pi1246 & w1022;
assign w2029 = ~w2027 & ~w2028;
assign w2030 = pi1014 & ~w2029;
assign w2031 = w1014 & w35896;
assign w2032 = pi1043 & ~pi1176;
assign w2033 = ~pi1043 & ~pi1316;
assign w2034 = w1010 & ~w2033;
assign w2035 = ~w2032 & w2034;
assign w2036 = w1039 & w35897;
assign w2037 = ~w2035 & w35898;
assign w2038 = ~w2030 & w2037;
assign w2039 = ~pi0976 & ~w2038;
assign w2040 = pi1134 & w1382;
assign w2041 = ~pi1043 & ~pi1190;
assign w2042 = (~w2041 & w2040) | (~w2041 & w35899) | (w2040 & w35899);
assign w2043 = pi1260 & w1022;
assign w2044 = pi1218 & w1039;
assign w2045 = ~w2043 & ~w2044;
assign w2046 = pi1106 & w1014;
assign w2047 = pi1162 & w1025;
assign w2048 = ~w2046 & ~w2047;
assign w2049 = w2045 & w2048;
assign w2050 = w1030 & ~w2049;
assign w2051 = pi1120 & w1037;
assign w2052 = pi1274 & w1678;
assign w2053 = ~w2051 & ~w2052;
assign w2054 = pi1288 & w1659;
assign w2055 = pi1232 & w1661;
assign w2056 = ~w2054 & ~w2055;
assign w2057 = w2053 & w2056;
assign w2058 = ~w2050 & w2057;
assign w2059 = ~w2042 & w2058;
assign w2060 = ~w2039 & w2059;
assign w2061 = w2059 & w35900;
assign w2062 = ~w2026 & ~w2061;
assign w2063 = (~pi2475 & ~w2059) | (~pi2475 & w35901) | (~w2059 & w35901);
assign w2064 = w2024 & w35902;
assign w2065 = ~w2063 & ~w2064;
assign w2066 = w2062 & w2065;
assign w2067 = ~pi2392 & pi2475;
assign w2068 = pi2373 & ~pi2476;
assign w2069 = ~w2067 & ~w2068;
assign w2070 = pi2374 & ~pi2478;
assign w2071 = pi2392 & ~pi2475;
assign w2072 = ~w2070 & ~w2071;
assign w2073 = w2069 & w2072;
assign w2074 = ~pi2013 & pi2481;
assign w2075 = pi2763 & ~w2074;
assign w2076 = ~pi2373 & pi2476;
assign w2077 = pi2010 & ~pi2477;
assign w2078 = ~w2076 & ~w2077;
assign w2079 = w2075 & w2078;
assign w2080 = w2073 & w2079;
assign w2081 = pi2011 & ~pi2479;
assign w2082 = ~pi2010 & pi2477;
assign w2083 = pi2376 & ~pi2485;
assign w2084 = ~w2082 & ~w2083;
assign w2085 = ~w2081 & w2084;
assign w2086 = ~pi2374 & pi2478;
assign w2087 = ~pi2376 & pi2485;
assign w2088 = ~w2086 & ~w2087;
assign w2089 = ~pi2015 & pi2483;
assign w2090 = ~pi2011 & pi2479;
assign w2091 = ~w2089 & ~w2090;
assign w2092 = w2088 & w2091;
assign w2093 = pi2013 & ~pi2481;
assign w2094 = ~pi2377 & pi2518;
assign w2095 = ~w2093 & ~w2094;
assign w2096 = pi2377 & ~pi2518;
assign w2097 = pi2015 & ~pi2483;
assign w2098 = ~w2096 & ~w2097;
assign w2099 = w2095 & w2098;
assign w2100 = w2092 & w2099;
assign w2101 = w2085 & w2100;
assign w2102 = w2080 & w2101;
assign w2103 = (~w2102 & ~w2066) | (~w2102 & w35903) | (~w2066 & w35903);
assign w2104 = (pi1014 & ~w1022) | (pi1014 & w35904) | (~w1022 & w35904);
assign w2105 = pi1306 & w1014;
assign w2106 = pi1152 & w1025;
assign w2107 = pi1208 & w1039;
assign w2108 = ~w2106 & ~w2107;
assign w2109 = w2108 & w35905;
assign w2110 = (~pi1014 & ~w1039) | (~pi1014 & w35906) | (~w1039 & w35906);
assign w2111 = pi1124 & w1014;
assign w2112 = pi1180 & w1025;
assign w2113 = pi1278 & w1022;
assign w2114 = ~w2112 & ~w2113;
assign w2115 = w2114 & w35907;
assign w2116 = ~w2109 & ~w2115;
assign w2117 = ~pi0976 & ~w2116;
assign w2118 = pi1264 & w1022;
assign w2119 = pi1222 & w1039;
assign w2120 = pi1166 & w1025;
assign w2121 = ~w2119 & ~w2120;
assign w2122 = w2121 & w35908;
assign w2123 = pi1194 & w1039;
assign w2124 = w1024 & ~w2123;
assign w2125 = pi1236 & w1022;
assign w2126 = pi1138 & w1025;
assign w2127 = pi1292 & w1014;
assign w2128 = ~w2126 & ~w2127;
assign w2129 = ~w2125 & w2128;
assign w2130 = w2124 & w2129;
assign w2131 = ~w2122 & ~w2130;
assign w2132 = ~w2117 & w2131;
assign w2133 = pi1110 & w1409;
assign w2134 = ~w2132 & ~w2133;
assign w2135 = ~w2132 & w35909;
assign w2136 = (~pi2479 & w2132) | (~pi2479 & w35910) | (w2132 & w35910);
assign w2137 = pi1233 & w1661;
assign w2138 = pi1261 & w1390;
assign w2139 = ~w2137 & ~w2138;
assign w2140 = pi1205 & w1046;
assign w2141 = pi1289 & w1659;
assign w2142 = ~w2140 & ~w2141;
assign w2143 = w2139 & w2142;
assign w2144 = pi1135 & w1382;
assign w2145 = pi1107 & w1409;
assign w2146 = pi1149 & w1388;
assign w2147 = ~w2145 & ~w2146;
assign w2148 = ~w2144 & w2147;
assign w2149 = w2143 & w2148;
assign w2150 = pi1275 & w1678;
assign w2151 = ~pi1043 & ~pi1121;
assign w2152 = (~w2151 & w2150) | (~w2151 & w35911) | (w2150 & w35911);
assign w2153 = pi1303 & w1416;
assign w2154 = pi1177 & w1385;
assign w2155 = pi1219 & w1043;
assign w2156 = ~w2154 & ~w2155;
assign w2157 = ~w2153 & w2156;
assign w2158 = pi1317 & w1040;
assign w2159 = pi1191 & w1687;
assign w2160 = ~w2158 & ~w2159;
assign w2161 = pi1163 & w1411;
assign w2162 = pi1247 & w1414;
assign w2163 = ~w2161 & ~w2162;
assign w2164 = w2160 & w2163;
assign w2165 = w2157 & w2164;
assign w2166 = ~w2152 & w2165;
assign w2167 = w2149 & w2166;
assign w2168 = w2166 & w35912;
assign w2169 = (~pi2476 & ~w2166) | (~pi2476 & w35913) | (~w2166 & w35913);
assign w2170 = ~w2168 & ~w2169;
assign w2171 = w2170 & w35914;
assign w2172 = ~pi2763 & ~w2171;
assign w2173 = ~w2103 & ~w2172;
assign w2174 = (w2173 & w1973) | (w2173 & w35915) | (w1973 & w35915);
assign w2175 = ~pi3190 & pi3291;
assign w2176 = ~pi2489 & w2175;
assign w2177 = (~pi2490 & ~w2175) | (~pi2490 & w35916) | (~w2175 & w35916);
assign w2178 = ~pi0134 & pi0152;
assign w2179 = pi0134 & ~pi0152;
assign w2180 = ~pi0149 & ~w2179;
assign w2181 = (pi2912 & ~w2180) | (pi2912 & w35917) | (~w2180 & w35917);
assign w2182 = ~pi0149 & ~pi2912;
assign w2183 = ~w2181 & w35918;
assign w2184 = ~pi2812 & ~pi2911;
assign w2185 = w2184 & w40096;
assign w2186 = ~w2183 & w2185;
assign w2187 = ~pi2912 & ~pi3633;
assign w2188 = ~pi2913 & w2187;
assign w2189 = pi2913 & ~w2187;
assign w2190 = ~pi0482 & pi2912;
assign w2191 = pi2812 & pi2911;
assign w2192 = ~w2190 & w2191;
assign w2193 = ~w2189 & w2192;
assign w2194 = (~pi0045 & ~w2193) | (~pi0045 & w35920) | (~w2193 & w35920);
assign w2195 = ~w2186 & w2194;
assign w2196 = (w2176 & w2186) | (w2176 & w35921) | (w2186 & w35921);
assign w2197 = w2180 & w35922;
assign w2198 = pi0149 & ~pi3267;
assign w2199 = ~pi3248 & w2198;
assign w2200 = pi3248 & ~w2198;
assign w2201 = ~w2199 & ~w2200;
assign w2202 = ~w2197 & w2201;
assign w2203 = ~pi3299 & ~w2202;
assign w2204 = ~pi3267 & pi3633;
assign w2205 = ~pi3248 & w2204;
assign w2206 = pi3248 & ~w2204;
assign w2207 = pi0482 & pi3267;
assign w2208 = pi3326 & ~w2207;
assign w2209 = ~w2206 & w2208;
assign w2210 = ~w2205 & w2209;
assign w2211 = ~w2203 & ~w2210;
assign w2212 = ~pi3299 & pi3326;
assign w2213 = (~w2212 & ~w2197) | (~w2212 & w35923) | (~w2197 & w35923);
assign w2214 = (~pi0038 & w2211) | (~pi0038 & w35924) | (w2211 & w35924);
assign w2215 = pi3268 & ~pi3426;
assign w2216 = pi2490 & ~w2215;
assign w2217 = (~pi3210 & ~w2215) | (~pi3210 & w35925) | (~w2215 & w35925);
assign w2218 = ~w2216 & w2217;
assign w2219 = w2218 & ~w2214;
assign w2220 = ~w2196 & w2219;
assign w2221 = (w2220 & w2174) | (w2220 & w35926) | (w2174 & w35926);
assign w2222 = w1971 & w2195;
assign w2223 = w2222 & w35927;
assign w2224 = (w2175 & ~w1966) | (w2175 & w35928) | (~w1966 & w35928);
assign w2225 = w2214 & ~w2215;
assign w2226 = ~w2224 & w2225;
assign w2227 = ~w2221 & ~w2226;
assign w2228 = ~pi0540 & ~w2227;
assign w2229 = ~pi3371 & ~pi3408;
assign w2230 = ~w2227 & w35929;
assign w2231 = ~pi0419 & ~pi0420;
assign w2232 = ~pi0403 & pi0418;
assign w2233 = w377 & w2232;
assign w2234 = w2231 & w2233;
assign w2235 = w2233 & w35930;
assign w2236 = ~pi0416 & pi0417;
assign w2237 = w378 & w2236;
assign w2238 = ~w2235 & ~w2237;
assign w2239 = ~w2235 & w35931;
assign w2240 = ~pi0422 & w2235;
assign w2241 = ~pi0418 & pi0419;
assign w2242 = ~pi0403 & w2236;
assign w2243 = ~w2241 & w2242;
assign w2244 = ~w2240 & ~w2243;
assign w2245 = ~w2240 & w35932;
assign w2246 = ~w2239 & ~w2245;
assign w2247 = w359 & w35933;
assign w2248 = ~pi0819 & ~pi3680;
assign w2249 = pi0909 & ~w2248;
assign w2250 = ~pi1422 & pi2515;
assign w2251 = w2249 & w2250;
assign w2252 = w2251 & w1324;
assign w2253 = w342 & w35935;
assign w2254 = ~w900 & ~w2253;
assign w2255 = ~w2252 & w2254;
assign w2256 = (w2255 & w2227) | (w2255 & w35936) | (w2227 & w35936);
assign w2257 = ~pi1422 & w2249;
assign w2258 = w2257 & w40097;
assign w2259 = ~w40129 & ~w2258;
assign w2260 = w341 & w35941;
assign w2261 = ~w358 & ~w370;
assign w2262 = (~w2260 & ~w2261) | (~w2260 & w35942) | (~w2261 & w35942);
assign w2263 = w2259 & w2262;
assign w2264 = (w2227 & w35943) | (w2227 & w35944) | (w35943 & w35944);
assign w2265 = w1351 & w40098;
assign w2266 = w1338 & w2265;
assign w2267 = ~w1344 & ~w1350;
assign w2268 = w2267 & w40098;
assign w2269 = w1338 & w2268;
assign w2270 = w1344 & w1350;
assign w2271 = w2270 & w40098;
assign w2272 = w1338 & w2271;
assign w2273 = w1344 & ~w1350;
assign w2274 = w2273 & w40098;
assign w2275 = w1338 & w2274;
assign w2276 = ~w1337 & w1331;
assign w2277 = w2265 & w2276;
assign w2278 = w2268 & w2276;
assign w2279 = w2271 & w2276;
assign w2280 = w2274 & w2276;
assign w2281 = (w342 & w35946) | (w342 & w35947) | (w35946 & w35947);
assign w2282 = ~w2262 & ~w2281;
assign w2283 = w2259 & ~w2282;
assign w2284 = ~w2283 & ~w1657;
assign w2285 = w1331 & w2284;
assign w2286 = ~pi3436 & ~pi3451;
assign w2287 = ~w367 & w35948;
assign w2288 = ~pi3392 & pi3398;
assign w2289 = w367 & w35949;
assign w2290 = (~pi3426 & w2289) | (~pi3426 & w35950) | (w2289 & w35950);
assign w2291 = ~w2287 & ~w2290;
assign w2292 = ~pi3551 & ~w2287;
assign w2293 = ~w333 & w35951;
assign w2294 = ~w2291 & ~w2293;
assign w2295 = w840 & w864;
assign w2296 = w2294 & w2295;
assign w2297 = w850 & w864;
assign w2298 = ~w367 & w35952;
assign w2299 = w354 & ~w2298;
assign w2300 = w850 & w35953;
assign w2301 = w367 & w35954;
assign w2302 = w367 & w35955;
assign w2303 = (~pi3426 & w2302) | (~pi3426 & w35956) | (w2302 & w35956);
assign w2304 = w2297 & w2303;
assign w2305 = (~w2300 & ~w2304) | (~w2300 & w35957) | (~w2304 & w35957);
assign w2306 = ~w2296 & w2305;
assign w2307 = pi3392 & pi3398;
assign w2308 = w367 & w35958;
assign w2309 = (~pi3426 & w2308) | (~pi3426 & w35959) | (w2308 & w35959);
assign w2310 = pi3436 & ~pi3451;
assign w2311 = ~w367 & w35960;
assign w2312 = ~w2309 & ~w2311;
assign w2313 = ~pi3551 & ~w2311;
assign w2314 = ~w333 & w35961;
assign w2315 = ~w2312 & ~w2314;
assign w2316 = w864 & w865;
assign w2317 = w2315 & w2316;
assign w2318 = ~w367 & w35962;
assign w2319 = (~pi0998 & ~w2301) | (~pi0998 & w35963) | (~w2301 & w35963);
assign w2320 = (~w2318 & w2319) | (~w2318 & w35964) | (w2319 & w35964);
assign w2321 = ~pi3551 & ~w2318;
assign w2322 = ~w333 & w35965;
assign w2323 = ~w2320 & ~w2322;
assign w2324 = w857 & w864;
assign w2325 = w2323 & w2324;
assign w2326 = ~w2317 & ~w2325;
assign w2327 = w2306 & w2326;
assign w2328 = ~w2290 & w35966;
assign w2329 = ~w2287 & w35967;
assign w2330 = ~w333 & w35968;
assign w2331 = ~w2328 & ~w2330;
assign w2332 = ~pi0414 & ~pi0415;
assign w2333 = ~w2298 & w2332;
assign w2334 = ~w2303 & w2333;
assign w2335 = ~w2298 & w35969;
assign w2336 = ~w333 & w35970;
assign w2337 = ~w2334 & ~w2336;
assign w2338 = w2331 & w2337;
assign w2339 = w397 & w2320;
assign w2340 = ~w2318 & w35971;
assign w2341 = ~w333 & w35972;
assign w2342 = ~w2339 & ~w2341;
assign w2343 = pi0414 & pi0415;
assign w2344 = ~w2309 & w35973;
assign w2345 = ~w2311 & w35974;
assign w2346 = ~w333 & w35975;
assign w2347 = ~w2344 & ~w2346;
assign w2348 = w2342 & w2347;
assign w2349 = w2338 & w2348;
assign w2350 = ~w354 & ~w2349;
assign w2351 = ~w2327 & ~w2350;
assign w2352 = pi3055 & ~pi3641;
assign w2353 = ~pi0403 & pi0416;
assign w2354 = ~pi0417 & w2353;
assign w2355 = ~w2352 & w2354;
assign w2356 = pi0416 & pi0417;
assign w2357 = (~w2356 & ~w2354) | (~w2356 & w35976) | (~w2354 & w35976);
assign w2358 = (~w375 & w2357) | (~w375 & w35977) | (w2357 & w35977);
assign w2359 = ~pi0692 & pi2789;
assign w2360 = (w2359 & ~w1212) | (w2359 & w35978) | (~w1212 & w35978);
assign w2361 = ~pi3426 & w2360;
assign w2362 = ~w2358 & ~w2361;
assign w2363 = w359 & w2362;
assign w2364 = (~w874 & ~w359) | (~w874 & w35979) | (~w359 & w35979);
assign w2365 = w359 & ~w2361;
assign w2366 = ~pi0830 & ~w2358;
assign w2367 = w359 & w35980;
assign w2368 = ~w2364 & ~w2367;
assign w2369 = ~w871 & w2368;
assign w2370 = ~w2351 & ~w2369;
assign w2371 = w421 & w35981;
assign w2372 = (w2358 & ~w870) | (w2358 & w35982) | (~w870 & w35982);
assign w2373 = ~w2371 & w2372;
assign w2374 = w2233 & w35983;
assign w2375 = pi0405 & w2374;
assign w2376 = pi0418 & ~w2357;
assign w2377 = ~w2375 & ~w2376;
assign w2378 = w874 & ~w2377;
assign w2379 = (w2358 & w2377) | (w2358 & w35984) | (w2377 & w35984);
assign w2380 = w359 & w35985;
assign w2381 = ~w2373 & w2380;
assign w2382 = ~pi2488 & w367;
assign w2383 = pi0830 & ~w2358;
assign w2384 = ~w2358 & w35986;
assign w2385 = ~w2327 & w35987;
assign w2386 = (~w363 & ~w2381) | (~w363 & w35988) | (~w2381 & w35988);
assign w2387 = ~w2370 & ~w2386;
assign w2388 = ~w871 & ~w2351;
assign w2389 = (~w354 & ~w359) | (~w354 & w35989) | (~w359 & w35989);
assign w2390 = w421 & w35990;
assign w2391 = w870 & w35991;
assign w2392 = ~w2390 & ~w2391;
assign w2393 = w874 & ~w2392;
assign w2394 = w2388 & ~w2393;
assign w2395 = ~w2358 & w35992;
assign w2396 = (~w363 & w2373) | (~w363 & w35994) | (w2373 & w35994);
assign w2397 = ~w2394 & ~w2396;
assign w2398 = ~w2387 & ~w2397;
assign w2399 = ~w680 & w688;
assign w2400 = ~w689 & ~w2399;
assign w2401 = (w2400 & w647) | (w2400 & w35995) | (w647 & w35995);
assign w2402 = ~w647 & w35996;
assign w2403 = w536 & w35997;
assign w2404 = ~w2402 & ~w2403;
assign w2405 = ~w2401 & w2404;
assign w2406 = w797 & w35998;
assign w2407 = ~w530 & w546;
assign w2408 = (w551 & w530) | (w551 & w35999) | (w530 & w35999);
assign w2409 = pi0505 & w40099;
assign w2410 = ~w2408 & ~w2409;
assign w2411 = pi0642 & ~w2410;
assign w2412 = ~w538 & w2410;
assign w2413 = ~w2411 & ~w2412;
assign w2414 = (~w2413 & ~w797) | (~w2413 & w36001) | (~w797 & w36001);
assign w2415 = ~w2406 & ~w2414;
assign w2416 = w2398 & ~w2415;
assign w2417 = w359 & w36002;
assign w2418 = ~w2373 & w2417;
assign w2419 = (~w363 & ~w359) | (~w363 & w36004) | (~w359 & w36004);
assign w2420 = ~w2418 & w2419;
assign w2421 = (w342 & w36005) | (w342 & w36006) | (w36005 & w36006);
assign w2422 = ~w2382 & ~w2421;
assign w2423 = ~w2327 & w36007;
assign w2424 = (~w2423 & ~w2388) | (~w2423 & w36008) | (~w2388 & w36008);
assign w2425 = ~w2420 & w2424;
assign w2426 = ~pi0670 & ~pi0671;
assign w2427 = ~pi0644 & ~pi0669;
assign w2428 = w2426 & w2427;
assign w2429 = ~pi0656 & ~pi0673;
assign w2430 = ~pi0674 & w2429;
assign w2431 = ~pi0657 & ~pi0672;
assign w2432 = w2430 & w2431;
assign w2433 = pi0674 & ~w2429;
assign w2434 = w2428 & ~w2433;
assign w2435 = ~w2432 & ~w2434;
assign w2436 = ~w2430 & ~w2431;
assign w2437 = pi0644 & pi0669;
assign w2438 = pi0645 & pi0646;
assign w2439 = pi0656 & pi0673;
assign w2440 = ~w2438 & ~w2439;
assign w2441 = ~w2437 & w2440;
assign w2442 = ~w2426 & ~w2427;
assign w2443 = pi0670 & pi0671;
assign w2444 = pi0657 & pi0672;
assign w2445 = ~w2443 & ~w2444;
assign w2446 = ~w2442 & w2445;
assign w2447 = w2441 & w2446;
assign w2448 = ~w2436 & w2447;
assign w2449 = ~w2435 & w2448;
assign w2450 = ~pi0645 & ~pi0646;
assign w2451 = ~pi0675 & w2450;
assign w2452 = w2450 & w36009;
assign w2453 = ~pi0668 & w2452;
assign w2454 = (w2453 & ~w2448) | (w2453 & w36010) | (~w2448 & w36010);
assign w2455 = w2428 & w2454;
assign w2456 = w2428 & w2432;
assign w2457 = ~w2453 & ~w2456;
assign w2458 = (pi0676 & ~w2450) | (pi0676 & w36011) | (~w2450 & w36011);
assign w2459 = (~pi0668 & w2450) | (~pi0668 & w36012) | (w2450 & w36012);
assign w2460 = ~w2452 & ~w2459;
assign w2461 = ~w2458 & ~w2460;
assign w2462 = w2449 & w36013;
assign w2463 = w2430 & w36014;
assign w2464 = w2462 & ~w2463;
assign w2465 = ~w2464 & w36015;
assign w2466 = ~pi0514 & ~w2465;
assign w2467 = pi0514 & w2465;
assign w2468 = ~w2456 & w2462;
assign w2469 = w2462 & w36016;
assign w2470 = ~pi0672 & w2428;
assign w2471 = w2454 & w2470;
assign w2472 = pi0515 & pi0704;
assign w2473 = (w2472 & ~w2454) | (w2472 & w36017) | (~w2454 & w36017);
assign w2474 = ~w2469 & w2473;
assign w2475 = ~w2467 & ~w2474;
assign w2476 = ~w2475 & w36018;
assign w2477 = ~pi0588 & ~pi0705;
assign w2478 = ~pi0657 & w2454;
assign w2479 = w2428 & w36019;
assign w2480 = (w2479 & w2468) | (w2479 & w36020) | (w2468 & w36020);
assign w2481 = ~w2477 & ~w2480;
assign w2482 = ~w2430 & w2462;
assign w2483 = ~pi0657 & ~pi0674;
assign w2484 = w2454 & w36021;
assign w2485 = ~w2482 & w36022;
assign w2486 = ~pi0516 & ~w2485;
assign w2487 = pi0521 & pi0707;
assign w2488 = ~pi0517 & ~w2487;
assign w2489 = ~w2488 & w40100;
assign w2490 = pi0517 & w2487;
assign w2491 = (w2490 & ~w2462) | (w2490 & w36024) | (~w2462 & w36024);
assign w2492 = ~w2489 & ~w2491;
assign w2493 = ~w2486 & ~w2492;
assign w2494 = pi0516 & w2485;
assign w2495 = (w2470 & w2468) | (w2470 & w36025) | (w2468 & w36025);
assign w2496 = pi0588 & pi0705;
assign w2497 = ~w2495 & w2496;
assign w2498 = ~w2494 & ~w2497;
assign w2499 = ~w2493 & w2498;
assign w2500 = w2481 & ~w2499;
assign w2501 = (pi0515 & w2469) | (pi0515 & w36026) | (w2469 & w36026);
assign w2502 = ~pi0515 & pi0704;
assign w2503 = ~w2469 & w36027;
assign w2504 = ~w2501 & ~w2503;
assign w2505 = ~w2466 & ~w2504;
assign w2506 = pi0513 & w2505;
assign w2507 = (~w2476 & ~w2500) | (~w2476 & w36028) | (~w2500 & w36028);
assign w2508 = ~pi0670 & w2454;
assign w2509 = (w2427 & w2468) | (w2427 & w36029) | (w2468 & w36029);
assign w2510 = pi0703 & ~w2509;
assign w2511 = w2505 & w2510;
assign w2512 = w2500 & w2511;
assign w2513 = (~pi0513 & w2475) | (~pi0513 & w36030) | (w2475 & w36030);
assign w2514 = w2510 & ~w2513;
assign w2515 = ~w2512 & ~w2514;
assign w2516 = w2462 & w36031;
assign w2517 = ~pi0644 & w2454;
assign w2518 = w2454 & w2427;
assign w2519 = ~w2516 & w36032;
assign w2520 = ~pi0587 & ~w2519;
assign w2521 = w2432 & w36033;
assign w2522 = (~w2454 & ~w2462) | (~w2454 & w36034) | (~w2462 & w36034);
assign w2523 = (~pi0511 & ~w2522) | (~pi0511 & w36035) | (~w2522 & w36035);
assign w2524 = ~w2468 & ~w2517;
assign w2525 = ~w2468 & w36036;
assign w2526 = ~pi0512 & ~w2525;
assign w2527 = (pi0520 & w2525) | (pi0520 & w36037) | (w2525 & w36037);
assign w2528 = ~w2523 & w2527;
assign w2529 = ~w2520 & w2528;
assign w2530 = (w2529 & ~w2515) | (w2529 & w36038) | (~w2515 & w36038);
assign w2531 = ~pi0676 & w2521;
assign w2532 = w2462 & ~w2531;
assign w2533 = (w2452 & ~w2449) | (w2452 & w36039) | (~w2449 & w36039);
assign w2534 = ~w2532 & w36040;
assign w2535 = w2522 & w36041;
assign w2536 = pi0520 & w2535;
assign w2537 = pi0587 & w2519;
assign w2538 = pi0512 & w2525;
assign w2539 = ~w2537 & ~w2538;
assign w2540 = w2528 & ~w2539;
assign w2541 = ~w2536 & ~w2540;
assign w2542 = ~w2540 & w36042;
assign w2543 = ~w2540 & w36043;
assign w2544 = ~w2530 & w2543;
assign w2545 = ~w2523 & ~w2535;
assign w2546 = ~w2526 & w2545;
assign w2547 = ~w2520 & w2546;
assign w2548 = (w2547 & ~w2515) | (w2547 & w36044) | (~w2515 & w36044);
assign w2549 = ~w2539 & w2546;
assign w2550 = (~pi0520 & ~w2522) | (~pi0520 & w36045) | (~w2522 & w36045);
assign w2551 = ~w2549 & w2550;
assign w2552 = ~w2549 & w36046;
assign w2553 = ~w2548 & w2552;
assign w2554 = ~w2544 & ~w2553;
assign w2555 = w2521 & w36047;
assign w2556 = (w2450 & ~w2521) | (w2450 & w36048) | (~w2521 & w36048);
assign w2557 = w2449 & w36049;
assign w2558 = pi0668 & ~w2451;
assign w2559 = w2557 & ~w2558;
assign w2560 = (~pi0675 & ~w2521) | (~pi0675 & w36050) | (~w2521 & w36050);
assign w2561 = (~w2556 & ~w2559) | (~w2556 & w36051) | (~w2559 & w36051);
assign w2562 = (~pi0589 & ~w2561) | (~pi0589 & w4488) | (~w2561 & w4488);
assign w2563 = w2557 & w36052;
assign w2564 = (pi0682 & w2557) | (pi0682 & w36053) | (w2557 & w36053);
assign w2565 = ~w2563 & w2564;
assign w2566 = ~w2562 & w2565;
assign w2567 = w2554 & w2566;
assign w2568 = ~w2548 & w2551;
assign w2569 = ~w2530 & w2542;
assign w2570 = ~w2568 & ~w2569;
assign w2571 = (w2561 & w36054) | (w2561 & w36055) | (w36054 & w36055);
assign w2572 = w2570 & w2571;
assign w2573 = ~w2567 & ~w2572;
assign w2574 = w2561 & w4491;
assign w2575 = (~w2555 & w2462) | (~w2555 & w36056) | (w2462 & w36056);
assign w2576 = pi0680 & ~w2575;
assign w2577 = (pi0518 & w2575) | (pi0518 & w36057) | (w2575 & w36057);
assign w2578 = ~w2574 & w2577;
assign w2579 = w2573 & w2578;
assign w2580 = pi0657 & pi0674;
assign w2581 = ~w2483 & ~w2580;
assign w2582 = w2481 & ~w2497;
assign w2583 = ~w2581 & w2582;
assign w2584 = w2581 & ~w2582;
assign w2585 = ~w2486 & ~w2494;
assign w2586 = ~w2584 & w2585;
assign w2587 = ~w2583 & w2586;
assign w2588 = ~pi0518 & pi0657;
assign w2589 = pi0518 & ~pi0657;
assign w2590 = ~w2588 & ~w2589;
assign w2591 = ~w2496 & w2590;
assign w2592 = w2470 & w2590;
assign w2593 = (w2592 & w2468) | (w2592 & w36058) | (w2468 & w36058);
assign w2594 = ~w2591 & ~w2593;
assign w2595 = w2481 & ~w2594;
assign w2596 = w2496 & ~w2590;
assign w2597 = ~w2495 & w2596;
assign w2598 = w2477 & ~w2590;
assign w2599 = w2479 & ~w2590;
assign w2600 = (w2599 & w2468) | (w2599 & w36059) | (w2468 & w36059);
assign w2601 = ~w2598 & ~w2600;
assign w2602 = ~w2597 & w2601;
assign w2603 = ~w2595 & w2602;
assign w2604 = w2494 & w2603;
assign w2605 = w2486 & ~w2603;
assign w2606 = ~w2604 & ~w2605;
assign w2607 = ~w2587 & w2606;
assign w2608 = ~pi0518 & pi0674;
assign w2609 = pi0518 & ~pi0674;
assign w2610 = ~w2608 & ~w2609;
assign w2611 = ~pi0516 & ~w2610;
assign w2612 = pi0516 & w2610;
assign w2613 = ~w2611 & ~w2612;
assign w2614 = ~w2485 & ~w2613;
assign w2615 = w2485 & w2613;
assign w2616 = ~w2614 & ~w2615;
assign w2617 = ~pi0518 & pi0673;
assign w2618 = pi0518 & ~pi0673;
assign w2619 = ~w2617 & ~w2618;
assign w2620 = ~pi0517 & ~w2619;
assign w2621 = pi0517 & w2619;
assign w2622 = ~w2620 & w40101;
assign w2623 = ~w2616 & ~w2622;
assign w2624 = w2616 & w2622;
assign w2625 = ~pi0518 & ~pi0656;
assign w2626 = w2487 & w2625;
assign w2627 = ~w2620 & ~w2621;
assign w2628 = ~w2627 & w40100;
assign w2629 = (w2462 & w36062) | (w2462 & w36063) | (w36062 & w36063);
assign w2630 = ~w2628 & ~w2629;
assign w2631 = ~pi0656 & ~pi0707;
assign w2632 = pi0521 & ~w2631;
assign w2633 = ~w2625 & ~w2632;
assign w2634 = ~w2626 & ~w2633;
assign w2635 = pi0656 & pi0707;
assign w2636 = (~w2634 & w2462) | (~w2634 & w36064) | (w2462 & w36064);
assign w2637 = ~w2630 & ~w2636;
assign w2638 = (~w2626 & w2630) | (~w2626 & w36065) | (w2630 & w36065);
assign w2639 = (w2638 & ~w2616) | (w2638 & w36066) | (~w2616 & w36066);
assign w2640 = ~w2623 & ~w2639;
assign w2641 = w2607 & w2640;
assign w2642 = (~w2612 & ~w2485) | (~w2612 & w36067) | (~w2485 & w36067);
assign w2643 = w2603 & ~w2642;
assign w2644 = ~w2469 & w36068;
assign w2645 = ~pi0515 & pi0518;
assign w2646 = pi0515 & ~pi0518;
assign w2647 = ~w2645 & ~w2646;
assign w2648 = ~pi0672 & w2647;
assign w2649 = pi0672 & ~w2647;
assign w2650 = ~w2648 & ~w2649;
assign w2651 = w2644 & ~w2650;
assign w2652 = ~w2644 & w2650;
assign w2653 = ~w2651 & ~w2652;
assign w2654 = ~w2497 & ~w2595;
assign w2655 = w2653 & ~w2654;
assign w2656 = ~w2643 & ~w2655;
assign w2657 = (w2656 & ~w2607) | (w2656 & w36069) | (~w2607 & w36069);
assign w2658 = ~w2497 & w2653;
assign w2659 = w2481 & ~w2653;
assign w2660 = ~w2658 & ~w2659;
assign w2661 = ~w2431 & ~w2444;
assign w2662 = w2504 & w2661;
assign w2663 = ~w2504 & ~w2661;
assign w2664 = w2582 & ~w2663;
assign w2665 = ~w2662 & w2664;
assign w2666 = ~w2660 & ~w2665;
assign w2667 = ~w2655 & ~w2666;
assign w2668 = ~pi0518 & pi0670;
assign w2669 = pi0518 & ~pi0670;
assign w2670 = ~w2668 & ~w2669;
assign w2671 = pi0513 & w2670;
assign w2672 = ~pi0513 & ~w2670;
assign w2673 = ~w2671 & ~w2672;
assign w2674 = ~w2509 & w36070;
assign w2675 = (~w2673 & w2509) | (~w2673 & w36071) | (w2509 & w36071);
assign w2676 = ~w2674 & ~w2675;
assign w2677 = ~pi0518 & pi0671;
assign w2678 = pi0518 & ~pi0671;
assign w2679 = ~w2677 & ~w2678;
assign w2680 = (~w2679 & ~w2465) | (~w2679 & w36072) | (~w2465 & w36072);
assign w2681 = ~w2466 & ~w2680;
assign w2682 = ~w2676 & ~w2681;
assign w2683 = ~w2520 & ~w2537;
assign w2684 = ~pi0518 & pi0669;
assign w2685 = pi0518 & ~pi0669;
assign w2686 = ~w2684 & ~w2685;
assign w2687 = ~w2671 & ~w2686;
assign w2688 = (w2687 & w2509) | (w2687 & w36073) | (w2509 & w36073);
assign w2689 = ~w2683 & w2688;
assign w2690 = ~w2671 & w2686;
assign w2691 = (w2690 & w2509) | (w2690 & w36074) | (w2509 & w36074);
assign w2692 = w2683 & w2691;
assign w2693 = ~w2689 & ~w2692;
assign w2694 = ~w2682 & w2693;
assign w2695 = pi0518 & pi0672;
assign w2696 = ~pi0518 & ~pi0672;
assign w2697 = ~w2695 & ~w2696;
assign w2698 = pi0515 & ~w2697;
assign w2699 = ~pi0672 & ~w2645;
assign w2700 = ~w2646 & ~w2695;
assign w2701 = (w2454 & w36076) | (w2454 & w36077) | (w36076 & w36077);
assign w2702 = ~w2469 & w36078;
assign w2703 = ~w2698 & ~w2702;
assign w2704 = ~w2466 & ~w2467;
assign w2705 = w2679 & ~w2704;
assign w2706 = ~w2679 & w2704;
assign w2707 = ~w2705 & ~w2706;
assign w2708 = w2703 & w2707;
assign w2709 = w2694 & ~w2708;
assign w2710 = ~w2667 & w2709;
assign w2711 = ~w2657 & w2710;
assign w2712 = w2676 & w2681;
assign w2713 = ~w2703 & ~w2707;
assign w2714 = (~w2712 & w2707) | (~w2712 & w36079) | (w2707 & w36079);
assign w2715 = w2694 & ~w2714;
assign w2716 = w2683 & w2686;
assign w2717 = (~w2671 & w2509) | (~w2671 & w36080) | (w2509 & w36080);
assign w2718 = (~w2717 & w2683) | (~w2717 & w36081) | (w2683 & w36081);
assign w2719 = ~w2716 & w2718;
assign w2720 = ~pi0512 & pi0518;
assign w2721 = pi0512 & ~pi0518;
assign w2722 = ~w2720 & ~w2721;
assign w2723 = pi0644 & ~w2722;
assign w2724 = ~pi0644 & w2722;
assign w2725 = ~w2723 & ~w2724;
assign w2726 = pi0512 & w2725;
assign w2727 = ~pi0644 & ~w2720;
assign w2728 = (~w2723 & w2454) | (~w2723 & w36082) | (w2454 & w36082);
assign w2729 = ~w2468 & w36083;
assign w2730 = ~w2726 & ~w2729;
assign w2731 = ~pi0518 & pi0668;
assign w2732 = pi0518 & ~pi0668;
assign w2733 = ~w2731 & ~w2732;
assign w2734 = ~w2545 & w2733;
assign w2735 = w2545 & ~w2733;
assign w2736 = ~w2734 & ~w2735;
assign w2737 = ~w2730 & ~w2736;
assign w2738 = (w2686 & w2519) | (w2686 & w36084) | (w2519 & w36084);
assign w2739 = ~w2537 & ~w2738;
assign w2740 = w2525 & ~w2725;
assign w2741 = ~w2525 & w2725;
assign w2742 = ~w2740 & ~w2741;
assign w2743 = ~w2739 & w2742;
assign w2744 = ~w2737 & ~w2743;
assign w2745 = ~w2719 & w2744;
assign w2746 = ~w2715 & w2745;
assign w2747 = ~pi0518 & pi0675;
assign w2748 = pi0518 & ~pi0675;
assign w2749 = ~w2747 & ~w2748;
assign w2750 = pi0519 & w2749;
assign w2751 = ~pi0519 & ~w2749;
assign w2752 = ~w2750 & ~w2751;
assign w2753 = w2565 & w2752;
assign w2754 = ~w2565 & ~w2752;
assign w2755 = ~w2753 & ~w2754;
assign w2756 = ~pi0518 & pi0676;
assign w2757 = pi0518 & ~pi0676;
assign w2758 = ~w2756 & ~w2757;
assign w2759 = ~pi0520 & ~w2758;
assign w2760 = pi0520 & w2758;
assign w2761 = (~w2759 & w2534) | (~w2759 & w36085) | (w2534 & w36085);
assign w2762 = ~w2755 & ~w2761;
assign w2763 = ~w2759 & ~w2760;
assign w2764 = w2534 & ~w2763;
assign w2765 = ~w2534 & w2763;
assign w2766 = ~w2764 & ~w2765;
assign w2767 = (w2522 & w36086) | (w2522 & w36087) | (w36086 & w36087);
assign w2768 = ~w2535 & ~w2767;
assign w2769 = ~w2766 & ~w2768;
assign w2770 = w2755 & w2761;
assign w2771 = ~w2769 & ~w2770;
assign w2772 = ~w2762 & ~w2771;
assign w2773 = (~w2750 & ~w2565) | (~w2750 & w36088) | (~w2565 & w36088);
assign w2774 = ~pi0518 & pi0646;
assign w2775 = pi0518 & ~pi0646;
assign w2776 = ~w2774 & ~w2775;
assign w2777 = ~pi0589 & w2776;
assign w2778 = pi0589 & ~w2776;
assign w2779 = ~w2777 & ~w2778;
assign w2780 = w2561 & w36089;
assign w2781 = (w2779 & ~w2561) | (w2779 & w36090) | (~w2561 & w36090);
assign w2782 = ~w2780 & ~w2781;
assign w2783 = ~w2773 & w2782;
assign w2784 = (~w2783 & w2771) | (~w2783 & w36091) | (w2771 & w36091);
assign w2785 = w2746 & w2784;
assign w2786 = ~w2711 & w2785;
assign w2787 = w2773 & ~w2782;
assign w2788 = w2739 & ~w2742;
assign w2789 = ~w2737 & w2788;
assign w2790 = w2730 & w2736;
assign w2791 = ~w2789 & ~w2790;
assign w2792 = w2766 & w2768;
assign w2793 = ~w2769 & ~w2792;
assign w2794 = ~w2762 & w2793;
assign w2795 = w2791 & w2794;
assign w2796 = (w2784 & ~w2791) | (w2784 & w36092) | (~w2791 & w36092);
assign w2797 = ~w2787 & ~w2796;
assign w2798 = (w2561 & w36093) | (w2561 & w36094) | (w36093 & w36094);
assign w2799 = ~w2574 & ~w2798;
assign w2800 = pi0645 & w2799;
assign w2801 = ~w2575 & w36095;
assign w2802 = (w2801 & ~w2799) | (w2801 & w36096) | (~w2799 & w36096);
assign w2803 = (w2802 & w2786) | (w2802 & w36097) | (w2786 & w36097);
assign w2804 = ~w2575 & w36098;
assign w2805 = (pi0645 & w2575) | (pi0645 & w36099) | (w2575 & w36099);
assign w2806 = ~w2804 & ~w2805;
assign w2807 = ~w2799 & w2806;
assign w2808 = w2784 & ~w2807;
assign w2809 = w2746 & w2808;
assign w2810 = ~w2711 & w2809;
assign w2811 = ~w2795 & w2808;
assign w2812 = w2799 & ~w2806;
assign w2813 = ~w2787 & ~w2812;
assign w2814 = ~w2807 & ~w2813;
assign w2815 = (~pi0518 & w2813) | (~pi0518 & w36100) | (w2813 & w36100);
assign w2816 = ~w2804 & w2815;
assign w2817 = (w2816 & w2795) | (w2816 & w36101) | (w2795 & w36101);
assign w2818 = ~w2810 & w2817;
assign w2819 = ~pi0645 & ~w2799;
assign w2820 = (w2801 & w2782) | (w2801 & w36102) | (w2782 & w36102);
assign w2821 = ~w2819 & w2820;
assign w2822 = ~w2796 & w2821;
assign w2823 = ~w2786 & w2822;
assign w2824 = ~w2818 & ~w2823;
assign w2825 = ~w2803 & w2824;
assign w2826 = ~w2579 & w2825;
assign w2827 = (pi0702 & w2516) | (pi0702 & w36103) | (w2516 & w36103);
assign w2828 = w2693 & ~w2719;
assign w2829 = ~w2827 & ~w2828;
assign w2830 = w2667 & ~w2713;
assign w2831 = w2656 & ~w2713;
assign w2832 = (~w2708 & w2641) | (~w2708 & w36104) | (w2641 & w36104);
assign w2833 = (~w2712 & ~w2832) | (~w2712 & w36105) | (~w2832 & w36105);
assign w2834 = ~w2682 & ~w2833;
assign w2835 = (w2829 & w2833) | (w2829 & w36106) | (w2833 & w36106);
assign w2836 = ~w2827 & w2828;
assign w2837 = ~w2833 & w36107;
assign w2838 = ~w2835 & ~w2837;
assign w2839 = ~w2826 & w2838;
assign w2840 = w2515 & w36108;
assign w2841 = (~w2683 & ~w2515) | (~w2683 & w36109) | (~w2515 & w36109);
assign w2842 = ~w2827 & ~w2841;
assign w2843 = ~w2840 & w2842;
assign w2844 = w2826 & ~w2843;
assign w2845 = ~w2839 & ~w2844;
assign w2846 = w2425 & w2845;
assign w2847 = ~w2416 & w2846;
assign w2848 = w2387 & ~w2397;
assign w2849 = w2425 & ~w2848;
assign w2850 = pi1977 & w1309;
assign w2851 = ~w414 & w36110;
assign w2852 = ~w2850 & ~w2851;
assign w2853 = pi2272 & w1316;
assign w2854 = pi2262 & w1314;
assign w2855 = ~w2853 & ~w2854;
assign w2856 = w2852 & w2855;
assign w2857 = ~w414 & w36111;
assign w2858 = ~w392 & w36112;
assign w2859 = ~w2857 & ~w2858;
assign w2860 = ~w371 & w36113;
assign w2861 = ~w405 & w36114;
assign w2862 = ~w2860 & ~w2861;
assign w2863 = w2859 & w2862;
assign w2864 = ~w354 & ~w2863;
assign w2865 = w2856 & ~w2864;
assign w2866 = (w2417 & w2864) | (w2417 & w36115) | (w2864 & w36115);
assign w2867 = (pi2454 & w2330) | (pi2454 & w36116) | (w2330 & w36116);
assign w2868 = pi3093 & ~w2342;
assign w2869 = ~w2867 & ~w2868;
assign w2870 = (pi2962 & w2346) | (pi2962 & w36117) | (w2346 & w36117);
assign w2871 = (pi2462 & w2336) | (pi2462 & w36118) | (w2336 & w36118);
assign w2872 = ~w2870 & ~w2871;
assign w2873 = w2869 & w2872;
assign w2874 = w2869 & w36119;
assign w2875 = (w341 & w36121) | (w341 & w36122) | (w36121 & w36122);
assign w2876 = w2297 & w2875;
assign w2877 = pi2462 & w2876;
assign w2878 = (pi2962 & w2314) | (pi2962 & w36123) | (w2314 & w36123);
assign w2879 = w2316 & w2878;
assign w2880 = w354 & ~w2879;
assign w2881 = ~w2323 & w2324;
assign w2882 = pi3093 & w2881;
assign w2883 = (pi2454 & w2293) | (pi2454 & w36124) | (w2293 & w36124);
assign w2884 = w2295 & w2883;
assign w2885 = ~w2882 & ~w2884;
assign w2886 = w2885 & w36125;
assign w2887 = ~w2874 & ~w2886;
assign w2888 = ~w2886 & w36126;
assign w2889 = ~pi2048 & ~pi2986;
assign w2890 = w892 & ~w893;
assign w2891 = ~w2889 & w2890;
assign w2892 = w904 & w2891;
assign w2893 = pi2990 & w2889;
assign w2894 = (~pi2986 & ~w2889) | (~pi2986 & w893) | (~w2889 & w893);
assign w2895 = pi3099 & w892;
assign w2896 = ~w2894 & w2895;
assign w2897 = w889 & w2896;
assign w2898 = ~w2892 & ~w2897;
assign w2899 = (~w2898 & ~w886) | (~w2898 & w36127) | (~w886 & w36127);
assign w2900 = w940 & w36128;
assign w2901 = pi0403 & w2236;
assign w2902 = w2236 & w36129;
assign w2903 = (~w2900 & ~w359) | (~w2900 & w36131) | (~w359 & w36131);
assign w2904 = ~w2899 & w2903;
assign w2905 = (w353 & w36133) | (w353 & w36134) | (w36133 & w36134);
assign w2906 = w2905 & w40102;
assign w2907 = w359 & w2361;
assign w2908 = w933 & ~w2907;
assign w2909 = (pi1031 & w2907) | (pi1031 & w36135) | (w2907 & w36135);
assign w2910 = ~w2906 & ~w2909;
assign w2911 = w2904 & w2910;
assign w2912 = ~w2888 & w2911;
assign w2913 = ~w2866 & w2912;
assign w2914 = ~pi0773 & w2899;
assign w2915 = (~w2914 & w2386) | (~w2914 & w36136) | (w2386 & w36136);
assign w2916 = ~w2913 & w2915;
assign w2917 = (pi2961 & w2346) | (pi2961 & w36137) | (w2346 & w36137);
assign w2918 = (pi2461 & w2336) | (pi2461 & w36138) | (w2336 & w36138);
assign w2919 = ~w2917 & ~w2918;
assign w2920 = (pi2453 & w2330) | (pi2453 & w36139) | (w2330 & w36139);
assign w2921 = pi3096 & ~w2342;
assign w2922 = ~w2920 & ~w2921;
assign w2923 = w2919 & w2922;
assign w2924 = w2922 & w36140;
assign w2925 = pi2461 & w2876;
assign w2926 = (pi2961 & w2314) | (pi2961 & w36141) | (w2314 & w36141);
assign w2927 = w2316 & w2926;
assign w2928 = w354 & ~w2927;
assign w2929 = pi3096 & w2881;
assign w2930 = (pi2453 & w2293) | (pi2453 & w36142) | (w2293 & w36142);
assign w2931 = w2295 & w2930;
assign w2932 = ~w2929 & ~w2931;
assign w2933 = w2932 & w36143;
assign w2934 = ~w2924 & ~w2933;
assign w2935 = ~w2386 & w36144;
assign w2936 = ~w2425 & ~w2935;
assign w2937 = ~w2916 & w2936;
assign w2938 = ~w2397 & ~w2937;
assign w2939 = (w2938 & ~w2415) | (w2938 & w36145) | (~w2415 & w36145);
assign w2940 = ~w2847 & w2939;
assign w2941 = w2387 & ~w2425;
assign w2942 = ~w2682 & ~w2712;
assign w2943 = pi0703 & w2509;
assign w2944 = w2942 & ~w2943;
assign w2945 = w2832 & w36146;
assign w2946 = ~w2942 & ~w2943;
assign w2947 = (w2946 & ~w2832) | (w2946 & w36147) | (~w2832 & w36147);
assign w2948 = ~w2945 & ~w2947;
assign w2949 = ~w2826 & ~w2948;
assign w2950 = ~w2499 & w36148;
assign w2951 = w2513 & ~w2950;
assign w2952 = w2507 & ~w2951;
assign w2953 = ~pi0703 & ~w2952;
assign w2954 = w2507 & ~w2515;
assign w2955 = ~w2953 & ~w2954;
assign w2956 = w2826 & ~w2955;
assign w2957 = ~w2949 & ~w2956;
assign w2958 = ~w2387 & w2425;
assign w2959 = w2865 & ~w2887;
assign w2960 = w2958 & ~w2959;
assign w2961 = ~w2387 & ~w2425;
assign w2962 = pi3866 & w983;
assign w2963 = w973 & w36149;
assign w2964 = w970 & w36150;
assign w2965 = w973 & w36151;
assign w2966 = ~w2964 & ~w2965;
assign w2967 = ~w2963 & w2966;
assign w2968 = w958 & w36152;
assign w2969 = w963 & w36153;
assign w2970 = w953 & w36154;
assign w2971 = ~w2969 & ~w2970;
assign w2972 = ~w2968 & w2971;
assign w2973 = w970 & w36155;
assign w2974 = w963 & w36156;
assign w2975 = ~w997 & ~w2974;
assign w2976 = ~w2973 & w2975;
assign w2977 = w2972 & w2976;
assign w2978 = w2967 & w2977;
assign w2979 = ~w2962 & w2978;
assign w2980 = w940 & w36157;
assign w2981 = (pi1331 & ~w1730) | (pi1331 & w36158) | (~w1730 & w36158);
assign w2982 = pi1053 & pi2409;
assign w2983 = pi0384 & pi1057;
assign w2984 = pi0914 & pi1358;
assign w2985 = ~w2983 & ~w2984;
assign w2986 = ~w2982 & w2985;
assign w2987 = pi3516 & ~w1054;
assign w2988 = pi1334 & pi3285;
assign w2989 = pi0571 & pi1359;
assign w2990 = ~w2988 & ~w2989;
assign w2991 = ~w2987 & w2990;
assign w2992 = w2986 & w2991;
assign w2993 = (pi0650 & w2981) | (pi0650 & w36159) | (w2981 & w36159);
assign w2994 = pi1339 & pi2245;
assign w2995 = pi1346 & pi2663;
assign w2996 = ~w2994 & ~w2995;
assign w2997 = pi1351 & pi2439;
assign w2998 = pi1348 & pi2688;
assign w2999 = ~w2997 & ~w2998;
assign w3000 = w2996 & w2999;
assign w3001 = pi1338 & pi2231;
assign w3002 = pi1353 & pi2276;
assign w3003 = ~w3001 & ~w3002;
assign w3004 = pi1347 & pi2677;
assign w3005 = pi1352 & pi2702;
assign w3006 = ~w3004 & ~w3005;
assign w3007 = w3003 & w3006;
assign w3008 = pi1350 & pi2699;
assign w3009 = pi1337 & pi2217;
assign w3010 = ~w3008 & ~w3009;
assign w3011 = pi1600 & pi2203;
assign w3012 = pi1345 & pi2649;
assign w3013 = ~w3011 & ~w3012;
assign w3014 = w3010 & w3013;
assign w3015 = w3007 & w3014;
assign w3016 = (pi0722 & ~w3015) | (pi0722 & w36160) | (~w3015 & w36160);
assign w3017 = pi1341 & pi2293;
assign w3018 = pi1055 & pi2531;
assign w3019 = ~w3017 & ~w3018;
assign w3020 = pi1355 & pi2453;
assign w3021 = pi1054 & pi2710;
assign w3022 = ~w3020 & ~w3021;
assign w3023 = w3019 & w3022;
assign w3024 = pi1340 & pi2281;
assign w3025 = pi1354 & pi2961;
assign w3026 = ~w3024 & ~w3025;
assign w3027 = pi1056 & pi2548;
assign w3028 = pi1343 & pi2316;
assign w3029 = ~w3027 & ~w3028;
assign w3030 = w3026 & w3029;
assign w3031 = pi1342 & pi2304;
assign w3032 = pi1357 & pi2461;
assign w3033 = ~w3031 & ~w3032;
assign w3034 = pi1349 & pi2729;
assign w3035 = pi1356 & pi3096;
assign w3036 = ~w3034 & ~w3035;
assign w3037 = w3033 & w3036;
assign w3038 = w3030 & w3037;
assign w3039 = (pi0539 & ~w3038) | (pi0539 & w36161) | (~w3038 & w36161);
assign w3040 = pi0247 & pi1336;
assign w3041 = pi1335 & pi2585;
assign w3042 = ~w3040 & ~w3041;
assign w3043 = pi1333 & pi1867;
assign w3044 = pi1332 & pi2569;
assign w3045 = ~w3043 & ~w3044;
assign w3046 = w3042 & w3045;
assign w3047 = pi0762 & ~w3046;
assign w3048 = ~w3039 & ~w3047;
assign w3049 = ~w3016 & w3048;
assign w3050 = pi0979 & pi3151;
assign w3051 = ~pi0979 & pi2862;
assign w3052 = ~w3050 & ~w3051;
assign w3053 = pi0763 & ~w3052;
assign w3054 = pi0979 & pi3125;
assign w3055 = ~pi0979 & pi3075;
assign w3056 = ~w3054 & ~w3055;
assign w3057 = pi0766 & ~w3056;
assign w3058 = pi0313 & ~pi0979;
assign w3059 = pi0312 & pi0979;
assign w3060 = ~w3058 & ~w3059;
assign w3061 = pi0721 & ~w3060;
assign w3062 = ~w3057 & ~w3061;
assign w3063 = ~w3053 & w3062;
assign w3064 = pi0979 & pi3160;
assign w3065 = ~pi0979 & pi2870;
assign w3066 = ~w3064 & ~w3065;
assign w3067 = pi0764 & ~w3066;
assign w3068 = ~w1144 & ~w3067;
assign w3069 = pi0979 & pi3169;
assign w3070 = ~pi0979 & pi2632;
assign w3071 = ~w3069 & ~w3070;
assign w3072 = pi0765 & ~w3071;
assign w3073 = pi0138 & ~pi0979;
assign w3074 = pi0136 & pi0979;
assign w3075 = ~w3073 & ~w3074;
assign w3076 = pi0720 & ~w3075;
assign w3077 = ~w3072 & ~w3076;
assign w3078 = w3068 & w3077;
assign w3079 = w3063 & w3078;
assign w3080 = pi0524 & ~w3079;
assign w3081 = pi0169 & ~pi0979;
assign w3082 = pi0155 & pi0979;
assign w3083 = ~w3081 & ~w3082;
assign w3084 = pi0586 & pi1360;
assign w3085 = (~w3084 & w3083) | (~w3084 & w36162) | (w3083 & w36162);
assign w3086 = pi0979 & pi1957;
assign w3087 = ~pi0979 & pi2422;
assign w3088 = ~w3086 & ~w3087;
assign w3089 = pi0768 & ~w3088;
assign w3090 = pi0979 & pi2179;
assign w3091 = ~pi0979 & pi2784;
assign w3092 = ~w3090 & ~w3091;
assign w3093 = pi0837 & ~w3092;
assign w3094 = ~w3089 & ~w3093;
assign w3095 = pi0979 & pi2146;
assign w3096 = ~pi0979 & pi2918;
assign w3097 = ~w3095 & ~w3096;
assign w3098 = pi0767 & ~w3097;
assign w3099 = pi0979 & pi2163;
assign w3100 = ~pi0979 & pi2932;
assign w3101 = ~w3099 & ~w3100;
assign w3102 = pi0836 & ~w3101;
assign w3103 = ~w3098 & ~w3102;
assign w3104 = w3094 & w3103;
assign w3105 = (pi0576 & ~w3104) | (pi0576 & w36163) | (~w3104 & w36163);
assign w3106 = pi0280 & ~pi0979;
assign w3107 = pi0279 & pi0979;
assign w3108 = ~w3106 & ~w3107;
assign w3109 = pi0716 & ~w3108;
assign w3110 = pi0253 & ~pi0979;
assign w3111 = pi0250 & pi0979;
assign w3112 = ~w3110 & ~w3111;
assign w3113 = pi0761 & ~w3112;
assign w3114 = pi0979 & pi2126;
assign w3115 = ~pi0979 & pi2843;
assign w3116 = ~w3114 & ~w3115;
assign w3117 = pi0717 & ~w3116;
assign w3118 = ~w3113 & ~w3117;
assign w3119 = ~w3109 & w3118;
assign w3120 = w1184 & w3119;
assign w3121 = (pi0538 & ~w3119) | (pi0538 & w35782) | (~w3119 & w35782);
assign w3122 = ~w3105 & ~w3121;
assign w3123 = ~w3080 & w3122;
assign w3124 = w3049 & w3123;
assign w3125 = ~w2993 & w3124;
assign w3126 = ~w941 & ~w3125;
assign w3127 = pi1033 & w1225;
assign w3128 = w1221 & w36164;
assign w3129 = w1216 & w36165;
assign w3130 = ~w3128 & ~w3129;
assign w3131 = w1221 & w36166;
assign w3132 = w1216 & w36167;
assign w3133 = ~w3131 & ~w3132;
assign w3134 = w3130 & w3133;
assign w3135 = pi0948 & w1291;
assign w3136 = pi1774 & w1258;
assign w3137 = ~w3135 & ~w3136;
assign w3138 = pi1830 & w1268;
assign w3139 = w1226 & w1257;
assign w3140 = pi1427 & w3139;
assign w3141 = ~w3138 & ~w3140;
assign w3142 = w3137 & w3141;
assign w3143 = pi0800 & w1234;
assign w3144 = ~pi1032 & w1256;
assign w3145 = w1226 & w3144;
assign w3146 = pi1938 & w3145;
assign w3147 = ~w3143 & ~w3146;
assign w3148 = w1226 & w1241;
assign w3149 = pi1452 & w3148;
assign w3150 = pi0876 & w1296;
assign w3151 = ~w3149 & ~w3150;
assign w3152 = w3147 & w3151;
assign w3153 = w3142 & w3152;
assign w3154 = pi2103 & w1275;
assign w3155 = pi1438 & w1280;
assign w3156 = ~w3154 & ~w3155;
assign w3157 = pi1020 & w1266;
assign w3158 = pi0956 & w1245;
assign w3159 = ~w3157 & ~w3158;
assign w3160 = w3156 & w3159;
assign w3161 = pi1921 & w1272;
assign w3162 = pi0496 & w1242;
assign w3163 = ~w3161 & ~w3162;
assign w3164 = pi2055 & w1238;
assign w3165 = pi0963 & w1288;
assign w3166 = ~w3164 & ~w3165;
assign w3167 = w3163 & w3166;
assign w3168 = w3160 & w3167;
assign w3169 = w3153 & w3168;
assign w3170 = w1221 & w36168;
assign w3171 = pi1706 & w1294;
assign w3172 = w1237 & w3144;
assign w3173 = pi1729 & w3172;
assign w3174 = ~w3171 & ~w3173;
assign w3175 = pi1857 & w1263;
assign w3176 = pi0880 & w1251;
assign w3177 = ~w3175 & ~w3176;
assign w3178 = w3174 & w3177;
assign w3179 = pi1751 & w1249;
assign w3180 = w1205 & w3144;
assign w3181 = ~w3179 & ~w3180;
assign w3182 = pi0742 & w1254;
assign w3183 = pi1884 & w1278;
assign w3184 = ~w3182 & ~w3183;
assign w3185 = w3181 & w3184;
assign w3186 = w3178 & w3185;
assign w3187 = ~w3170 & w3186;
assign w3188 = w3169 & w3187;
assign w3189 = (pi1934 & ~w3188) | (pi1934 & w36169) | (~w3188 & w36169);
assign w3190 = ~w3126 & ~w3189;
assign w3191 = ~w3126 & w36170;
assign w3192 = pi1787 & pi2826;
assign w3193 = w958 & w36171;
assign w3194 = (w3193 & w3191) | (w3193 & w36172) | (w3191 & w36172);
assign w3195 = ~w2979 & ~w3194;
assign w3196 = w2961 & w3195;
assign w3197 = w940 & w36173;
assign w3198 = w1221 & w36174;
assign w3199 = w1216 & w36175;
assign w3200 = ~w3198 & ~w3199;
assign w3201 = w1216 & w36176;
assign w3202 = w1221 & w36177;
assign w3203 = ~w3201 & ~w3202;
assign w3204 = w3200 & w3203;
assign w3205 = pi1453 & w3148;
assign w3206 = pi1730 & w3172;
assign w3207 = ~w3205 & ~w3206;
assign w3208 = pi1099 & w1266;
assign w3209 = pi1716 & w1294;
assign w3210 = ~w3208 & ~w3209;
assign w3211 = w3207 & w3210;
assign w3212 = pi1752 & w1249;
assign w3213 = pi0577 & w1242;
assign w3214 = ~w3212 & ~w3213;
assign w3215 = pi0904 & w1296;
assign w3216 = pi1831 & w1268;
assign w3217 = ~w3215 & ~w3216;
assign w3218 = w3214 & w3217;
assign w3219 = w3211 & w3218;
assign w3220 = pi1885 & w1278;
assign w3221 = pi0801 & w1234;
assign w3222 = ~w3220 & ~w3221;
assign w3223 = pi1428 & w3139;
assign w3224 = pi0743 & w1254;
assign w3225 = ~w3223 & ~w3224;
assign w3226 = w3222 & w3225;
assign w3227 = pi1775 & w1258;
assign w3228 = pi1939 & w3145;
assign w3229 = ~w3227 & ~w3228;
assign w3230 = pi1763 & w1263;
assign w3231 = pi1922 & w1272;
assign w3232 = ~w3230 & ~w3231;
assign w3233 = w3229 & w3232;
assign w3234 = w3226 & w3233;
assign w3235 = w3219 & w3234;
assign w3236 = w1221 & w36178;
assign w3237 = pi0954 & w1245;
assign w3238 = pi0964 & w1288;
assign w3239 = ~w3237 & ~w3238;
assign w3240 = pi1899 & w1238;
assign w3241 = pi0881 & w1251;
assign w3242 = ~w3240 & ~w3241;
assign w3243 = w3239 & w3242;
assign w3244 = pi0949 & w1291;
assign w3245 = ~w3180 & ~w3244;
assign w3246 = pi2104 & w1275;
assign w3247 = pi1439 & w1280;
assign w3248 = ~w3246 & ~w3247;
assign w3249 = w3245 & w3248;
assign w3250 = w3243 & w3249;
assign w3251 = ~w3236 & w3250;
assign w3252 = w3235 & w3251;
assign w3253 = (pi1934 & ~w3252) | (pi1934 & w36179) | (~w3252 & w36179);
assign w3254 = pi0572 & pi1359;
assign w3255 = pi1053 & pi2473;
assign w3256 = ~w3254 & ~w3255;
assign w3257 = pi0915 & pi1358;
assign w3258 = pi0385 & pi1057;
assign w3259 = ~w3257 & ~w3258;
assign w3260 = w3256 & w3259;
assign w3261 = pi3517 & ~w1054;
assign w3262 = pi0826 & pi1344;
assign w3263 = pi1334 & pi2767;
assign w3264 = ~w3262 & ~w3263;
assign w3265 = ~w3261 & w3264;
assign w3266 = w3260 & w3265;
assign w3267 = (w3266 & w1808) | (w3266 & w36180) | (w1808 & w36180);
assign w3268 = pi0650 & ~w3267;
assign w3269 = pi1343 & pi2317;
assign w3270 = pi1054 & pi2711;
assign w3271 = ~w3269 & ~w3270;
assign w3272 = pi1349 & pi2730;
assign w3273 = pi1356 & pi3093;
assign w3274 = ~w3272 & ~w3273;
assign w3275 = w3271 & w3274;
assign w3276 = pi1355 & pi2454;
assign w3277 = pi1342 & pi2305;
assign w3278 = ~w3276 & ~w3277;
assign w3279 = pi1055 & pi2528;
assign w3280 = pi1354 & pi2962;
assign w3281 = ~w3279 & ~w3280;
assign w3282 = w3278 & w3281;
assign w3283 = pi1357 & pi2462;
assign w3284 = pi1341 & pi2294;
assign w3285 = ~w3283 & ~w3284;
assign w3286 = pi1340 & pi2282;
assign w3287 = pi1056 & pi2740;
assign w3288 = ~w3286 & ~w3287;
assign w3289 = w3285 & w3288;
assign w3290 = w3282 & w3289;
assign w3291 = (pi0539 & ~w3290) | (pi0539 & w36181) | (~w3290 & w36181);
assign w3292 = pi1353 & pi1977;
assign w3293 = pi1351 & pi2262;
assign w3294 = ~w3292 & ~w3293;
assign w3295 = pi1352 & pi2272;
assign w3296 = pi1348 & pi2563;
assign w3297 = ~w3295 & ~w3296;
assign w3298 = w3294 & w3297;
assign w3299 = pi1600 & pi2204;
assign w3300 = pi1345 & pi2650;
assign w3301 = ~w3299 & ~w3300;
assign w3302 = pi1338 & pi2232;
assign w3303 = pi1346 & pi2664;
assign w3304 = ~w3302 & ~w3303;
assign w3305 = w3301 & w3304;
assign w3306 = pi1350 & pi2258;
assign w3307 = pi1337 & pi2218;
assign w3308 = ~w3306 & ~w3307;
assign w3309 = pi1339 & pi2246;
assign w3310 = pi1347 & pi2678;
assign w3311 = ~w3309 & ~w3310;
assign w3312 = w3308 & w3311;
assign w3313 = w3305 & w3312;
assign w3314 = (pi0722 & ~w3313) | (pi0722 & w36182) | (~w3313 & w36182);
assign w3315 = pi0248 & pi1336;
assign w3316 = pi1332 & pi2570;
assign w3317 = ~w3315 & ~w3316;
assign w3318 = pi0368 & pi1333;
assign w3319 = pi1335 & pi2586;
assign w3320 = ~w3318 & ~w3319;
assign w3321 = w3317 & w3320;
assign w3322 = pi0762 & ~w3321;
assign w3323 = ~w3314 & ~w3322;
assign w3324 = ~w3291 & w3323;
assign w3325 = pi0979 & pi3161;
assign w3326 = ~pi0979 & pi2871;
assign w3327 = ~w3325 & ~w3326;
assign w3328 = pi0764 & ~w3327;
assign w3329 = pi0979 & pi3152;
assign w3330 = ~pi0979 & pi2863;
assign w3331 = ~w3329 & ~w3330;
assign w3332 = pi0763 & ~w3331;
assign w3333 = pi0054 & ~pi0979;
assign w3334 = pi0052 & pi0979;
assign w3335 = ~w3333 & ~w3334;
assign w3336 = pi0719 & ~w3335;
assign w3337 = ~w3332 & ~w3336;
assign w3338 = ~w3328 & w3337;
assign w3339 = pi0979 & pi3178;
assign w3340 = ~pi0979 & pi2890;
assign w3341 = ~w3339 & ~w3340;
assign w3342 = pi0766 & ~w3341;
assign w3343 = pi0979 & pi3133;
assign w3344 = ~pi0979 & pi2633;
assign w3345 = ~w3343 & ~w3344;
assign w3346 = pi0765 & ~w3345;
assign w3347 = ~w3342 & ~w3346;
assign w3348 = pi0131 & ~pi0979;
assign w3349 = pi0130 & pi0979;
assign w3350 = ~w3348 & ~w3349;
assign w3351 = pi0720 & ~w3350;
assign w3352 = pi0328 & ~pi0979;
assign w3353 = pi0327 & pi0979;
assign w3354 = ~w3352 & ~w3353;
assign w3355 = pi0721 & ~w3354;
assign w3356 = ~w3351 & ~w3355;
assign w3357 = w3347 & w3356;
assign w3358 = w3338 & w3357;
assign w3359 = pi0524 & ~w3358;
assign w3360 = pi0979 & pi1958;
assign w3361 = ~pi0979 & pi2423;
assign w3362 = ~w3360 & ~w3361;
assign w3363 = pi1360 & ~pi3633;
assign w3364 = (~w3363 & w3362) | (~w3363 & w36183) | (w3362 & w36183);
assign w3365 = pi0170 & ~pi0979;
assign w3366 = pi0156 & pi0979;
assign w3367 = ~w3365 & ~w3366;
assign w3368 = pi0838 & ~w3367;
assign w3369 = pi0979 & pi2180;
assign w3370 = ~pi0979 & pi2941;
assign w3371 = ~w3369 & ~w3370;
assign w3372 = pi0837 & ~w3371;
assign w3373 = ~w3368 & ~w3372;
assign w3374 = pi0979 & pi2164;
assign w3375 = ~pi0979 & pi2808;
assign w3376 = ~w3374 & ~w3375;
assign w3377 = pi0836 & ~w3376;
assign w3378 = pi0979 & pi2147;
assign w3379 = ~pi0979 & pi2919;
assign w3380 = ~w3378 & ~w3379;
assign w3381 = pi0767 & ~w3380;
assign w3382 = ~w3377 & ~w3381;
assign w3383 = w3373 & w3382;
assign w3384 = (pi0576 & ~w3383) | (pi0576 & w36184) | (~w3383 & w36184);
assign w3385 = pi0290 & ~pi0979;
assign w3386 = pi0287 & pi0979;
assign w3387 = ~w3385 & ~w3386;
assign w3388 = pi0761 & ~w3387;
assign w3389 = ~w1179 & ~w3388;
assign w3390 = pi0487 & ~pi0979;
assign w3391 = pi0484 & pi0979;
assign w3392 = ~w3390 & ~w3391;
assign w3393 = pi0718 & ~w3392;
assign w3394 = pi0264 & ~pi0979;
assign w3395 = pi0260 & pi0979;
assign w3396 = ~w3394 & ~w3395;
assign w3397 = pi0716 & ~w3396;
assign w3398 = pi0979 & pi2127;
assign w3399 = ~pi0979 & pi2844;
assign w3400 = ~w3398 & ~w3399;
assign w3401 = pi0717 & ~w3400;
assign w3402 = ~w3397 & ~w3401;
assign w3403 = ~w3393 & w3402;
assign w3404 = w3389 & w3403;
assign w3405 = (pi0538 & ~w3403) | (pi0538 & w36185) | (~w3403 & w36185);
assign w3406 = ~w3384 & ~w3405;
assign w3407 = ~w3359 & w3406;
assign w3408 = w3324 & w3407;
assign w3409 = ~w3268 & w3408;
assign w3410 = ~w941 & ~w3409;
assign w3411 = ~w3253 & ~w3410;
assign w3412 = ~w3410 & w36186;
assign w3413 = pi1787 & pi2819;
assign w3414 = w958 & w36187;
assign w3415 = pi3865 & w983;
assign w3416 = w973 & w36189;
assign w3417 = w973 & w36190;
assign w3418 = w970 & w36191;
assign w3419 = ~w3417 & ~w3418;
assign w3420 = ~w3416 & w3419;
assign w3421 = w958 & w36192;
assign w3422 = w953 & w36193;
assign w3423 = w963 & w36194;
assign w3424 = ~w3422 & ~w3423;
assign w3425 = ~w3421 & w3424;
assign w3426 = w970 & w36195;
assign w3427 = w963 & w36196;
assign w3428 = ~w997 & ~w3427;
assign w3429 = ~w3426 & w3428;
assign w3430 = w3425 & w3429;
assign w3431 = w3420 & w3430;
assign w3432 = ~w3415 & w3431;
assign w3433 = w2387 & w2425;
assign w3434 = w40134 & w3433;
assign w3435 = ~w3196 & ~w3434;
assign w3436 = ~w2960 & w3435;
assign w3437 = (w3436 & ~w2957) | (w3436 & w36199) | (~w2957 & w36199);
assign w3438 = w2397 & ~w3437;
assign w3439 = ~w2940 & ~w3438;
assign w3440 = w2397 & w2941;
assign w3441 = w2573 & ~w2574;
assign w3442 = (w2573 & w36201) | (w2573 & w36202) | (w36201 & w36202);
assign w3443 = w2746 & ~w2772;
assign w3444 = ~w2711 & w3443;
assign w3445 = (~w2772 & ~w2791) | (~w2772 & w36203) | (~w2791 & w36203);
assign w3446 = ~w2787 & ~w2800;
assign w3447 = (~pi0518 & w2799) | (~pi0518 & w36205) | (w2799 & w36205);
assign w3448 = w2783 & ~w2800;
assign w3449 = w3447 & ~w3448;
assign w3450 = (w3449 & w3444) | (w3449 & w36206) | (w3444 & w36206);
assign w3451 = (~pi0680 & w3441) | (~pi0680 & w36207) | (w3441 & w36207);
assign w3452 = ~w3442 & ~w3451;
assign w3453 = ~w2800 & ~w2819;
assign w3454 = pi0518 & ~w3453;
assign w3455 = ~pi0680 & ~w3447;
assign w3456 = ~w3453 & w3455;
assign w3457 = w2802 & ~w2819;
assign w3458 = ~w3456 & ~w3457;
assign w3459 = ~w2786 & w36209;
assign w3460 = (w2573 & w36210) | (w2573 & w36211) | (w36210 & w36211);
assign w3461 = ~w2579 & w3453;
assign w3462 = ~w2801 & ~w3453;
assign w3463 = (~w3462 & w2786) | (~w3462 & w36212) | (w2786 & w36212);
assign w3464 = (~w3460 & w3461) | (~w3460 & w36213) | (w3461 & w36213);
assign w3465 = ~w3452 & w3464;
assign w3466 = w3440 & ~w3465;
assign w3467 = pi3859 & w983;
assign w3468 = w973 & w36214;
assign w3469 = w970 & w36215;
assign w3470 = w973 & w36216;
assign w3471 = ~w3469 & ~w3470;
assign w3472 = ~w3468 & w3471;
assign w3473 = w958 & w36217;
assign w3474 = w963 & w36218;
assign w3475 = w953 & w36219;
assign w3476 = ~w3474 & ~w3475;
assign w3477 = ~w3473 & w3476;
assign w3478 = w970 & w36220;
assign w3479 = w963 & w36221;
assign w3480 = ~w997 & ~w3479;
assign w3481 = ~w3478 & w3480;
assign w3482 = w3477 & w3481;
assign w3483 = w3472 & w3482;
assign w3484 = ~w3467 & w3483;
assign w3485 = w940 & w36222;
assign w3486 = pi0393 & pi1057;
assign w3487 = pi0979 & pi1344;
assign w3488 = ~w3486 & ~w3487;
assign w3489 = pi0980 & pi1358;
assign w3490 = pi0585 & pi1359;
assign w3491 = ~w3489 & ~w3490;
assign w3492 = w3488 & w3491;
assign w3493 = pi3520 & ~w1054;
assign w3494 = pi1053 & pi2408;
assign w3495 = pi1047 & pi1334;
assign w3496 = ~w3494 & ~w3495;
assign w3497 = pi1059 & pi2981;
assign w3498 = pi1058 & pi3361;
assign w3499 = ~w3497 & ~w3498;
assign w3500 = w3496 & w3499;
assign w3501 = ~w3493 & w3500;
assign w3502 = w3492 & w3501;
assign w3503 = (w3502 & w1770) | (w3502 & w36223) | (w1770 & w36223);
assign w3504 = pi0650 & ~w3503;
assign w3505 = pi1339 & pi2256;
assign w3506 = pi1352 & pi2447;
assign w3507 = ~w3505 & ~w3506;
assign w3508 = pi1347 & pi2603;
assign w3509 = pi1600 & pi2214;
assign w3510 = ~w3508 & ~w3509;
assign w3511 = w3507 & w3510;
assign w3512 = pi1351 & pi2270;
assign w3513 = pi1350 & pi2437;
assign w3514 = ~w3512 & ~w3513;
assign w3515 = pi1337 & pi2228;
assign w3516 = pi1345 & pi2660;
assign w3517 = ~w3515 & ~w3516;
assign w3518 = w3514 & w3517;
assign w3519 = pi1348 & pi2562;
assign w3520 = pi1338 & pi2242;
assign w3521 = ~w3519 & ~w3520;
assign w3522 = pi1353 & pi1985;
assign w3523 = pi1346 & pi2674;
assign w3524 = ~w3522 & ~w3523;
assign w3525 = w3521 & w3524;
assign w3526 = w3518 & w3525;
assign w3527 = (pi0722 & ~w3526) | (pi0722 & w36224) | (~w3526 & w36224);
assign w3528 = pi1343 & pi2327;
assign w3529 = pi1055 & pi2727;
assign w3530 = ~w3528 & ~w3529;
assign w3531 = pi1357 & pi2470;
assign w3532 = pi1349 & pi2552;
assign w3533 = ~w3531 & ~w3532;
assign w3534 = w3530 & w3533;
assign w3535 = pi1355 & pi2524;
assign w3536 = pi1354 & pi2964;
assign w3537 = ~w3535 & ~w3536;
assign w3538 = pi1056 & pi2542;
assign w3539 = pi1356 & pi2968;
assign w3540 = ~w3538 & ~w3539;
assign w3541 = w3537 & w3540;
assign w3542 = pi1054 & pi2532;
assign w3543 = pi1341 & pi2302;
assign w3544 = ~w3542 & ~w3543;
assign w3545 = pi1340 & pi2291;
assign w3546 = pi1342 & pi2313;
assign w3547 = ~w3545 & ~w3546;
assign w3548 = w3544 & w3547;
assign w3549 = w3541 & w3548;
assign w3550 = (pi0539 & ~w3549) | (pi0539 & w36225) | (~w3549 & w36225);
assign w3551 = pi0128 & pi1333;
assign w3552 = pi0479 & pi1336;
assign w3553 = ~w3551 & ~w3552;
assign w3554 = pi1332 & pi2582;
assign w3555 = pi1335 & pi2597;
assign w3556 = ~w3554 & ~w3555;
assign w3557 = w3553 & w3556;
assign w3558 = pi0762 & ~w3557;
assign w3559 = ~w3550 & ~w3558;
assign w3560 = ~w3527 & w3559;
assign w3561 = pi0208 & ~pi0979;
assign w3562 = pi0205 & pi0979;
assign w3563 = ~w3561 & ~w3562;
assign w3564 = pi1599 & ~w3563;
assign w3565 = pi0333 & ~pi0979;
assign w3566 = pi0332 & pi0979;
assign w3567 = ~w3565 & ~w3566;
assign w3568 = pi0718 & ~w3567;
assign w3569 = ~w3564 & ~w3568;
assign w3570 = pi0979 & pi2139;
assign w3571 = ~pi0979 & pi2856;
assign w3572 = ~w3570 & ~w3571;
assign w3573 = pi0717 & ~w3572;
assign w3574 = pi0266 & ~pi0979;
assign w3575 = pi0262 & pi0979;
assign w3576 = ~w3574 & ~w3575;
assign w3577 = pi0716 & ~w3576;
assign w3578 = pi0311 & ~pi0979;
assign w3579 = pi0309 & pi0979;
assign w3580 = ~w3578 & ~w3579;
assign w3581 = pi0761 & ~w3580;
assign w3582 = ~w3577 & ~w3581;
assign w3583 = ~w3573 & w3582;
assign w3584 = w3569 & w3583;
assign w3585 = (pi0538 & ~w3583) | (pi0538 & w36226) | (~w3583 & w36226);
assign w3586 = pi0182 & ~pi0979;
assign w3587 = pi0174 & pi0979;
assign w3588 = ~w3586 & ~w3587;
assign w3589 = pi0149 & pi1360;
assign w3590 = (~w3589 & w3588) | (~w3589 & w36227) | (w3588 & w36227);
assign w3591 = pi0144 & ~pi0979;
assign w3592 = pi0129 & pi0979;
assign w3593 = ~w3591 & ~w3592;
assign w3594 = pi0768 & ~w3593;
assign w3595 = pi0979 & pi2192;
assign w3596 = ~pi0979 & pi2950;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = pi0837 & ~w3597;
assign w3599 = ~w3594 & ~w3598;
assign w3600 = pi0979 & pi2176;
assign w3601 = ~pi0979 & pi2938;
assign w3602 = ~w3600 & ~w3601;
assign w3603 = pi0836 & ~w3602;
assign w3604 = pi0979 & pi2158;
assign w3605 = ~pi0979 & pi2929;
assign w3606 = ~w3604 & ~w3605;
assign w3607 = pi0767 & ~w3606;
assign w3608 = ~w3603 & ~w3607;
assign w3609 = w3599 & w3608;
assign w3610 = (pi0576 & ~w3609) | (pi0576 & w36228) | (~w3609 & w36228);
assign w3611 = pi0088 & ~pi0979;
assign w3612 = pi0086 & pi0979;
assign w3613 = ~w3611 & ~w3612;
assign w3614 = pi0720 & ~w3613;
assign w3615 = pi0979 & pi3166;
assign w3616 = ~pi0979 & pi2879;
assign w3617 = ~w3615 & ~w3616;
assign w3618 = pi0764 & ~w3617;
assign w3619 = pi0979 & pi3202;
assign w3620 = ~pi0979 & pi2897;
assign w3621 = ~w3619 & ~w3620;
assign w3622 = pi0766 & ~w3621;
assign w3623 = ~w3618 & ~w3622;
assign w3624 = ~w3614 & w3623;
assign w3625 = pi0050 & ~pi0979;
assign w3626 = pi0049 & pi0979;
assign w3627 = ~w3625 & ~w3626;
assign w3628 = pi0719 & ~w3627;
assign w3629 = pi0751 & ~pi0979;
assign w3630 = pi0750 & pi0979;
assign w3631 = ~w3629 & ~w3630;
assign w3632 = pi0721 & ~w3631;
assign w3633 = ~w3628 & ~w3632;
assign w3634 = pi0979 & pi3127;
assign w3635 = ~pi0979 & pi2537;
assign w3636 = ~w3634 & ~w3635;
assign w3637 = pi0765 & ~w3636;
assign w3638 = pi0979 & pi3159;
assign w3639 = ~pi0979 & pi3084;
assign w3640 = ~w3638 & ~w3639;
assign w3641 = pi0763 & ~w3640;
assign w3642 = ~w3637 & ~w3641;
assign w3643 = w3633 & w3642;
assign w3644 = w3624 & w3643;
assign w3645 = pi0524 & ~w3644;
assign w3646 = ~w3645 & w36229;
assign w3647 = w3560 & w3646;
assign w3648 = ~w3504 & w3647;
assign w3649 = ~w941 & ~w3648;
assign w3650 = w1221 & w36230;
assign w3651 = w1216 & w36231;
assign w3652 = ~w3650 & ~w3651;
assign w3653 = w1221 & w36232;
assign w3654 = w1216 & w36233;
assign w3655 = ~w3653 & ~w3654;
assign w3656 = w3652 & w3655;
assign w3657 = pi1907 & w1238;
assign w3658 = pi1738 & w3172;
assign w3659 = ~w3657 & ~w3658;
assign w3660 = pi0849 & w1242;
assign w3661 = pi1726 & w1294;
assign w3662 = ~w3660 & ~w3661;
assign w3663 = w3659 & w3662;
assign w3664 = pi1786 & w1258;
assign w3665 = pi0741 & w1251;
assign w3666 = ~w3664 & ~w3665;
assign w3667 = pi0873 & w1296;
assign w3668 = pi1461 & w3148;
assign w3669 = ~w3667 & ~w3668;
assign w3670 = w3666 & w3669;
assign w3671 = w3663 & w3670;
assign w3672 = pi2110 & w1275;
assign w3673 = pi0967 & w1288;
assign w3674 = ~w3672 & ~w3673;
assign w3675 = pi0795 & w1245;
assign w3676 = pi1447 & w1280;
assign w3677 = ~w3675 & ~w3676;
assign w3678 = w3674 & w3677;
assign w3679 = pi1873 & w1278;
assign w3680 = pi1760 & w1249;
assign w3681 = ~w3679 & ~w3680;
assign w3682 = pi1434 & w3139;
assign w3683 = pi1769 & w1263;
assign w3684 = ~w3682 & ~w3683;
assign w3685 = w3681 & w3684;
assign w3686 = w3678 & w3685;
assign w3687 = w3671 & w3686;
assign w3688 = w1221 & w36234;
assign w3689 = pi1933 & w1272;
assign w3690 = pi0953 & w1291;
assign w3691 = ~w3689 & ~w3690;
assign w3692 = pi0805 & w1234;
assign w3693 = pi1945 & w3145;
assign w3694 = ~w3692 & ~w3693;
assign w3695 = w3691 & w3694;
assign w3696 = pi1839 & w1268;
assign w3697 = ~w3180 & ~w3696;
assign w3698 = pi1103 & w1266;
assign w3699 = pi0748 & w1254;
assign w3700 = ~w3698 & ~w3699;
assign w3701 = w3697 & w3700;
assign w3702 = w3695 & w3701;
assign w3703 = ~w3688 & w3702;
assign w3704 = w3687 & w3703;
assign w3705 = (pi1934 & ~w3704) | (pi1934 & w36235) | (~w3704 & w36235);
assign w3706 = ~w3649 & ~w3705;
assign w3707 = ~w3649 & w36236;
assign w3708 = pi1787 & pi2836;
assign w3709 = w958 & w36237;
assign w3710 = (w3709 & w3707) | (w3709 & w36238) | (w3707 & w36238);
assign w3711 = ~w3484 & ~w3710;
assign w3712 = w2961 & w3711;
assign w3713 = w1639 & w2425;
assign w3714 = w2387 & w3713;
assign w3715 = (pi2458 & w2330) | (pi2458 & w36239) | (w2330 & w36239);
assign w3716 = pi2530 & ~w2342;
assign w3717 = ~w3715 & ~w3716;
assign w3718 = (pi2748 & w2346) | (pi2748 & w36240) | (w2346 & w36240);
assign w3719 = (pi2410 & w2336) | (pi2410 & w36241) | (w2336 & w36241);
assign w3720 = ~w3718 & ~w3719;
assign w3721 = w3717 & w3720;
assign w3722 = w3717 & w36242;
assign w3723 = pi2410 & w2876;
assign w3724 = (pi2458 & w2293) | (pi2458 & w36243) | (w2293 & w36243);
assign w3725 = w2295 & w3724;
assign w3726 = w354 & ~w3725;
assign w3727 = (pi2748 & w2314) | (pi2748 & w36244) | (w2314 & w36244);
assign w3728 = w2316 & w3727;
assign w3729 = pi2530 & w2881;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = w3730 & w36245;
assign w3732 = ~w3722 & ~w3731;
assign w3733 = ~w354 & ~w1377;
assign w3734 = w1653 & ~w3733;
assign w3735 = ~w3732 & w3734;
assign w3736 = w2425 & ~w3735;
assign w3737 = ~w2387 & w3736;
assign w3738 = ~w3714 & ~w3737;
assign w3739 = (w2397 & ~w3738) | (w2397 & w36246) | (~w3738 & w36246);
assign w3740 = ~w2377 & ~w3734;
assign w3741 = ~w3731 & w36247;
assign w3742 = ~w1643 & ~w2899;
assign w3743 = w1642 & w40102;
assign w3744 = (pi1035 & w2907) | (pi1035 & w36248) | (w2907 & w36248);
assign w3745 = ~w3744 & w36249;
assign w3746 = pi0421 & w2901;
assign w3747 = w3745 & ~w3746;
assign w3748 = ~w3741 & w3747;
assign w3749 = ~w3740 & w3748;
assign w3750 = ~pi0752 & w2899;
assign w3751 = (~w3750 & ~w3745) | (~w3750 & w36250) | (~w3745 & w36250);
assign w3752 = ~w3749 & w3751;
assign w3753 = ~w2387 & ~w3752;
assign w3754 = ~w2397 & ~w2425;
assign w3755 = (pi2524 & w2330) | (pi2524 & w36251) | (w2330 & w36251);
assign w3756 = (pi2964 & w2346) | (pi2964 & w36252) | (w2346 & w36252);
assign w3757 = ~w3755 & ~w3756;
assign w3758 = (pi2470 & w2336) | (pi2470 & w36253) | (w2336 & w36253);
assign w3759 = pi2968 & ~w2342;
assign w3760 = ~w3758 & ~w3759;
assign w3761 = w3757 & w3760;
assign w3762 = w3760 & w36254;
assign w3763 = pi2470 & w2875;
assign w3764 = w2297 & w3763;
assign w3765 = (pi2964 & w2314) | (pi2964 & w36255) | (w2314 & w36255);
assign w3766 = w2316 & w3765;
assign w3767 = w354 & ~w3766;
assign w3768 = (pi2968 & w2322) | (pi2968 & w36256) | (w2322 & w36256);
assign w3769 = w2324 & w3768;
assign w3770 = (pi2524 & w2293) | (pi2524 & w36257) | (w2293 & w36257);
assign w3771 = w2295 & w3770;
assign w3772 = ~w3769 & ~w3771;
assign w3773 = w3767 & w3772;
assign w3774 = ~w3764 & w3773;
assign w3775 = ~w3762 & ~w3774;
assign w3776 = ~w2386 & w36258;
assign w3777 = w3754 & ~w3776;
assign w3778 = ~w3753 & w3777;
assign w3779 = ~w1367 & ~w3778;
assign w3780 = ~w3739 & w3779;
assign w3781 = (w3780 & w797) | (w3780 & w36259) | (w797 & w36259);
assign w3782 = ~w2397 & w2958;
assign w3783 = ~w3778 & ~w3782;
assign w3784 = ~w3739 & w3783;
assign w3785 = (~w3784 & w1357) | (~w3784 & w36260) | (w1357 & w36260);
assign w3786 = ~w2397 & w3433;
assign w3787 = ~pi0521 & ~pi0707;
assign w3788 = ~w2487 & ~w3787;
assign w3789 = pi0518 & w3788;
assign w3790 = (w3789 & ~w2573) | (w3789 & w36261) | (~w2573 & w36261);
assign w3791 = pi0656 & ~w3788;
assign w3792 = w2573 & w36262;
assign w3793 = ~w2810 & w36263;
assign w3794 = pi0518 & pi0645;
assign w3795 = (~w3794 & w2575) | (~w3794 & w36264) | (w2575 & w36264);
assign w3796 = (~w3788 & ~w2462) | (~w3788 & w36265) | (~w2462 & w36265);
assign w3797 = w3795 & w3796;
assign w3798 = ~pi0518 & pi0656;
assign w3799 = (w3798 & ~w3795) | (w3798 & w36266) | (~w3795 & w36266);
assign w3800 = ~w3793 & w3799;
assign w3801 = w3788 & ~w3795;
assign w3802 = (w2575 & w36267) | (w2575 & w36268) | (w36267 & w36268);
assign w3803 = (w2575 & w36271) | (w2575 & w36272) | (w36271 & w36272);
assign w3804 = ~w3802 & w3803;
assign w3805 = ~w3797 & ~w3804;
assign w3806 = (~w3801 & w3805) | (~w3801 & w36273) | (w3805 & w36273);
assign w3807 = w2815 & ~w3806;
assign w3808 = ~w2810 & w36274;
assign w3809 = ~pi0656 & w3788;
assign w3810 = (~w3809 & ~w2462) | (~w3809 & w36275) | (~w2462 & w36275);
assign w3811 = ~w3808 & w3810;
assign w3812 = ~w3800 & w3811;
assign w3813 = ~w3792 & w3812;
assign w3814 = ~w3790 & w3813;
assign w3815 = (w3786 & ~w3813) | (w3786 & w36276) | (~w3813 & w36276);
assign w3816 = ~w3785 & ~w3815;
assign w3817 = ~w3466 & w3816;
assign w3818 = (~w565 & w561) | (~w565 & w36277) | (w561 & w36277);
assign w3819 = pi0660 & w486;
assign w3820 = (~w3819 & w561) | (~w3819 & w36278) | (w561 & w36278);
assign w3821 = ~w3818 & w3820;
assign w3822 = (w3821 & ~w797) | (w3821 & w36279) | (~w797 & w36279);
assign w3823 = ~w659 & ~w719;
assign w3824 = ~w677 & ~w717;
assign w3825 = ~w677 & w702;
assign w3826 = (~w3824 & w647) | (~w3824 & w36280) | (w647 & w36280);
assign w3827 = w3823 & w3826;
assign w3828 = (~w3819 & w3826) | (~w3819 & w36281) | (w3826 & w36281);
assign w3829 = ~w3827 & w3828;
assign w3830 = w797 & w36282;
assign w3831 = ~w3822 & ~w3830;
assign w3832 = w2958 & w3831;
assign w3833 = (~w2472 & w2644) | (~w2472 & w36283) | (w2644 & w36283);
assign w3834 = ~w2500 & w3833;
assign w3835 = (pi0704 & w2469) | (pi0704 & w36284) | (w2469 & w36284);
assign w3836 = (~w3833 & w2500) | (~w3833 & w36285) | (w2500 & w36285);
assign w3837 = ~w3834 & ~w3836;
assign w3838 = w2826 & ~w3837;
assign w3839 = w2826 & w36286;
assign w3840 = w2666 & w40104;
assign w3841 = (w2607 & w36288) | (w2607 & w36289) | (w36288 & w36289);
assign w3842 = ~w3835 & ~w3841;
assign w3843 = ~w3840 & w3842;
assign w3844 = (w3433 & ~w3842) | (w3433 & w36290) | (~w3842 & w36290);
assign w3845 = (pi2452 & w2330) | (pi2452 & w36291) | (w2330 & w36291);
assign w3846 = (pi2413 & w2336) | (pi2413 & w36292) | (w2336 & w36292);
assign w3847 = ~w3845 & ~w3846;
assign w3848 = (pi2960 & w2346) | (pi2960 & w36293) | (w2346 & w36293);
assign w3849 = pi2965 & ~w2342;
assign w3850 = ~w3848 & ~w3849;
assign w3851 = w3847 & w3850;
assign w3852 = w3850 & w36294;
assign w3853 = pi2413 & w2875;
assign w3854 = w2297 & w3853;
assign w3855 = (pi2452 & w2293) | (pi2452 & w36295) | (w2293 & w36295);
assign w3856 = w2295 & w3855;
assign w3857 = w354 & ~w3856;
assign w3858 = (pi2960 & w2314) | (pi2960 & w36296) | (w2314 & w36296);
assign w3859 = w2316 & w3858;
assign w3860 = pi2965 & w2881;
assign w3861 = ~w3859 & ~w3860;
assign w3862 = w3861 & w36297;
assign w3863 = ~w3852 & ~w3862;
assign w3864 = ~w3862 & w36298;
assign w3865 = pi2261 & w1314;
assign w3866 = ~w414 & w36299;
assign w3867 = ~w3865 & ~w3866;
assign w3868 = pi2271 & w1316;
assign w3869 = pi1976 & w1309;
assign w3870 = ~w3868 & ~w3869;
assign w3871 = w3867 & w3870;
assign w3872 = ~w371 & w36300;
assign w3873 = ~w392 & w36301;
assign w3874 = ~w3872 & ~w3873;
assign w3875 = ~w414 & w36302;
assign w3876 = ~w405 & w36303;
assign w3877 = ~w3875 & ~w3876;
assign w3878 = w3874 & w3877;
assign w3879 = (~w354 & ~w3877) | (~w354 & w36304) | (~w3877 & w36304);
assign w3880 = w3871 & ~w3879;
assign w3881 = w2236 & w36305;
assign w3882 = (~w3881 & w3880) | (~w3881 & w36306) | (w3880 & w36306);
assign w3883 = (w2365 & ~w3882) | (w2365 & w36307) | (~w3882 & w36307);
assign w3884 = pi2448 & w941;
assign w3885 = ~w2899 & ~w3884;
assign w3886 = (w353 & w36308) | (w353 & w36309) | (w36308 & w36309);
assign w3887 = w3886 & w40102;
assign w3888 = (pi1028 & w2907) | (pi1028 & w36310) | (w2907 & w36310);
assign w3889 = ~w3888 & w36311;
assign w3890 = ~w3883 & w3889;
assign w3891 = ~pi0845 & w2899;
assign w3892 = w2961 & w36312;
assign w3893 = pi2455 & ~w2331;
assign w3894 = (pi2963 & w2346) | (pi2963 & w36313) | (w2346 & w36313);
assign w3895 = ~w3893 & ~w3894;
assign w3896 = (pi2464 & w2336) | (pi2464 & w36314) | (w2336 & w36314);
assign w3897 = pi2966 & ~w2342;
assign w3898 = ~w3896 & ~w3897;
assign w3899 = w3895 & w3898;
assign w3900 = ~w354 & w3899;
assign w3901 = pi2464 & w2875;
assign w3902 = w2297 & w3901;
assign w3903 = (pi2455 & w2293) | (pi2455 & w36315) | (w2293 & w36315);
assign w3904 = w2295 & w3903;
assign w3905 = w354 & ~w3904;
assign w3906 = pi2966 & w2881;
assign w3907 = ~w2315 & w2316;
assign w3908 = pi2963 & w3907;
assign w3909 = ~w3906 & ~w3908;
assign w3910 = w3909 & w36316;
assign w3911 = ~w3900 & ~w3910;
assign w3912 = (~w2397 & ~w2941) | (~w2397 & w36317) | (~w2941 & w36317);
assign w3913 = ~w3892 & w3912;
assign w3914 = (w3913 & w2826) | (w3913 & w36318) | (w2826 & w36318);
assign w3915 = ~w3839 & w3914;
assign w3916 = ~w3832 & w3915;
assign w3917 = ~w2715 & ~w2719;
assign w3918 = ~w2743 & ~w2788;
assign w3919 = ~w2711 & w36319;
assign w3920 = ~w2737 & ~w2790;
assign w3921 = ~w2788 & ~w3920;
assign w3922 = ~w3919 & w3921;
assign w3923 = (~w2789 & w2711) | (~w2789 & w36320) | (w2711 & w36320);
assign w3924 = pi0701 & ~w2522;
assign w3925 = (~w3924 & w3923) | (~w3924 & w36321) | (w3923 & w36321);
assign w3926 = ~w3922 & w3925;
assign w3927 = ~w2826 & w3926;
assign w3928 = (~w2520 & ~w2515) | (~w2520 & w36322) | (~w2515 & w36322);
assign w3929 = (~w2526 & w3928) | (~w2526 & w36323) | (w3928 & w36323);
assign w3930 = ~w2545 & w3929;
assign w3931 = (w3928 & w36326) | (w3928 & w36327) | (w36326 & w36327);
assign w3932 = ~w3930 & w3931;
assign w3933 = w2826 & w3932;
assign w3934 = ~w3927 & ~w3933;
assign w3935 = ~w3863 & w3880;
assign w3936 = (w2397 & ~w2958) | (w2397 & w36328) | (~w2958 & w36328);
assign w3937 = pi3868 & w983;
assign w3938 = w970 & w36329;
assign w3939 = w973 & w36330;
assign w3940 = w973 & w36331;
assign w3941 = ~w3939 & ~w3940;
assign w3942 = ~w3938 & w3941;
assign w3943 = w958 & w36332;
assign w3944 = w963 & w36333;
assign w3945 = w953 & w36334;
assign w3946 = ~w3944 & ~w3945;
assign w3947 = ~w3943 & w3946;
assign w3948 = w970 & w36335;
assign w3949 = w963 & w36336;
assign w3950 = ~w997 & ~w3949;
assign w3951 = ~w3948 & w3950;
assign w3952 = w3947 & w3951;
assign w3953 = w3942 & w3952;
assign w3954 = ~w3937 & w3953;
assign w3955 = w940 & w36337;
assign w3956 = (pi1331 & ~w2059) | (pi1331 & w36338) | (~w2059 & w36338);
assign w3957 = pi3514 & ~w1054;
assign w3958 = pi0382 & pi1057;
assign w3959 = pi0912 & pi1358;
assign w3960 = pi0590 & pi1359;
assign w3961 = ~w3959 & ~w3960;
assign w3962 = ~w3958 & w3961;
assign w3963 = ~w3957 & w3962;
assign w3964 = (pi0650 & w3956) | (pi0650 & w36339) | (w3956 & w36339);
assign w3965 = pi1351 & pi2261;
assign w3966 = pi1348 & pi2602;
assign w3967 = ~w3965 & ~w3966;
assign w3968 = pi1338 & pi2229;
assign w3969 = pi1346 & pi2661;
assign w3970 = ~w3968 & ~w3969;
assign w3971 = w3967 & w3970;
assign w3972 = pi1600 & pi2201;
assign w3973 = pi1347 & pi2675;
assign w3974 = ~w3972 & ~w3973;
assign w3975 = pi1337 & pi2215;
assign w3976 = pi1350 & pi2257;
assign w3977 = ~w3975 & ~w3976;
assign w3978 = w3974 & w3977;
assign w3979 = pi1339 & pi2243;
assign w3980 = pi1353 & pi1976;
assign w3981 = ~w3979 & ~w3980;
assign w3982 = pi1352 & pi2271;
assign w3983 = pi1345 & pi2550;
assign w3984 = ~w3982 & ~w3983;
assign w3985 = w3981 & w3984;
assign w3986 = w3978 & w3985;
assign w3987 = (pi0722 & ~w3986) | (pi0722 & w36340) | (~w3986 & w36340);
assign w3988 = pi1355 & pi2452;
assign w3989 = pi1054 & pi2708;
assign w3990 = ~w3988 & ~w3989;
assign w3991 = pi1356 & pi2965;
assign w3992 = pi1341 & pi2292;
assign w3993 = ~w3991 & ~w3992;
assign w3994 = w3990 & w3993;
assign w3995 = pi1357 & pi2413;
assign w3996 = pi1055 & pi2719;
assign w3997 = ~w3995 & ~w3996;
assign w3998 = pi1354 & pi2960;
assign w3999 = pi1340 & pi2279;
assign w4000 = ~w3998 & ~w3999;
assign w4001 = w3997 & w4000;
assign w4002 = pi1349 & pi2728;
assign w4003 = pi1343 & pi2314;
assign w4004 = ~w4002 & ~w4003;
assign w4005 = pi1342 & pi2303;
assign w4006 = pi1056 & pi2738;
assign w4007 = ~w4005 & ~w4006;
assign w4008 = w4004 & w4007;
assign w4009 = w4001 & w4008;
assign w4010 = (pi0539 & ~w4009) | (pi0539 & w36341) | (~w4009 & w36341);
assign w4011 = pi1333 & pi1742;
assign w4012 = pi1332 & pi2768;
assign w4013 = ~w4011 & ~w4012;
assign w4014 = pi0237 & pi1336;
assign w4015 = pi1335 & pi2583;
assign w4016 = ~w4014 & ~w4015;
assign w4017 = w4013 & w4016;
assign w4018 = pi0762 & ~w4017;
assign w4019 = ~w4010 & ~w4018;
assign w4020 = ~w3987 & w4019;
assign w4021 = pi0137 & ~pi0979;
assign w4022 = pi0135 & pi0979;
assign w4023 = ~w4021 & ~w4022;
assign w4024 = pi0720 & ~w4023;
assign w4025 = pi0979 & pi3126;
assign w4026 = ~pi0979 & pi2888;
assign w4027 = ~w4025 & ~w4026;
assign w4028 = pi0766 & ~w4027;
assign w4029 = pi0979 & pi3167;
assign w4030 = ~pi0979 & pi2630;
assign w4031 = ~w4029 & ~w4030;
assign w4032 = pi0765 & ~w4031;
assign w4033 = ~w4028 & ~w4032;
assign w4034 = ~w4024 & w4033;
assign w4035 = pi0979 & pi2618;
assign w4036 = ~pi0979 & pi2624;
assign w4037 = ~w4035 & ~w4036;
assign w4038 = pi0764 & ~w4037;
assign w4039 = ~w1144 & ~w4038;
assign w4040 = pi0268 & ~pi0979;
assign w4041 = pi0267 & pi0979;
assign w4042 = ~w4040 & ~w4041;
assign w4043 = pi0721 & ~w4042;
assign w4044 = pi0979 & pi2605;
assign w4045 = ~pi0979 & pi2611;
assign w4046 = ~w4044 & ~w4045;
assign w4047 = pi0763 & ~w4046;
assign w4048 = ~w4043 & ~w4047;
assign w4049 = w4039 & w4048;
assign w4050 = w4034 & w4049;
assign w4051 = pi0524 & ~w4050;
assign w4052 = pi0837 & pi2939;
assign w4053 = pi0767 & pi2916;
assign w4054 = pi0836 & pi2931;
assign w4055 = ~w4053 & ~w4054;
assign w4056 = (~pi0979 & ~w4055) | (~pi0979 & w36342) | (~w4055 & w36342);
assign w4057 = pi0837 & pi2177;
assign w4058 = pi0767 & pi2144;
assign w4059 = pi0836 & pi2161;
assign w4060 = ~w4058 & ~w4059;
assign w4061 = (pi0979 & ~w4060) | (pi0979 & w36343) | (~w4060 & w36343);
assign w4062 = pi0167 & ~pi0979;
assign w4063 = pi0153 & pi0979;
assign w4064 = ~w4062 & ~w4063;
assign w4065 = pi0838 & ~w4064;
assign w4066 = pi0979 & pi1955;
assign w4067 = ~pi0979 & pi2420;
assign w4068 = ~w4066 & ~w4067;
assign w4069 = pi0768 & ~w4068;
assign w4070 = ~w4065 & ~w4069;
assign w4071 = w4070 & w36344;
assign w4072 = pi0576 & ~w4071;
assign w4073 = pi0252 & ~pi0979;
assign w4074 = pi0249 & pi0979;
assign w4075 = ~w4073 & ~w4074;
assign w4076 = pi0761 & ~w4075;
assign w4077 = pi0979 & pi2124;
assign w4078 = ~pi0979 & pi2841;
assign w4079 = ~w4077 & ~w4078;
assign w4080 = pi0717 & ~w4079;
assign w4081 = pi0198 & ~pi0979;
assign w4082 = pi0197 & pi0979;
assign w4083 = ~w4081 & ~w4082;
assign w4084 = pi0716 & ~w4083;
assign w4085 = ~w4080 & ~w4084;
assign w4086 = ~w4076 & w4085;
assign w4087 = (pi0538 & ~w4086) | (pi0538 & w35782) | (~w4086 & w35782);
assign w4088 = ~w4072 & ~w4087;
assign w4089 = ~w4051 & w4088;
assign w4090 = w4020 & w4089;
assign w4091 = ~w3964 & w4090;
assign w4092 = ~w941 & ~w4091;
assign w4093 = w1221 & w36345;
assign w4094 = w1216 & w36346;
assign w4095 = ~w4093 & ~w4094;
assign w4096 = w1221 & w36347;
assign w4097 = w1216 & w36348;
assign w4098 = ~w4096 & ~w4097;
assign w4099 = w4095 & w4098;
assign w4100 = pi1450 & w3148;
assign w4101 = pi1772 & w1258;
assign w4102 = ~w4100 & ~w4101;
assign w4103 = pi0738 & w1251;
assign w4104 = pi1877 & w1294;
assign w4105 = ~w4103 & ~w4104;
assign w4106 = w4102 & w4105;
assign w4107 = pi1727 & w3172;
assign w4108 = pi0792 & w1245;
assign w4109 = ~w4107 & ~w4108;
assign w4110 = pi2057 & w1238;
assign w4111 = pi1436 & w1280;
assign w4112 = ~w4110 & ~w4111;
assign w4113 = w4109 & w4112;
assign w4114 = pi1828 & w1268;
assign w4115 = pi1918 & w1272;
assign w4116 = ~w4114 & ~w4115;
assign w4117 = pi0869 & w1254;
assign w4118 = pi0977 & w1234;
assign w4119 = ~w4117 & ~w4118;
assign w4120 = w4116 & w4119;
assign w4121 = w4113 & w4120;
assign w4122 = w4106 & w4121;
assign w4123 = w1221 & w36349;
assign w4124 = pi1952 & w1278;
assign w4125 = ~w3180 & ~w4124;
assign w4126 = pi0902 & w1296;
assign w4127 = pi0398 & w1242;
assign w4128 = ~w4126 & ~w4127;
assign w4129 = w4125 & w4128;
assign w4130 = w1288 & w36350;
assign w4131 = w1291 & w36351;
assign w4132 = ~w4130 & ~w4131;
assign w4133 = w4129 & w36352;
assign w4134 = w4122 & w36353;
assign w4135 = pi1934 & ~w4134;
assign w4136 = ~w4092 & ~w4135;
assign w4137 = ~w4092 & w36354;
assign w4138 = pi1787 & pi3149;
assign w4139 = w958 & w36355;
assign w4140 = (w4139 & w4137) | (w4139 & w36356) | (w4137 & w36356);
assign w4141 = ~w3954 & ~w4140;
assign w4142 = w3433 & w4141;
assign w4143 = pi3863 & w983;
assign w4144 = w970 & w36357;
assign w4145 = w973 & w36358;
assign w4146 = w973 & w36359;
assign w4147 = ~w4145 & ~w4146;
assign w4148 = ~w4144 & w4147;
assign w4149 = w958 & w36360;
assign w4150 = w963 & w36361;
assign w4151 = w953 & w36362;
assign w4152 = ~w4150 & ~w4151;
assign w4153 = ~w4149 & w4152;
assign w4154 = w970 & w36363;
assign w4155 = w963 & w36364;
assign w4156 = ~w997 & ~w4155;
assign w4157 = ~w4154 & w4156;
assign w4158 = w4153 & w4157;
assign w4159 = w4148 & w4158;
assign w4160 = ~w4143 & w4159;
assign w4161 = w940 & w36365;
assign w4162 = w1221 & w36366;
assign w4163 = w1221 & w36367;
assign w4164 = ~w4162 & ~w4163;
assign w4165 = w1216 & w36368;
assign w4166 = w1216 & w36369;
assign w4167 = ~w4165 & ~w4166;
assign w4168 = w4164 & w4167;
assign w4169 = pi1455 & w3148;
assign w4170 = pi1777 & w1258;
assign w4171 = ~w4169 & ~w4170;
assign w4172 = pi1732 & w3172;
assign w4173 = pi0745 & w1254;
assign w4174 = ~w4172 & ~w4173;
assign w4175 = w4171 & w4174;
assign w4176 = pi0900 & w1288;
assign w4177 = pi0883 & w1251;
assign w4178 = ~w4176 & ~w4177;
assign w4179 = pi0850 & w1234;
assign w4180 = pi0906 & w1296;
assign w4181 = ~w4179 & ~w4180;
assign w4182 = w4178 & w4181;
assign w4183 = w4175 & w4182;
assign w4184 = pi1924 & w1272;
assign w4185 = pi1017 & w1245;
assign w4186 = ~w4184 & ~w4185;
assign w4187 = pi1754 & w1249;
assign w4188 = pi0863 & w1242;
assign w4189 = ~w4187 & ~w4188;
assign w4190 = w4186 & w4189;
assign w4191 = pi1441 & w1280;
assign w4192 = pi1100 & w1266;
assign w4193 = ~w4191 & ~w4192;
assign w4194 = pi1765 & w1263;
assign w4195 = pi1886 & w1278;
assign w4196 = ~w4194 & ~w4195;
assign w4197 = w4193 & w4196;
assign w4198 = w4190 & w4197;
assign w4199 = w4183 & w4198;
assign w4200 = w1221 & w36370;
assign w4201 = pi1833 & w1268;
assign w4202 = pi0951 & w1291;
assign w4203 = ~w4201 & ~w4202;
assign w4204 = pi1430 & w3139;
assign w4205 = pi1900 & w1238;
assign w4206 = ~w4204 & ~w4205;
assign w4207 = w4203 & w4206;
assign w4208 = pi1941 & w3145;
assign w4209 = ~w3180 & ~w4208;
assign w4210 = pi2106 & w1275;
assign w4211 = pi1718 & w1294;
assign w4212 = ~w4210 & ~w4211;
assign w4213 = w4209 & w4212;
assign w4214 = w4207 & w4213;
assign w4215 = ~w4200 & w4214;
assign w4216 = w4199 & w4215;
assign w4217 = (pi1934 & ~w4216) | (pi1934 & w36371) | (~w4216 & w36371);
assign w4218 = pi1053 & pi2405;
assign w4219 = pi0387 & pi1057;
assign w4220 = pi0917 & pi1358;
assign w4221 = ~w4219 & ~w4220;
assign w4222 = ~w4218 & w4221;
assign w4223 = pi3509 & ~w1054;
assign w4224 = pi0591 & pi1359;
assign w4225 = pi1058 & pi3293;
assign w4226 = ~w4224 & ~w4225;
assign w4227 = pi1334 & pi2380;
assign w4228 = pi0868 & pi1344;
assign w4229 = ~w4227 & ~w4228;
assign w4230 = w4226 & w4229;
assign w4231 = ~w4223 & w4230;
assign w4232 = w4222 & w4231;
assign w4233 = (w4232 & w1918) | (w4232 & w36372) | (w1918 & w36372);
assign w4234 = pi0650 & ~w4233;
assign w4235 = pi1341 & pi2296;
assign w4236 = pi1356 & pi2966;
assign w4237 = ~w4235 & ~w4236;
assign w4238 = pi1056 & pi2546;
assign w4239 = pi1054 & pi2712;
assign w4240 = ~w4238 & ~w4239;
assign w4241 = w4237 & w4240;
assign w4242 = pi1355 & pi2455;
assign w4243 = pi1357 & pi2464;
assign w4244 = ~w4242 & ~w4243;
assign w4245 = pi1340 & pi2284;
assign w4246 = pi1349 & pi2732;
assign w4247 = ~w4245 & ~w4246;
assign w4248 = w4244 & w4247;
assign w4249 = pi1354 & pi2963;
assign w4250 = pi1343 & pi2319;
assign w4251 = ~w4249 & ~w4250;
assign w4252 = pi1342 & pi2087;
assign w4253 = pi1055 & pi2722;
assign w4254 = ~w4252 & ~w4253;
assign w4255 = w4251 & w4254;
assign w4256 = w4248 & w4255;
assign w4257 = (pi0539 & ~w4256) | (pi0539 & w36373) | (~w4256 & w36373);
assign w4258 = pi1600 & pi2206;
assign w4259 = pi1350 & pi2259;
assign w4260 = ~w4258 & ~w4259;
assign w4261 = pi1345 & pi2652;
assign w4262 = pi1348 & pi2690;
assign w4263 = ~w4261 & ~w4262;
assign w4264 = w4260 & w4263;
assign w4265 = pi1353 & pi1979;
assign w4266 = pi1351 & pi2264;
assign w4267 = ~w4265 & ~w4266;
assign w4268 = pi1339 & pi2248;
assign w4269 = pi1347 & pi2680;
assign w4270 = ~w4268 & ~w4269;
assign w4271 = w4267 & w4270;
assign w4272 = pi1346 & pi2666;
assign w4273 = pi1338 & pi2234;
assign w4274 = ~w4272 & ~w4273;
assign w4275 = pi1337 & pi2220;
assign w4276 = pi1352 & pi2273;
assign w4277 = ~w4275 & ~w4276;
assign w4278 = w4274 & w4277;
assign w4279 = w4271 & w4278;
assign w4280 = (pi0722 & ~w4279) | (pi0722 & w36374) | (~w4279 & w36374);
assign w4281 = pi1332 & pi2572;
assign w4282 = pi1335 & pi2587;
assign w4283 = ~w4281 & ~w4282;
assign w4284 = pi0330 & pi1333;
assign w4285 = pi0329 & pi1336;
assign w4286 = ~w4284 & ~w4285;
assign w4287 = w4283 & w4286;
assign w4288 = pi0762 & ~w4287;
assign w4289 = ~w4280 & ~w4288;
assign w4290 = ~w4257 & w4289;
assign w4291 = pi0172 & ~pi0979;
assign w4292 = pi0158 & pi0979;
assign w4293 = ~w4291 & ~w4292;
assign w4294 = pi0659 & pi1360;
assign w4295 = (~w4294 & w4293) | (~w4294 & w36375) | (w4293 & w36375);
assign w4296 = pi0979 & pi1960;
assign w4297 = ~pi0979 & pi2425;
assign w4298 = ~w4296 & ~w4297;
assign w4299 = pi0768 & ~w4298;
assign w4300 = pi0979 & pi2148;
assign w4301 = ~pi0979 & pi2920;
assign w4302 = ~w4300 & ~w4301;
assign w4303 = pi0767 & ~w4302;
assign w4304 = ~w4299 & ~w4303;
assign w4305 = pi0979 & pi2166;
assign w4306 = ~pi0979 & pi2933;
assign w4307 = ~w4305 & ~w4306;
assign w4308 = pi0836 & ~w4307;
assign w4309 = pi0979 & pi2182;
assign w4310 = ~pi0979 & pi2943;
assign w4311 = ~w4309 & ~w4310;
assign w4312 = pi0837 & ~w4311;
assign w4313 = ~w4308 & ~w4312;
assign w4314 = w4304 & w4313;
assign w4315 = (pi0576 & ~w4314) | (pi0576 & w36376) | (~w4314 & w36376);
assign w4316 = pi0979 & pi2129;
assign w4317 = ~pi0979 & pi2846;
assign w4318 = ~w4316 & ~w4317;
assign w4319 = pi0717 & ~w4318;
assign w4320 = ~w1179 & ~w4319;
assign w4321 = pi0270 & ~pi0979;
assign w4322 = pi0269 & pi0979;
assign w4323 = ~w4321 & ~w4322;
assign w4324 = pi0716 & ~w4323;
assign w4325 = pi0495 & ~pi0979;
assign w4326 = pi0494 & pi0979;
assign w4327 = ~w4325 & ~w4326;
assign w4328 = pi0718 & ~w4327;
assign w4329 = pi0319 & ~pi0979;
assign w4330 = pi0317 & pi0979;
assign w4331 = ~w4329 & ~w4330;
assign w4332 = pi0761 & ~w4331;
assign w4333 = ~w4328 & ~w4332;
assign w4334 = ~w4324 & w4333;
assign w4335 = w4320 & w4334;
assign w4336 = (pi0538 & ~w4334) | (pi0538 & w36377) | (~w4334 & w36377);
assign w4337 = pi0186 & ~pi0979;
assign w4338 = pi0185 & pi0979;
assign w4339 = ~w4337 & ~w4338;
assign w4340 = pi0720 & ~w4339;
assign w4341 = pi0979 & pi3180;
assign w4342 = ~pi0979 & pi3059;
assign w4343 = ~w4341 & ~w4342;
assign w4344 = pi0766 & ~w4343;
assign w4345 = pi0979 & pi3132;
assign w4346 = ~pi0979 & pi2635;
assign w4347 = ~w4345 & ~w4346;
assign w4348 = pi0765 & ~w4347;
assign w4349 = ~w4344 & ~w4348;
assign w4350 = ~w4340 & w4349;
assign w4351 = pi0979 & pi3154;
assign w4352 = ~pi0979 & pi2782;
assign w4353 = ~w4351 & ~w4352;
assign w4354 = pi0763 & ~w4353;
assign w4355 = pi0345 & ~pi0979;
assign w4356 = pi0344 & pi0979;
assign w4357 = ~w4355 & ~w4356;
assign w4358 = pi0721 & ~w4357;
assign w4359 = ~w4354 & ~w4358;
assign w4360 = pi0979 & pi3201;
assign w4361 = ~pi0979 & pi2873;
assign w4362 = ~w4360 & ~w4361;
assign w4363 = pi0764 & ~w4362;
assign w4364 = pi0065 & ~pi0979;
assign w4365 = pi0063 & pi0979;
assign w4366 = ~w4364 & ~w4365;
assign w4367 = pi0719 & ~w4366;
assign w4368 = ~w4363 & ~w4367;
assign w4369 = w4359 & w4368;
assign w4370 = w4350 & w4369;
assign w4371 = pi0524 & ~w4370;
assign w4372 = ~w4371 & w36378;
assign w4373 = w4290 & w4372;
assign w4374 = (~w941 & w4234) | (~w941 & w36379) | (w4234 & w36379);
assign w4375 = ~w4217 & ~w4374;
assign w4376 = ~w4374 & w36380;
assign w4377 = pi1787 & pi2828;
assign w4378 = w958 & w36381;
assign w4379 = (w4378 & w4376) | (w4378 & w36382) | (w4376 & w36382);
assign w4380 = ~w4160 & ~w4379;
assign w4381 = w2961 & w4380;
assign w4382 = ~w4142 & ~w4381;
assign w4383 = w3936 & w4382;
assign w4384 = (w4383 & ~w3934) | (w4383 & w36383) | (~w3934 & w36383);
assign w4385 = ~w3916 & ~w4384;
assign w4386 = ~w3817 & w4385;
assign w4387 = ~w3439 & w4386;
assign w4388 = ~w674 & w40105;
assign w4389 = w539 & w706;
assign w4390 = ~w713 & ~w4389;
assign w4391 = w4390 & w40106;
assign w4392 = ~w4388 & ~w4391;
assign w4393 = w707 & ~w711;
assign w4394 = ~w674 & ~w4389;
assign w4395 = ~w4393 & ~w4394;
assign w4396 = ~w674 & w4393;
assign w4397 = ~w4395 & ~w4396;
assign w4398 = ~w647 & w36387;
assign w4399 = ~w4392 & ~w4398;
assign w4400 = w797 & w36388;
assign w4401 = ~w550 & ~w2408;
assign w4402 = ~w553 & ~w567;
assign w4403 = ~w4401 & ~w4402;
assign w4404 = w4401 & w4402;
assign w4405 = ~w4403 & ~w4404;
assign w4406 = pi0755 & w552;
assign w4407 = (w797 & w36390) | (w797 & w36391) | (w36390 & w36391);
assign w4408 = ~w4400 & w4407;
assign w4409 = ~w2933 & w36392;
assign w4410 = pi2702 & w1316;
assign w4411 = ~w414 & w36393;
assign w4412 = ~w4410 & ~w4411;
assign w4413 = pi2276 & w1309;
assign w4414 = pi2439 & w1314;
assign w4415 = ~w4413 & ~w4414;
assign w4416 = w4412 & w4415;
assign w4417 = ~w371 & w36394;
assign w4418 = ~w392 & w36395;
assign w4419 = ~w4417 & ~w4418;
assign w4420 = ~w414 & w36396;
assign w4421 = ~w405 & w36397;
assign w4422 = ~w4420 & ~w4421;
assign w4423 = w4419 & w4422;
assign w4424 = (~w354 & ~w4422) | (~w354 & w36398) | (~w4422 & w36398);
assign w4425 = w4416 & ~w4424;
assign w4426 = w2236 & w36399;
assign w4427 = (~w4426 & w4425) | (~w4426 & w36400) | (w4425 & w36400);
assign w4428 = (w2365 & ~w4427) | (w2365 & w36401) | (~w4427 & w36401);
assign w4429 = pi2449 & w941;
assign w4430 = ~w2899 & ~w4429;
assign w4431 = (w353 & w36402) | (w353 & w36403) | (w36402 & w36403);
assign w4432 = w4431 & w40102;
assign w4433 = (pi1030 & w2907) | (pi1030 & w36404) | (w2907 & w36404);
assign w4434 = ~w4433 & w36405;
assign w4435 = ~w4428 & w4434;
assign w4436 = ~pi0861 & w2899;
assign w4437 = w2398 & w36406;
assign w4438 = w2961 & w36407;
assign w4439 = ~w3782 & ~w4438;
assign w4440 = ~w4437 & w4439;
assign w4441 = (~w4440 & ~w4408) | (~w4440 & w36408) | (~w4408 & w36408);
assign w4442 = ~w2425 & ~w2887;
assign w4443 = w2848 & ~w4442;
assign w4444 = (w4443 & w2957) | (w4443 & w36409) | (w2957 & w36409);
assign w4445 = ~w2934 & w4425;
assign w4446 = w2958 & ~w4445;
assign w4447 = w3195 & w3433;
assign w4448 = ~w4446 & ~w4447;
assign w4449 = w2397 & ~w4448;
assign w4450 = (~w4449 & w2845) | (~w4449 & w36410) | (w2845 & w36410);
assign w4451 = ~w4444 & w4450;
assign w4452 = ~w4441 & w4451;
assign w4453 = (w2487 & ~w2462) | (w2487 & w36411) | (~w2462 & w36411);
assign w4454 = ~pi0517 & ~w4453;
assign w4455 = (~pi0679 & w4454) | (~pi0679 & w36412) | (w4454 & w36412);
assign w4456 = w2489 & ~w2490;
assign w4457 = ~w4455 & ~w4456;
assign w4458 = w2826 & ~w4457;
assign w4459 = w2462 & w36413;
assign w4460 = w2630 & w2636;
assign w4461 = ~w2637 & ~w4460;
assign w4462 = ~w4459 & ~w4461;
assign w4463 = ~w2826 & w4462;
assign w4464 = ~w4458 & ~w4463;
assign w4465 = (pi2457 & w2330) | (pi2457 & w36414) | (w2330 & w36414);
assign w4466 = pi2754 & ~w2342;
assign w4467 = ~w4465 & ~w4466;
assign w4468 = (pi2747 & w2346) | (pi2747 & w36415) | (w2346 & w36415);
assign w4469 = (pi2466 & w2336) | (pi2466 & w36416) | (w2336 & w36416);
assign w4470 = ~w4468 & ~w4469;
assign w4471 = w4467 & w4470;
assign w4472 = w4467 & w36417;
assign w4473 = pi2466 & w2876;
assign w4474 = (pi2457 & w2293) | (pi2457 & w36418) | (w2293 & w36418);
assign w4475 = w2295 & w4474;
assign w4476 = w354 & ~w4475;
assign w4477 = pi2747 & w3907;
assign w4478 = pi2754 & w2881;
assign w4479 = ~w4477 & ~w4478;
assign w4480 = w4479 & w36419;
assign w4481 = ~w4472 & ~w4480;
assign w4482 = ~w2425 & ~w4481;
assign w4483 = w2848 & ~w4482;
assign w4484 = (w4483 & w4464) | (w4483 & w36420) | (w4464 & w36420);
assign w4485 = pi0519 & w2570;
assign w4486 = w2554 & w2565;
assign w4487 = ~w4485 & ~w4486;
assign w4488 = ~pi0589 & ~pi0681;
assign w4489 = (~w4488 & ~w2561) | (~w4488 & w36421) | (~w2561 & w36421);
assign w4490 = w4487 & w4489;
assign w4491 = pi0589 & pi0681;
assign w4492 = (w2561 & w36422) | (w2561 & w36421) | (w36422 & w36421);
assign w4493 = ~w4487 & ~w4492;
assign w4494 = ~w4490 & ~w4493;
assign w4495 = w2826 & ~w4494;
assign w4496 = ~w2783 & ~w2787;
assign w4497 = (w4496 & w3444) | (w4496 & w36423) | (w3444 & w36423);
assign w4498 = pi0681 & ~w2561;
assign w4499 = (~w4498 & w3444) | (~w4498 & w36425) | (w3444 & w36425);
assign w4500 = ~w4497 & w4499;
assign w4501 = ~w2826 & ~w4500;
assign w4502 = ~w4495 & ~w4501;
assign w4503 = w3440 & ~w4502;
assign w4504 = (w3782 & w818) | (w3782 & w36426) | (w818 & w36426);
assign w4505 = w1308 & w3433;
assign w4506 = pi3860 & w983;
assign w4507 = w973 & w36427;
assign w4508 = w970 & w36428;
assign w4509 = w973 & w36429;
assign w4510 = ~w4508 & ~w4509;
assign w4511 = ~w4507 & w4510;
assign w4512 = w958 & w36430;
assign w4513 = w963 & w36431;
assign w4514 = w953 & w36432;
assign w4515 = ~w4513 & ~w4514;
assign w4516 = ~w4512 & w4515;
assign w4517 = w970 & w36433;
assign w4518 = w963 & w36434;
assign w4519 = ~w997 & ~w4518;
assign w4520 = ~w4517 & w4519;
assign w4521 = w4516 & w4520;
assign w4522 = w4511 & w4521;
assign w4523 = ~w4506 & w4522;
assign w4524 = w1221 & w36435;
assign w4525 = w1221 & w36436;
assign w4526 = ~w4524 & ~w4525;
assign w4527 = w1216 & w36437;
assign w4528 = w1216 & w36438;
assign w4529 = ~w4527 & ~w4528;
assign w4530 = w4526 & w4529;
assign w4531 = pi1458 & w3148;
assign w4532 = pi0804 & w1234;
assign w4533 = ~w4531 & ~w4532;
assign w4534 = pi1757 & w1249;
assign w4535 = pi0793 & w1245;
assign w4536 = ~w4534 & ~w4535;
assign w4537 = w4533 & w4536;
assign w4538 = pi0699 & w1242;
assign w4539 = pi2052 & w1238;
assign w4540 = ~w4538 & ~w4539;
assign w4541 = pi1444 & w1280;
assign w4542 = pi0908 & w1296;
assign w4543 = ~w4541 & ~w4542;
assign w4544 = w4540 & w4543;
assign w4545 = w4537 & w4544;
assign w4546 = pi1853 & w1268;
assign w4547 = pi1862 & w1278;
assign w4548 = ~w4546 & ~w4547;
assign w4549 = pi0966 & w1288;
assign w4550 = pi1023 & w1266;
assign w4551 = ~w4549 & ~w4550;
assign w4552 = w4548 & w4551;
assign w4553 = pi1721 & w1294;
assign w4554 = pi1944 & w3145;
assign w4555 = ~w4553 & ~w4554;
assign w4556 = pi1767 & w1263;
assign w4557 = pi1735 & w3172;
assign w4558 = ~w4556 & ~w4557;
assign w4559 = w4555 & w4558;
assign w4560 = w4552 & w4559;
assign w4561 = w4545 & w4560;
assign w4562 = w1221 & w36439;
assign w4563 = pi0747 & w1254;
assign w4564 = pi2108 & w1275;
assign w4565 = ~w4563 & ~w4564;
assign w4566 = pi1780 & w1258;
assign w4567 = pi1927 & w1272;
assign w4568 = ~w4566 & ~w4567;
assign w4569 = w4565 & w4568;
assign w4570 = pi1433 & w3139;
assign w4571 = ~w3180 & ~w4570;
assign w4572 = pi0739 & w1251;
assign w4573 = pi0952 & w1291;
assign w4574 = ~w4572 & ~w4573;
assign w4575 = w4571 & w4574;
assign w4576 = w4569 & w4575;
assign w4577 = ~w4562 & w4576;
assign w4578 = w4561 & w4577;
assign w4579 = (pi1934 & ~w4578) | (pi1934 & w36440) | (~w4578 & w36440);
assign w4580 = pi0830 & pi1344;
assign w4581 = pi1334 & pi2766;
assign w4582 = ~w4580 & ~w4581;
assign w4583 = pi0390 & pi1057;
assign w4584 = pi0919 & pi1358;
assign w4585 = ~w4583 & ~w4584;
assign w4586 = w4582 & w4585;
assign w4587 = pi3511 & ~w1054;
assign w4588 = pi1058 & pi3360;
assign w4589 = pi0632 & pi1359;
assign w4590 = ~w4588 & ~w4589;
assign w4591 = pi1059 & pi2980;
assign w4592 = pi1053 & pi2400;
assign w4593 = ~w4591 & ~w4592;
assign w4594 = w4590 & w4593;
assign w4595 = ~w4587 & w4594;
assign w4596 = w4586 & w4595;
assign w4597 = (w4596 & w1693) | (w4596 & w36441) | (w1693 & w36441);
assign w4598 = pi0650 & ~w4597;
assign w4599 = pi1350 & pi2434;
assign w4600 = pi1347 & pi2683;
assign w4601 = ~w4599 & ~w4600;
assign w4602 = pi1339 & pi2251;
assign w4603 = pi1346 & pi2669;
assign w4604 = ~w4602 & ~w4603;
assign w4605 = w4601 & w4604;
assign w4606 = pi1353 & pi1982;
assign w4607 = pi1352 & pi2444;
assign w4608 = ~w4606 & ~w4607;
assign w4609 = pi1600 & pi2209;
assign w4610 = pi1348 & pi2693;
assign w4611 = ~w4609 & ~w4610;
assign w4612 = w4608 & w4611;
assign w4613 = pi1351 & pi2267;
assign w4614 = pi1338 & pi2237;
assign w4615 = ~w4613 & ~w4614;
assign w4616 = pi1337 & pi2223;
assign w4617 = pi1345 & pi2655;
assign w4618 = ~w4616 & ~w4617;
assign w4619 = w4615 & w4618;
assign w4620 = w4612 & w4619;
assign w4621 = (pi0722 & ~w4620) | (pi0722 & w36442) | (~w4620 & w36442);
assign w4622 = pi1340 & pi2068;
assign w4623 = pi1054 & pi2715;
assign w4624 = ~w4622 & ~w4623;
assign w4625 = pi1355 & pi2457;
assign w4626 = pi1349 & pi2734;
assign w4627 = ~w4625 & ~w4626;
assign w4628 = w4624 & w4627;
assign w4629 = pi1056 & pi2743;
assign w4630 = pi1343 & pi2322;
assign w4631 = ~w4629 & ~w4630;
assign w4632 = pi1342 & pi2308;
assign w4633 = pi1354 & pi2747;
assign w4634 = ~w4632 & ~w4633;
assign w4635 = w4631 & w4634;
assign w4636 = pi1356 & pi2754;
assign w4637 = pi1341 & pi2299;
assign w4638 = ~w4636 & ~w4637;
assign w4639 = pi1357 & pi2466;
assign w4640 = pi1055 & pi2773;
assign w4641 = ~w4639 & ~w4640;
assign w4642 = w4638 & w4641;
assign w4643 = w4635 & w4642;
assign w4644 = (pi0539 & ~w4643) | (pi0539 & w36443) | (~w4643 & w36443);
assign w4645 = pi0370 & pi1336;
assign w4646 = pi1335 & pi2590;
assign w4647 = ~w4645 & ~w4646;
assign w4648 = pi0073 & pi1333;
assign w4649 = pi1332 & pi2575;
assign w4650 = ~w4648 & ~w4649;
assign w4651 = w4647 & w4650;
assign w4652 = pi0762 & ~w4651;
assign w4653 = ~w4644 & ~w4652;
assign w4654 = ~w4621 & w4653;
assign w4655 = pi0292 & ~pi0979;
assign w4656 = pi0289 & pi0979;
assign w4657 = ~w4655 & ~w4656;
assign w4658 = pi0761 & ~w4657;
assign w4659 = pi0307 & ~pi0979;
assign w4660 = pi0305 & pi0979;
assign w4661 = ~w4659 & ~w4660;
assign w4662 = pi0716 & ~w4661;
assign w4663 = ~w4658 & ~w4662;
assign w4664 = pi0979 & pi2132;
assign w4665 = ~pi0979 & pi2849;
assign w4666 = ~w4664 & ~w4665;
assign w4667 = pi0717 & ~w4666;
assign w4668 = pi0395 & ~pi0979;
assign w4669 = pi0394 & pi0979;
assign w4670 = ~w4668 & ~w4669;
assign w4671 = pi0718 & ~w4670;
assign w4672 = pi0206 & ~pi0979;
assign w4673 = pi0202 & pi0979;
assign w4674 = ~w4672 & ~w4673;
assign w4675 = pi1599 & ~w4674;
assign w4676 = ~w4671 & ~w4675;
assign w4677 = ~w4667 & w4676;
assign w4678 = (pi0538 & ~w4677) | (pi0538 & w36444) | (~w4677 & w36444);
assign w4679 = pi0979 & pi3157;
assign w4680 = ~pi0979 & pi2781;
assign w4681 = ~w4679 & ~w4680;
assign w4682 = pi0763 & ~w4681;
assign w4683 = pi0584 & ~pi0979;
assign w4684 = pi0583 & pi0979;
assign w4685 = ~w4683 & ~w4684;
assign w4686 = pi0721 & ~w4685;
assign w4687 = pi0047 & ~pi0979;
assign w4688 = pi0046 & pi0979;
assign w4689 = ~w4687 & ~w4688;
assign w4690 = pi0719 & ~w4689;
assign w4691 = ~w4686 & ~w4690;
assign w4692 = ~w4682 & w4691;
assign w4693 = pi0210 & ~pi0979;
assign w4694 = pi0209 & pi0979;
assign w4695 = ~w4693 & ~w4694;
assign w4696 = pi0720 & ~w4695;
assign w4697 = pi0979 & pi3123;
assign w4698 = ~pi0979 & pi2893;
assign w4699 = ~w4697 & ~w4698;
assign w4700 = pi0766 & ~w4699;
assign w4701 = ~w4696 & ~w4700;
assign w4702 = pi0979 & pi3128;
assign w4703 = ~pi0979 & pi2637;
assign w4704 = ~w4702 & ~w4703;
assign w4705 = pi0765 & ~w4704;
assign w4706 = pi0979 & pi3165;
assign w4707 = ~pi0979 & pi2876;
assign w4708 = ~w4706 & ~w4707;
assign w4709 = pi0764 & ~w4708;
assign w4710 = ~w4705 & ~w4709;
assign w4711 = w4701 & w4710;
assign w4712 = w4692 & w4711;
assign w4713 = pi0524 & ~w4712;
assign w4714 = pi0979 & pi1790;
assign w4715 = ~pi0979 & pi2159;
assign w4716 = ~w4714 & ~w4715;
assign w4717 = pi0134 & pi1360;
assign w4718 = (~w4717 & w4716) | (~w4717 & w36445) | (w4716 & w36445);
assign w4719 = pi0176 & ~pi0979;
assign w4720 = pi0161 & pi0979;
assign w4721 = ~w4719 & ~w4720;
assign w4722 = pi0838 & ~w4721;
assign w4723 = pi0979 & pi2169;
assign w4724 = ~pi0979 & pi2935;
assign w4725 = ~w4723 & ~w4724;
assign w4726 = pi0836 & ~w4725;
assign w4727 = ~w4722 & ~w4726;
assign w4728 = pi0979 & pi2185;
assign w4729 = ~pi0979 & pi2783;
assign w4730 = ~w4728 & ~w4729;
assign w4731 = pi0837 & ~w4730;
assign w4732 = pi0979 & pi2151;
assign w4733 = ~pi0979 & pi2923;
assign w4734 = ~w4732 & ~w4733;
assign w4735 = pi0767 & ~w4734;
assign w4736 = ~w4731 & ~w4735;
assign w4737 = w4727 & w4736;
assign w4738 = w4718 & w4737;
assign w4739 = (pi0576 & ~w4737) | (pi0576 & w36446) | (~w4737 & w36446);
assign w4740 = ~w4713 & w36447;
assign w4741 = w4654 & w4740;
assign w4742 = (~w941 & w4598) | (~w941 & w36448) | (w4598 & w36448);
assign w4743 = ~w4579 & ~w4742;
assign w4744 = w940 & w36449;
assign w4745 = ~w4742 & w36450;
assign w4746 = pi1787 & pi2831;
assign w4747 = w958 & w36451;
assign w4748 = (w4747 & w4745) | (w4747 & w36452) | (w4745 & w36452);
assign w4749 = ~w4523 & ~w4748;
assign w4750 = w2961 & w4749;
assign w4751 = (pi2467 & w2336) | (pi2467 & w36453) | (w2336 & w36453);
assign w4752 = pi2755 & ~w2342;
assign w4753 = ~w4751 & ~w4752;
assign w4754 = (pi2525 & w2330) | (pi2525 & w36454) | (w2330 & w36454);
assign w4755 = (pi2533 & w2346) | (pi2533 & w36455) | (w2346 & w36455);
assign w4756 = ~w4754 & ~w4755;
assign w4757 = w4753 & w4756;
assign w4758 = w4753 & w36456;
assign w4759 = pi2467 & w2875;
assign w4760 = w2297 & w4759;
assign w4761 = (pi2533 & w2314) | (pi2533 & w36457) | (w2314 & w36457);
assign w4762 = w2316 & w4761;
assign w4763 = w354 & ~w4762;
assign w4764 = (pi2755 & w2322) | (pi2755 & w36458) | (w2322 & w36458);
assign w4765 = w2324 & w4764;
assign w4766 = (pi2525 & w2293) | (pi2525 & w36459) | (w2293 & w36459);
assign w4767 = w2295 & w4766;
assign w4768 = ~w4765 & ~w4767;
assign w4769 = w4763 & w4768;
assign w4770 = ~w4760 & w4769;
assign w4771 = ~w4758 & ~w4770;
assign w4772 = (~w354 & ~w879) | (~w354 & w36460) | (~w879 & w36460);
assign w4773 = w1319 & ~w4772;
assign w4774 = ~w4771 & w4773;
assign w4775 = w2958 & ~w4774;
assign w4776 = ~w4750 & ~w4775;
assign w4777 = (w2397 & ~w4776) | (w2397 & w36461) | (~w4776 & w36461);
assign w4778 = pi0405 & w2901;
assign w4779 = ~w4770 & w36462;
assign w4780 = (w2365 & w4779) | (w2365 & w36463) | (w4779 & w36463);
assign w4781 = w2417 & ~w4773;
assign w4782 = ~w942 & ~w2899;
assign w4783 = w939 & w40102;
assign w4784 = (pi1036 & w2907) | (pi1036 & w36464) | (w2907 & w36464);
assign w4785 = ~w4784 & w36465;
assign w4786 = ~w4781 & w4785;
assign w4787 = ~w4780 & w4786;
assign w4788 = ~pi0779 & w2899;
assign w4789 = ~w2425 & ~w4788;
assign w4790 = w2398 & w4789;
assign w4791 = ~w4787 & w4790;
assign w4792 = ~w4777 & ~w4791;
assign w4793 = ~w4504 & w4792;
assign w4794 = ~w4503 & w4793;
assign w4795 = ~w4484 & w4794;
assign w4796 = ~w4452 & ~w4795;
assign w4797 = w4387 & w4796;
assign w4798 = ~w474 & w36467;
assign w4799 = ~w720 & ~w4798;
assign w4800 = w4799 & w40107;
assign w4801 = w491 & ~w494;
assign w4802 = (w4801 & w561) | (w4801 & w36468) | (w561 & w36468);
assign w4803 = ~w4800 & ~w4802;
assign w4804 = (w4803 & ~w797) | (w4803 & w36469) | (~w797 & w36469);
assign w4805 = ~w659 & ~w731;
assign w4806 = (w4805 & ~w3826) | (w4805 & w36470) | (~w3826 & w36470);
assign w4807 = ~w718 & w732;
assign w4808 = ~w704 & w4807;
assign w4809 = (~w4798 & w704) | (~w4798 & w36471) | (w704 & w36471);
assign w4810 = ~w4806 & w4809;
assign w4811 = w797 & w36472;
assign w4812 = ~w4804 & ~w4811;
assign w4813 = pi2441 & w1314;
assign w4814 = ~w414 & w36473;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = pi2751 & w1316;
assign w4817 = pi2278 & w1309;
assign w4818 = ~w4816 & ~w4817;
assign w4819 = w4815 & w4818;
assign w4820 = ~w414 & w36474;
assign w4821 = ~w405 & w36475;
assign w4822 = ~w4820 & ~w4821;
assign w4823 = ~w371 & w36476;
assign w4824 = ~w392 & w36477;
assign w4825 = ~w4823 & ~w4824;
assign w4826 = w4822 & w4825;
assign w4827 = (~w354 & ~w4822) | (~w354 & w36478) | (~w4822 & w36478);
assign w4828 = w4819 & ~w4827;
assign w4829 = (pi2460 & w2330) | (pi2460 & w36479) | (w2330 & w36479);
assign w4830 = (pi2469 & w2336) | (pi2469 & w36480) | (w2336 & w36480);
assign w4831 = ~w4829 & ~w4830;
assign w4832 = (pi2750 & w2346) | (pi2750 & w36481) | (w2346 & w36481);
assign w4833 = pi2756 & ~w2342;
assign w4834 = ~w4832 & ~w4833;
assign w4835 = w4831 & w4834;
assign w4836 = w4834 & w36482;
assign w4837 = pi2469 & w2875;
assign w4838 = w2297 & w4837;
assign w4839 = (pi2460 & w2293) | (pi2460 & w36483) | (w2293 & w36483);
assign w4840 = w2295 & w4839;
assign w4841 = w354 & ~w4840;
assign w4842 = pi2750 & w3907;
assign w4843 = pi2756 & w2881;
assign w4844 = ~w4842 & ~w4843;
assign w4845 = w4844 & w36484;
assign w4846 = ~w4836 & ~w4845;
assign w4847 = w4828 & ~w4846;
assign w4848 = w2958 & ~w4847;
assign w4849 = pi3869 & w983;
assign w4850 = w973 & w36485;
assign w4851 = w973 & w36486;
assign w4852 = w970 & w36487;
assign w4853 = ~w4851 & ~w4852;
assign w4854 = ~w4850 & w4853;
assign w4855 = w958 & w36488;
assign w4856 = w963 & w36489;
assign w4857 = w953 & w36490;
assign w4858 = ~w4856 & ~w4857;
assign w4859 = ~w4855 & w4858;
assign w4860 = w970 & w36491;
assign w4861 = w963 & w36492;
assign w4862 = ~w997 & ~w4861;
assign w4863 = ~w4860 & w4862;
assign w4864 = w4859 & w4863;
assign w4865 = w4854 & w4864;
assign w4866 = ~w4849 & w4865;
assign w4867 = w940 & w36493;
assign w4868 = pi3504 & ~w1054;
assign w4869 = pi0392 & pi1057;
assign w4870 = pi0594 & pi1359;
assign w4871 = ~w4869 & ~w4870;
assign w4872 = ~w4868 & w4871;
assign w4873 = (w4872 & w1845) | (w4872 & w36494) | (w1845 & w36494);
assign w4874 = pi0650 & ~w4873;
assign w4875 = pi1355 & pi2460;
assign w4876 = pi1356 & pi2756;
assign w4877 = ~w4875 & ~w4876;
assign w4878 = pi1343 & pi2326;
assign w4879 = pi1357 & pi2469;
assign w4880 = ~w4878 & ~w4879;
assign w4881 = w4877 & w4880;
assign w4882 = pi1341 & pi2301;
assign w4883 = pi1349 & pi2737;
assign w4884 = ~w4882 & ~w4883;
assign w4885 = pi1054 & pi2718;
assign w4886 = pi1056 & pi2745;
assign w4887 = ~w4885 & ~w4886;
assign w4888 = w4884 & w4887;
assign w4889 = pi1055 & pi2726;
assign w4890 = pi1340 & pi2290;
assign w4891 = ~w4889 & ~w4890;
assign w4892 = pi1342 & pi2312;
assign w4893 = pi1354 & pi2750;
assign w4894 = ~w4892 & ~w4893;
assign w4895 = w4891 & w4894;
assign w4896 = w4888 & w4895;
assign w4897 = (pi0539 & ~w4896) | (pi0539 & w36495) | (~w4896 & w36495);
assign w4898 = pi1348 & pi2697;
assign w4899 = pi1351 & pi2441;
assign w4900 = ~w4898 & ~w4899;
assign w4901 = pi1346 & pi2673;
assign w4902 = pi1600 & pi2213;
assign w4903 = ~w4901 & ~w4902;
assign w4904 = w4900 & w4903;
assign w4905 = pi1339 & pi2255;
assign w4906 = pi1337 & pi2227;
assign w4907 = ~w4905 & ~w4906;
assign w4908 = pi1352 & pi2751;
assign w4909 = pi1347 & pi2686;
assign w4910 = ~w4908 & ~w4909;
assign w4911 = w4907 & w4910;
assign w4912 = pi1345 & pi2659;
assign w4913 = pi1338 & pi2241;
assign w4914 = ~w4912 & ~w4913;
assign w4915 = pi1353 & pi2278;
assign w4916 = pi1350 & pi2700;
assign w4917 = ~w4915 & ~w4916;
assign w4918 = w4914 & w4917;
assign w4919 = w4911 & w4918;
assign w4920 = (pi0722 & ~w4919) | (pi0722 & w36496) | (~w4919 & w36496);
assign w4921 = pi0225 & pi1336;
assign w4922 = pi1333 & pi1745;
assign w4923 = ~w4921 & ~w4922;
assign w4924 = pi1332 & pi2581;
assign w4925 = pi1335 & pi2596;
assign w4926 = ~w4924 & ~w4925;
assign w4927 = w4923 & w4926;
assign w4928 = pi0762 & ~w4927;
assign w4929 = ~w4920 & ~w4928;
assign w4930 = ~w4897 & w4929;
assign w4931 = pi0284 & ~pi0979;
assign w4932 = pi0282 & pi0979;
assign w4933 = ~w4931 & ~w4932;
assign w4934 = pi0761 & ~w4933;
assign w4935 = pi0979 & pi2138;
assign w4936 = ~pi0979 & pi2855;
assign w4937 = ~w4935 & ~w4936;
assign w4938 = pi0717 & ~w4937;
assign w4939 = pi0227 & ~pi0979;
assign w4940 = pi0226 & pi0979;
assign w4941 = ~w4939 & ~w4940;
assign w4942 = pi0716 & ~w4941;
assign w4943 = ~w4938 & ~w4942;
assign w4944 = ~w4934 & w4943;
assign w4945 = w1184 & w4944;
assign w4946 = (pi0538 & ~w4944) | (pi0538 & w35782) | (~w4944 & w35782);
assign w4947 = pi0979 & pi1967;
assign w4948 = ~pi0979 & pi2431;
assign w4949 = ~w4947 & ~w4948;
assign w4950 = pi0768 & ~w4949;
assign w4951 = pi0979 & pi2175;
assign w4952 = ~pi0979 & pi2937;
assign w4953 = ~w4951 & ~w4952;
assign w4954 = pi0836 & ~w4953;
assign w4955 = ~w4950 & ~w4954;
assign w4956 = pi0979 & pi2157;
assign w4957 = ~pi0979 & pi2928;
assign w4958 = ~w4956 & ~w4957;
assign w4959 = pi0767 & ~w4958;
assign w4960 = pi0181 & ~pi0979;
assign w4961 = pi0166 & pi0979;
assign w4962 = ~w4960 & ~w4961;
assign w4963 = pi0838 & ~w4962;
assign w4964 = pi0979 & pi2191;
assign w4965 = ~pi0979 & pi3113;
assign w4966 = ~w4964 & ~w4965;
assign w4967 = pi0837 & ~w4966;
assign w4968 = ~w4963 & ~w4967;
assign w4969 = ~w4959 & w4968;
assign w4970 = (pi0576 & ~w4969) | (pi0576 & w36497) | (~w4969 & w36497);
assign w4971 = pi0258 & ~pi0979;
assign w4972 = pi0256 & pi0979;
assign w4973 = ~w4971 & ~w4972;
assign w4974 = pi0721 & ~w4973;
assign w4975 = pi0069 & ~pi0979;
assign w4976 = pi0068 & pi0979;
assign w4977 = ~w4975 & ~w4976;
assign w4978 = pi0720 & ~w4977;
assign w4979 = pi0979 & pi3176;
assign w4980 = ~pi0979 & pi2642;
assign w4981 = ~w4979 & ~w4980;
assign w4982 = pi0765 & ~w4981;
assign w4983 = ~w4978 & ~w4982;
assign w4984 = ~w4974 & w4983;
assign w4985 = pi0979 & pi2610;
assign w4986 = ~pi0979 & pi2617;
assign w4987 = ~w4985 & ~w4986;
assign w4988 = pi0763 & ~w4987;
assign w4989 = ~w1144 & ~w4988;
assign w4990 = pi0979 & pi2623;
assign w4991 = ~pi0979 & pi2629;
assign w4992 = ~w4990 & ~w4991;
assign w4993 = pi0764 & ~w4992;
assign w4994 = pi0979 & pi3185;
assign w4995 = ~pi0979 & pi2840;
assign w4996 = ~w4994 & ~w4995;
assign w4997 = pi0766 & ~w4996;
assign w4998 = ~w4993 & ~w4997;
assign w4999 = w4989 & w4998;
assign w5000 = w4984 & w4999;
assign w5001 = pi0524 & ~w5000;
assign w5002 = ~w5001 & w36498;
assign w5003 = w4930 & w5002;
assign w5004 = ~w4874 & w5003;
assign w5005 = ~w941 & ~w5004;
assign w5006 = w1221 & w36499;
assign w5007 = w1216 & w36500;
assign w5008 = ~w5006 & ~w5007;
assign w5009 = w1221 & w36501;
assign w5010 = w1216 & w36502;
assign w5011 = ~w5009 & ~w5010;
assign w5012 = w5008 & w5011;
assign w5013 = pi0367 & w1242;
assign w5014 = pi0871 & w1254;
assign w5015 = pi1891 & w1278;
assign w5016 = ~w5014 & ~w5015;
assign w5017 = ~w5013 & w5016;
assign w5018 = pi0978 & w1234;
assign w5019 = pi1785 & w1258;
assign w5020 = ~w5018 & ~w5019;
assign w5021 = pi1932 & w1272;
assign w5022 = pi1460 & w3148;
assign w5023 = ~w5021 & ~w5022;
assign w5024 = w5020 & w5023;
assign w5025 = pi1725 & w1294;
assign w5026 = pi2051 & w1238;
assign w5027 = ~w5025 & ~w5026;
assign w5028 = pi0794 & w1245;
assign w5029 = pi1737 & w3172;
assign w5030 = ~w5028 & ~w5029;
assign w5031 = w5027 & w5030;
assign w5032 = w5024 & w5031;
assign w5033 = w5017 & w5032;
assign w5034 = w1221 & w36503;
assign w5035 = pi0740 & w1251;
assign w5036 = pi0910 & w1296;
assign w5037 = ~w5035 & ~w5036;
assign w5038 = pi1705 & w1268;
assign w5039 = pi1446 & w1280;
assign w5040 = ~w5038 & ~w5039;
assign w5041 = w5037 & w5040;
assign w5042 = w1291 & w36504;
assign w5043 = w1288 & w36505;
assign w5044 = ~w5042 & ~w5043;
assign w5045 = w5041 & w36506;
assign w5046 = w5033 & w36507;
assign w5047 = pi1934 & ~w5046;
assign w5048 = ~w5005 & ~w5047;
assign w5049 = ~w5005 & w36508;
assign w5050 = pi1787 & pi2835;
assign w5051 = w958 & w36509;
assign w5052 = (w5051 & w5049) | (w5051 & w36510) | (w5049 & w36510);
assign w5053 = ~w4866 & ~w5052;
assign w5054 = w3433 & w5053;
assign w5055 = ~w4848 & ~w5054;
assign w5056 = w2397 & ~w5055;
assign w5057 = (w2425 & w5055) | (w2425 & w36511) | (w5055 & w36511);
assign w5058 = ~pi0781 & w2899;
assign w5059 = w2417 & ~w4828;
assign w5060 = ~w4845 & w36512;
assign w5061 = w940 & w36513;
assign w5062 = w2236 & w36514;
assign w5063 = (~w5061 & ~w359) | (~w5061 & w36516) | (~w359 & w36516);
assign w5064 = ~w2899 & w5063;
assign w5065 = (w353 & w36517) | (w353 & w36518) | (w36517 & w36518);
assign w5066 = w5065 & w40102;
assign w5067 = (pi1038 & w2907) | (pi1038 & w36519) | (w2907 & w36519);
assign w5068 = ~w5066 & ~w5067;
assign w5069 = w5064 & w5068;
assign w5070 = ~w5060 & w5069;
assign w5071 = ~w5059 & w5070;
assign w5072 = ~w5058 & ~w5071;
assign w5073 = ~w2425 & ~w5072;
assign w5074 = w2398 & ~w5073;
assign w5075 = pi3862 & w983;
assign w5076 = w973 & w36520;
assign w5077 = w973 & w36521;
assign w5078 = w970 & w36522;
assign w5079 = ~w5077 & ~w5078;
assign w5080 = ~w5076 & w5079;
assign w5081 = w958 & w36523;
assign w5082 = w963 & w36524;
assign w5083 = w953 & w36525;
assign w5084 = ~w5082 & ~w5083;
assign w5085 = ~w5081 & w5084;
assign w5086 = w970 & w36526;
assign w5087 = w963 & w36527;
assign w5088 = ~w997 & ~w5087;
assign w5089 = ~w5086 & w5088;
assign w5090 = w5085 & w5089;
assign w5091 = w5080 & w5090;
assign w5092 = ~w5075 & w5091;
assign w5093 = w940 & w36528;
assign w5094 = (pi1331 & ~w2024) | (pi1331 & w36529) | (~w2024 & w36529);
assign w5095 = pi0388 & pi1057;
assign w5096 = pi0603 & pi1359;
assign w5097 = ~w5095 & ~w5096;
assign w5098 = pi0828 & pi1344;
assign w5099 = pi0708 & pi1358;
assign w5100 = ~w5098 & ~w5099;
assign w5101 = w5097 & w5100;
assign w5102 = pi3521 & ~w1054;
assign w5103 = pi1334 & pi3204;
assign w5104 = pi1053 & pi2472;
assign w5105 = ~w5103 & ~w5104;
assign w5106 = pi1059 & pi2978;
assign w5107 = pi1058 & pi3407;
assign w5108 = ~w5106 & ~w5107;
assign w5109 = w5105 & w5108;
assign w5110 = ~w5102 & w5109;
assign w5111 = w5101 & w5110;
assign w5112 = (pi0650 & w5094) | (pi0650 & w36530) | (w5094 & w36530);
assign w5113 = pi0979 & pi3131;
assign w5114 = ~pi0979 & pi2541;
assign w5115 = ~w5113 & ~w5114;
assign w5116 = pi0765 & ~w5115;
assign w5117 = pi0041 & ~pi0979;
assign w5118 = pi0039 & pi0979;
assign w5119 = ~w5117 & ~w5118;
assign w5120 = pi0719 & ~w5119;
assign w5121 = pi0218 & ~pi0979;
assign w5122 = pi0215 & pi0979;
assign w5123 = ~w5121 & ~w5122;
assign w5124 = pi0720 & ~w5123;
assign w5125 = ~w5120 & ~w5124;
assign w5126 = ~w5116 & w5125;
assign w5127 = pi0397 & ~pi0979;
assign w5128 = pi0396 & pi0979;
assign w5129 = ~w5127 & ~w5128;
assign w5130 = pi0721 & ~w5129;
assign w5131 = pi0979 & pi3181;
assign w5132 = ~pi0979 & pi2891;
assign w5133 = ~w5131 & ~w5132;
assign w5134 = pi0766 & ~w5133;
assign w5135 = ~w5130 & ~w5134;
assign w5136 = pi0979 & pi3155;
assign w5137 = ~pi0979 & pi2865;
assign w5138 = ~w5136 & ~w5137;
assign w5139 = pi0763 & ~w5138;
assign w5140 = pi0979 & pi3163;
assign w5141 = ~pi0979 & pi2874;
assign w5142 = ~w5140 & ~w5141;
assign w5143 = pi0764 & ~w5142;
assign w5144 = ~w5139 & ~w5143;
assign w5145 = w5135 & w5144;
assign w5146 = w5126 & w5145;
assign w5147 = pi0524 & ~w5146;
assign w5148 = pi1338 & pi2235;
assign w5149 = pi1352 & pi2443;
assign w5150 = ~w5148 & ~w5149;
assign w5151 = pi1353 & pi1980;
assign w5152 = pi1337 & pi2221;
assign w5153 = ~w5151 & ~w5152;
assign w5154 = w5150 & w5153;
assign w5155 = pi1347 & pi2681;
assign w5156 = pi1345 & pi2653;
assign w5157 = ~w5155 & ~w5156;
assign w5158 = pi1600 & pi2207;
assign w5159 = pi1346 & pi2667;
assign w5160 = ~w5158 & ~w5159;
assign w5161 = w5157 & w5160;
assign w5162 = pi1348 & pi2691;
assign w5163 = pi1339 & pi2249;
assign w5164 = ~w5162 & ~w5163;
assign w5165 = pi1350 & pi2260;
assign w5166 = pi1351 & pi2265;
assign w5167 = ~w5165 & ~w5166;
assign w5168 = w5164 & w5167;
assign w5169 = w5161 & w5168;
assign w5170 = (pi0722 & ~w5169) | (pi0722 & w36531) | (~w5169 & w36531);
assign w5171 = ~w5147 & ~w5170;
assign w5172 = pi0196 & pi1360;
assign w5173 = pi0979 & pi2183;
assign w5174 = ~pi0979 & pi2944;
assign w5175 = ~w5173 & ~w5174;
assign w5176 = (~w5172 & w5175) | (~w5172 & w36532) | (w5175 & w36532);
assign w5177 = pi0173 & ~pi0979;
assign w5178 = pi0159 & pi0979;
assign w5179 = ~w5177 & ~w5178;
assign w5180 = pi0838 & ~w5179;
assign w5181 = pi0979 & pi1961;
assign w5182 = ~pi0979 & pi2426;
assign w5183 = ~w5181 & ~w5182;
assign w5184 = pi0768 & ~w5183;
assign w5185 = ~w5180 & ~w5184;
assign w5186 = pi0979 & pi2167;
assign w5187 = ~pi0979 & pi2793;
assign w5188 = ~w5186 & ~w5187;
assign w5189 = pi0836 & ~w5188;
assign w5190 = pi0979 & pi2149;
assign w5191 = ~pi0979 & pi2921;
assign w5192 = ~w5190 & ~w5191;
assign w5193 = pi0767 & ~w5192;
assign w5194 = ~w5189 & ~w5193;
assign w5195 = w5185 & w5194;
assign w5196 = w5176 & w5195;
assign w5197 = (pi0576 & ~w5195) | (pi0576 & w36533) | (~w5195 & w36533);
assign w5198 = pi0324 & ~pi0979;
assign w5199 = pi0323 & pi0979;
assign w5200 = ~w5198 & ~w5199;
assign w5201 = pi0761 & ~w5200;
assign w5202 = pi0306 & ~pi0979;
assign w5203 = pi0304 & pi0979;
assign w5204 = ~w5202 & ~w5203;
assign w5205 = pi0716 & ~w5204;
assign w5206 = ~w5201 & ~w5205;
assign w5207 = pi0481 & ~pi0979;
assign w5208 = pi0480 & pi0979;
assign w5209 = ~w5207 & ~w5208;
assign w5210 = pi0718 & ~w5209;
assign w5211 = pi0979 & pi2130;
assign w5212 = ~pi0979 & pi2847;
assign w5213 = ~w5211 & ~w5212;
assign w5214 = pi0717 & ~w5213;
assign w5215 = pi0204 & ~pi0979;
assign w5216 = pi0200 & pi0979;
assign w5217 = ~w5215 & ~w5216;
assign w5218 = pi1599 & ~w5217;
assign w5219 = ~w5214 & ~w5218;
assign w5220 = ~w5210 & w5219;
assign w5221 = (pi0538 & ~w5220) | (pi0538 & w36534) | (~w5220 & w36534);
assign w5222 = ~w5197 & ~w5221;
assign w5223 = w5171 & w5222;
assign w5224 = ~w5112 & w5223;
assign w5225 = ~w941 & ~w5224;
assign w5226 = w1221 & w36535;
assign w5227 = w1216 & w36536;
assign w5228 = ~w5226 & ~w5227;
assign w5229 = w1221 & w36537;
assign w5230 = w1216 & w36538;
assign w5231 = ~w5229 & ~w5230;
assign w5232 = w5228 & w5231;
assign w5233 = pi1456 & w3148;
assign w5234 = pi2107 & w1275;
assign w5235 = ~w5233 & ~w5234;
assign w5236 = pi1022 & w1266;
assign w5237 = pi1431 & w3139;
assign w5238 = ~w5236 & ~w5237;
assign w5239 = w5235 & w5238;
assign w5240 = pi0797 & w1288;
assign w5241 = pi1442 & w1280;
assign w5242 = ~w5240 & ~w5241;
assign w5243 = pi1733 & w3172;
assign w5244 = pi0874 & w1296;
assign w5245 = ~w5243 & ~w5244;
assign w5246 = w5242 & w5245;
assign w5247 = w5239 & w5246;
assign w5248 = pi1719 & w1294;
assign w5249 = pi1901 & w1238;
assign w5250 = ~w5248 & ~w5249;
assign w5251 = pi1942 & w3145;
assign w5252 = pi1852 & w1268;
assign w5253 = ~w5251 & ~w5252;
assign w5254 = w5250 & w5253;
assign w5255 = pi1858 & w1263;
assign w5256 = pi0884 & w1251;
assign w5257 = ~w5255 & ~w5256;
assign w5258 = pi1887 & w1278;
assign w5259 = pi1755 & w1249;
assign w5260 = ~w5258 & ~w5259;
assign w5261 = w5257 & w5260;
assign w5262 = w5254 & w5261;
assign w5263 = w5247 & w5262;
assign w5264 = w1221 & w36539;
assign w5265 = pi0803 & w1234;
assign w5266 = pi0822 & w1242;
assign w5267 = ~w5265 & ~w5266;
assign w5268 = pi1925 & w1272;
assign w5269 = pi0957 & w1245;
assign w5270 = ~w5268 & ~w5269;
assign w5271 = w5267 & w5270;
assign w5272 = pi0746 & w1254;
assign w5273 = ~w3180 & ~w5272;
assign w5274 = pi1778 & w1258;
assign w5275 = pi0891 & w1291;
assign w5276 = ~w5274 & ~w5275;
assign w5277 = w5273 & w5276;
assign w5278 = w5271 & w5277;
assign w5279 = ~w5264 & w5278;
assign w5280 = w5263 & w5279;
assign w5281 = pi1332 & pi2573;
assign w5282 = pi1335 & pi2588;
assign w5283 = ~w5281 & ~w5282;
assign w5284 = pi0072 & pi1333;
assign w5285 = pi0331 & pi1336;
assign w5286 = ~w5284 & ~w5285;
assign w5287 = w5283 & w5286;
assign w5288 = w1607 & ~w5287;
assign w5289 = (pi0539 & ~w940) | (pi0539 & w36541) | (~w940 & w36541);
assign w5290 = pi1342 & pi2306;
assign w5291 = pi1356 & pi2810;
assign w5292 = ~w5290 & ~w5291;
assign w5293 = pi1341 & pi2297;
assign w5294 = pi1056 & pi2742;
assign w5295 = ~w5293 & ~w5294;
assign w5296 = w5292 & w5295;
assign w5297 = pi1355 & pi2456;
assign w5298 = pi1354 & pi2780;
assign w5299 = ~w5297 & ~w5298;
assign w5300 = pi1055 & pi2723;
assign w5301 = pi1054 & pi2713;
assign w5302 = ~w5300 & ~w5301;
assign w5303 = w5299 & w5302;
assign w5304 = pi1349 & pi2733;
assign w5305 = pi1340 & pi2285;
assign w5306 = ~w5304 & ~w5305;
assign w5307 = pi1343 & pi2320;
assign w5308 = pi1357 & pi2465;
assign w5309 = ~w5307 & ~w5308;
assign w5310 = w5306 & w5309;
assign w5311 = w5303 & w5310;
assign w5312 = (w5289 & ~w5311) | (w5289 & w36542) | (~w5311 & w36542);
assign w5313 = ~w5288 & ~w5312;
assign w5314 = (w5280 & w36543) | (w5280 & w36544) | (w36543 & w36544);
assign w5315 = ~w5225 & w5314;
assign w5316 = ~w5225 & w36545;
assign w5317 = pi1787 & pi2829;
assign w5318 = w958 & w36546;
assign w5319 = (w5318 & w5316) | (w5318 & w36547) | (w5316 & w36547);
assign w5320 = ~w5092 & ~w5319;
assign w5321 = w2961 & w36548;
assign w5322 = ~w5074 & ~w5321;
assign w5323 = ~w5056 & w5322;
assign w5324 = (~w5323 & ~w4812) | (~w5323 & w36549) | (~w4812 & w36549);
assign w5325 = ~w2493 & w36550;
assign w5326 = (pi0588 & w2493) | (pi0588 & w36551) | (w2493 & w36551);
assign w5327 = ~w5325 & ~w5326;
assign w5328 = ~pi0705 & w5327;
assign w5329 = pi0705 & w2495;
assign w5330 = (~w5329 & w5327) | (~w5329 & w36552) | (w5327 & w36552);
assign w5331 = ~w5328 & w5330;
assign w5332 = (~w5331 & w2810) | (~w5331 & w36553) | (w2810 & w36553);
assign w5333 = (w5332 & ~w2573) | (w5332 & w36554) | (~w2573 & w36554);
assign w5334 = ~w2607 & ~w2640;
assign w5335 = ~w2641 & ~w5334;
assign w5336 = ~w5329 & ~w5335;
assign w5337 = (w2578 & w5335) | (w2578 & w36555) | (w5335 & w36555);
assign w5338 = w2573 & w5337;
assign w5339 = w2818 & ~w5336;
assign w5340 = ~w5338 & ~w5339;
assign w5341 = ~w5333 & w5340;
assign w5342 = w5340 & w36556;
assign w5343 = (pi2456 & w2330) | (pi2456 & w36557) | (w2330 & w36557);
assign w5344 = (pi2780 & w2346) | (pi2780 & w36558) | (w2346 & w36558);
assign w5345 = ~w5343 & ~w5344;
assign w5346 = (pi2465 & w2336) | (pi2465 & w36559) | (w2336 & w36559);
assign w5347 = pi2810 & ~w2342;
assign w5348 = ~w5346 & ~w5347;
assign w5349 = w5345 & w5348;
assign w5350 = w5348 & w36560;
assign w5351 = pi2465 & w2875;
assign w5352 = w2297 & w5351;
assign w5353 = (pi2456 & w2293) | (pi2456 & w36561) | (w2293 & w36561);
assign w5354 = w2295 & w5353;
assign w5355 = w354 & ~w5354;
assign w5356 = pi2810 & w2881;
assign w5357 = pi2780 & w3907;
assign w5358 = ~w5356 & ~w5357;
assign w5359 = w5358 & w36562;
assign w5360 = ~w5350 & ~w5359;
assign w5361 = ~w2425 & ~w5360;
assign w5362 = w2848 & ~w5361;
assign w5363 = ~w5342 & w5362;
assign w5364 = (pi0683 & w2532) | (pi0683 & w36563) | (w2532 & w36563);
assign w5365 = w2791 & w2793;
assign w5366 = (w5365 & w2711) | (w5365 & w36564) | (w2711 & w36564);
assign w5367 = (w2791 & w2711) | (w2791 & w36565) | (w2711 & w36565);
assign w5368 = ~w2793 & ~w5367;
assign w5369 = (~w5364 & w5368) | (~w5364 & w36566) | (w5368 & w36566);
assign w5370 = ~w2826 & w5369;
assign w5371 = ~w2530 & w2541;
assign w5372 = ~w2568 & w5371;
assign w5373 = ~pi0683 & ~w5372;
assign w5374 = w2534 & w5372;
assign w5375 = ~w5373 & ~w5374;
assign w5376 = w2826 & ~w5375;
assign w5377 = ~w5370 & ~w5376;
assign w5378 = w3440 & w5377;
assign w5379 = ~w5378 & w36567;
assign w5380 = ~w5366 & w36568;
assign w5381 = ~pi0682 & ~w2752;
assign w5382 = (~w5381 & ~w2565) | (~w5381 & w36570) | (~w2565 & w36570);
assign w5383 = w5382 & w40108;
assign w5384 = ~w5380 & w5383;
assign w5385 = pi0682 & w2752;
assign w5386 = (~w5385 & w2565) | (~w5385 & w36571) | (w2565 & w36571);
assign w5387 = w2761 & ~w5386;
assign w5388 = ~w5366 & w36572;
assign w5389 = ~w2761 & ~w5386;
assign w5390 = (w5389 & w5366) | (w5389 & w36573) | (w5366 & w36573);
assign w5391 = ~w5388 & ~w5390;
assign w5392 = ~w2826 & w36574;
assign w5393 = ~w4485 & w36575;
assign w5394 = (pi0682 & w4485) | (pi0682 & w36576) | (w4485 & w36576);
assign w5395 = ~w5393 & ~w5394;
assign w5396 = w2826 & w5395;
assign w5397 = ~w5392 & ~w5396;
assign w5398 = w3440 & w5397;
assign w5399 = w491 & ~w493;
assign w5400 = (w5399 & w561) | (w5399 & w36577) | (w561 & w36577);
assign w5401 = ~w493 & w495;
assign w5402 = ~w475 & w36578;
assign w5403 = ~w5401 & ~w5402;
assign w5404 = ~w497 & w5403;
assign w5405 = (w5404 & w561) | (w5404 & w36579) | (w561 & w36579);
assign w5406 = ~w5400 & w5405;
assign w5407 = (w5406 & ~w797) | (w5406 & w36580) | (~w797 & w36580);
assign w5408 = (~w729 & w704) | (~w729 & w36581) | (w704 & w36581);
assign w5409 = w782 & ~w5402;
assign w5410 = ~w5408 & w5409;
assign w5411 = ~w782 & w36582;
assign w5412 = ~w4808 & w5411;
assign w5413 = ~w5410 & ~w5412;
assign w5414 = w798 & ~w5413;
assign w5415 = ~w5407 & ~w5414;
assign w5416 = ~w5414 & w36583;
assign w5417 = ~pi0516 & w2492;
assign w5418 = pi0516 & ~w2492;
assign w5419 = ~w5417 & ~w5418;
assign w5420 = pi0706 & ~w5419;
assign w5421 = ~w2485 & w5419;
assign w5422 = ~w5420 & ~w5421;
assign w5423 = w2826 & ~w5422;
assign w5424 = w2826 & w36584;
assign w5425 = ~w2623 & ~w2624;
assign w5426 = w2638 & w5425;
assign w5427 = (pi0706 & w2482) | (pi0706 & w36585) | (w2482 & w36585);
assign w5428 = (~w5427 & w5425) | (~w5427 & w36586) | (w5425 & w36586);
assign w5429 = ~w5426 & w5428;
assign w5430 = w3433 & w36587;
assign w5431 = pi3870 & w983;
assign w5432 = w973 & w36588;
assign w5433 = w970 & w36589;
assign w5434 = w973 & w36590;
assign w5435 = ~w5433 & ~w5434;
assign w5436 = ~w5432 & w5435;
assign w5437 = w958 & w36591;
assign w5438 = w963 & w36592;
assign w5439 = w953 & w36593;
assign w5440 = ~w5438 & ~w5439;
assign w5441 = ~w5437 & w5440;
assign w5442 = w970 & w36594;
assign w5443 = w963 & w36595;
assign w5444 = ~w997 & ~w5443;
assign w5445 = ~w5442 & w5444;
assign w5446 = w5441 & w5445;
assign w5447 = w5436 & w5446;
assign w5448 = ~w5431 & w5447;
assign w5449 = w1221 & w36596;
assign w5450 = w1216 & w36597;
assign w5451 = ~w5449 & ~w5450;
assign w5452 = w1221 & w36598;
assign w5453 = w1216 & w36599;
assign w5454 = ~w5452 & ~w5453;
assign w5455 = w5451 & w5454;
assign w5456 = pi1459 & w3148;
assign w5457 = pi1838 & w1268;
assign w5458 = ~w5456 & ~w5457;
assign w5459 = pi1931 & w1272;
assign w5460 = pi0971 & w1234;
assign w5461 = ~w5459 & ~w5460;
assign w5462 = w5458 & w5461;
assign w5463 = pi0336 & w1242;
assign w5464 = pi0791 & w1251;
assign w5465 = ~w5463 & ~w5464;
assign w5466 = pi1736 & w3172;
assign w5467 = pi1892 & w1278;
assign w5468 = ~w5466 & ~w5467;
assign w5469 = w5465 & w5468;
assign w5470 = pi0872 & w1254;
assign w5471 = pi1784 & w1258;
assign w5472 = ~w5470 & ~w5471;
assign w5473 = pi1724 & w1294;
assign w5474 = pi1445 & w1280;
assign w5475 = ~w5473 & ~w5474;
assign w5476 = w5472 & w5475;
assign w5477 = w5469 & w5476;
assign w5478 = w5462 & w5477;
assign w5479 = w1221 & w36600;
assign w5480 = pi1906 & w1238;
assign w5481 = ~w3180 & ~w5480;
assign w5482 = pi0820 & w1296;
assign w5483 = pi0899 & w1245;
assign w5484 = ~w5482 & ~w5483;
assign w5485 = w5481 & w5484;
assign w5486 = w1288 & w36601;
assign w5487 = w1291 & w36602;
assign w5488 = ~w5486 & ~w5487;
assign w5489 = w5485 & w36603;
assign w5490 = w5478 & w36604;
assign w5491 = pi1934 & ~w5490;
assign w5492 = pi3513 & ~w1054;
assign w5493 = pi0391 & pi1057;
assign w5494 = pi0595 & pi1359;
assign w5495 = ~w5493 & ~w5494;
assign w5496 = ~w5492 & w5495;
assign w5497 = (w5496 & w1879) | (w5496 & w36605) | (w1879 & w36605);
assign w5498 = pi0650 & ~w5497;
assign w5499 = pi1600 & pi2212;
assign w5500 = pi1350 & pi2539;
assign w5501 = ~w5499 & ~w5500;
assign w5502 = pi1338 & pi2240;
assign w5503 = pi1346 & pi2672;
assign w5504 = ~w5502 & ~w5503;
assign w5505 = w5501 & w5504;
assign w5506 = pi1337 & pi2226;
assign w5507 = pi1348 & pi2696;
assign w5508 = ~w5506 & ~w5507;
assign w5509 = pi1351 & pi2440;
assign w5510 = pi1347 & pi2615;
assign w5511 = ~w5509 & ~w5510;
assign w5512 = w5508 & w5511;
assign w5513 = pi1353 & pi2277;
assign w5514 = pi1345 & pi2658;
assign w5515 = ~w5513 & ~w5514;
assign w5516 = pi1339 & pi2254;
assign w5517 = pi1352 & pi2703;
assign w5518 = ~w5516 & ~w5517;
assign w5519 = w5515 & w5518;
assign w5520 = w5512 & w5519;
assign w5521 = (pi0722 & ~w5520) | (pi0722 & w36606) | (~w5520 & w36606);
assign w5522 = pi1356 & pi2544;
assign w5523 = pi1056 & pi2545;
assign w5524 = ~w5522 & ~w5523;
assign w5525 = pi1054 & pi2534;
assign w5526 = pi1055 & pi2565;
assign w5527 = ~w5525 & ~w5526;
assign w5528 = w5524 & w5527;
assign w5529 = pi1343 & pi2325;
assign w5530 = pi1342 & pi2311;
assign w5531 = ~w5529 & ~w5530;
assign w5532 = pi1355 & pi2459;
assign w5533 = pi1357 & pi2468;
assign w5534 = ~w5532 & ~w5533;
assign w5535 = w5531 & w5534;
assign w5536 = pi1349 & pi2736;
assign w5537 = pi1340 & pi2289;
assign w5538 = ~w5536 & ~w5537;
assign w5539 = pi1341 & pi2088;
assign w5540 = pi1354 & pi2749;
assign w5541 = ~w5539 & ~w5540;
assign w5542 = w5538 & w5541;
assign w5543 = w5535 & w5542;
assign w5544 = (pi0539 & ~w5543) | (pi0539 & w36607) | (~w5543 & w36607);
assign w5545 = pi1333 & pi1714;
assign w5546 = pi1332 & pi2580;
assign w5547 = ~w5545 & ~w5546;
assign w5548 = pi0224 & pi1336;
assign w5549 = pi1335 & pi2595;
assign w5550 = ~w5548 & ~w5549;
assign w5551 = w5547 & w5550;
assign w5552 = (~w941 & w5551) | (~w941 & w36608) | (w5551 & w36608);
assign w5553 = ~w5544 & w5552;
assign w5554 = ~w5521 & w5553;
assign w5555 = pi0979 & pi1966;
assign w5556 = ~pi0979 & pi2511;
assign w5557 = ~w5555 & ~w5556;
assign w5558 = pi0768 & ~w5557;
assign w5559 = pi0979 & pi2156;
assign w5560 = ~pi0979 & pi2778;
assign w5561 = ~w5559 & ~w5560;
assign w5562 = pi0767 & ~w5561;
assign w5563 = ~w5558 & ~w5562;
assign w5564 = pi0180 & ~pi0979;
assign w5565 = pi0165 & pi0979;
assign w5566 = ~w5564 & ~w5565;
assign w5567 = pi0838 & ~w5566;
assign w5568 = pi0979 & pi2174;
assign w5569 = ~pi0979 & pi2801;
assign w5570 = ~w5568 & ~w5569;
assign w5571 = pi0836 & ~w5570;
assign w5572 = pi0979 & pi2190;
assign w5573 = ~pi0979 & pi3079;
assign w5574 = ~w5572 & ~w5573;
assign w5575 = pi0837 & ~w5574;
assign w5576 = ~w5571 & ~w5575;
assign w5577 = ~w5567 & w5576;
assign w5578 = w5563 & w5577;
assign w5579 = (pi0576 & ~w5577) | (pi0576 & w36609) | (~w5577 & w36609);
assign w5580 = pi0979 & pi2622;
assign w5581 = ~pi0979 & pi2628;
assign w5582 = ~w5580 & ~w5581;
assign w5583 = pi0764 & ~w5582;
assign w5584 = pi0979 & pi3184;
assign w5585 = ~pi0979 & pi2896;
assign w5586 = ~w5584 & ~w5585;
assign w5587 = pi0766 & ~w5586;
assign w5588 = pi0087 & ~pi0979;
assign w5589 = pi0085 & pi0979;
assign w5590 = ~w5588 & ~w5589;
assign w5591 = pi0720 & ~w5590;
assign w5592 = ~w5587 & ~w5591;
assign w5593 = ~w5583 & w5592;
assign w5594 = pi0979 & pi3175;
assign w5595 = ~pi0979 & pi2538;
assign w5596 = ~w5594 & ~w5595;
assign w5597 = pi0765 & ~w5596;
assign w5598 = ~w1144 & ~w5597;
assign w5599 = pi0979 & pi2609;
assign w5600 = ~pi0979 & pi2616;
assign w5601 = ~w5599 & ~w5600;
assign w5602 = pi0763 & ~w5601;
assign w5603 = pi0257 & ~pi0979;
assign w5604 = pi0255 & pi0979;
assign w5605 = ~w5603 & ~w5604;
assign w5606 = pi0721 & ~w5605;
assign w5607 = ~w5602 & ~w5606;
assign w5608 = w5598 & w5607;
assign w5609 = w5593 & w5608;
assign w5610 = pi0524 & ~w5609;
assign w5611 = pi0234 & ~pi0979;
assign w5612 = pi0233 & pi0979;
assign w5613 = ~w5611 & ~w5612;
assign w5614 = pi0716 & ~w5613;
assign w5615 = pi0283 & ~pi0979;
assign w5616 = pi0281 & pi0979;
assign w5617 = ~w5615 & ~w5616;
assign w5618 = pi0761 & ~w5617;
assign w5619 = pi0979 & pi2137;
assign w5620 = ~pi0979 & pi2854;
assign w5621 = ~w5619 & ~w5620;
assign w5622 = pi0717 & ~w5621;
assign w5623 = ~w5618 & ~w5622;
assign w5624 = ~w5614 & w5623;
assign w5625 = (pi0538 & ~w5624) | (pi0538 & w35782) | (~w5624 & w35782);
assign w5626 = ~w5610 & w36610;
assign w5627 = w5554 & w5626;
assign w5628 = ~w5498 & w5627;
assign w5629 = ~w941 & ~w5628;
assign w5630 = ~w5491 & ~w5629;
assign w5631 = pi3295 & ~w5628;
assign w5632 = (~pi1787 & ~w5630) | (~pi1787 & w36611) | (~w5630 & w36611);
assign w5633 = pi1787 & pi2834;
assign w5634 = w958 & w36612;
assign w5635 = (~w5448 & w5632) | (~w5448 & w36613) | (w5632 & w36613);
assign w5636 = w3433 & w5635;
assign w5637 = pi2440 & w1314;
assign w5638 = ~w414 & w36614;
assign w5639 = ~w5637 & ~w5638;
assign w5640 = pi2703 & w1316;
assign w5641 = pi2277 & w1309;
assign w5642 = ~w5640 & ~w5641;
assign w5643 = w5639 & w5642;
assign w5644 = ~w414 & w36615;
assign w5645 = ~w405 & w36616;
assign w5646 = ~w5644 & ~w5645;
assign w5647 = ~w371 & w36617;
assign w5648 = ~w392 & w36618;
assign w5649 = ~w5647 & ~w5648;
assign w5650 = w5646 & w5649;
assign w5651 = (~w354 & ~w5646) | (~w354 & w36619) | (~w5646 & w36619);
assign w5652 = w5643 & ~w5651;
assign w5653 = (pi2749 & w2346) | (pi2749 & w36620) | (w2346 & w36620);
assign w5654 = (pi2468 & w2336) | (pi2468 & w36621) | (w2336 & w36621);
assign w5655 = ~w5653 & ~w5654;
assign w5656 = (pi2459 & w2330) | (pi2459 & w36622) | (w2330 & w36622);
assign w5657 = pi2544 & ~w2342;
assign w5658 = ~w5656 & ~w5657;
assign w5659 = w5655 & w5658;
assign w5660 = w5658 & w36623;
assign w5661 = pi2468 & w2875;
assign w5662 = w2297 & w5661;
assign w5663 = (pi2459 & w2293) | (pi2459 & w36624) | (w2293 & w36624);
assign w5664 = w2295 & w5663;
assign w5665 = w354 & ~w5664;
assign w5666 = pi2749 & w3907;
assign w5667 = pi2544 & w2881;
assign w5668 = ~w5666 & ~w5667;
assign w5669 = w5668 & w36625;
assign w5670 = ~w5660 & ~w5669;
assign w5671 = w5652 & ~w5670;
assign w5672 = w2958 & ~w5671;
assign w5673 = w940 & w36626;
assign w5674 = (pi1331 & ~w1956) | (pi1331 & w36627) | (~w1956 & w36627);
assign w5675 = pi0685 & pi1334;
assign w5676 = pi1053 & pi2514;
assign w5677 = ~w5675 & ~w5676;
assign w5678 = pi0592 & pi1359;
assign w5679 = pi1058 & pi3328;
assign w5680 = ~w5678 & ~w5679;
assign w5681 = w5677 & w5680;
assign w5682 = pi3510 & ~w1054;
assign w5683 = pi0918 & pi1358;
assign w5684 = pi0829 & pi1344;
assign w5685 = ~w5683 & ~w5684;
assign w5686 = pi1059 & pi2979;
assign w5687 = pi0389 & pi1057;
assign w5688 = ~w5686 & ~w5687;
assign w5689 = w5685 & w5688;
assign w5690 = ~w5682 & w5689;
assign w5691 = w5681 & w5690;
assign w5692 = (pi0650 & w5674) | (pi0650 & w36628) | (w5674 & w36628);
assign w5693 = pi0042 & ~pi0979;
assign w5694 = pi0040 & pi0979;
assign w5695 = ~w5693 & ~w5694;
assign w5696 = pi0719 & ~w5695;
assign w5697 = pi0979 & pi3170;
assign w5698 = ~pi0979 & pi2636;
assign w5699 = ~w5697 & ~w5698;
assign w5700 = pi0765 & ~w5699;
assign w5701 = pi0490 & ~pi0979;
assign w5702 = pi0489 & pi0979;
assign w5703 = ~w5701 & ~w5702;
assign w5704 = pi0721 & ~w5703;
assign w5705 = ~w5700 & ~w5704;
assign w5706 = ~w5696 & w5705;
assign w5707 = pi0979 & pi3122;
assign w5708 = ~pi0979 & pi2892;
assign w5709 = ~w5707 & ~w5708;
assign w5710 = pi0766 & ~w5709;
assign w5711 = pi0979 & pi3156;
assign w5712 = ~pi0979 & pi2866;
assign w5713 = ~w5711 & ~w5712;
assign w5714 = pi0763 & ~w5713;
assign w5715 = ~w5710 & ~w5714;
assign w5716 = pi0217 & ~pi0979;
assign w5717 = pi0216 & pi0979;
assign w5718 = ~w5716 & ~w5717;
assign w5719 = pi0720 & ~w5718;
assign w5720 = pi0979 & pi3164;
assign w5721 = ~pi0979 & pi2875;
assign w5722 = ~w5720 & ~w5721;
assign w5723 = pi0764 & ~w5722;
assign w5724 = ~w5719 & ~w5723;
assign w5725 = w5715 & w5724;
assign w5726 = w5706 & w5725;
assign w5727 = pi0524 & ~w5726;
assign w5728 = pi1347 & pi2682;
assign w5729 = pi1339 & pi2250;
assign w5730 = ~w5728 & ~w5729;
assign w5731 = pi1352 & pi2274;
assign w5732 = pi1346 & pi2668;
assign w5733 = ~w5731 & ~w5732;
assign w5734 = w5730 & w5733;
assign w5735 = pi1600 & pi2208;
assign w5736 = pi1353 & pi1981;
assign w5737 = ~w5735 & ~w5736;
assign w5738 = pi1348 & pi2692;
assign w5739 = pi1338 & pi2236;
assign w5740 = ~w5738 & ~w5739;
assign w5741 = w5737 & w5740;
assign w5742 = pi1350 & pi2433;
assign w5743 = pi1337 & pi2222;
assign w5744 = ~w5742 & ~w5743;
assign w5745 = pi1345 & pi2654;
assign w5746 = pi1351 & pi2266;
assign w5747 = ~w5745 & ~w5746;
assign w5748 = w5744 & w5747;
assign w5749 = w5741 & w5748;
assign w5750 = (pi0722 & ~w5749) | (pi0722 & w36629) | (~w5749 & w36629);
assign w5751 = ~w5727 & ~w5750;
assign w5752 = pi0207 & ~pi0979;
assign w5753 = pi0201 & pi0979;
assign w5754 = ~w5752 & ~w5753;
assign w5755 = pi1599 & ~w5754;
assign w5756 = pi0300 & ~pi0979;
assign w5757 = pi0299 & pi0979;
assign w5758 = ~w5756 & ~w5757;
assign w5759 = pi0761 & ~w5758;
assign w5760 = ~w5755 & ~w5759;
assign w5761 = pi0400 & ~pi0979;
assign w5762 = pi0399 & pi0979;
assign w5763 = ~w5761 & ~w5762;
assign w5764 = pi0718 & ~w5763;
assign w5765 = pi0316 & ~pi0979;
assign w5766 = pi0315 & pi0979;
assign w5767 = ~w5765 & ~w5766;
assign w5768 = pi0716 & ~w5767;
assign w5769 = pi0979 & pi2131;
assign w5770 = ~pi0979 & pi2848;
assign w5771 = ~w5769 & ~w5770;
assign w5772 = pi0717 & ~w5771;
assign w5773 = ~w5768 & ~w5772;
assign w5774 = ~w5764 & w5773;
assign w5775 = (pi0538 & ~w5774) | (pi0538 & w36630) | (~w5774 & w36630);
assign w5776 = pi0979 & pi1962;
assign w5777 = ~pi0979 & pi2427;
assign w5778 = ~w5776 & ~w5777;
assign w5779 = pi0152 & pi1360;
assign w5780 = (~w5779 & w5778) | (~w5779 & w36631) | (w5778 & w36631);
assign w5781 = pi0175 & ~pi0979;
assign w5782 = pi0160 & pi0979;
assign w5783 = ~w5781 & ~w5782;
assign w5784 = pi0838 & ~w5783;
assign w5785 = pi0979 & pi2150;
assign w5786 = ~pi0979 & pi2922;
assign w5787 = ~w5785 & ~w5786;
assign w5788 = pi0767 & ~w5787;
assign w5789 = ~w5784 & ~w5788;
assign w5790 = pi0979 & pi2184;
assign w5791 = ~pi0979 & pi2945;
assign w5792 = ~w5790 & ~w5791;
assign w5793 = pi0837 & ~w5792;
assign w5794 = pi0979 & pi2168;
assign w5795 = ~pi0979 & pi2934;
assign w5796 = ~w5794 & ~w5795;
assign w5797 = pi0836 & ~w5796;
assign w5798 = ~w5793 & ~w5797;
assign w5799 = w5789 & w5798;
assign w5800 = (pi0576 & ~w5799) | (pi0576 & w36632) | (~w5799 & w36632);
assign w5801 = ~w5775 & ~w5800;
assign w5802 = w5751 & w5801;
assign w5803 = ~w5692 & w5802;
assign w5804 = ~w941 & ~w5803;
assign w5805 = w1216 & w36633;
assign w5806 = w1221 & w36634;
assign w5807 = w1221 & w36635;
assign w5808 = ~w5806 & ~w5807;
assign w5809 = ~w5805 & w5808;
assign w5810 = pi1943 & w3145;
assign w5811 = pi1032 & ~pi1432;
assign w5812 = (~w5811 & w5810) | (~w5811 & w36636) | (w5810 & w36636);
assign w5813 = pi1902 & w1238;
assign w5814 = pi1834 & w1268;
assign w5815 = ~w5813 & ~w5814;
assign w5816 = pi1443 & w1280;
assign w5817 = pi0846 & w1234;
assign w5818 = ~w5816 & ~w5817;
assign w5819 = w5815 & w5818;
assign w5820 = pi1101 & w1266;
assign w5821 = pi0737 & w1254;
assign w5822 = ~w5820 & ~w5821;
assign w5823 = pi0892 & w1291;
assign w5824 = pi1888 & w1278;
assign w5825 = ~w5823 & ~w5824;
assign w5826 = w5822 & w5825;
assign w5827 = w5819 & w5826;
assign w5828 = ~w5812 & w5827;
assign w5829 = pi2141 & w1275;
assign w5830 = ~w3180 & ~w5829;
assign w5831 = pi1734 & w3172;
assign w5832 = pi1756 & w1249;
assign w5833 = ~w5831 & ~w5832;
assign w5834 = pi0798 & w1288;
assign w5835 = pi1779 & w1258;
assign w5836 = ~w5834 & ~w5835;
assign w5837 = w5833 & w5836;
assign w5838 = w5830 & w5837;
assign w5839 = pi0907 & w1296;
assign w5840 = pi1457 & w3148;
assign w5841 = ~w5839 & ~w5840;
assign w5842 = pi0728 & w1242;
assign w5843 = pi1926 & w1272;
assign w5844 = ~w5842 & ~w5843;
assign w5845 = w5841 & w5844;
assign w5846 = pi1766 & w1263;
assign w5847 = pi1009 & w1245;
assign w5848 = ~w5846 & ~w5847;
assign w5849 = pi1720 & w1294;
assign w5850 = pi0885 & w1251;
assign w5851 = ~w5849 & ~w5850;
assign w5852 = w5848 & w5851;
assign w5853 = w5845 & w5852;
assign w5854 = w5838 & w5853;
assign w5855 = w1216 & w36637;
assign w5856 = w1221 & w36638;
assign w5857 = ~w5855 & ~w5856;
assign w5858 = w5854 & w5857;
assign w5859 = w5858 & w36639;
assign w5860 = pi1357 & pi2411;
assign w5861 = pi1349 & pi2560;
assign w5862 = ~w5860 & ~w5861;
assign w5863 = pi1355 & pi2526;
assign w5864 = pi1054 & pi2714;
assign w5865 = ~w5863 & ~w5864;
assign w5866 = w5862 & w5865;
assign w5867 = pi1342 & pi2307;
assign w5868 = pi1055 & pi2724;
assign w5869 = ~w5867 & ~w5868;
assign w5870 = pi1354 & pi2776;
assign w5871 = pi1340 & pi2286;
assign w5872 = ~w5870 & ~w5871;
assign w5873 = w5869 & w5872;
assign w5874 = pi1056 & pi2547;
assign w5875 = pi1343 & pi2321;
assign w5876 = ~w5874 & ~w5875;
assign w5877 = pi1341 & pi2298;
assign w5878 = pi1356 & pi2967;
assign w5879 = ~w5877 & ~w5878;
assign w5880 = w5876 & w5879;
assign w5881 = w5873 & w5880;
assign w5882 = (w5289 & ~w5881) | (w5289 & w36640) | (~w5881 & w36640);
assign w5883 = pi1332 & pi2574;
assign w5884 = pi1335 & pi2589;
assign w5885 = ~w5883 & ~w5884;
assign w5886 = pi0127 & pi1333;
assign w5887 = pi0350 & pi1336;
assign w5888 = ~w5886 & ~w5887;
assign w5889 = w5885 & w5888;
assign w5890 = w1607 & ~w5889;
assign w5891 = ~w5882 & ~w5890;
assign w5892 = (w5891 & w5859) | (w5891 & w36641) | (w5859 & w36641);
assign w5893 = ~w5804 & w5892;
assign w5894 = pi1787 & pi2830;
assign w5895 = w958 & w36643;
assign w5896 = pi3861 & w983;
assign w5897 = w973 & w36646;
assign w5898 = w970 & w36647;
assign w5899 = w970 & w36648;
assign w5900 = ~w5898 & ~w5899;
assign w5901 = ~w5897 & w5900;
assign w5902 = w963 & w36649;
assign w5903 = w953 & w36650;
assign w5904 = w958 & w36651;
assign w5905 = ~w5903 & ~w5904;
assign w5906 = ~w5902 & w5905;
assign w5907 = w973 & w36652;
assign w5908 = w963 & w36653;
assign w5909 = ~w997 & ~w5908;
assign w5910 = ~w5907 & w5909;
assign w5911 = w5906 & w5910;
assign w5912 = w5901 & w5911;
assign w5913 = ~w5896 & w5912;
assign w5914 = ~w5913 & w40109;
assign w5915 = w2961 & w5914;
assign w5916 = ~w5672 & ~w5915;
assign w5917 = (w2397 & ~w5916) | (w2397 & w36656) | (~w5916 & w36656);
assign w5918 = w2417 & ~w5652;
assign w5919 = ~w5669 & w36657;
assign w5920 = (w353 & w36658) | (w353 & w36659) | (w36658 & w36659);
assign w5921 = w5920 & w40102;
assign w5922 = (pi1037 & w2907) | (pi1037 & w36660) | (w2907 & w36660);
assign w5923 = w940 & w36661;
assign w5924 = w2236 & w36662;
assign w5925 = (~w5923 & ~w359) | (~w5923 & w36664) | (~w359 & w36664);
assign w5926 = ~w5922 & w36665;
assign w5927 = ~w5919 & w5926;
assign w5928 = ~w5918 & w5927;
assign w5929 = ~w2899 & ~w5928;
assign w5930 = pi0780 & w2899;
assign w5931 = (~w5930 & w2386) | (~w5930 & w36666) | (w2386 & w36666);
assign w5932 = ~w5929 & w5931;
assign w5933 = (pi2526 & w2330) | (pi2526 & w36667) | (w2330 & w36667);
assign w5934 = (pi2411 & w2336) | (pi2411 & w36668) | (w2336 & w36668);
assign w5935 = ~w5933 & ~w5934;
assign w5936 = (pi2776 & w2346) | (pi2776 & w36669) | (w2346 & w36669);
assign w5937 = pi2967 & ~w2342;
assign w5938 = ~w5936 & ~w5937;
assign w5939 = w5935 & w5938;
assign w5940 = w5938 & w36670;
assign w5941 = pi2411 & w2875;
assign w5942 = w2297 & w5941;
assign w5943 = (pi2526 & w2293) | (pi2526 & w36671) | (w2293 & w36671);
assign w5944 = w2295 & w5943;
assign w5945 = w354 & ~w5944;
assign w5946 = pi2967 & w2881;
assign w5947 = pi2776 & w3907;
assign w5948 = ~w5946 & ~w5947;
assign w5949 = w5948 & w36672;
assign w5950 = ~w5940 & ~w5949;
assign w5951 = ~w2386 & w36673;
assign w5952 = w3754 & ~w5951;
assign w5953 = ~w5932 & w5952;
assign w5954 = ~w5917 & ~w5953;
assign w5955 = (w5954 & w2826) | (w5954 & w36674) | (w2826 & w36674);
assign w5956 = ~w5424 & w5955;
assign w5957 = ~w5416 & w5956;
assign w5958 = ~w5398 & w5957;
assign w5959 = ~w5379 & ~w5958;
assign w5960 = pi0661 & w541;
assign w5961 = (~w544 & w530) | (~w544 & w36675) | (w530 & w36675);
assign w5962 = ~w2407 & ~w5961;
assign w5963 = ~w5960 & ~w5962;
assign w5964 = (w5963 & ~w797) | (w5963 & w36676) | (~w797 & w36676);
assign w5965 = (~w645 & w634) | (~w645 & w36677) | (w634 & w36677);
assign w5966 = ~w647 & ~w5960;
assign w5967 = ~w5965 & w5966;
assign w5968 = w797 & w36678;
assign w5969 = ~w5964 & ~w5968;
assign w5970 = pi3867 & w983;
assign w5971 = w970 & w36679;
assign w5972 = w973 & w36680;
assign w5973 = w970 & w36681;
assign w5974 = ~w5972 & ~w5973;
assign w5975 = ~w5971 & w5974;
assign w5976 = w963 & w36682;
assign w5977 = w953 & w36683;
assign w5978 = w963 & w36684;
assign w5979 = ~w5977 & ~w5978;
assign w5980 = ~w5976 & w5979;
assign w5981 = w973 & w36685;
assign w5982 = w958 & w36686;
assign w5983 = ~w997 & ~w5982;
assign w5984 = ~w5981 & w5983;
assign w5985 = w5980 & w5984;
assign w5986 = w5975 & w5985;
assign w5987 = ~w5970 & w5986;
assign w5988 = w940 & w36687;
assign w5989 = (pi1331 & ~w2166) | (pi1331 & w36688) | (~w2166 & w36688);
assign w5990 = pi3518 & ~w1054;
assign w5991 = pi0383 & pi1057;
assign w5992 = pi0602 & pi1359;
assign w5993 = pi0913 & pi1358;
assign w5994 = ~w5992 & ~w5993;
assign w5995 = ~w5991 & w5994;
assign w5996 = ~w5990 & w5995;
assign w5997 = (pi0650 & w5989) | (pi0650 & w36689) | (w5989 & w36689);
assign w5998 = pi1054 & pi2709;
assign w5999 = pi1055 & pi2720;
assign w6000 = ~w5998 & ~w5999;
assign w6001 = pi1355 & pi2520;
assign w6002 = pi1356 & pi2752;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = w6000 & w6003;
assign w6005 = pi1340 & pi2280;
assign w6006 = pi1354 & pi2535;
assign w6007 = ~w6005 & ~w6006;
assign w6008 = pi1357 & pi2412;
assign w6009 = pi1056 & pi2739;
assign w6010 = ~w6008 & ~w6009;
assign w6011 = w6007 & w6010;
assign w6012 = pi1349 & pi2566;
assign w6013 = pi1342 & pi2089;
assign w6014 = ~w6012 & ~w6013;
assign w6015 = pi1341 & pi2067;
assign w6016 = pi1343 & pi2315;
assign w6017 = ~w6015 & ~w6016;
assign w6018 = w6014 & w6017;
assign w6019 = w6011 & w6018;
assign w6020 = (pi0539 & ~w6019) | (pi0539 & w36690) | (~w6019 & w36690);
assign w6021 = pi1600 & pi2202;
assign w6022 = pi1348 & pi2687;
assign w6023 = ~w6021 & ~w6022;
assign w6024 = pi1339 & pi2244;
assign w6025 = pi1352 & pi2701;
assign w6026 = ~w6024 & ~w6025;
assign w6027 = w6023 & w6026;
assign w6028 = pi1345 & pi2648;
assign w6029 = pi1346 & pi2662;
assign w6030 = ~w6028 & ~w6029;
assign w6031 = pi1337 & pi2216;
assign w6032 = pi1353 & pi2275;
assign w6033 = ~w6031 & ~w6032;
assign w6034 = w6030 & w6033;
assign w6035 = pi1350 & pi2698;
assign w6036 = pi1351 & pi2438;
assign w6037 = ~w6035 & ~w6036;
assign w6038 = pi1338 & pi2230;
assign w6039 = pi1347 & pi2676;
assign w6040 = ~w6038 & ~w6039;
assign w6041 = w6037 & w6040;
assign w6042 = w6034 & w6041;
assign w6043 = (pi0722 & ~w6042) | (pi0722 & w36691) | (~w6042 & w36691);
assign w6044 = pi0232 & pi1336;
assign w6045 = pi1335 & pi2584;
assign w6046 = ~w6044 & ~w6045;
assign w6047 = pi1333 & pi1741;
assign w6048 = pi1332 & pi2568;
assign w6049 = ~w6047 & ~w6048;
assign w6050 = w6046 & w6049;
assign w6051 = pi0762 & ~w6050;
assign w6052 = ~w6043 & ~w6051;
assign w6053 = ~w6020 & w6052;
assign w6054 = pi0294 & ~pi0979;
assign w6055 = pi0293 & pi0979;
assign w6056 = ~w6054 & ~w6055;
assign w6057 = pi0721 & ~w6056;
assign w6058 = pi0146 & ~pi0979;
assign w6059 = pi0145 & pi0979;
assign w6060 = ~w6058 & ~w6059;
assign w6061 = pi0720 & ~w6060;
assign w6062 = pi0979 & pi3168;
assign w6063 = ~pi0979 & pi2631;
assign w6064 = ~w6062 & ~w6063;
assign w6065 = pi0765 & ~w6064;
assign w6066 = ~w6061 & ~w6065;
assign w6067 = ~w6057 & w6066;
assign w6068 = pi0979 & pi3177;
assign w6069 = ~pi0979 & pi2889;
assign w6070 = ~w6068 & ~w6069;
assign w6071 = pi0766 & ~w6070;
assign w6072 = ~w1144 & ~w6071;
assign w6073 = pi0979 & pi2619;
assign w6074 = ~pi0979 & pi2625;
assign w6075 = ~w6073 & ~w6074;
assign w6076 = pi0764 & ~w6075;
assign w6077 = pi0979 & pi2606;
assign w6078 = ~pi0979 & pi2612;
assign w6079 = ~w6077 & ~w6078;
assign w6080 = pi0763 & ~w6079;
assign w6081 = ~w6076 & ~w6080;
assign w6082 = w6072 & w6081;
assign w6083 = w6067 & w6082;
assign w6084 = pi0524 & ~w6083;
assign w6085 = pi0239 & ~pi0979;
assign w6086 = pi0238 & pi0979;
assign w6087 = ~w6085 & ~w6086;
assign w6088 = pi0716 & ~w6087;
assign w6089 = pi0236 & ~pi0979;
assign w6090 = pi0235 & pi0979;
assign w6091 = ~w6089 & ~w6090;
assign w6092 = pi0761 & ~w6091;
assign w6093 = pi0979 & pi2125;
assign w6094 = ~pi0979 & pi2842;
assign w6095 = ~w6093 & ~w6094;
assign w6096 = pi0717 & ~w6095;
assign w6097 = ~w6092 & ~w6096;
assign w6098 = ~w6088 & w6097;
assign w6099 = (pi0538 & ~w6098) | (pi0538 & w35782) | (~w6098 & w35782);
assign w6100 = pi0979 & pi2178;
assign w6101 = ~pi0979 & pi2940;
assign w6102 = ~w6100 & ~w6101;
assign w6103 = pi0837 & ~w6102;
assign w6104 = pi0979 & pi2145;
assign w6105 = ~pi0979 & pi2917;
assign w6106 = ~w6104 & ~w6105;
assign w6107 = pi0767 & ~w6106;
assign w6108 = ~w6103 & ~w6107;
assign w6109 = pi0168 & ~pi0979;
assign w6110 = pi0154 & pi0979;
assign w6111 = ~w6109 & ~w6110;
assign w6112 = pi0838 & ~w6111;
assign w6113 = pi0979 & pi1956;
assign w6114 = ~pi0979 & pi2421;
assign w6115 = ~w6113 & ~w6114;
assign w6116 = pi0768 & ~w6115;
assign w6117 = pi0979 & pi2162;
assign w6118 = ~pi0979 & pi2809;
assign w6119 = ~w6117 & ~w6118;
assign w6120 = pi0836 & ~w6119;
assign w6121 = ~w6116 & ~w6120;
assign w6122 = ~w6112 & w6121;
assign w6123 = (pi0576 & ~w6122) | (pi0576 & w36692) | (~w6122 & w36692);
assign w6124 = ~w6099 & ~w6123;
assign w6125 = ~w6084 & w6124;
assign w6126 = w6053 & w6125;
assign w6127 = ~w5997 & w6126;
assign w6128 = ~w941 & ~w6127;
assign w6129 = w1221 & w36693;
assign w6130 = w1216 & w36694;
assign w6131 = ~w6129 & ~w6130;
assign w6132 = w1221 & w36695;
assign w6133 = w1216 & w36696;
assign w6134 = ~w6132 & ~w6133;
assign w6135 = w6131 & w6134;
assign w6136 = pi1451 & w3148;
assign w6137 = pi1898 & w1238;
assign w6138 = ~w6136 & ~w6137;
assign w6139 = pi1883 & w1278;
assign w6140 = pi1773 & w1258;
assign w6141 = ~w6139 & ~w6140;
assign w6142 = w6138 & w6141;
assign w6143 = pi1437 & w1280;
assign w6144 = pi1728 & w3172;
assign w6145 = ~w6143 & ~w6144;
assign w6146 = pi1919 & w1272;
assign w6147 = pi1878 & w1294;
assign w6148 = ~w6146 & ~w6147;
assign w6149 = w6145 & w6148;
assign w6150 = pi0790 & w1251;
assign w6151 = pi0458 & w1242;
assign w6152 = ~w6150 & ~w6151;
assign w6153 = pi0968 & w1234;
assign w6154 = pi0894 & w1254;
assign w6155 = ~w6153 & ~w6154;
assign w6156 = w6152 & w6155;
assign w6157 = w6149 & w6156;
assign w6158 = w6142 & w6157;
assign w6159 = w1221 & w36697;
assign w6160 = pi1829 & w1268;
assign w6161 = ~w3180 & ~w6160;
assign w6162 = pi0903 & w1296;
assign w6163 = pi0941 & w1245;
assign w6164 = ~w6162 & ~w6163;
assign w6165 = w6161 & w6164;
assign w6166 = w1291 & w36698;
assign w6167 = w1288 & w36699;
assign w6168 = ~w6166 & ~w6167;
assign w6169 = w6165 & w36700;
assign w6170 = w6158 & w36701;
assign w6171 = pi1934 & ~w6170;
assign w6172 = ~w6128 & ~w6171;
assign w6173 = ~w6128 & w36702;
assign w6174 = pi1787 & pi3150;
assign w6175 = w958 & w36703;
assign w6176 = (w6175 & w6173) | (w6175 & w36704) | (w6173 & w36704);
assign w6177 = ~w5987 & ~w6176;
assign w6178 = w2961 & w6177;
assign w6179 = pi3864 & w983;
assign w6180 = w970 & w36705;
assign w6181 = w973 & w36706;
assign w6182 = w970 & w36707;
assign w6183 = ~w6181 & ~w6182;
assign w6184 = ~w6180 & w6183;
assign w6185 = w958 & w36708;
assign w6186 = w963 & w36709;
assign w6187 = w953 & w36710;
assign w6188 = ~w6186 & ~w6187;
assign w6189 = ~w6185 & w6188;
assign w6190 = w973 & w36711;
assign w6191 = w963 & w36712;
assign w6192 = ~w997 & ~w6191;
assign w6193 = ~w6190 & w6192;
assign w6194 = w6189 & w6193;
assign w6195 = w6184 & w6194;
assign w6196 = ~w6179 & w6195;
assign w6197 = pi1334 & pi2379;
assign w6198 = pi1053 & pi2404;
assign w6199 = ~w6197 & ~w6198;
assign w6200 = pi0386 & pi1057;
assign w6201 = pi0827 & pi1344;
assign w6202 = ~w6200 & ~w6201;
assign w6203 = w6199 & w6202;
assign w6204 = pi3508 & ~w1054;
assign w6205 = pi0916 & pi1358;
assign w6206 = pi0578 & pi1359;
assign w6207 = ~w6205 & ~w6206;
assign w6208 = ~w6204 & w6207;
assign w6209 = w6203 & w6208;
assign w6210 = w6209 & w40110;
assign w6211 = pi0650 & ~w6210;
assign w6212 = pi1342 & pi2084;
assign w6213 = pi1056 & pi2741;
assign w6214 = ~w6212 & ~w6213;
assign w6215 = pi1355 & pi2527;
assign w6216 = pi1349 & pi2731;
assign w6217 = ~w6215 & ~w6216;
assign w6218 = w6214 & w6217;
assign w6219 = pi1341 & pi2295;
assign w6220 = pi1357 & pi2463;
assign w6221 = ~w6219 & ~w6220;
assign w6222 = pi1054 & pi2536;
assign w6223 = pi1055 & pi2721;
assign w6224 = ~w6222 & ~w6223;
assign w6225 = w6221 & w6224;
assign w6226 = pi1356 & pi2753;
assign w6227 = pi1340 & pi2283;
assign w6228 = ~w6226 & ~w6227;
assign w6229 = pi1343 & pi2318;
assign w6230 = pi1354 & pi2746;
assign w6231 = ~w6229 & ~w6230;
assign w6232 = w6228 & w6231;
assign w6233 = w6225 & w6232;
assign w6234 = (pi0539 & ~w6233) | (pi0539 & w36714) | (~w6233 & w36714);
assign w6235 = pi1337 & pi2219;
assign w6236 = pi1348 & pi2689;
assign w6237 = ~w6235 & ~w6236;
assign w6238 = pi1350 & pi2432;
assign w6239 = pi1352 & pi2442;
assign w6240 = ~w6238 & ~w6239;
assign w6241 = w6237 & w6240;
assign w6242 = pi1600 & pi2205;
assign w6243 = pi1345 & pi2651;
assign w6244 = ~w6242 & ~w6243;
assign w6245 = pi1339 & pi2247;
assign w6246 = pi1347 & pi2679;
assign w6247 = ~w6245 & ~w6246;
assign w6248 = w6244 & w6247;
assign w6249 = pi1351 & pi2263;
assign w6250 = pi1353 & pi1978;
assign w6251 = ~w6249 & ~w6250;
assign w6252 = pi1338 & pi2233;
assign w6253 = pi1346 & pi2665;
assign w6254 = ~w6252 & ~w6253;
assign w6255 = w6251 & w6254;
assign w6256 = w6248 & w6255;
assign w6257 = (pi0722 & ~w6256) | (pi0722 & w36715) | (~w6256 & w36715);
assign w6258 = pi0314 & pi1333;
assign w6259 = pi1335 & pi2764;
assign w6260 = ~w6258 & ~w6259;
assign w6261 = pi0278 & pi1336;
assign w6262 = pi1332 & pi2571;
assign w6263 = ~w6261 & ~w6262;
assign w6264 = w6260 & w6263;
assign w6265 = (~w941 & w6264) | (~w941 & w36608) | (w6264 & w36608);
assign w6266 = ~w6257 & w6265;
assign w6267 = ~w6234 & w6266;
assign w6268 = pi0171 & ~pi0979;
assign w6269 = pi0157 & pi0979;
assign w6270 = ~w6268 & ~w6269;
assign w6271 = pi0143 & pi1360;
assign w6272 = (~w6271 & w6270) | (~w6271 & w36716) | (w6270 & w36716);
assign w6273 = pi0979 & pi1959;
assign w6274 = ~pi0979 & pi2424;
assign w6275 = ~w6273 & ~w6274;
assign w6276 = pi0768 & ~w6275;
assign w6277 = pi0979 & pi2181;
assign w6278 = ~pi0979 & pi2942;
assign w6279 = ~w6277 & ~w6278;
assign w6280 = pi0837 & ~w6279;
assign w6281 = ~w6276 & ~w6280;
assign w6282 = pi0979 & pi2085;
assign w6283 = ~pi0979 & pi2787;
assign w6284 = ~w6282 & ~w6283;
assign w6285 = pi0767 & ~w6284;
assign w6286 = pi0979 & pi2165;
assign w6287 = ~pi0979 & pi2807;
assign w6288 = ~w6286 & ~w6287;
assign w6289 = pi0836 & ~w6288;
assign w6290 = ~w6285 & ~w6289;
assign w6291 = w6281 & w6290;
assign w6292 = (pi0576 & ~w6291) | (pi0576 & w36717) | (~w6291 & w36717);
assign w6293 = pi0488 & ~pi0979;
assign w6294 = pi0485 & pi0979;
assign w6295 = ~w6293 & ~w6294;
assign w6296 = pi0718 & ~w6295;
assign w6297 = ~w1179 & ~w6296;
assign w6298 = pi0979 & pi2128;
assign w6299 = ~pi0979 & pi2845;
assign w6300 = ~w6298 & ~w6299;
assign w6301 = pi0717 & ~w6300;
assign w6302 = pi0263 & ~pi0979;
assign w6303 = pi0259 & pi0979;
assign w6304 = ~w6302 & ~w6303;
assign w6305 = pi0716 & ~w6304;
assign w6306 = pi0291 & ~pi0979;
assign w6307 = pi0288 & pi0979;
assign w6308 = ~w6306 & ~w6307;
assign w6309 = pi0761 & ~w6308;
assign w6310 = ~w6305 & ~w6309;
assign w6311 = ~w6301 & w6310;
assign w6312 = w6297 & w6311;
assign w6313 = (pi0538 & ~w6311) | (pi0538 & w36718) | (~w6311 & w36718);
assign w6314 = pi0064 & ~pi0979;
assign w6315 = pi0062 & pi0979;
assign w6316 = ~w6314 & ~w6315;
assign w6317 = pi0719 & ~w6316;
assign w6318 = pi0335 & ~pi0979;
assign w6319 = pi0334 & pi0979;
assign w6320 = ~w6318 & ~w6319;
assign w6321 = pi0721 & ~w6320;
assign w6322 = pi0979 & pi3153;
assign w6323 = ~pi0979 & pi2864;
assign w6324 = ~w6322 & ~w6323;
assign w6325 = pi0763 & ~w6324;
assign w6326 = ~w6321 & ~w6325;
assign w6327 = ~w6317 & w6326;
assign w6328 = pi0191 & ~pi0979;
assign w6329 = pi0190 & pi0979;
assign w6330 = ~w6328 & ~w6329;
assign w6331 = pi0720 & ~w6330;
assign w6332 = pi0979 & pi3179;
assign w6333 = ~pi0979 & pi3074;
assign w6334 = ~w6332 & ~w6333;
assign w6335 = pi0766 & ~w6334;
assign w6336 = ~w6331 & ~w6335;
assign w6337 = pi0979 & pi3134;
assign w6338 = ~pi0979 & pi2634;
assign w6339 = ~w6337 & ~w6338;
assign w6340 = pi0765 & ~w6339;
assign w6341 = pi0979 & pi3162;
assign w6342 = ~pi0979 & pi2872;
assign w6343 = ~w6341 & ~w6342;
assign w6344 = pi0764 & ~w6343;
assign w6345 = ~w6340 & ~w6344;
assign w6346 = w6336 & w6345;
assign w6347 = w6327 & w6346;
assign w6348 = pi0524 & ~w6347;
assign w6349 = ~w6348 & w36719;
assign w6350 = w6267 & w6349;
assign w6351 = ~w6211 & w6350;
assign w6352 = w940 & w36720;
assign w6353 = ~w6351 & ~w6352;
assign w6354 = w1221 & w36721;
assign w6355 = pi2522 & w1227;
assign w6356 = ~w6354 & ~w6355;
assign w6357 = w1221 & w36722;
assign w6358 = pi1603 & w1217;
assign w6359 = ~w6357 & ~w6358;
assign w6360 = w6356 & w6359;
assign w6361 = pi1454 & w3148;
assign w6362 = pi1717 & w1294;
assign w6363 = ~w6361 & ~w6362;
assign w6364 = pi0653 & w1242;
assign w6365 = pi1776 & w1258;
assign w6366 = ~w6364 & ~w6365;
assign w6367 = w6363 & w6366;
assign w6368 = pi0950 & w1291;
assign w6369 = pi1429 & w3139;
assign w6370 = ~w6368 & ~w6369;
assign w6371 = pi0955 & w1245;
assign w6372 = pi0905 & w1296;
assign w6373 = ~w6371 & ~w6372;
assign w6374 = w6370 & w6373;
assign w6375 = w6367 & w6374;
assign w6376 = pi2105 & w1275;
assign w6377 = pi1440 & w1280;
assign w6378 = ~w6376 & ~w6377;
assign w6379 = pi1940 & w3145;
assign w6380 = pi2054 & w1238;
assign w6381 = ~w6379 & ~w6380;
assign w6382 = w6378 & w6381;
assign w6383 = pi1753 & w1249;
assign w6384 = pi0882 & w1251;
assign w6385 = ~w6383 & ~w6384;
assign w6386 = pi1764 & w1263;
assign w6387 = pi0965 & w1288;
assign w6388 = ~w6386 & ~w6387;
assign w6389 = w6385 & w6388;
assign w6390 = w6382 & w6389;
assign w6391 = w6375 & w6390;
assign w6392 = w1221 & w36723;
assign w6393 = pi1920 & w1278;
assign w6394 = pi0744 & w1254;
assign w6395 = ~w6393 & ~w6394;
assign w6396 = pi1832 & w1268;
assign w6397 = pi1731 & w3172;
assign w6398 = ~w6396 & ~w6397;
assign w6399 = w6395 & w6398;
assign w6400 = pi1923 & w1272;
assign w6401 = ~w3180 & ~w6400;
assign w6402 = pi0802 & w1234;
assign w6403 = pi1021 & w1266;
assign w6404 = ~w6402 & ~w6403;
assign w6405 = w6401 & w6404;
assign w6406 = w6399 & w6405;
assign w6407 = ~w6392 & w6406;
assign w6408 = w6391 & w6407;
assign w6409 = (pi1934 & ~w6408) | (pi1934 & w36724) | (~w6408 & w36724);
assign w6410 = (~pi1787 & w6353) | (~pi1787 & w36725) | (w6353 & w36725);
assign w6411 = pi1787 & pi2827;
assign w6412 = w958 & w36726;
assign w6413 = (~w6196 & w6410) | (~w6196 & w36727) | (w6410 & w36727);
assign w6414 = w3433 & w6413;
assign w6415 = (pi2746 & w2346) | (pi2746 & w36728) | (w2346 & w36728);
assign w6416 = pi2753 & ~w2342;
assign w6417 = ~w6415 & ~w6416;
assign w6418 = (pi2527 & w2330) | (pi2527 & w36729) | (w2330 & w36729);
assign w6419 = (pi2463 & w2336) | (pi2463 & w36730) | (w2336 & w36730);
assign w6420 = ~w6418 & ~w6419;
assign w6421 = w6417 & w6420;
assign w6422 = w6417 & w36731;
assign w6423 = pi2463 & w2875;
assign w6424 = w2297 & w6423;
assign w6425 = (pi2527 & w2293) | (pi2527 & w36732) | (w2293 & w36732);
assign w6426 = w2295 & w6425;
assign w6427 = w354 & ~w6426;
assign w6428 = pi2746 & w3907;
assign w6429 = pi2753 & w2881;
assign w6430 = ~w6428 & ~w6429;
assign w6431 = w6430 & w36733;
assign w6432 = ~w6422 & ~w6431;
assign w6433 = pi1978 & w1309;
assign w6434 = ~w414 & w36734;
assign w6435 = ~w6433 & ~w6434;
assign w6436 = pi2442 & w1316;
assign w6437 = pi2263 & w1314;
assign w6438 = ~w6436 & ~w6437;
assign w6439 = w6435 & w6438;
assign w6440 = ~w371 & w36735;
assign w6441 = ~w392 & w36736;
assign w6442 = ~w6440 & ~w6441;
assign w6443 = ~w414 & w36737;
assign w6444 = ~w405 & w36738;
assign w6445 = ~w6443 & ~w6444;
assign w6446 = w6442 & w6445;
assign w6447 = (~w354 & ~w6445) | (~w354 & w36739) | (~w6445 & w36739);
assign w6448 = w6439 & ~w6447;
assign w6449 = ~w6432 & w6448;
assign w6450 = w2958 & ~w6449;
assign w6451 = ~w6414 & ~w6450;
assign w6452 = (w2397 & ~w6451) | (w2397 & w36740) | (~w6451 & w36740);
assign w6453 = ~pi0774 & w2899;
assign w6454 = w2236 & w36741;
assign w6455 = ~w6431 & w36742;
assign w6456 = (w2365 & w6455) | (w2365 & w36743) | (w6455 & w36743);
assign w6457 = w2417 & ~w6448;
assign w6458 = w940 & w36744;
assign w6459 = ~w2899 & ~w6458;
assign w6460 = (w353 & w36745) | (w353 & w36746) | (w36745 & w36746);
assign w6461 = w6460 & w40102;
assign w6462 = (pi1013 & w2907) | (pi1013 & w36747) | (w2907 & w36747);
assign w6463 = ~w6462 & w36748;
assign w6464 = ~w6457 & w6463;
assign w6465 = (~w6453 & ~w6464) | (~w6453 & w36749) | (~w6464 & w36749);
assign w6466 = ~w2387 & ~w6465;
assign w6467 = (pi2535 & w2346) | (pi2535 & w36750) | (w2346 & w36750);
assign w6468 = pi2752 & ~w2342;
assign w6469 = ~w6467 & ~w6468;
assign w6470 = (pi2520 & w2330) | (pi2520 & w36751) | (w2330 & w36751);
assign w6471 = (pi2412 & w2336) | (pi2412 & w36752) | (w2336 & w36752);
assign w6472 = ~w6470 & ~w6471;
assign w6473 = w6469 & w6472;
assign w6474 = w6469 & w36753;
assign w6475 = pi2412 & w2875;
assign w6476 = w2297 & w6475;
assign w6477 = (pi2520 & w2293) | (pi2520 & w36754) | (w2293 & w36754);
assign w6478 = w2295 & w6477;
assign w6479 = w354 & ~w6478;
assign w6480 = (pi2535 & w2314) | (pi2535 & w36755) | (w2314 & w36755);
assign w6481 = w2316 & w6480;
assign w6482 = pi2752 & w2881;
assign w6483 = ~w6481 & ~w6482;
assign w6484 = w6483 & w36756;
assign w6485 = ~w6474 & ~w6484;
assign w6486 = ~w2386 & w36757;
assign w6487 = w3754 & ~w6486;
assign w6488 = ~w6466 & w6487;
assign w6489 = ~w6452 & ~w6488;
assign w6490 = (w6489 & ~w5969) | (w6489 & w36758) | (~w5969 & w36758);
assign w6491 = ~w2657 & ~w2667;
assign w6492 = ~w2708 & ~w2713;
assign w6493 = (w6492 & w2657) | (w6492 & w36759) | (w2657 & w36759);
assign w6494 = (pi0678 & w2464) | (pi0678 & w36760) | (w2464 & w36760);
assign w6495 = (~w6494 & ~w6491) | (~w6494 & w36761) | (~w6491 & w36761);
assign w6496 = ~w6493 & w6495;
assign w6497 = ~w2826 & ~w6496;
assign w6498 = (~w2474 & w2499) | (~w2474 & w36763) | (w2499 & w36763);
assign w6499 = ~pi0514 & w6498;
assign w6500 = pi0514 & ~w6498;
assign w6501 = ~w6499 & ~w6500;
assign w6502 = pi0678 & ~w6501;
assign w6503 = ~w2465 & w6501;
assign w6504 = ~w6502 & ~w6503;
assign w6505 = w2826 & ~w6504;
assign w6506 = ~w6497 & ~w6505;
assign w6507 = w3440 & ~w6506;
assign w6508 = ~w3928 & w36764;
assign w6509 = (pi0512 & w3928) | (pi0512 & w36765) | (w3928 & w36765);
assign w6510 = ~w6508 & ~w6509;
assign w6511 = pi0677 & ~w6510;
assign w6512 = ~w2525 & w6510;
assign w6513 = ~w6511 & ~w6512;
assign w6514 = w2826 & w6513;
assign w6515 = (~w3918 & w2711) | (~w3918 & w36766) | (w2711 & w36766);
assign w6516 = pi0677 & ~w2524;
assign w6517 = ~w3919 & ~w6516;
assign w6518 = ~w6515 & w6517;
assign w6519 = ~w2826 & w6518;
assign w6520 = ~w6514 & ~w6519;
assign w6521 = w3786 & w6520;
assign w6522 = ~w6507 & ~w6521;
assign w6523 = w6490 & w6522;
assign w6524 = (w2397 & ~w2961) | (w2397 & w36767) | (~w2961 & w36767);
assign w6525 = pi2438 & w1314;
assign w6526 = ~w414 & w36768;
assign w6527 = ~w6525 & ~w6526;
assign w6528 = pi2701 & w1316;
assign w6529 = pi2275 & w1309;
assign w6530 = ~w6528 & ~w6529;
assign w6531 = w6527 & w6530;
assign w6532 = ~w371 & w36769;
assign w6533 = ~w392 & w36770;
assign w6534 = ~w6532 & ~w6533;
assign w6535 = ~w414 & w36771;
assign w6536 = ~w405 & w36772;
assign w6537 = ~w6535 & ~w6536;
assign w6538 = w6534 & w6537;
assign w6539 = (~w354 & ~w6537) | (~w354 & w36773) | (~w6537 & w36773);
assign w6540 = w6531 & ~w6539;
assign w6541 = ~w6485 & w6540;
assign w6542 = w2958 & ~w6541;
assign w6543 = w3433 & w6177;
assign w6544 = ~w6542 & ~w6543;
assign w6545 = w6524 & w6544;
assign w6546 = (w6545 & ~w6520) | (w6545 & w36774) | (~w6520 & w36774);
assign w6547 = pi0566 & ~pi0754;
assign w6548 = (~w553 & w4401) | (~w553 & w36775) | (w4401 & w36775);
assign w6549 = ~w6547 & w6548;
assign w6550 = ~pi0566 & ~pi0754;
assign w6551 = ~w6550 & ~w6548;
assign w6552 = ~w6549 & ~w6551;
assign w6553 = ~w555 & w36777;
assign w6554 = w6548 & w6553;
assign w6555 = w566 & ~w6548;
assign w6556 = ~w6554 & ~w6555;
assign w6557 = ~w6554 & w36778;
assign w6558 = w6557 & w40111;
assign w6559 = w3433 & ~w6504;
assign w6560 = ~w6484 & w36779;
assign w6561 = w2236 & w36780;
assign w6562 = (~w6561 & w6540) | (~w6561 & w36781) | (w6540 & w36781);
assign w6563 = (w2365 & ~w6562) | (w2365 & w36782) | (~w6562 & w36782);
assign w6564 = pi2415 & w941;
assign w6565 = ~w2899 & ~w6564;
assign w6566 = (w353 & w36783) | (w353 & w36784) | (w36783 & w36784);
assign w6567 = w6566 & w40102;
assign w6568 = (pi1029 & w2907) | (pi1029 & w36785) | (w2907 & w36785);
assign w6569 = ~w6568 & w36786;
assign w6570 = ~w6563 & w6569;
assign w6571 = ~pi0862 & w2899;
assign w6572 = w2961 & w36787;
assign w6573 = (~w2397 & ~w2941) | (~w2397 & w36788) | (~w2941 & w36788);
assign w6574 = ~w6572 & w6573;
assign w6575 = (w6574 & ~w2826) | (w6574 & w36789) | (~w2826 & w36789);
assign w6576 = ~w6558 & w6575;
assign w6577 = ~w2826 & w36790;
assign w6578 = ~pi0658 & w660;
assign w6579 = pi0658 & ~w660;
assign w6580 = ~w6578 & ~w6579;
assign w6581 = w667 & ~w4402;
assign w6582 = pi0636 & w4402;
assign w6583 = ~w6581 & ~w6582;
assign w6584 = w6580 & ~w6583;
assign w6585 = ~w6580 & w6583;
assign w6586 = ~w6584 & ~w6585;
assign w6587 = w6586 & w40112;
assign w6588 = (w647 & w36792) | (w647 & w36793) | (w36792 & w36793);
assign w6589 = pi0754 & w555;
assign w6590 = ~w6588 & ~w6589;
assign w6591 = ~w6587 & w6590;
assign w6592 = w797 & w36794;
assign w6593 = w2958 & w6592;
assign w6594 = ~w6577 & ~w6593;
assign w6595 = w6576 & w6594;
assign w6596 = ~w6546 & ~w6595;
assign w6597 = ~w6523 & w6596;
assign w6598 = w5959 & w6597;
assign w6599 = w4797 & w6598;
assign w6600 = w886 & w36795;
assign w6601 = w2374 & w36796;
assign w6602 = w2236 & w36797;
assign w6603 = w2354 & w36798;
assign w6604 = ~w6602 & ~w6603;
assign w6605 = ~w6601 & w6604;
assign w6606 = ~w375 & w6605;
assign w6607 = w359 & w36799;
assign w6608 = w342 & w36801;
assign w6609 = pi1422 & pi2515;
assign w6610 = (w353 & w36802) | (w353 & w36803) | (w36802 & w36803);
assign w6611 = (~w6610 & ~w342) | (~w6610 & w36804) | (~w342 & w36804);
assign w6612 = (w6611 & w2227) | (w6611 & w36805) | (w2227 & w36805);
assign w6613 = ~w828 & ~w830;
assign w6614 = ~w2897 & w6613;
assign w6615 = ~w6600 & w40113;
assign w6616 = pi1422 & pi2769;
assign w6617 = (w353 & w36810) | (w353 & w36811) | (w36810 & w36811);
assign w6618 = (~w6617 & ~w904) | (~w6617 & w36812) | (~w904 & w36812);
assign w6619 = ~w822 & ~w825;
assign w6620 = w6618 & w6619;
assign w6621 = (~w6620 & ~w886) | (~w6620 & w36813) | (~w886 & w36813);
assign w6622 = w341 & w36814;
assign w6623 = (~w6622 & ~w2261) | (~w6622 & w36815) | (~w2261 & w36815);
assign w6624 = ~w6621 & w6623;
assign w6625 = (w2227 & w36816) | (w2227 & w36817) | (w36816 & w36817);
assign w6626 = ~w3817 & ~w6625;
assign w6627 = ~w6599 & w6626;
assign w6628 = pi1452 & w1324;
assign w6629 = ~pi2978 & ~w889;
assign w6630 = ~pi2495 & w889;
assign w6631 = ~w6629 & ~w6630;
assign w6632 = (w886 & w36818) | (w886 & w36819) | (w36818 & w36819);
assign w6633 = ~w6628 & ~w6632;
assign w6634 = pi1453 & w1324;
assign w6635 = ~pi2979 & ~w889;
assign w6636 = ~pi2496 & w889;
assign w6637 = ~w6635 & ~w6636;
assign w6638 = (w886 & w36820) | (w886 & w36821) | (w36820 & w36821);
assign w6639 = ~w6634 & ~w6638;
assign w6640 = pi1455 & w1324;
assign w6641 = ~pi2981 & ~w889;
assign w6642 = ~pi2513 & w889;
assign w6643 = ~w6641 & ~w6642;
assign w6644 = (w886 & w36823) | (w886 & w36824) | (w36823 & w36824);
assign w6645 = ~w6640 & ~w6644;
assign w6646 = w3817 & w36825;
assign w6647 = pi1454 & w1324;
assign w6648 = ~pi2980 & ~w889;
assign w6649 = ~pi2497 & w889;
assign w6650 = ~w6648 & ~w6649;
assign w6651 = (w886 & w36826) | (w886 & w36827) | (w36826 & w36827);
assign w6652 = ~w6647 & ~w6651;
assign w6653 = w6652 & ~w6625;
assign w6654 = w6646 & w6653;
assign w6655 = w3817 & w36828;
assign w6656 = w6653 & w6655;
assign w6657 = ~w6652 & ~w6625;
assign w6658 = w6646 & w6657;
assign w6659 = w6655 & w6657;
assign w6660 = w3817 & w36829;
assign w6661 = w6645 & w6660;
assign w6662 = w6653 & w6661;
assign w6663 = w3817 & w36830;
assign w6664 = w6653 & w6663;
assign w6665 = w6657 & w6661;
assign w6666 = w6657 & w6663;
assign w6667 = w3817 & ~w6633;
assign w6668 = (~pi3426 & ~w341) | (~pi3426 & w35945) | (~w341 & w35945);
assign w6669 = (w341 & w35946) | (w341 & w35947) | (w35946 & w35947);
assign w6670 = (~w6621 & w6623) | (~w6621 & w36831) | (w6623 & w36831);
assign w6671 = ~w6667 & ~w6670;
assign w6672 = ~w6599 & w6671;
assign w6673 = w2352 & w2354;
assign w6674 = (~pi3390 & ~w2354) | (~pi3390 & w36832) | (~w2354 & w36832);
assign w6675 = pi3505 & ~pi3515;
assign w6676 = (pi0404 & w6675) | (pi0404 & w36833) | (w6675 & w36833);
assign w6677 = ~pi0684 & w6676;
assign w6678 = (pi0684 & w6675) | (pi0684 & w36834) | (w6675 & w36834);
assign w6679 = pi3236 & pi3547;
assign w6680 = (~w6679 & w909) | (~w6679 & w36835) | (w909 & w36835);
assign w6681 = ~w6678 & w6680;
assign w6682 = ~w6677 & w6681;
assign w6683 = w342 & w6682;
assign w6684 = w342 & w36836;
assign w6685 = w6674 & ~w6684;
assign w6686 = ~w358 & w6685;
assign w6687 = w347 & w36837;
assign w6688 = pi2489 & ~w2214;
assign w6689 = w2175 & ~w6688;
assign w6690 = ~w6688 & w36838;
assign w6691 = (w6690 & w2227) | (w6690 & w36839) | (w2227 & w36839);
assign w6692 = ~pi0684 & ~pi3481;
assign w6693 = ~pi3236 & w6692;
assign w6694 = ~pi0007 & pi3432;
assign w6695 = ~pi0005 & pi3454;
assign w6696 = ~w6694 & ~w6695;
assign w6697 = pi0006 & ~pi3453;
assign w6698 = pi0005 & ~pi3454;
assign w6699 = ~w6697 & ~w6698;
assign w6700 = w6696 & w6699;
assign w6701 = ~pi0006 & pi3453;
assign w6702 = pi0002 & ~w6701;
assign w6703 = pi0011 & ~pi3458;
assign w6704 = pi0010 & ~pi3450;
assign w6705 = ~w6703 & ~w6704;
assign w6706 = w6702 & w6705;
assign w6707 = w6700 & w6706;
assign w6708 = pi0009 & ~pi3478;
assign w6709 = ~pi0004 & pi3455;
assign w6710 = ~pi0010 & pi3450;
assign w6711 = ~w6709 & ~w6710;
assign w6712 = ~w6708 & w6711;
assign w6713 = ~pi0003 & pi3434;
assign w6714 = pi0004 & ~pi3455;
assign w6715 = ~w6713 & ~w6714;
assign w6716 = pi0007 & ~pi3432;
assign w6717 = ~pi0009 & pi3478;
assign w6718 = ~w6716 & ~w6717;
assign w6719 = w6715 & w6718;
assign w6720 = pi0003 & ~pi3434;
assign w6721 = ~pi0008 & pi3459;
assign w6722 = ~w6720 & ~w6721;
assign w6723 = pi0008 & ~pi3459;
assign w6724 = ~pi0011 & pi3458;
assign w6725 = ~w6723 & ~w6724;
assign w6726 = w6722 & w6725;
assign w6727 = w6719 & w6726;
assign w6728 = w6712 & w6727;
assign w6729 = w6707 & w6728;
assign w6730 = pi3332 & ~pi3460;
assign w6731 = pi3352 & ~pi3457;
assign w6732 = ~pi3332 & pi3460;
assign w6733 = ~w6731 & ~w6732;
assign w6734 = ~w6730 & w6733;
assign w6735 = ~pi3331 & pi3433;
assign w6736 = ~pi3347 & pi3437;
assign w6737 = ~w6735 & ~w6736;
assign w6738 = ~pi3352 & pi3457;
assign w6739 = pi3354 & ~pi3456;
assign w6740 = ~w6738 & ~w6739;
assign w6741 = w6737 & w6740;
assign w6742 = pi3331 & ~pi3433;
assign w6743 = pi3423 & ~w6742;
assign w6744 = ~pi3354 & pi3456;
assign w6745 = pi3347 & ~pi3437;
assign w6746 = ~w6744 & ~w6745;
assign w6747 = w6743 & w6746;
assign w6748 = w6741 & w6747;
assign w6749 = (pi1930 & ~w6748) | (pi1930 & w36840) | (~w6748 & w36840);
assign w6750 = pi0001 & w6749;
assign w6751 = pi0000 & w6749;
assign w6752 = ~w6750 & ~w6751;
assign w6753 = w6729 & ~w6752;
assign w6754 = ~pi1798 & pi2073;
assign w6755 = pi1798 & pi2075;
assign w6756 = pi1713 & ~w6755;
assign w6757 = ~w6754 & w6756;
assign w6758 = ~pi1713 & ~pi1798;
assign w6759 = ~pi2389 & w6758;
assign w6760 = ~pi1713 & pi1798;
assign w6761 = ~pi1998 & w6760;
assign w6762 = ~w6759 & ~w6761;
assign w6763 = ~w6757 & w6762;
assign w6764 = pi3434 & ~w6763;
assign w6765 = ~pi1798 & pi2346;
assign w6766 = pi1798 & pi2330;
assign w6767 = pi1713 & ~w6766;
assign w6768 = ~w6765 & w6767;
assign w6769 = ~pi2368 & w6758;
assign w6770 = ~pi2005 & w6760;
assign w6771 = ~w6769 & ~w6770;
assign w6772 = ~w6768 & w6771;
assign w6773 = pi3459 & ~w6772;
assign w6774 = ~w6764 & ~w6773;
assign w6775 = ~pi1798 & pi2336;
assign w6776 = pi1798 & pi1987;
assign w6777 = pi1713 & ~w6776;
assign w6778 = ~w6775 & w6777;
assign w6779 = ~pi2359 & w6758;
assign w6780 = ~pi2351 & w6760;
assign w6781 = ~w6779 & ~w6780;
assign w6782 = ~w6778 & w6781;
assign w6783 = ~pi3456 & w6782;
assign w6784 = ~pi1798 & pi2339;
assign w6785 = pi1798 & pi1991;
assign w6786 = pi1713 & ~w6785;
assign w6787 = ~w6784 & w6786;
assign w6788 = ~pi2363 & w6758;
assign w6789 = ~pi2002 & w6760;
assign w6790 = ~w6788 & ~w6789;
assign w6791 = ~w6787 & w6790;
assign w6792 = ~pi2514 & w6791;
assign w6793 = ~w6783 & ~w6792;
assign w6794 = w6774 & w6793;
assign w6795 = ~pi1798 & pi2337;
assign w6796 = pi1798 & pi1986;
assign w6797 = pi1713 & ~w6796;
assign w6798 = ~w6795 & w6797;
assign w6799 = ~pi2360 & w6758;
assign w6800 = ~pi2352 & w6760;
assign w6801 = ~w6799 & ~w6800;
assign w6802 = ~w6798 & w6801;
assign w6803 = ~pi3457 & w6802;
assign w6804 = ~pi1798 & pi2349;
assign w6805 = pi1798 & pi2333;
assign w6806 = pi1713 & ~w6805;
assign w6807 = ~w6804 & w6806;
assign w6808 = ~pi2371 & w6758;
assign w6809 = ~pi2007 & w6760;
assign w6810 = ~w6808 & ~w6809;
assign w6811 = ~w6807 & w6810;
assign w6812 = ~pi3454 & w6811;
assign w6813 = ~w6803 & ~w6812;
assign w6814 = ~pi3434 & w6763;
assign w6815 = pi3457 & ~w6802;
assign w6816 = ~w6814 & ~w6815;
assign w6817 = w6813 & w6816;
assign w6818 = w6794 & w6817;
assign w6819 = ~pi1798 & pi1996;
assign w6820 = pi1798 & pi1799;
assign w6821 = pi1713 & ~w6820;
assign w6822 = ~w6819 & w6821;
assign w6823 = ~pi2008 & w6758;
assign w6824 = ~pi1800 & w6760;
assign w6825 = ~w6823 & ~w6824;
assign w6826 = ~w6822 & w6825;
assign w6827 = pi3437 & ~w6826;
assign w6828 = ~pi1798 & pi1997;
assign w6829 = pi1798 & pi1989;
assign w6830 = pi1713 & ~w6829;
assign w6831 = ~w6828 & w6830;
assign w6832 = ~pi2009 & w6758;
assign w6833 = ~pi2000 & w6760;
assign w6834 = ~w6832 & ~w6833;
assign w6835 = ~w6831 & w6834;
assign w6836 = pi3460 & ~w6835;
assign w6837 = ~pi1798 & pi2350;
assign w6838 = pi1798 & pi2334;
assign w6839 = pi1713 & ~w6838;
assign w6840 = ~w6837 & w6839;
assign w6841 = ~pi2388 & w6760;
assign w6842 = ~pi2372 & w6758;
assign w6843 = ~w6841 & ~w6842;
assign w6844 = ~w6840 & w6843;
assign w6845 = pi3455 & ~w6844;
assign w6846 = ~w6836 & ~w6845;
assign w6847 = ~w6827 & w6846;
assign w6848 = ~pi1798 & pi2070;
assign w6849 = pi1798 & pi2077;
assign w6850 = pi1713 & ~w6849;
assign w6851 = ~w6848 & w6850;
assign w6852 = ~pi2390 & w6760;
assign w6853 = ~pi2076 & w6758;
assign w6854 = ~w6852 & ~w6853;
assign w6855 = ~w6851 & w6854;
assign w6856 = pi2472 & ~w6855;
assign w6857 = ~pi1798 & pi2347;
assign w6858 = pi1798 & pi2331;
assign w6859 = pi1713 & ~w6858;
assign w6860 = ~w6857 & w6859;
assign w6861 = ~pi2369 & w6758;
assign w6862 = ~pi2357 & w6760;
assign w6863 = ~w6861 & ~w6862;
assign w6864 = ~w6860 & w6863;
assign w6865 = ~pi3432 & w6864;
assign w6866 = ~w6856 & ~w6865;
assign w6867 = ~pi1798 & pi2341;
assign w6868 = pi1798 & pi1992;
assign w6869 = pi1713 & ~w6868;
assign w6870 = ~w6867 & w6869;
assign w6871 = ~pi2391 & w6760;
assign w6872 = ~pi2365 & w6758;
assign w6873 = ~w6871 & ~w6872;
assign w6874 = ~w6870 & w6873;
assign w6875 = ~pi2400 & w6874;
assign w6876 = ~pi1798 & pi2342;
assign w6877 = pi1798 & pi2074;
assign w6878 = pi1713 & ~w6877;
assign w6879 = ~w6876 & w6878;
assign w6880 = ~pi2355 & w6760;
assign w6881 = ~pi2072 & w6758;
assign w6882 = ~w6880 & ~w6881;
assign w6883 = ~w6879 & w6882;
assign w6884 = pi2408 & ~w6883;
assign w6885 = ~w6875 & ~w6884;
assign w6886 = w6866 & w6885;
assign w6887 = w6847 & w6886;
assign w6888 = w6818 & w6887;
assign w6889 = ~pi1798 & pi2343;
assign w6890 = pi1798 & pi1993;
assign w6891 = pi1713 & ~w6890;
assign w6892 = ~w6889 & w6891;
assign w6893 = ~pi2366 & w6758;
assign w6894 = ~pi2003 & w6760;
assign w6895 = ~w6893 & ~w6894;
assign w6896 = ~w6892 & w6895;
assign w6897 = (~pi1797 & ~w6896) | (~pi1797 & w36841) | (~w6896 & w36841);
assign w6898 = ~pi3460 & w6835;
assign w6899 = ~pi3459 & w6772;
assign w6900 = ~w6898 & ~w6899;
assign w6901 = pi2514 & ~w6791;
assign w6902 = pi3456 & ~w6782;
assign w6903 = ~w6901 & ~w6902;
assign w6904 = w6900 & w6903;
assign w6905 = w6897 & w6904;
assign w6906 = ~pi3455 & w6844;
assign w6907 = ~pi1798 & pi2071;
assign w6908 = pi1798 & pi1988;
assign w6909 = pi1713 & ~w6908;
assign w6910 = ~w6907 & w6909;
assign w6911 = ~pi2361 & w6758;
assign w6912 = ~pi1999 & w6760;
assign w6913 = ~w6911 & ~w6912;
assign w6914 = ~w6910 & w6913;
assign w6915 = pi3433 & ~w6914;
assign w6916 = ~w6906 & ~w6915;
assign w6917 = ~pi1798 & pi2348;
assign w6918 = pi1798 & pi2332;
assign w6919 = pi1713 & ~w6918;
assign w6920 = ~w6917 & w6919;
assign w6921 = ~pi2370 & w6758;
assign w6922 = ~pi2006 & w6760;
assign w6923 = ~w6921 & ~w6922;
assign w6924 = ~w6920 & w6923;
assign w6925 = pi3453 & ~w6924;
assign w6926 = ~pi3437 & w6826;
assign w6927 = ~w6925 & ~w6926;
assign w6928 = w6916 & w6927;
assign w6929 = ~pi3433 & w6914;
assign w6930 = pi2400 & ~w6874;
assign w6931 = ~w6929 & ~w6930;
assign w6932 = pi3432 & ~w6864;
assign w6933 = ~pi2408 & w6883;
assign w6934 = ~w6932 & ~w6933;
assign w6935 = w6931 & w6934;
assign w6936 = w6928 & w6935;
assign w6937 = ~pi1798 & pi2344;
assign w6938 = pi1798 & pi1994;
assign w6939 = pi1713 & ~w6938;
assign w6940 = ~w6937 & w6939;
assign w6941 = ~pi2367 & w6758;
assign w6942 = ~pi2356 & w6760;
assign w6943 = ~w6941 & ~w6942;
assign w6944 = ~w6940 & w6943;
assign w6945 = pi3450 & ~w6944;
assign w6946 = ~pi1798 & pi2345;
assign w6947 = pi1798 & pi1995;
assign w6948 = pi1713 & ~w6947;
assign w6949 = ~w6946 & w6948;
assign w6950 = ~pi2069 & w6758;
assign w6951 = ~pi2004 & w6760;
assign w6952 = ~w6950 & ~w6951;
assign w6953 = ~w6949 & w6952;
assign w6954 = ~pi3478 & w6953;
assign w6955 = ~w6945 & ~w6954;
assign w6956 = ~pi3450 & w6944;
assign w6957 = pi3478 & ~w6953;
assign w6958 = ~w6956 & ~w6957;
assign w6959 = w6955 & w6958;
assign w6960 = ~pi3453 & w6924;
assign w6961 = pi3458 & ~w6896;
assign w6962 = ~w6960 & ~w6961;
assign w6963 = pi3454 & ~w6811;
assign w6964 = ~pi2472 & w6855;
assign w6965 = ~w6963 & ~w6964;
assign w6966 = w6962 & w6965;
assign w6967 = w6959 & w6966;
assign w6968 = w6936 & w6967;
assign w6969 = w6905 & w6968;
assign w6970 = w6888 & w6969;
assign w6971 = pi0419 & ~pi0420;
assign w6972 = ~pi3641 & w6971;
assign w6973 = (pi0405 & ~w6971) | (pi0405 & w36842) | (~w6971 & w36842);
assign w6974 = w380 & w6973;
assign w6975 = w380 & w36843;
assign w6976 = pi2193 & w6975;
assign w6977 = w6969 & w36844;
assign w6978 = (w6693 & w6977) | (w6693 & w36845) | (w6977 & w36845);
assign w6979 = w2228 & w6978;
assign w6980 = (w6687 & w6979) | (w6687 & w36846) | (w6979 & w36846);
assign w6981 = ~w1052 & w6980;
assign w6982 = w909 & w6693;
assign w6983 = w6969 & w36848;
assign w6984 = ~w2227 & w36849;
assign w6985 = pi0976 & ~w1016;
assign w6986 = (w1045 & ~w1034) | (w1045 & w36850) | (~w1034 & w36850);
assign w6987 = pi1144 & w1037;
assign w6988 = pi1043 & w1036;
assign w6989 = ~w1020 & w6988;
assign w6990 = pi1242 & w1040;
assign w6991 = ~w6989 & ~w6990;
assign w6992 = ~w6987 & w6991;
assign w6993 = pi1326 & w1043;
assign w6994 = pi1214 & w1687;
assign w6995 = ~w6993 & ~w6994;
assign w6996 = pi1130 & w1409;
assign w6997 = pi1228 & w1046;
assign w6998 = ~w6996 & ~w6997;
assign w6999 = w6995 & w6998;
assign w7000 = w6992 & w6999;
assign w7001 = w7000 & w36851;
assign w7002 = w6984 & ~w7001;
assign w7003 = w6687 & w6688;
assign w7004 = pi2763 & ~w2214;
assign w7005 = w1052 & ~w7004;
assign w7006 = ~pi2376 & w7004;
assign w7007 = ~w7005 & ~w7006;
assign w7008 = w2227 & w36852;
assign w7009 = ~w6688 & w36853;
assign w7010 = pi0540 & ~w7009;
assign w7011 = pi0032 & ~pi3453;
assign w7012 = pi0031 & ~pi3454;
assign w7013 = ~w7011 & ~w7012;
assign w7014 = ~pi0036 & pi3450;
assign w7015 = pi0029 & ~pi3434;
assign w7016 = ~w7014 & ~w7015;
assign w7017 = w7013 & w7016;
assign w7018 = pi0033 & ~pi3432;
assign w7019 = pi0028 & ~w7018;
assign w7020 = pi0037 & ~pi3458;
assign w7021 = ~pi0029 & pi3434;
assign w7022 = ~w7020 & ~w7021;
assign w7023 = w7019 & w7022;
assign w7024 = w7017 & w7023;
assign w7025 = ~pi0032 & pi3453;
assign w7026 = ~pi0031 & pi3454;
assign w7027 = pi0036 & ~pi3450;
assign w7028 = ~w7026 & ~w7027;
assign w7029 = ~w7025 & w7028;
assign w7030 = ~pi0033 & pi3432;
assign w7031 = pi0030 & ~pi3455;
assign w7032 = ~w7030 & ~w7031;
assign w7033 = ~pi0030 & pi3455;
assign w7034 = pi0035 & ~pi3478;
assign w7035 = ~w7033 & ~w7034;
assign w7036 = w7032 & w7035;
assign w7037 = ~pi0037 & pi3458;
assign w7038 = ~pi0034 & pi3459;
assign w7039 = ~w7037 & ~w7038;
assign w7040 = pi0034 & ~pi3459;
assign w7041 = ~pi0035 & pi3478;
assign w7042 = ~w7040 & ~w7041;
assign w7043 = w7039 & w7042;
assign w7044 = w7036 & w7043;
assign w7045 = w7029 & w7044;
assign w7046 = w7024 & w7045;
assign w7047 = pi0012 & w6749;
assign w7048 = pi0013 & w6749;
assign w7049 = ~w7047 & ~w7048;
assign w7050 = w7046 & ~w7049;
assign w7051 = ~w6753 & ~w7050;
assign w7052 = w6982 & w7051;
assign w7053 = ~w6970 & w36854;
assign w7054 = pi3437 & pi3460;
assign w7055 = pi3433 & w7054;
assign w7056 = w7054 & w36855;
assign w7057 = pi3456 & w7056;
assign w7058 = w7056 & w36856;
assign w7059 = w7056 & w36857;
assign w7060 = pi3454 & w7059;
assign w7061 = w7059 & w36858;
assign w7062 = w7059 & w36859;
assign w7063 = w7059 & w36860;
assign w7064 = pi3478 & w7063;
assign w7065 = w7063 & w36861;
assign w7066 = (~pi3450 & ~w7063) | (~pi3450 & w36862) | (~w7063 & w36862);
assign w7067 = ~w7065 & ~w7066;
assign w7068 = pi3236 & w6687;
assign w7069 = w6687 & w36864;
assign w7070 = (~w7069 & w2227) | (~w7069 & w36865) | (w2227 & w36865);
assign w7071 = ~w7008 & w7070;
assign w7072 = ~w7002 & w7071;
assign w7073 = ~w2227 & w36866;
assign w7074 = pi0026 & w7073;
assign w7075 = ~w6688 & ~w6690;
assign w7076 = w2227 & w7075;
assign w7077 = ~pi3481 & w40114;
assign w7078 = pi3400 & pi3403;
assign w7079 = pi3402 & w7078;
assign w7080 = w7078 & w36869;
assign w7081 = pi3414 & w7080;
assign w7082 = w7080 & w36870;
assign w7083 = w7080 & w36871;
assign w7084 = pi3406 & w7083;
assign w7085 = w7083 & w36872;
assign w7086 = w7083 & w36873;
assign w7087 = w7083 & w36874;
assign w7088 = pi3422 & w7087;
assign w7089 = w7087 & w36875;
assign w7090 = (~pi3421 & ~w7087) | (~pi3421 & w36876) | (~w7087 & w36876);
assign w7091 = ~w7089 & ~w7090;
assign w7092 = (w7076 & w36877) | (w7076 & w36878) | (w36877 & w36878);
assign w7093 = ~w7074 & ~w7092;
assign w7094 = w7072 & w7093;
assign w7095 = ~w6981 & w7094;
assign w7096 = pi0779 & w889;
assign w7097 = ~w939 & ~w7096;
assign w7098 = ~w350 & w36879;
assign w7099 = (pi0405 & ~w342) | (pi0405 & w36880) | (~w342 & w36880);
assign w7100 = w342 & w36881;
assign w7101 = ~w7099 & ~w7100;
assign w7102 = ~w6674 & w7101;
assign w7103 = ~pi3450 & w6674;
assign w7104 = ~w6685 & w36882;
assign w7105 = ~w7102 & w7104;
assign w7106 = ~w7098 & ~w7105;
assign w7107 = (w7106 & w7095) | (w7106 & w36883) | (w7095 & w36883);
assign w7108 = pi3680 & ~w7107;
assign w7109 = ~w1422 & w6980;
assign w7110 = ~w2227 & w36884;
assign w7111 = (~pi3458 & ~w7063) | (~pi3458 & w36885) | (~w7063 & w36885);
assign w7112 = w7063 & w36886;
assign w7113 = ~w7111 & ~w7112;
assign w7114 = ~w2227 & w36887;
assign w7115 = w1422 & ~w7004;
assign w7116 = ~pi2375 & w7004;
assign w7117 = ~w7115 & ~w7116;
assign w7118 = w6687 & w36889;
assign w7119 = (~w7118 & ~w2227) | (~w7118 & w36890) | (~w2227 & w36890);
assign w7120 = ~w7114 & w7119;
assign w7121 = ~w7110 & w7120;
assign w7122 = pi1157 & w1382;
assign w7123 = pi1255 & w1661;
assign w7124 = pi1171 & w1388;
assign w7125 = ~w7123 & ~w7124;
assign w7126 = pi1311 & w1659;
assign w7127 = pi1297 & w1678;
assign w7128 = ~w7126 & ~w7127;
assign w7129 = w7125 & w7128;
assign w7130 = ~w7122 & w7129;
assign w7131 = (w1030 & ~w1398) | (w1030 & w36891) | (~w1398 & w36891);
assign w7132 = pi1213 & w1687;
assign w7133 = pi1199 & w1385;
assign w7134 = ~w7132 & ~w7133;
assign w7135 = pi1241 & w1040;
assign w7136 = pi1185 & w1411;
assign w7137 = ~w7135 & ~w7136;
assign w7138 = w7134 & w7137;
assign w7139 = pi1143 & w1037;
assign w7140 = pi1269 & w1414;
assign w7141 = ~w7139 & ~w7140;
assign w7142 = pi1227 & w1046;
assign w7143 = pi1115 & w1416;
assign w7144 = ~w7142 & ~w7143;
assign w7145 = w7141 & w7144;
assign w7146 = w7138 & w7145;
assign w7147 = ~w7131 & w7146;
assign w7148 = w7130 & w7147;
assign w7149 = ~w2227 & w36892;
assign w7150 = w7087 & w36893;
assign w7151 = (~pi3430 & ~w7087) | (~pi3430 & w36894) | (~w7087 & w36894);
assign w7152 = ~w7150 & ~w7151;
assign w7153 = (w7076 & w36895) | (w7076 & w36896) | (w36895 & w36896);
assign w7154 = ~w7149 & ~w7153;
assign w7155 = w7121 & w7154;
assign w7156 = ~w7109 & w7155;
assign w7157 = pi0752 & w889;
assign w7158 = ~w1642 & ~w7157;
assign w7159 = ~w350 & w36897;
assign w7160 = (pi0421 & ~w342) | (pi0421 & w36898) | (~w342 & w36898);
assign w7161 = w342 & w36899;
assign w7162 = ~w7160 & ~w7161;
assign w7163 = ~w6674 & w7162;
assign w7164 = ~pi3458 & w6674;
assign w7165 = ~w6685 & w36900;
assign w7166 = ~w7163 & w7165;
assign w7167 = ~w7159 & ~w7166;
assign w7168 = (w7167 & w7156) | (w7167 & w36901) | (w7156 & w36901);
assign w7169 = pi3523 & ~w338;
assign w7170 = ~pi3547 & ~w6675;
assign w7171 = pi3190 & w327;
assign w7172 = ~w7170 & w7171;
assign w7173 = ~w7169 & ~w7172;
assign w7174 = w6682 & w7173;
assign w7175 = w930 & w36902;
assign w7176 = w887 & w7175;
assign w7177 = pi3586 & pi3591;
assign w7178 = ~w889 & ~w7177;
assign w7179 = w7178 & w36903;
assign w7180 = (~pi3682 & w7173) | (~pi3682 & w36904) | (w7173 & w36904);
assign w7181 = ~w7179 & w7180;
assign w7182 = ~w7176 & w7181;
assign w7183 = (w7156 & w36905) | (w7156 & w36906) | (w36905 & w36906);
assign w7184 = ~w7108 & w7183;
assign w7185 = ~pi1456 & w1324;
assign w7186 = pi2472 & ~w889;
assign w7187 = pi2498 & w889;
assign w7188 = ~w7186 & ~w7187;
assign w7189 = (w886 & w36907) | (w886 & w36908) | (w36907 & w36908);
assign w7190 = ~w7185 & ~w7189;
assign w7191 = pi1458 & w1324;
assign w7192 = ~pi2400 & ~w889;
assign w7193 = ~pi2499 & w889;
assign w7194 = ~w7192 & ~w7193;
assign w7195 = (w886 & w36909) | (w886 & w36910) | (w36909 & w36910);
assign w7196 = ~w7191 & ~w7195;
assign w7197 = w7182 & w36911;
assign w7198 = pi1461 & w1324;
assign w7199 = ~pi2408 & ~w889;
assign w7200 = ~pi2502 & w889;
assign w7201 = ~w7199 & ~w7200;
assign w7202 = (w886 & w36912) | (w886 & w36913) | (w36912 & w36913);
assign w7203 = ~w7198 & ~w7202;
assign w7204 = w7197 & w7203;
assign w7205 = w7107 & ~w7168;
assign w7206 = ~pi3680 & w7205;
assign w7207 = ~w7107 & w7168;
assign w7208 = pi3680 & w7207;
assign w7209 = ~w7206 & ~w7208;
assign w7210 = ~pi1457 & w1324;
assign w7211 = pi2514 & ~w889;
assign w7212 = pi2512 & w889;
assign w7213 = ~w7211 & ~w7212;
assign w7214 = (w886 & w36914) | (w886 & w36915) | (w36914 & w36915);
assign w7215 = ~w7210 & ~w7214;
assign w7216 = ~w7209 & ~w7215;
assign w7217 = w7204 & w7216;
assign w7218 = w7197 & ~w7203;
assign w7219 = w7216 & w7218;
assign w7220 = w7182 & w36916;
assign w7221 = w7203 & w7220;
assign w7222 = w7216 & w7221;
assign w7223 = ~w7203 & w7220;
assign w7224 = w7216 & w7223;
assign w7225 = ~w7209 & w7215;
assign w7226 = w7204 & w7225;
assign w7227 = w7218 & w7225;
assign w7228 = w7221 & w7225;
assign w7229 = w7223 & w7225;
assign w7230 = (~pi1422 & w2248) | (~pi1422 & w36917) | (w2248 & w36917);
assign w7231 = w7230 & w40097;
assign w7232 = pi1840 & ~w891;
assign w7233 = w895 & w7232;
assign w7234 = w904 & w7233;
assign w7235 = (w7234 & ~w886) | (w7234 & w36918) | (~w886 & w36918);
assign w7236 = ~w7231 & ~w7235;
assign w7237 = w7173 & ~w7236;
assign w7238 = (w6673 & ~w342) | (w6673 & w36919) | (~w342 & w36919);
assign w7239 = (pi0418 & w7169) | (pi0418 & w36920) | (w7169 & w36920);
assign w7240 = w7239 & w7238;
assign w7241 = ~w7237 & ~w7240;
assign w7242 = (w178 & w36921) | (w178 & w36922) | (w36921 & w36922);
assign w7243 = (w178 & w36923) | (w178 & w36924) | (w36923 & w36924);
assign w7244 = w110 & w36926;
assign w7245 = (~pi3496 & ~w110) | (~pi3496 & w36927) | (~w110 & w36927);
assign w7246 = pi3350 & ~w7245;
assign w7247 = ~w7244 & w7246;
assign w7248 = ~w7247 & w40115;
assign w7249 = ~w7243 & w7248;
assign w7250 = (pi3626 & ~w7249) | (pi3626 & w36928) | (~w7249 & w36928);
assign w7251 = pi2059 & ~pi3626;
assign w7252 = ~w7250 & ~w7251;
assign w7253 = (w178 & w36929) | (w178 & w36930) | (w36929 & w36930);
assign w7254 = (w178 & w36931) | (w178 & w36932) | (w36931 & w36932);
assign w7255 = (~pi3497 & ~w110) | (~pi3497 & w36934) | (~w110 & w36934);
assign w7256 = w110 & w36935;
assign w7257 = pi3350 & ~w7256;
assign w7258 = ~w7255 & w7257;
assign w7259 = ~w7258 & w40116;
assign w7260 = ~w7254 & w7259;
assign w7261 = (pi3626 & ~w7260) | (pi3626 & w36936) | (~w7260 & w36936);
assign w7262 = pi2061 & ~pi3626;
assign w7263 = ~w7261 & ~w7262;
assign w7264 = (w178 & w36937) | (w178 & w36938) | (w36937 & w36938);
assign w7265 = (w178 & w36939) | (w178 & w36940) | (w36939 & w36940);
assign w7266 = w110 & w36942;
assign w7267 = (~pi3495 & ~w110) | (~pi3495 & w36943) | (~w110 & w36943);
assign w7268 = pi3350 & ~w7267;
assign w7269 = ~w7266 & w7268;
assign w7270 = ~w7269 & w40117;
assign w7271 = ~w7265 & w7270;
assign w7272 = (pi3626 & ~w7271) | (pi3626 & w36944) | (~w7271 & w36944);
assign w7273 = pi2058 & ~pi3626;
assign w7274 = ~w7272 & ~w7273;
assign w7275 = (w178 & w36945) | (w178 & w36946) | (w36945 & w36946);
assign w7276 = (w178 & w36947) | (w178 & w36948) | (w36947 & w36948);
assign w7277 = w110 & w36950;
assign w7278 = (~pi3500 & ~w110) | (~pi3500 & w36951) | (~w110 & w36951);
assign w7279 = pi3350 & ~w7278;
assign w7280 = ~w7277 & w7279;
assign w7281 = ~w7280 & w40118;
assign w7282 = ~w7276 & w7281;
assign w7283 = (pi3626 & ~w7282) | (pi3626 & w36952) | (~w7282 & w36952);
assign w7284 = pi1841 & ~pi3626;
assign w7285 = ~w7283 & ~w7284;
assign w7286 = (w178 & w36953) | (w178 & w36954) | (w36953 & w36954);
assign w7287 = (w178 & w36955) | (w178 & w36956) | (w36955 & w36956);
assign w7288 = w110 & w36958;
assign w7289 = (~pi3499 & ~w110) | (~pi3499 & w36959) | (~w110 & w36959);
assign w7290 = pi3350 & ~w7289;
assign w7291 = ~w7288 & w7290;
assign w7292 = ~w7291 & w40119;
assign w7293 = ~w7287 & w7292;
assign w7294 = (pi3626 & ~w7293) | (pi3626 & w36960) | (~w7293 & w36960);
assign w7295 = pi1467 & ~pi3626;
assign w7296 = ~w7294 & ~w7295;
assign w7297 = (w178 & w36961) | (w178 & w36962) | (w36961 & w36962);
assign w7298 = (w178 & w36963) | (w178 & w36964) | (w36963 & w36964);
assign w7299 = w110 & w36966;
assign w7300 = (~pi3503 & ~w110) | (~pi3503 & w36967) | (~w110 & w36967);
assign w7301 = pi3350 & ~w7300;
assign w7302 = ~w7299 & w7301;
assign w7303 = ~w7302 & w40120;
assign w7304 = ~w7298 & w7303;
assign w7305 = (pi3626 & ~w7304) | (pi3626 & w36968) | (~w7304 & w36968);
assign w7306 = pi1603 & ~pi3626;
assign w7307 = ~w7305 & ~w7306;
assign w7308 = (w178 & w36969) | (w178 & w36970) | (w36969 & w36970);
assign w7309 = (w178 & w36971) | (w178 & w36972) | (w36971 & w36972);
assign w7310 = (~pi3489 & ~w110) | (~pi3489 & w36974) | (~w110 & w36974);
assign w7311 = w110 & w36975;
assign w7312 = pi3350 & ~w7311;
assign w7313 = ~w7310 & w7312;
assign w7314 = ~w7313 & w40121;
assign w7315 = ~w7309 & w7314;
assign w7316 = (pi3626 & ~w7315) | (pi3626 & w36976) | (~w7315 & w36976);
assign w7317 = pi1474 & ~pi3626;
assign w7318 = ~w7316 & ~w7317;
assign w7319 = (w178 & w36977) | (w178 & w36978) | (w36977 & w36978);
assign w7320 = (w178 & w36979) | (w178 & w36980) | (w36979 & w36980);
assign w7321 = (~pi3492 & ~w110) | (~pi3492 & w36982) | (~w110 & w36982);
assign w7322 = w110 & w36983;
assign w7323 = pi3350 & ~w7322;
assign w7324 = ~w7321 & w7323;
assign w7325 = ~w7324 & w40122;
assign w7326 = ~w7320 & w7325;
assign w7327 = (pi3626 & ~w7326) | (pi3626 & w36984) | (~w7326 & w36984);
assign w7328 = pi1602 & ~pi3626;
assign w7329 = ~w7327 & ~w7328;
assign w7330 = (w178 & w36985) | (w178 & w36986) | (w36985 & w36986);
assign w7331 = (w178 & w36987) | (w178 & w36988) | (w36987 & w36988);
assign w7332 = pi3350 & pi3501;
assign w7333 = ~w7332 & w40123;
assign w7334 = ~w7331 & w7333;
assign w7335 = (pi3626 & ~w7334) | (pi3626 & w36990) | (~w7334 & w36990);
assign w7336 = pi0928 & ~pi3626;
assign w7337 = ~w7335 & ~w7336;
assign w7338 = (w178 & w36991) | (w178 & w36992) | (w36991 & w36992);
assign w7339 = (w178 & w36993) | (w178 & w36994) | (w36993 & w36994);
assign w7340 = pi3350 & pi3491;
assign w7341 = ~w7340 & w40124;
assign w7342 = ~w7339 & w7341;
assign w7343 = (pi3626 & ~w7342) | (pi3626 & w36996) | (~w7342 & w36996);
assign w7344 = pi1066 & ~pi3626;
assign w7345 = ~w7343 & ~w7344;
assign w7346 = (w178 & w36997) | (w178 & w36998) | (w36997 & w36998);
assign w7347 = (w178 & w36999) | (w178 & w37000) | (w36999 & w37000);
assign w7348 = pi3350 & pi3494;
assign w7349 = ~w7348 & w40125;
assign w7350 = ~w7347 & w7349;
assign w7351 = (pi3626 & ~w7350) | (pi3626 & w37002) | (~w7350 & w37002);
assign w7352 = pi1090 & ~pi3626;
assign w7353 = ~w7351 & ~w7352;
assign w7354 = (w178 & w37003) | (w178 & w37004) | (w37003 & w37004);
assign w7355 = pi3350 & pi3498;
assign w7356 = ~w7355 & w40126;
assign w7357 = ~w7354 & w7356;
assign w7358 = pi3626 & ~w7357;
assign w7359 = pi0930 & ~pi3626;
assign w7360 = ~w7358 & ~w7359;
assign w7361 = pi2400 & pi2514;
assign w7362 = ~pi2472 & ~w7361;
assign w7363 = (w7205 & w37007) | (w7205 & w37008) | (w37007 & w37008);
assign w7364 = ~pi2400 & ~pi2514;
assign w7365 = (~pi3449 & w7364) | (~pi3449 & w37009) | (w7364 & w37009);
assign w7366 = ~pi2408 & ~pi2472;
assign w7367 = ~w7365 & w7366;
assign w7368 = w7207 & w7367;
assign w7369 = ~w7363 & ~w7368;
assign w7370 = pi3350 & pi3626;
assign w7371 = (w7370 & ~w7205) | (w7370 & w37011) | (~w7205 & w37011);
assign w7372 = ~w7369 & w7371;
assign w7373 = pi0688 & ~pi3626;
assign w7374 = (w178 & w37012) | (w178 & w37013) | (w37012 & w37013);
assign w7375 = ~pi2405 & ~pi3680;
assign w7376 = ~pi2529 & pi3680;
assign w7377 = ~w7375 & ~w7376;
assign w7378 = (w7377 & w184) | (w7377 & w37014) | (w184 & w37014);
assign w7379 = ~w7374 & ~w7378;
assign w7380 = (~w7373 & w7379) | (~w7373 & w37015) | (w7379 & w37015);
assign w7381 = ~w7372 & w7380;
assign w7382 = ~pi0929 & ~pi3626;
assign w7383 = ~pi2472 & pi3350;
assign w7384 = pi2400 & pi2408;
assign w7385 = ~pi2400 & ~pi2408;
assign w7386 = ~w7384 & ~w7385;
assign w7387 = w7207 & w37016;
assign w7388 = w7205 & w37017;
assign w7389 = ~w7387 & ~w7388;
assign w7390 = (w178 & w37018) | (w178 & w37019) | (w37018 & w37019);
assign w7391 = ~pi2404 & ~pi3680;
assign w7392 = ~pi2405 & pi3680;
assign w7393 = ~w7391 & ~w7392;
assign w7394 = pi3626 & w40127;
assign w7395 = ~w7390 & w7394;
assign w7396 = (w7395 & w7389) | (w7395 & w37021) | (w7389 & w37021);
assign w7397 = ~w7382 & ~w7396;
assign w7398 = pi2980 & w181;
assign w7399 = ~pi2473 & ~pi3680;
assign w7400 = ~pi2404 & pi3680;
assign w7401 = ~w7399 & ~w7400;
assign w7402 = pi3626 & w40128;
assign w7403 = ~w7398 & w37024;
assign w7404 = (w7403 & ~w7205) | (w7403 & w37025) | (~w7205 & w37025);
assign w7405 = pi2514 & w7384;
assign w7406 = ~pi2514 & ~w7384;
assign w7407 = w7383 & ~w7406;
assign w7408 = ~w7405 & w7407;
assign w7409 = w7207 & w7408;
assign w7410 = pi3350 & ~pi3680;
assign w7411 = ~w7398 & w37026;
assign w7412 = ~pi3101 & ~pi3626;
assign w7413 = (~w7412 & w7409) | (~w7412 & w37027) | (w7409 & w37027);
assign w7414 = ~w7404 & w7413;
assign w7415 = pi0942 & w203;
assign w7416 = pi3625 & ~w183;
assign w7417 = (pi3624 & w184) | (pi3624 & w37028) | (w184 & w37028);
assign w7418 = (~w7417 & w183) | (~w7417 & w37029) | (w183 & w37029);
assign w7419 = pi0393 & w7418;
assign w7420 = pi0523 & ~w3644;
assign w7421 = (pi0574 & ~w3609) | (pi0574 & w37030) | (~w3609 & w37030);
assign w7422 = pi0537 & ~w3584;
assign w7423 = ~w7421 & ~w7422;
assign w7424 = (~w941 & ~w7423) | (~w941 & w37031) | (~w7423 & w37031);
assign w7425 = pi2121 & pi2419;
assign w7426 = ~pi3380 & ~pi3381;
assign w7427 = ~pi3383 & ~pi3384;
assign w7428 = w7426 & w7427;
assign w7429 = ~pi3369 & ~pi3379;
assign w7430 = ~pi3366 & ~pi3368;
assign w7431 = w7429 & w7430;
assign w7432 = w7428 & w7431;
assign w7433 = ~w7425 & w7432;
assign w7434 = w7427 & w7431;
assign w7435 = pi3380 & ~pi3381;
assign w7436 = w7431 & w37033;
assign w7437 = pi3366 & ~pi3368;
assign w7438 = w7428 & w37034;
assign w7439 = ~pi3380 & pi3381;
assign w7440 = w7431 & w37035;
assign w7441 = ~w7438 & ~w7440;
assign w7442 = ~w7436 & w7441;
assign w7443 = ~pi3366 & pi3368;
assign w7444 = w7428 & w37036;
assign w7445 = pi3383 & ~pi3384;
assign w7446 = w7426 & w7445;
assign w7447 = w7431 & w7446;
assign w7448 = ~w7444 & ~w7447;
assign w7449 = ~pi3369 & pi3379;
assign w7450 = w7428 & w37037;
assign w7451 = pi3369 & ~pi3379;
assign w7452 = w7428 & w37038;
assign w7453 = ~w7450 & ~w7452;
assign w7454 = w7448 & w7453;
assign w7455 = w7442 & w7454;
assign w7456 = pi3715 & w7455;
assign w7457 = pi3779 & w7444;
assign w7458 = pi3747 & w7447;
assign w7459 = ~pi3381 & pi3811;
assign w7460 = pi3380 & ~w7459;
assign w7461 = pi3381 & ~pi3795;
assign w7462 = ~w7460 & ~w7461;
assign w7463 = w7434 & w7462;
assign w7464 = ~w7458 & ~w7463;
assign w7465 = ~w7457 & w7464;
assign w7466 = pi3763 & w7452;
assign w7467 = pi3827 & w7450;
assign w7468 = pi3731 & w7438;
assign w7469 = ~w7467 & ~w7468;
assign w7470 = ~w7466 & w7469;
assign w7471 = w7465 & w7470;
assign w7472 = ~w7456 & w7471;
assign w7473 = (w7424 & w37039) | (w7424 & w37040) | (w37039 & w37040);
assign w7474 = w7417 & w7473;
assign w7475 = (~w7474 & ~w7416) | (~w7474 & w37041) | (~w7416 & w37041);
assign w7476 = ~w7419 & w7475;
assign w7477 = w201 & ~w7476;
assign w7478 = ~w7415 & ~w7477;
assign w7479 = pi0927 & w203;
assign w7480 = pi0390 & w7418;
assign w7481 = pi3716 & w7455;
assign w7482 = pi3732 & w7438;
assign w7483 = pi3828 & w7450;
assign w7484 = pi3812 & w7436;
assign w7485 = ~w7483 & ~w7484;
assign w7486 = ~w7482 & w7485;
assign w7487 = pi3764 & w7452;
assign w7488 = pi3748 & w7447;
assign w7489 = ~w7432 & ~w7488;
assign w7490 = ~w7487 & w7489;
assign w7491 = pi3796 & w7440;
assign w7492 = pi3780 & w7444;
assign w7493 = ~w7491 & ~w7492;
assign w7494 = w7490 & w7493;
assign w7495 = w7486 & w7494;
assign w7496 = ~w7481 & w7495;
assign w7497 = (pi0537 & ~w4677) | (pi0537 & w37042) | (~w4677 & w37042);
assign w7498 = pi0574 & ~w4738;
assign w7499 = pi0523 & ~w4712;
assign w7500 = ~w7498 & ~w7499;
assign w7501 = (~w941 & ~w7500) | (~w941 & w37043) | (~w7500 & w37043);
assign w7502 = pi2120 & pi2419;
assign w7503 = w7432 & ~w7502;
assign w7504 = (w7503 & ~w7501) | (w7503 & w37044) | (~w7501 & w37044);
assign w7505 = ~w7496 & ~w7504;
assign w7506 = (w184 & w37045) | (w184 & w37046) | (w37045 & w37046);
assign w7507 = (~w7506 & ~w7416) | (~w7506 & w37047) | (~w7416 & w37047);
assign w7508 = ~w7480 & w7507;
assign w7509 = w201 & ~w7508;
assign w7510 = ~w7479 & ~w7509;
assign w7511 = pi0926 & w203;
assign w7512 = pi0389 & w7418;
assign w7513 = pi3717 & w7455;
assign w7514 = pi3829 & w7450;
assign w7515 = pi3733 & w7438;
assign w7516 = pi3813 & w7436;
assign w7517 = ~w7515 & ~w7516;
assign w7518 = ~w7514 & w7517;
assign w7519 = pi3765 & w7452;
assign w7520 = pi3749 & w7447;
assign w7521 = ~w7432 & ~w7520;
assign w7522 = ~w7519 & w7521;
assign w7523 = pi3797 & w7440;
assign w7524 = pi3781 & w7444;
assign w7525 = ~w7523 & ~w7524;
assign w7526 = w7522 & w7525;
assign w7527 = w7518 & w7526;
assign w7528 = ~w7513 & w7527;
assign w7529 = (pi0537 & ~w5774) | (pi0537 & w37048) | (~w5774 & w37048);
assign w7530 = pi0523 & ~w5726;
assign w7531 = (pi0574 & ~w5799) | (pi0574 & w37049) | (~w5799 & w37049);
assign w7532 = ~w7530 & w37050;
assign w7533 = ~w941 & ~w7532;
assign w7534 = pi2119 & pi2419;
assign w7535 = w7432 & ~w7534;
assign w7536 = (w7535 & w7532) | (w7535 & w37052) | (w7532 & w37052);
assign w7537 = ~w7528 & ~w7536;
assign w7538 = (w184 & w37053) | (w184 & w37054) | (w37053 & w37054);
assign w7539 = ~w183 & w37055;
assign w7540 = ~w7538 & ~w7539;
assign w7541 = ~w7512 & w7540;
assign w7542 = w201 & ~w7541;
assign w7543 = ~w7511 & ~w7542;
assign w7544 = pi0925 & w203;
assign w7545 = pi0388 & w7418;
assign w7546 = pi3718 & w7455;
assign w7547 = pi3766 & w7452;
assign w7548 = pi3830 & w7450;
assign w7549 = pi3734 & w7438;
assign w7550 = ~w7548 & ~w7549;
assign w7551 = ~w7547 & w7550;
assign w7552 = pi3814 & w7436;
assign w7553 = pi3750 & w7447;
assign w7554 = ~w7432 & ~w7553;
assign w7555 = ~w7552 & w7554;
assign w7556 = pi3798 & w7440;
assign w7557 = pi3782 & w7444;
assign w7558 = ~w7556 & ~w7557;
assign w7559 = w7555 & w7558;
assign w7560 = w7551 & w7559;
assign w7561 = ~w7546 & w7560;
assign w7562 = (pi0537 & ~w5220) | (pi0537 & w37056) | (~w5220 & w37056);
assign w7563 = pi0574 & ~w5196;
assign w7564 = pi0523 & ~w5146;
assign w7565 = ~w7563 & ~w7564;
assign w7566 = (~w941 & ~w7565) | (~w941 & w37057) | (~w7565 & w37057);
assign w7567 = pi2118 & pi2419;
assign w7568 = w7432 & ~w7567;
assign w7569 = (w7568 & ~w7566) | (w7568 & w37058) | (~w7566 & w37058);
assign w7570 = ~w7561 & ~w7569;
assign w7571 = (w184 & w37059) | (w184 & w37060) | (w37059 & w37060);
assign w7572 = (~w7571 & ~w7416) | (~w7571 & w37061) | (~w7416 & w37061);
assign w7573 = ~w7545 & w7572;
assign w7574 = w201 & ~w7573;
assign w7575 = ~w7544 & ~w7574;
assign w7576 = pi0943 & w203;
assign w7577 = pi0387 & w7418;
assign w7578 = pi3719 & w7455;
assign w7579 = pi3799 & w7440;
assign w7580 = pi3831 & w7450;
assign w7581 = pi3815 & w7436;
assign w7582 = ~w7580 & ~w7581;
assign w7583 = ~w7579 & w7582;
assign w7584 = pi3783 & w7444;
assign w7585 = pi3751 & w7447;
assign w7586 = ~w7432 & ~w7585;
assign w7587 = ~w7584 & w7586;
assign w7588 = pi3735 & w7438;
assign w7589 = pi3767 & w7452;
assign w7590 = ~w7588 & ~w7589;
assign w7591 = w7587 & w7590;
assign w7592 = w7583 & w7591;
assign w7593 = ~w7578 & w7592;
assign w7594 = (pi0574 & ~w4314) | (pi0574 & w37062) | (~w4314 & w37062);
assign w7595 = pi0537 & ~w4335;
assign w7596 = pi0523 & ~w4370;
assign w7597 = ~w7595 & ~w7596;
assign w7598 = (~w941 & ~w7597) | (~w941 & w37063) | (~w7597 & w37063);
assign w7599 = pi2117 & pi2419;
assign w7600 = w7432 & ~w7599;
assign w7601 = (w7600 & ~w7598) | (w7600 & w37064) | (~w7598 & w37064);
assign w7602 = ~w7593 & ~w7601;
assign w7603 = (w184 & w37065) | (w184 & w37066) | (w37065 & w37066);
assign w7604 = (~w7603 & ~w7416) | (~w7603 & w37067) | (~w7416 & w37067);
assign w7605 = ~w7577 & w7604;
assign w7606 = w201 & ~w7605;
assign w7607 = ~w7576 & ~w7606;
assign w7608 = pi0924 & w203;
assign w7609 = pi0386 & w7418;
assign w7610 = ~w183 & w37068;
assign w7611 = pi3720 & w7455;
assign w7612 = pi3800 & w7440;
assign w7613 = pi3768 & w7452;
assign w7614 = pi3816 & w7436;
assign w7615 = ~w7613 & ~w7614;
assign w7616 = ~w7612 & w7615;
assign w7617 = pi3784 & w7444;
assign w7618 = pi3752 & w7447;
assign w7619 = ~w7432 & ~w7618;
assign w7620 = ~w7617 & w7619;
assign w7621 = pi3832 & w7450;
assign w7622 = pi3736 & w7438;
assign w7623 = ~w7621 & ~w7622;
assign w7624 = w7620 & w7623;
assign w7625 = w7616 & w7624;
assign w7626 = ~w7611 & w7625;
assign w7627 = pi0523 & ~w6347;
assign w7628 = (pi0574 & ~w6291) | (pi0574 & w37069) | (~w6291 & w37069);
assign w7629 = pi0537 & ~w6312;
assign w7630 = ~w7628 & ~w7629;
assign w7631 = (~w941 & ~w7630) | (~w941 & w37070) | (~w7630 & w37070);
assign w7632 = pi2078 & pi2419;
assign w7633 = w7432 & ~w7632;
assign w7634 = (w7633 & ~w7631) | (w7633 & w37071) | (~w7631 & w37071);
assign w7635 = ~w7626 & ~w7634;
assign w7636 = (w184 & w37072) | (w184 & w37073) | (w37072 & w37073);
assign w7637 = ~w7610 & ~w7636;
assign w7638 = ~w7609 & w7637;
assign w7639 = w201 & ~w7638;
assign w7640 = ~w7608 & ~w7639;
assign w7641 = pi0923 & w203;
assign w7642 = pi0385 & w7418;
assign w7643 = ~w183 & w37074;
assign w7644 = pi3721 & w7455;
assign w7645 = pi3801 & w7440;
assign w7646 = pi3769 & w7452;
assign w7647 = pi3817 & w7436;
assign w7648 = ~w7646 & ~w7647;
assign w7649 = ~w7645 & w7648;
assign w7650 = pi3785 & w7444;
assign w7651 = pi3753 & w7447;
assign w7652 = ~w7432 & ~w7651;
assign w7653 = ~w7650 & w7652;
assign w7654 = pi3833 & w7450;
assign w7655 = pi3737 & w7438;
assign w7656 = ~w7654 & ~w7655;
assign w7657 = w7653 & w7656;
assign w7658 = w7649 & w7657;
assign w7659 = ~w7644 & w7658;
assign w7660 = pi0523 & ~w3358;
assign w7661 = (pi0574 & ~w3383) | (pi0574 & w37075) | (~w3383 & w37075);
assign w7662 = pi0537 & ~w3404;
assign w7663 = ~w7661 & ~w7662;
assign w7664 = (~w941 & ~w7663) | (~w941 & w37076) | (~w7663 & w37076);
assign w7665 = pi2116 & pi2419;
assign w7666 = w7432 & ~w7665;
assign w7667 = (w7666 & ~w7664) | (w7666 & w37077) | (~w7664 & w37077);
assign w7668 = ~w7659 & ~w7667;
assign w7669 = (w184 & w37078) | (w184 & w37079) | (w37078 & w37079);
assign w7670 = ~w7643 & ~w7669;
assign w7671 = ~w7642 & w7670;
assign w7672 = w201 & ~w7671;
assign w7673 = ~w7641 & ~w7672;
assign w7674 = pi0922 & w203;
assign w7675 = pi0384 & w7418;
assign w7676 = pi3722 & w7455;
assign w7677 = pi3834 & w7450;
assign w7678 = pi3770 & w7452;
assign w7679 = pi3818 & w7436;
assign w7680 = ~w7678 & ~w7679;
assign w7681 = ~w7677 & w7680;
assign w7682 = pi3802 & w7440;
assign w7683 = pi3754 & w7447;
assign w7684 = ~w7432 & ~w7683;
assign w7685 = ~w7682 & w7684;
assign w7686 = pi3738 & w7438;
assign w7687 = pi3786 & w7444;
assign w7688 = ~w7686 & ~w7687;
assign w7689 = w7685 & w7688;
assign w7690 = w7681 & w7689;
assign w7691 = ~w7676 & w7690;
assign w7692 = (pi0574 & ~w3104) | (pi0574 & w37080) | (~w3104 & w37080);
assign w7693 = pi0537 & ~w3120;
assign w7694 = pi0523 & ~w3079;
assign w7695 = ~w7693 & ~w7694;
assign w7696 = (~w941 & ~w7695) | (~w941 & w37081) | (~w7695 & w37081);
assign w7697 = pi2115 & pi2419;
assign w7698 = w7432 & ~w7697;
assign w7699 = (w7698 & ~w7696) | (w7698 & w37082) | (~w7696 & w37082);
assign w7700 = ~w7691 & ~w7699;
assign w7701 = (w184 & w37083) | (w184 & w37084) | (w37083 & w37084);
assign w7702 = (~w7701 & ~w7416) | (~w7701 & w37085) | (~w7416 & w37085);
assign w7703 = ~w7675 & w7702;
assign w7704 = w201 & ~w7703;
assign w7705 = ~w7674 & ~w7704;
assign w7706 = pi3107 & ~pi3626;
assign w7707 = pi0383 & w7418;
assign w7708 = pi3723 & w7455;
assign w7709 = pi3803 & w7440;
assign w7710 = pi3771 & w7452;
assign w7711 = pi3819 & w7436;
assign w7712 = ~w7710 & ~w7711;
assign w7713 = ~w7709 & w7712;
assign w7714 = pi3787 & w7444;
assign w7715 = pi3755 & w7447;
assign w7716 = ~w7432 & ~w7715;
assign w7717 = ~w7714 & w7716;
assign w7718 = pi3739 & w7438;
assign w7719 = pi3835 & w7450;
assign w7720 = ~w7718 & ~w7719;
assign w7721 = w7717 & w7720;
assign w7722 = w7713 & w7721;
assign w7723 = ~w7708 & w7722;
assign w7724 = (pi0574 & ~w6122) | (pi0574 & w37086) | (~w6122 & w37086);
assign w7725 = pi0523 & ~w6083;
assign w7726 = (pi0537 & ~w6098) | (pi0537 & w37087) | (~w6098 & w37087);
assign w7727 = ~w7725 & w37088;
assign w7728 = ~w941 & ~w7727;
assign w7729 = pi2414 & pi2419;
assign w7730 = w7432 & ~w7729;
assign w7731 = (w7730 & w7727) | (w7730 & w37089) | (w7727 & w37089);
assign w7732 = ~w7723 & ~w7731;
assign w7733 = (w184 & w37090) | (w184 & w37091) | (w37090 & w37091);
assign w7734 = (~w7733 & ~w7416) | (~w7733 & w37092) | (~w7416 & w37092);
assign w7735 = ~w7707 & w7734;
assign w7736 = w201 & ~w7735;
assign w7737 = ~w7706 & ~w7736;
assign w7738 = pi3063 & ~pi3626;
assign w7739 = pi0382 & w7418;
assign w7740 = pi3724 & w7455;
assign w7741 = pi3740 & w7438;
assign w7742 = pi3788 & w7444;
assign w7743 = pi3820 & w7436;
assign w7744 = ~w7742 & ~w7743;
assign w7745 = ~w7741 & w7744;
assign w7746 = pi3772 & w7452;
assign w7747 = pi3756 & w7447;
assign w7748 = ~w7432 & ~w7747;
assign w7749 = ~w7746 & w7748;
assign w7750 = pi3836 & w7450;
assign w7751 = pi3804 & w7440;
assign w7752 = ~w7750 & ~w7751;
assign w7753 = w7749 & w7752;
assign w7754 = w7745 & w7753;
assign w7755 = ~w7740 & w7754;
assign w7756 = pi0574 & ~w4071;
assign w7757 = (pi0537 & ~w4086) | (pi0537 & w37087) | (~w4086 & w37087);
assign w7758 = pi0523 & ~w4050;
assign w7759 = ~w7758 & w37093;
assign w7760 = ~w941 & ~w7759;
assign w7761 = pi2418 & pi2419;
assign w7762 = w7432 & ~w7761;
assign w7763 = (w7762 & w7759) | (w7762 & w37094) | (w7759 & w37094);
assign w7764 = ~w7755 & ~w7763;
assign w7765 = (w184 & w37095) | (w184 & w37096) | (w37095 & w37096);
assign w7766 = (~w7765 & ~w7416) | (~w7765 & w37097) | (~w7416 & w37097);
assign w7767 = ~w7739 & w7766;
assign w7768 = w201 & ~w7767;
assign w7769 = ~w7738 & ~w7768;
assign w7770 = pi3091 & ~pi3626;
assign w7771 = pi0392 & w7418;
assign w7772 = pi3725 & w7455;
assign w7773 = pi3805 & w7440;
assign w7774 = pi3773 & w7452;
assign w7775 = pi3821 & w7436;
assign w7776 = ~w7774 & ~w7775;
assign w7777 = ~w7773 & w7776;
assign w7778 = pi3789 & w7444;
assign w7779 = pi3757 & w7447;
assign w7780 = ~w7432 & ~w7779;
assign w7781 = ~w7778 & w7780;
assign w7782 = pi3837 & w7450;
assign w7783 = pi3741 & w7438;
assign w7784 = ~w7782 & ~w7783;
assign w7785 = w7781 & w7784;
assign w7786 = w7777 & w7785;
assign w7787 = ~w7772 & w7786;
assign w7788 = pi0523 & ~w5000;
assign w7789 = (pi0574 & ~w4969) | (pi0574 & w37098) | (~w4969 & w37098);
assign w7790 = pi0537 & ~w4945;
assign w7791 = ~w7789 & ~w7790;
assign w7792 = (~w941 & ~w7791) | (~w941 & w37099) | (~w7791 & w37099);
assign w7793 = pi1951 & pi2419;
assign w7794 = w7432 & ~w7793;
assign w7795 = (w7794 & ~w7792) | (w7794 & w37100) | (~w7792 & w37100);
assign w7796 = ~w7787 & ~w7795;
assign w7797 = (w184 & w37101) | (w184 & w37102) | (w37101 & w37102);
assign w7798 = (~w7797 & ~w7416) | (~w7797 & w37103) | (~w7416 & w37103);
assign w7799 = ~w7771 & w7798;
assign w7800 = w201 & ~w7799;
assign w7801 = ~w7770 & ~w7800;
assign w7802 = pi2989 & ~pi3626;
assign w7803 = pi0391 & w7418;
assign w7804 = pi3726 & w7455;
assign w7805 = pi3806 & w7440;
assign w7806 = pi3838 & w7450;
assign w7807 = pi3822 & w7436;
assign w7808 = ~w7806 & ~w7807;
assign w7809 = ~w7805 & w7808;
assign w7810 = pi3790 & w7444;
assign w7811 = pi3758 & w7447;
assign w7812 = ~w7432 & ~w7811;
assign w7813 = ~w7810 & w7812;
assign w7814 = pi3742 & w7438;
assign w7815 = pi3774 & w7452;
assign w7816 = ~w7814 & ~w7815;
assign w7817 = w7813 & w7816;
assign w7818 = w7809 & w7817;
assign w7819 = ~w7804 & w7818;
assign w7820 = (pi0537 & ~w5624) | (pi0537 & w37087) | (~w5624 & w37087);
assign w7821 = pi0574 & ~w5578;
assign w7822 = pi0523 & ~w5609;
assign w7823 = ~w7821 & ~w7822;
assign w7824 = (~w941 & ~w7823) | (~w941 & w37104) | (~w7823 & w37104);
assign w7825 = pi1950 & pi2419;
assign w7826 = w7432 & ~w7825;
assign w7827 = (w7826 & ~w7824) | (w7826 & w37105) | (~w7824 & w37105);
assign w7828 = ~w7819 & ~w7827;
assign w7829 = (w184 & w37106) | (w184 & w37107) | (w37106 & w37107);
assign w7830 = (~w7829 & ~w7416) | (~w7829 & w37108) | (~w7416 & w37108);
assign w7831 = ~w7803 & w7830;
assign w7832 = w201 & ~w7831;
assign w7833 = ~w7802 & ~w7832;
assign w7834 = pi2988 & ~pi3626;
assign w7835 = pi0381 & w7418;
assign w7836 = pi3727 & w7455;
assign w7837 = pi3839 & w7450;
assign w7838 = pi3775 & w7452;
assign w7839 = pi3823 & w7436;
assign w7840 = ~w7838 & ~w7839;
assign w7841 = ~w7837 & w7840;
assign w7842 = pi3807 & w7440;
assign w7843 = pi3759 & w7447;
assign w7844 = ~w7432 & ~w7843;
assign w7845 = ~w7842 & w7844;
assign w7846 = pi3743 & w7438;
assign w7847 = pi3791 & w7444;
assign w7848 = ~w7846 & ~w7847;
assign w7849 = w7845 & w7848;
assign w7850 = w7841 & w7849;
assign w7851 = ~w7836 & w7850;
assign w7852 = (pi0574 & ~w1139) | (pi0574 & w37109) | (~w1139 & w37109);
assign w7853 = pi0523 & ~w1174;
assign w7854 = (pi0537 & ~w1198) | (pi0537 & w37087) | (~w1198 & w37087);
assign w7855 = ~w7853 & w37110;
assign w7856 = ~w941 & ~w7855;
assign w7857 = pi1949 & pi2419;
assign w7858 = w7432 & ~w7857;
assign w7859 = (w7858 & w7855) | (w7858 & w37111) | (w7855 & w37111);
assign w7860 = ~w7851 & ~w7859;
assign w7861 = (w184 & w37112) | (w184 & w37113) | (w37112 & w37113);
assign w7862 = (~w7861 & ~w7416) | (~w7861 & w37114) | (~w7416 & w37114);
assign w7863 = ~w7835 & w7862;
assign w7864 = w201 & ~w7863;
assign w7865 = ~w7834 & ~w7864;
assign w7866 = pi2987 & ~pi3626;
assign w7867 = pi0378 & w7418;
assign w7868 = pi3728 & w7455;
assign w7869 = pi3808 & w7440;
assign w7870 = pi3840 & w7450;
assign w7871 = pi3824 & w7436;
assign w7872 = ~w7870 & ~w7871;
assign w7873 = ~w7869 & w7872;
assign w7874 = pi3792 & w7444;
assign w7875 = pi3760 & w7447;
assign w7876 = ~w7432 & ~w7875;
assign w7877 = ~w7874 & w7876;
assign w7878 = pi3744 & w7438;
assign w7879 = pi3776 & w7452;
assign w7880 = ~w7878 & ~w7879;
assign w7881 = w7877 & w7880;
assign w7882 = w7873 & w7881;
assign w7883 = ~w7868 & w7882;
assign w7884 = pi0523 & ~w1536;
assign w7885 = (pi0537 & ~w1551) | (pi0537 & w37087) | (~w1551 & w37087);
assign w7886 = pi0574 & ~w1453;
assign w7887 = ~w7885 & ~w7886;
assign w7888 = (~w941 & ~w7887) | (~w941 & w37115) | (~w7887 & w37115);
assign w7889 = pi1948 & pi2419;
assign w7890 = w7432 & ~w7889;
assign w7891 = (w7890 & ~w7888) | (w7890 & w37116) | (~w7888 & w37116);
assign w7892 = ~w7883 & ~w7891;
assign w7893 = (w184 & w37117) | (w184 & w37118) | (w37117 & w37118);
assign w7894 = ~w183 & w37119;
assign w7895 = ~w7893 & ~w7894;
assign w7896 = ~w7867 & w7895;
assign w7897 = w201 & ~w7896;
assign w7898 = ~w7866 & ~w7897;
assign w7899 = pi3097 & ~pi3626;
assign w7900 = pi0377 & w7418;
assign w7901 = pi3729 & w7455;
assign w7902 = pi3809 & w7440;
assign w7903 = pi3841 & w7450;
assign w7904 = pi3825 & w7436;
assign w7905 = ~w7903 & ~w7904;
assign w7906 = ~w7902 & w7905;
assign w7907 = pi3793 & w7444;
assign w7908 = pi3761 & w7447;
assign w7909 = ~w7432 & ~w7908;
assign w7910 = ~w7907 & w7909;
assign w7911 = pi3745 & w7438;
assign w7912 = pi3777 & w7452;
assign w7913 = ~w7911 & ~w7912;
assign w7914 = w7910 & w7913;
assign w7915 = w7906 & w7914;
assign w7916 = ~w7901 & w7915;
assign w7917 = pi0979 & pi2861;
assign w7918 = ~pi0979 & pi2868;
assign w7919 = ~w7917 & ~w7918;
assign w7920 = pi0763 & ~w7919;
assign w7921 = pi0979 & pi3172;
assign w7922 = ~pi0979 & pi2639;
assign w7923 = ~w7921 & ~w7922;
assign w7924 = pi0765 & ~w7923;
assign w7925 = pi0212 & ~pi0979;
assign w7926 = pi0211 & pi0979;
assign w7927 = ~w7925 & ~w7926;
assign w7928 = pi0721 & ~w7927;
assign w7929 = ~w7924 & ~w7928;
assign w7930 = ~w7920 & w7929;
assign w7931 = pi0979 & pi3183;
assign w7932 = ~pi0979 & pi2914;
assign w7933 = ~w7931 & ~w7932;
assign w7934 = pi0766 & ~w7933;
assign w7935 = ~w1144 & ~w7934;
assign w7936 = pi0979 & pi2869;
assign w7937 = ~pi0979 & pi2878;
assign w7938 = ~w7936 & ~w7937;
assign w7939 = pi0764 & ~w7938;
assign w7940 = pi0119 & ~pi0979;
assign w7941 = pi0115 & pi0979;
assign w7942 = ~w7940 & ~w7941;
assign w7943 = pi0720 & ~w7942;
assign w7944 = ~w7939 & ~w7943;
assign w7945 = w7935 & w7944;
assign w7946 = w7930 & w7945;
assign w7947 = pi0523 & ~w7946;
assign w7948 = pi0298 & ~pi0979;
assign w7949 = pi0297 & pi0979;
assign w7950 = ~w7948 & ~w7949;
assign w7951 = pi0716 & ~w7950;
assign w7952 = pi0979 & pi2134;
assign w7953 = ~pi0979 & pi2851;
assign w7954 = ~w7952 & ~w7953;
assign w7955 = pi0717 & ~w7954;
assign w7956 = pi0320 & ~pi0979;
assign w7957 = pi0318 & pi0979;
assign w7958 = ~w7956 & ~w7957;
assign w7959 = pi0761 & ~w7958;
assign w7960 = ~w7955 & ~w7959;
assign w7961 = ~w7951 & w7960;
assign w7962 = (pi0537 & ~w7961) | (pi0537 & w37087) | (~w7961 & w37087);
assign w7963 = pi0979 & pi1791;
assign w7964 = ~pi0979 & pi2160;
assign w7965 = ~w7963 & ~w7964;
assign w7966 = pi0768 & ~w7965;
assign w7967 = pi0979 & pi2187;
assign w7968 = ~pi0979 & pi2947;
assign w7969 = ~w7967 & ~w7968;
assign w7970 = pi0837 & ~w7969;
assign w7971 = ~w7966 & ~w7970;
assign w7972 = pi0979 & pi2171;
assign w7973 = ~pi0979 & pi2804;
assign w7974 = ~w7972 & ~w7973;
assign w7975 = pi0836 & ~w7974;
assign w7976 = pi0979 & pi2153;
assign w7977 = ~pi0979 & pi2925;
assign w7978 = ~w7976 & ~w7977;
assign w7979 = pi0767 & ~w7978;
assign w7980 = pi0177 & ~pi0979;
assign w7981 = pi0162 & pi0979;
assign w7982 = ~w7980 & ~w7981;
assign w7983 = pi0838 & ~w7982;
assign w7984 = ~w7979 & ~w7983;
assign w7985 = ~w7975 & w7984;
assign w7986 = w7971 & w7985;
assign w7987 = (pi0574 & ~w7985) | (pi0574 & w37120) | (~w7985 & w37120);
assign w7988 = ~w7962 & ~w7987;
assign w7989 = ~w7947 & w7988;
assign w7990 = ~w941 & ~w7989;
assign w7991 = pi1947 & pi2419;
assign w7992 = w7432 & ~w7991;
assign w7993 = (w7992 & w7989) | (w7992 & w37121) | (w7989 & w37121);
assign w7994 = ~w7916 & ~w7993;
assign w7995 = (w184 & w37122) | (w184 & w37123) | (w37122 & w37123);
assign w7996 = pi3873 & w983;
assign w7997 = w970 & w37124;
assign w7998 = w973 & w37125;
assign w7999 = w970 & w37126;
assign w8000 = ~w7998 & ~w7999;
assign w8001 = ~w7997 & w8000;
assign w8002 = w963 & w37127;
assign w8003 = w953 & w37128;
assign w8004 = w958 & w37129;
assign w8005 = ~w8003 & ~w8004;
assign w8006 = ~w8002 & w8005;
assign w8007 = w973 & w37130;
assign w8008 = w963 & w37131;
assign w8009 = ~w997 & ~w8008;
assign w8010 = ~w8007 & w8009;
assign w8011 = w8006 & w8010;
assign w8012 = w8001 & w8011;
assign w8013 = ~w7996 & w8012;
assign w8014 = w940 & w37132;
assign w8015 = pi1854 & w1263;
assign w8016 = pi1723 & w1294;
assign w8017 = ~w8015 & ~w8016;
assign w8018 = pi1869 & w1278;
assign w8019 = pi1904 & w1238;
assign w8020 = ~w8018 & ~w8019;
assign w8021 = w8017 & w8020;
assign w8022 = pi1792 & w1268;
assign w8023 = pi1929 & w1272;
assign w8024 = ~w8022 & ~w8023;
assign w8025 = pi3680 & w3180;
assign w8026 = pi0887 & w1251;
assign w8027 = ~w8025 & ~w8026;
assign w8028 = w8024 & w8027;
assign w8029 = pi1102 & w1266;
assign w8030 = pi0896 & w1254;
assign w8031 = ~w8029 & ~w8030;
assign w8032 = pi2123 & w1275;
assign w8033 = pi1759 & w1249;
assign w8034 = ~w8032 & ~w8033;
assign w8035 = w8031 & w8034;
assign w8036 = w8028 & w8035;
assign w8037 = w8021 & w8036;
assign w8038 = w1216 & w37133;
assign w8039 = pi0959 & w1245;
assign w8040 = pi0246 & w1242;
assign w8041 = ~w8039 & ~w8040;
assign w8042 = pi0970 & w1234;
assign w8043 = pi1917 & w1280;
assign w8044 = ~w8042 & ~w8043;
assign w8045 = w8041 & w8044;
assign w8046 = ~w1289 & ~w1292;
assign w8047 = pi1422 & w1296;
assign w8048 = pi1781 & w1258;
assign w8049 = ~w8047 & ~w8048;
assign w8050 = w8046 & w8049;
assign w8051 = w8045 & w8050;
assign w8052 = ~w8038 & w8051;
assign w8053 = w8037 & w8052;
assign w8054 = pi1934 & ~w8053;
assign w8055 = pi0524 & ~w7946;
assign w8056 = pi0607 & pi1336;
assign w8057 = pi1335 & pi2592;
assign w8058 = ~w8056 & ~w8057;
assign w8059 = pi1332 & pi2577;
assign w8060 = pi1333 & pi1866;
assign w8061 = ~w8059 & ~w8060;
assign w8062 = w8058 & w8061;
assign w8063 = pi0762 & ~w8062;
assign w8064 = pi3233 & pi3396;
assign w8065 = pi0377 & pi1057;
assign w8066 = pi3329 & pi3519;
assign w8067 = ~w8065 & ~w8066;
assign w8068 = (pi0650 & ~w8067) | (pi0650 & w37134) | (~w8067 & w37134);
assign w8069 = ~w8063 & ~w8068;
assign w8070 = w1487 & w8069;
assign w8071 = ~w8055 & w8070;
assign w8072 = (pi0538 & ~w7961) | (pi0538 & w35782) | (~w7961 & w35782);
assign w8073 = pi0576 & ~w7986;
assign w8074 = ~w8072 & ~w8073;
assign w8075 = w8071 & w8074;
assign w8076 = ~w941 & ~w8075;
assign w8077 = ~w8054 & ~w8076;
assign w8078 = pi1787 & pi2832;
assign w8079 = w958 & w37136;
assign w8080 = (w8077 & w37137) | (w8077 & w37138) | (w37137 & w37138);
assign w8081 = ~w8013 & ~w8080;
assign w8082 = ~w183 & w37139;
assign w8083 = ~w7995 & ~w8082;
assign w8084 = ~w7900 & w8083;
assign w8085 = w201 & ~w8084;
assign w8086 = ~w7899 & ~w8085;
assign w8087 = pi0376 & w7418;
assign w8088 = pi3874 & w983;
assign w8089 = w970 & w37140;
assign w8090 = w973 & w37141;
assign w8091 = w970 & w37142;
assign w8092 = ~w8090 & ~w8091;
assign w8093 = ~w8089 & w8092;
assign w8094 = w963 & w37143;
assign w8095 = w953 & w37144;
assign w8096 = w963 & w37145;
assign w8097 = ~w8095 & ~w8096;
assign w8098 = ~w8094 & w8097;
assign w8099 = w973 & w37146;
assign w8100 = w958 & w37147;
assign w8101 = ~w997 & ~w8100;
assign w8102 = ~w8099 & w8101;
assign w8103 = w8098 & w8102;
assign w8104 = w8093 & w8103;
assign w8105 = ~w8088 & w8104;
assign w8106 = w940 & w37148;
assign w8107 = pi0895 & w1254;
assign w8108 = pi0958 & w1245;
assign w8109 = pi1758 & w1249;
assign w8110 = ~w8108 & ~w8109;
assign w8111 = ~w8107 & w8110;
assign w8112 = pi0969 & w1234;
assign w8113 = pi1889 & w1278;
assign w8114 = ~w8112 & ~w8113;
assign w8115 = pi0886 & w1251;
assign w8116 = pi2109 & w1275;
assign w8117 = ~w8115 & ~w8116;
assign w8118 = w8114 & w8117;
assign w8119 = pi0893 & w1291;
assign w8120 = pi0223 & w1242;
assign w8121 = ~w8119 & ~w8120;
assign w8122 = pi1722 & w1294;
assign w8123 = pi1928 & w1272;
assign w8124 = ~w8122 & ~w8123;
assign w8125 = w8121 & w8124;
assign w8126 = w8118 & w8125;
assign w8127 = w8111 & w8126;
assign w8128 = w1216 & w37149;
assign w8129 = pi1835 & w1268;
assign w8130 = pi0799 & w1288;
assign w8131 = ~w8129 & ~w8130;
assign w8132 = pi2385 & w3180;
assign w8133 = pi1768 & w1263;
assign w8134 = ~w8132 & ~w8133;
assign w8135 = w8131 & w8134;
assign w8136 = pi1908 & w1280;
assign w8137 = pi1903 & w1238;
assign w8138 = ~w8136 & ~w8137;
assign w8139 = pi1024 & w1266;
assign w8140 = pi1426 & w3139;
assign w8141 = ~w8139 & ~w8140;
assign w8142 = w8138 & w8141;
assign w8143 = w8135 & w8142;
assign w8144 = ~w8128 & w8143;
assign w8145 = w8127 & w8144;
assign w8146 = pi1934 & ~w8145;
assign w8147 = pi0979 & pi3140;
assign w8148 = ~pi0979 & pi2877;
assign w8149 = ~w8147 & ~w8148;
assign w8150 = pi0764 & ~w8149;
assign w8151 = pi0979 & pi3182;
assign w8152 = ~pi0979 & pi2894;
assign w8153 = ~w8151 & ~w8152;
assign w8154 = pi0766 & ~w8153;
assign w8155 = pi0059 & ~pi0979;
assign w8156 = pi0058 & pi0979;
assign w8157 = ~w8155 & ~w8156;
assign w8158 = pi0720 & ~w8157;
assign w8159 = ~w8154 & ~w8158;
assign w8160 = ~w8150 & w8159;
assign w8161 = pi0979 & pi3158;
assign w8162 = ~pi0979 & pi2867;
assign w8163 = ~w8161 & ~w8162;
assign w8164 = pi0763 & ~w8163;
assign w8165 = ~w1144 & ~w8164;
assign w8166 = pi0979 & pi3171;
assign w8167 = ~pi0979 & pi2638;
assign w8168 = ~w8166 & ~w8167;
assign w8169 = pi0765 & ~w8168;
assign w8170 = pi0193 & ~pi0979;
assign w8171 = pi0192 & pi0979;
assign w8172 = ~w8170 & ~w8171;
assign w8173 = pi0721 & ~w8172;
assign w8174 = ~w8169 & ~w8173;
assign w8175 = w8165 & w8174;
assign w8176 = w8160 & w8175;
assign w8177 = pi0524 & ~w8176;
assign w8178 = pi1333 & pi1897;
assign w8179 = pi1335 & pi2591;
assign w8180 = ~w8178 & ~w8179;
assign w8181 = pi0605 & pi1336;
assign w8182 = pi1332 & pi2576;
assign w8183 = ~w8181 & ~w8182;
assign w8184 = w8180 & w8183;
assign w8185 = pi0762 & ~w8184;
assign w8186 = pi3233 & pi3393;
assign w8187 = pi0376 & pi1057;
assign w8188 = ~w8066 & ~w8187;
assign w8189 = (pi0650 & ~w8188) | (pi0650 & w37150) | (~w8188 & w37150);
assign w8190 = ~w8185 & ~w8189;
assign w8191 = w1487 & w8190;
assign w8192 = ~w8177 & w8191;
assign w8193 = pi0286 & ~pi0979;
assign w8194 = pi0285 & pi0979;
assign w8195 = ~w8193 & ~w8194;
assign w8196 = pi0716 & ~w8195;
assign w8197 = pi0979 & pi2133;
assign w8198 = ~pi0979 & pi2850;
assign w8199 = ~w8197 & ~w8198;
assign w8200 = pi0717 & ~w8199;
assign w8201 = pi0254 & ~pi0979;
assign w8202 = pi0251 & pi0979;
assign w8203 = ~w8201 & ~w8202;
assign w8204 = pi0761 & ~w8203;
assign w8205 = ~w8200 & ~w8204;
assign w8206 = ~w8196 & w8205;
assign w8207 = w1184 & w8206;
assign w8208 = (pi0538 & ~w8206) | (pi0538 & w35782) | (~w8206 & w35782);
assign w8209 = pi0979 & pi1963;
assign w8210 = ~pi0979 & pi2428;
assign w8211 = ~w8209 & ~w8210;
assign w8212 = pi0768 & ~w8211;
assign w8213 = pi0979 & pi2170;
assign w8214 = ~pi0979 & pi2805;
assign w8215 = ~w8213 & ~w8214;
assign w8216 = pi0836 & ~w8215;
assign w8217 = ~w8212 & ~w8216;
assign w8218 = pi0151 & ~pi0979;
assign w8219 = pi0150 & pi0979;
assign w8220 = ~w8218 & ~w8219;
assign w8221 = pi0838 & ~w8220;
assign w8222 = pi0979 & pi2186;
assign w8223 = ~pi0979 & pi2946;
assign w8224 = ~w8222 & ~w8223;
assign w8225 = pi0837 & ~w8224;
assign w8226 = pi0979 & pi2152;
assign w8227 = ~pi0979 & pi2924;
assign w8228 = ~w8226 & ~w8227;
assign w8229 = pi0767 & ~w8228;
assign w8230 = ~w8225 & ~w8229;
assign w8231 = ~w8221 & w8230;
assign w8232 = (pi0576 & ~w8231) | (pi0576 & w37151) | (~w8231 & w37151);
assign w8233 = ~w8208 & ~w8232;
assign w8234 = (~w941 & ~w8192) | (~w941 & w37152) | (~w8192 & w37152);
assign w8235 = ~w8146 & ~w8234;
assign w8236 = ~w8146 & w37153;
assign w8237 = pi1787 & pi2816;
assign w8238 = w958 & w37154;
assign w8239 = (w8238 & w8236) | (w8238 & w37155) | (w8236 & w37155);
assign w8240 = ~w8105 & ~w8239;
assign w8241 = ~w183 & w37156;
assign w8242 = pi3730 & w7455;
assign w8243 = pi3810 & w7440;
assign w8244 = pi3778 & w7452;
assign w8245 = pi3826 & w7436;
assign w8246 = ~w8244 & ~w8245;
assign w8247 = ~w8243 & w8246;
assign w8248 = pi3794 & w7444;
assign w8249 = pi3762 & w7447;
assign w8250 = ~w7432 & ~w8249;
assign w8251 = ~w8248 & w8250;
assign w8252 = pi3842 & w7450;
assign w8253 = pi3746 & w7438;
assign w8254 = ~w8252 & ~w8253;
assign w8255 = w8251 & w8254;
assign w8256 = w8247 & w8255;
assign w8257 = ~w8242 & w8256;
assign w8258 = pi0523 & ~w8176;
assign w8259 = (pi0574 & ~w8231) | (pi0574 & w37157) | (~w8231 & w37157);
assign w8260 = pi0537 & ~w8207;
assign w8261 = ~w8259 & ~w8260;
assign w8262 = (~w941 & ~w8261) | (~w941 & w37158) | (~w8261 & w37158);
assign w8263 = pi1946 & pi2419;
assign w8264 = w7432 & ~w8263;
assign w8265 = (w8264 & ~w8262) | (w8264 & w37159) | (~w8262 & w37159);
assign w8266 = ~w8257 & ~w8265;
assign w8267 = (w184 & w37160) | (w184 & w37161) | (w37160 & w37161);
assign w8268 = ~w8241 & ~w8267;
assign w8269 = ~w8087 & w8268;
assign w8270 = ~pi1422 & ~pi1856;
assign w8271 = ~pi0366 & ~w8270;
assign w8272 = (pi3641 & ~w8270) | (pi3641 & w37162) | (~w8270 & w37162);
assign w8273 = ~w8271 & w8272;
assign w8274 = ~pi0359 & ~w8270;
assign w8275 = (pi3641 & ~w8270) | (pi3641 & w37163) | (~w8270 & w37163);
assign w8276 = ~w8274 & w8275;
assign w8277 = pi0432 & w8270;
assign w8278 = (pi3641 & w8270) | (pi3641 & w37164) | (w8270 & w37164);
assign w8279 = ~w8277 & w8278;
assign w8280 = ~pi0357 & ~w8270;
assign w8281 = (pi3641 & ~w8270) | (pi3641 & w37165) | (~w8270 & w37165);
assign w8282 = ~w8280 & w8281;
assign w8283 = ~pi0356 & ~w8270;
assign w8284 = (pi3641 & ~w8270) | (pi3641 & w37166) | (~w8270 & w37166);
assign w8285 = ~w8283 & w8284;
assign w8286 = pi0429 & w8270;
assign w8287 = (pi3641 & w8270) | (pi3641 & w37167) | (w8270 & w37167);
assign w8288 = ~w8286 & w8287;
assign w8289 = ~pi0354 & ~w8270;
assign w8290 = (pi3641 & ~w8270) | (pi3641 & w37168) | (~w8270 & w37168);
assign w8291 = ~w8289 & w8290;
assign w8292 = pi0435 & w8270;
assign w8293 = (pi3641 & w8270) | (pi3641 & w37169) | (w8270 & w37169);
assign w8294 = ~w8292 & w8293;
assign w8295 = pi3641 & ~w8270;
assign w8296 = pi0352 & w8295;
assign w8297 = pi0351 & w8295;
assign w8298 = pi0365 & ~w8270;
assign w8299 = pi3641 & ~w8298;
assign w8300 = pi0364 & w8295;
assign w8301 = pi0363 & w8295;
assign w8302 = pi0362 & ~w8270;
assign w8303 = pi3641 & ~w8302;
assign w8304 = pi0361 & w8295;
assign w8305 = pi0360 & ~w8270;
assign w8306 = pi3641 & ~w8305;
assign w8307 = ~w3485 & ~w7424;
assign w8308 = w2259 & w8307;
assign w8309 = ~pi1092 & w40129;
assign w8310 = ~pi0366 & w40130;
assign w8311 = ~w8309 & ~w8310;
assign w8312 = ~w8308 & w8311;
assign w8313 = (w7500 & w37170) | (w7500 & w37171) | (w37170 & w37171);
assign w8314 = w2259 & w8313;
assign w8315 = ~pi1060 & w40129;
assign w8316 = ~pi0359 & w40130;
assign w8317 = ~w8315 & ~w8316;
assign w8318 = ~w8314 & w8317;
assign w8319 = (~w5673 & w7532) | (~w5673 & w37172) | (w7532 & w37172);
assign w8320 = w2259 & w8319;
assign w8321 = ~pi1089 & w40129;
assign w8322 = ~pi0358 & w40130;
assign w8323 = ~w8321 & ~w8322;
assign w8324 = ~w8320 & w8323;
assign w8325 = (w7565 & w37173) | (w7565 & w37174) | (w37173 & w37174);
assign w8326 = w2259 & w8325;
assign w8327 = ~pi1065 & w40129;
assign w8328 = ~pi0357 & w40130;
assign w8329 = ~w8327 & ~w8328;
assign w8330 = ~w8326 & w8329;
assign w8331 = (w7597 & w37175) | (w7597 & w37176) | (w37175 & w37176);
assign w8332 = w2259 & w8331;
assign w8333 = ~pi1064 & w40129;
assign w8334 = ~pi0356 & w40130;
assign w8335 = ~w8333 & ~w8334;
assign w8336 = ~w8332 & w8335;
assign w8337 = w940 & w37177;
assign w8338 = ~w7631 & ~w8337;
assign w8339 = w2259 & w8338;
assign w8340 = ~pi1063 & w40129;
assign w8341 = ~pi0355 & w40130;
assign w8342 = ~w8340 & ~w8341;
assign w8343 = ~w8339 & w8342;
assign w8344 = ~w3197 & ~w7664;
assign w8345 = w2259 & w8344;
assign w8346 = ~pi1062 & w40129;
assign w8347 = ~pi0354 & w40130;
assign w8348 = ~w8346 & ~w8347;
assign w8349 = ~w8345 & w8348;
assign w8350 = (w7695 & w37178) | (w7695 & w37179) | (w37178 & w37179);
assign w8351 = w2259 & w8350;
assign w8352 = ~pi1061 & w40129;
assign w8353 = ~pi0353 & w40130;
assign w8354 = ~w8352 & ~w8353;
assign w8355 = ~w8351 & w8354;
assign w8356 = (~w5988 & w7727) | (~w5988 & w37180) | (w7727 & w37180);
assign w8357 = w2259 & w8356;
assign w8358 = ~pi3106 & w40129;
assign w8359 = ~pi0352 & w40130;
assign w8360 = ~w8358 & ~w8359;
assign w8361 = ~w8357 & w8360;
assign w8362 = (~w3955 & w7759) | (~w3955 & w37181) | (w7759 & w37181);
assign w8363 = w2259 & w8362;
assign w8364 = ~pi3105 & w40129;
assign w8365 = ~pi0351 & w40130;
assign w8366 = ~w8364 & ~w8365;
assign w8367 = ~w8363 & w8366;
assign w8368 = ~w4867 & ~w7792;
assign w8369 = w2259 & w8368;
assign w8370 = ~pi3104 & w40129;
assign w8371 = ~pi0365 & w40130;
assign w8372 = ~w8370 & ~w8371;
assign w8373 = ~w8369 & w8372;
assign w8374 = w940 & w37182;
assign w8375 = (w7823 & w37183) | (w7823 & w37184) | (w37183 & w37184);
assign w8376 = w2259 & w8375;
assign w8377 = ~pi0364 & w40130;
assign w8378 = ~pi2985 & w40129;
assign w8379 = ~w8377 & ~w8378;
assign w8380 = ~w8376 & w8379;
assign w8381 = (~w1003 & w7855) | (~w1003 & w37185) | (w7855 & w37185);
assign w8382 = w2259 & w8381;
assign w8383 = ~pi3102 & w40129;
assign w8384 = ~pi0363 & w40130;
assign w8385 = ~w8383 & ~w8384;
assign w8386 = ~w8382 & w8385;
assign w8387 = ~w1380 & ~w7888;
assign w8388 = w2259 & w8387;
assign w8389 = ~pi3109 & w40129;
assign w8390 = ~pi0362 & w40130;
assign w8391 = ~w8389 & ~w8390;
assign w8392 = ~w8388 & w8391;
assign w8393 = (~w8014 & w7989) | (~w8014 & w37186) | (w7989 & w37186);
assign w8394 = w2259 & w8393;
assign w8395 = ~pi3111 & w40129;
assign w8396 = ~pi0361 & w40130;
assign w8397 = ~w8395 & ~w8396;
assign w8398 = ~w8394 & w8397;
assign w8399 = ~w8106 & ~w8262;
assign w8400 = w2259 & w8399;
assign w8401 = ~pi3112 & w40129;
assign w8402 = ~pi0360 & w40130;
assign w8403 = ~w8401 & ~w8402;
assign w8404 = ~w8400 & w8403;
assign w8405 = pi0366 & w40131;
assign w8406 = w342 & w346;
assign w8407 = (w825 & ~w342) | (w825 & w37187) | (~w342 & w37187);
assign w8408 = pi0479 & w8407;
assign w8409 = (w822 & ~w342) | (w822 & w37188) | (~w342 & w37188);
assign w8410 = pi2597 & w8409;
assign w8411 = ~w8408 & ~w8410;
assign w8412 = ~w8405 & w8411;
assign w8413 = w342 & w37189;
assign w8414 = w6621 & ~w8413;
assign w8415 = w2891 & w40094;
assign w8416 = pi0844 & w8415;
assign w8417 = (~w8416 & w3707) | (~w8416 & w37190) | (w3707 & w37190);
assign w8418 = w8412 & w8417;
assign w8419 = pi0359 & w40131;
assign w8420 = pi0370 & w8407;
assign w8421 = pi2590 & w8409;
assign w8422 = ~w8420 & ~w8421;
assign w8423 = ~w8419 & w8422;
assign w8424 = pi0843 & w40132;
assign w8425 = (~w8424 & w4745) | (~w8424 & w37191) | (w4745 & w37191);
assign w8426 = w8423 & w8425;
assign w8427 = pi0358 & w40131;
assign w8428 = pi0350 & w8407;
assign w8429 = pi2589 & w8409;
assign w8430 = ~w8428 & ~w8429;
assign w8431 = ~w8427 & w8430;
assign w8432 = pi0842 & w8415;
assign w8433 = (w5893 & w37193) | (w5893 & w37194) | (w37193 & w37194);
assign w8434 = w8431 & w8433;
assign w8435 = pi0357 & w40131;
assign w8436 = pi0331 & w8407;
assign w8437 = pi2588 & w8409;
assign w8438 = ~w8436 & ~w8437;
assign w8439 = ~w8435 & w8438;
assign w8440 = pi0864 & w40132;
assign w8441 = (~w8440 & w5316) | (~w8440 & w37195) | (w5316 & w37195);
assign w8442 = w8439 & w8441;
assign w8443 = pi0356 & w40131;
assign w8444 = pi0329 & w8407;
assign w8445 = pi2587 & w8409;
assign w8446 = ~w8444 & ~w8445;
assign w8447 = ~w8443 & w8446;
assign w8448 = pi0841 & w40132;
assign w8449 = (~w8448 & w4376) | (~w8448 & w37196) | (w4376 & w37196);
assign w8450 = w8447 & w8449;
assign w8451 = pi0355 & w40131;
assign w8452 = pi0278 & w8407;
assign w8453 = pi2764 & w8409;
assign w8454 = ~w8452 & ~w8453;
assign w8455 = ~w8451 & w8454;
assign w8456 = (~w8414 & w6353) | (~w8414 & w37197) | (w6353 & w37197);
assign w8457 = pi0865 & w8415;
assign w8458 = ~w8456 & ~w8457;
assign w8459 = w8455 & w8458;
assign w8460 = pi0354 & w40131;
assign w8461 = pi0248 & w8407;
assign w8462 = pi2586 & w8409;
assign w8463 = ~w8461 & ~w8462;
assign w8464 = ~w8460 & w8463;
assign w8465 = pi0840 & w40132;
assign w8466 = (~w8465 & w3412) | (~w8465 & w37198) | (w3412 & w37198);
assign w8467 = w8464 & w8466;
assign w8468 = pi0353 & w40131;
assign w8469 = pi0247 & w8407;
assign w8470 = pi2585 & w8409;
assign w8471 = ~w8469 & ~w8470;
assign w8472 = ~w8468 & w8471;
assign w8473 = pi0839 & w40132;
assign w8474 = (~w8473 & w3191) | (~w8473 & w37199) | (w3191 & w37199);
assign w8475 = w8472 & w8474;
assign w8476 = pi0352 & w40131;
assign w8477 = pi0232 & w8407;
assign w8478 = pi2584 & w8409;
assign w8479 = ~w8477 & ~w8478;
assign w8480 = ~w8476 & w8479;
assign w8481 = pi1092 & w40132;
assign w8482 = (~w8481 & w6173) | (~w8481 & w37200) | (w6173 & w37200);
assign w8483 = w8480 & w8482;
assign w8484 = pi0351 & w40131;
assign w8485 = pi0237 & w8407;
assign w8486 = pi2583 & w8409;
assign w8487 = ~w8485 & ~w8486;
assign w8488 = ~w8484 & w8487;
assign w8489 = pi1060 & w40132;
assign w8490 = (~w8489 & w4137) | (~w8489 & w37201) | (w4137 & w37201);
assign w8491 = w8488 & w8490;
assign w8492 = pi0365 & w40131;
assign w8493 = pi0225 & w8407;
assign w8494 = pi2596 & w8409;
assign w8495 = ~w8493 & ~w8494;
assign w8496 = ~w8492 & w8495;
assign w8497 = pi1089 & w40132;
assign w8498 = (~w8497 & w5049) | (~w8497 & w37202) | (w5049 & w37202);
assign w8499 = w8496 & w8498;
assign w8500 = pi0364 & w40131;
assign w8501 = pi0224 & w8407;
assign w8502 = pi2595 & w8409;
assign w8503 = ~w8501 & ~w8502;
assign w8504 = ~w8500 & w8503;
assign w8505 = (~w8414 & ~w5630) | (~w8414 & w37203) | (~w5630 & w37203);
assign w8506 = pi1065 & w8415;
assign w8507 = ~w8505 & ~w8506;
assign w8508 = w8504 & w8507;
assign w8509 = pi0363 & w40131;
assign w8510 = pi0189 & w8407;
assign w8511 = pi2594 & w8409;
assign w8512 = ~w8510 & ~w8511;
assign w8513 = ~w8509 & w8512;
assign w8514 = pi1064 & w40132;
assign w8515 = (~w8514 & w1304) | (~w8514 & w37204) | (w1304 & w37204);
assign w8516 = w8513 & w8515;
assign w8517 = pi0362 & w40131;
assign w8518 = pi0606 & w8407;
assign w8519 = pi2593 & w8409;
assign w8520 = ~w8518 & ~w8519;
assign w8521 = ~w8517 & w8520;
assign w8522 = pi1063 & w40132;
assign w8523 = (~w8522 & w1618) | (~w8522 & w37205) | (w1618 & w37205);
assign w8524 = w8521 & w8523;
assign w8525 = pi0361 & w40131;
assign w8526 = pi0607 & w8407;
assign w8527 = pi2592 & w8409;
assign w8528 = ~w8526 & ~w8527;
assign w8529 = ~w8525 & w8528;
assign w8530 = pi1062 & w8415;
assign w8531 = (w8077 & w37207) | (w8077 & w37208) | (w37207 & w37208);
assign w8532 = w8529 & w8531;
assign w8533 = pi0360 & w40131;
assign w8534 = pi0605 & w8407;
assign w8535 = pi2591 & w8409;
assign w8536 = ~w8534 & ~w8535;
assign w8537 = ~w8533 & w8536;
assign w8538 = pi1061 & w40132;
assign w8539 = (~w8538 & w8236) | (~w8538 & w37209) | (w8236 & w37209);
assign w8540 = w8537 & w8539;
assign w8541 = (w788 & w704) | (w788 & w37210) | (w704 & w37210);
assign w8542 = ~w764 & ~w8541;
assign w8543 = ~pi0569 & ~pi0667;
assign w8544 = (~w8543 & ~w463) | (~w8543 & w37211) | (~w463 & w37211);
assign w8545 = ~w502 & w8544;
assign w8546 = (~pi0568 & ~w501) | (~pi0568 & w37212) | (~w501 & w37212);
assign w8547 = (w8546 & ~w8545) | (w8546 & w37213) | (~w8545 & w37213);
assign w8548 = ~w8542 & w8547;
assign w8549 = (w8545 & w770) | (w8545 & w37214) | (w770 & w37214);
assign w8550 = ~w8548 & ~w8549;
assign w8551 = pi0667 & w463;
assign w8552 = ~w501 & ~w8543;
assign w8553 = pi0568 & ~w8552;
assign w8554 = (~w8551 & w574) | (~w8551 & w37215) | (w574 & w37215);
assign w8555 = (pi0641 & ~w8550) | (pi0641 & w37216) | (~w8550 & w37216);
assign w8556 = (~w501 & w575) | (~w501 & w37217) | (w575 & w37217);
assign w8557 = (~w8543 & ~w8550) | (~w8543 & w37218) | (~w8550 & w37218);
assign w8558 = ~w8555 & ~w8557;
assign w8559 = (w874 & w3710) | (w874 & w37219) | (w3710 & w37219);
assign w8560 = (~w8559 & ~w8558) | (~w8559 & w37220) | (~w8558 & w37220);
assign w8561 = ~w371 & w37221;
assign w8562 = ~w414 & w37222;
assign w8563 = ~w8561 & ~w8562;
assign w8564 = ~w392 & w37223;
assign w8565 = ~w405 & w37224;
assign w8566 = ~w8564 & ~w8565;
assign w8567 = w8563 & w8566;
assign w8568 = w423 & ~w8567;
assign w8569 = w873 & ~w8568;
assign w8570 = (w8569 & ~w8560) | (w8569 & w37225) | (~w8560 & w37225);
assign w8571 = pi2540 & ~w935;
assign w8572 = (w353 & w37226) | (w353 & w37227) | (w37226 & w37227);
assign w8573 = w940 & w37230;
assign w8574 = (w342 & w37231) | (w342 & w37232) | (w37231 & w37232);
assign w8575 = ~w8571 & w37233;
assign w8576 = ~pi0749 & ~w905;
assign w8577 = (~w8576 & w423) | (~w8576 & w37234) | (w423 & w37234);
assign w8578 = ~w8575 & w8577;
assign w8579 = pi2447 & w1316;
assign w8580 = ~w414 & w37235;
assign w8581 = ~w8579 & ~w8580;
assign w8582 = pi1985 & w1309;
assign w8583 = pi2270 & w1314;
assign w8584 = ~w8582 & ~w8583;
assign w8585 = w8581 & w8584;
assign w8586 = w424 & ~w8585;
assign w8587 = ~w873 & ~w8586;
assign w8588 = ~w8578 & w8587;
assign w8589 = ~w8570 & ~w8588;
assign w8590 = ~w600 & ~w609;
assign w8591 = (~w8590 & w463) | (~w8590 & w37237) | (w463 & w37237);
assign w8592 = w597 & ~w8591;
assign w8593 = (w463 & w37238) | (w463 & w37239) | (w37238 & w37239);
assign w8594 = ~w8592 & w37240;
assign w8595 = (pi0665 & w8592) | (pi0665 & w37241) | (w8592 & w37241);
assign w8596 = ~w8594 & ~w8595;
assign w8597 = w797 & w37242;
assign w8598 = (pi0665 & w503) | (pi0665 & w37243) | (w503 & w37243);
assign w8599 = ~w503 & w506;
assign w8600 = ~w8598 & ~w8599;
assign w8601 = (w8600 & ~w797) | (w8600 & w37244) | (~w797 & w37244);
assign w8602 = ~w8597 & ~w8601;
assign w8603 = ~w371 & w37245;
assign w8604 = ~w392 & w37246;
assign w8605 = ~w8603 & ~w8604;
assign w8606 = ~w414 & w37247;
assign w8607 = ~w405 & w37248;
assign w8608 = ~w8606 & ~w8607;
assign w8609 = w8605 & w8608;
assign w8610 = ~w424 & w8609;
assign w8611 = w876 & ~w8610;
assign w8612 = (w8611 & w8602) | (w8611 & w37249) | (w8602 & w37249);
assign w8613 = pi1982 & w1309;
assign w8614 = ~w414 & w37250;
assign w8615 = ~w8613 & ~w8614;
assign w8616 = pi2444 & w1316;
assign w8617 = pi2267 & w1314;
assign w8618 = ~w8616 & ~w8617;
assign w8619 = w8615 & w8618;
assign w8620 = w424 & ~w8619;
assign w8621 = ~pi0778 & ~w905;
assign w8622 = (pi2549 & w934) | (pi2549 & w37251) | (w934 & w37251);
assign w8623 = (w353 & w37252) | (w353 & w37253) | (w37252 & w37253);
assign w8624 = w940 & w37256;
assign w8625 = (w342 & w37257) | (w342 & w37258) | (w37257 & w37258);
assign w8626 = ~w8622 & w37259;
assign w8627 = ~w424 & w37260;
assign w8628 = ~w8620 & ~w8627;
assign w8629 = ~w873 & ~w8628;
assign w8630 = w948 & w4749;
assign w8631 = ~w8629 & ~w8630;
assign w8632 = ~w8612 & w8631;
assign w8633 = (w353 & w37261) | (w353 & w37262) | (w37261 & w37262);
assign w8634 = w8633 & w937;
assign w8635 = (pi2646 & w934) | (pi2646 & w37263) | (w934 & w37263);
assign w8636 = w940 & w37264;
assign w8637 = ~w8635 & w37265;
assign w8638 = w905 & w8637;
assign w8639 = ~pi0777 & ~w905;
assign w8640 = (~w8639 & w423) | (~w8639 & w37266) | (w423 & w37266);
assign w8641 = ~w8638 & w8640;
assign w8642 = pi1981 & w1309;
assign w8643 = ~w414 & w37267;
assign w8644 = ~w8642 & ~w8643;
assign w8645 = pi2274 & w1316;
assign w8646 = pi2266 & w1314;
assign w8647 = ~w8645 & ~w8646;
assign w8648 = w8644 & w8647;
assign w8649 = w424 & ~w8648;
assign w8650 = ~w873 & ~w8649;
assign w8651 = ~w8641 & w8650;
assign w8652 = (pi0664 & w508) | (pi0664 & w37268) | (w508 & w37268);
assign w8653 = w508 & ~w514;
assign w8654 = ~w516 & ~w8653;
assign w8655 = ~w8652 & ~w8654;
assign w8656 = (w8655 & ~w797) | (w8655 & w37269) | (~w797 & w37269);
assign w8657 = ~w613 & ~w628;
assign w8658 = ~w624 & ~w629;
assign w8659 = ~w626 & ~w8658;
assign w8660 = w8657 & w8659;
assign w8661 = pi0664 & ~w514;
assign w8662 = (~w8661 & w8657) | (~w8661 & w37270) | (w8657 & w37270);
assign w8663 = ~w8660 & w8662;
assign w8664 = w797 & w37271;
assign w8665 = ~w8656 & ~w8664;
assign w8666 = w874 & w40133;
assign w8667 = (~w8666 & ~w8665) | (~w8666 & w37272) | (~w8665 & w37272);
assign w8668 = ~w414 & w37273;
assign w8669 = ~w405 & w37274;
assign w8670 = ~w8668 & ~w8669;
assign w8671 = ~w371 & w37275;
assign w8672 = ~w392 & w37276;
assign w8673 = ~w8671 & ~w8672;
assign w8674 = w8670 & w8673;
assign w8675 = w423 & ~w8674;
assign w8676 = w873 & ~w8675;
assign w8677 = (w8676 & w8667) | (w8676 & w37277) | (w8667 & w37277);
assign w8678 = ~w8651 & ~w8677;
assign w8679 = ~w517 & ~w528;
assign w8680 = (w797 & w37279) | (w797 & w37280) | (w37279 & w37280);
assign w8681 = (w522 & w798) | (w522 & w37281) | (w798 & w37281);
assign w8682 = (w505 & w37282) | (w505 & w37283) | (w37282 & w37283);
assign w8683 = (~w8682 & w604) | (~w8682 & w37284) | (w604 & w37284);
assign w8684 = (w505 & w37287) | (w505 & w37288) | (w37287 & w37288);
assign w8685 = w514 & w8684;
assign w8686 = ~w8683 & w8685;
assign w8687 = w622 & ~w612;
assign w8688 = ~w604 & w37289;
assign w8689 = ~w8688 & w37290;
assign w8690 = ~w8682 & ~w8687;
assign w8691 = (~w8690 & w613) | (~w8690 & w37291) | (w613 & w37291);
assign w8692 = ~w8691 & w37292;
assign w8693 = ~w617 & w8692;
assign w8694 = w617 & ~w8692;
assign w8695 = ~w8693 & ~w8694;
assign w8696 = w797 & w37293;
assign w8697 = (~w8696 & w8681) | (~w8696 & w37294) | (w8681 & w37294);
assign w8698 = (w874 & w5319) | (w874 & w37295) | (w5319 & w37295);
assign w8699 = (~w8698 & ~w8697) | (~w8698 & w37296) | (~w8697 & w37296);
assign w8700 = ~w371 & w37297;
assign w8701 = ~w392 & w37298;
assign w8702 = ~w8700 & ~w8701;
assign w8703 = ~w414 & w37299;
assign w8704 = (pi1980 & w848) | (pi1980 & w37300) | (w848 & w37300);
assign w8705 = w409 & w8704;
assign w8706 = ~w8703 & ~w8705;
assign w8707 = w8702 & w8706;
assign w8708 = w423 & ~w8707;
assign w8709 = w873 & ~w8708;
assign w8710 = (w8709 & ~w8699) | (w8709 & w37301) | (~w8699 & w37301);
assign w8711 = pi2551 & ~w935;
assign w8712 = (w353 & w37302) | (w353 & w37303) | (w37302 & w37303);
assign w8713 = w940 & w37306;
assign w8714 = (w342 & w37307) | (w342 & w37308) | (w37307 & w37308);
assign w8715 = ~w8711 & w37309;
assign w8716 = ~pi0776 & ~w905;
assign w8717 = (~w8716 & w423) | (~w8716 & w37310) | (w423 & w37310);
assign w8718 = ~w8715 & w8717;
assign w8719 = pi2265 & w1314;
assign w8720 = ~w414 & w37311;
assign w8721 = ~w8719 & ~w8720;
assign w8722 = pi2443 & w1316;
assign w8723 = pi1980 & w1309;
assign w8724 = ~w8722 & ~w8723;
assign w8725 = w8721 & w8724;
assign w8726 = w424 & ~w8725;
assign w8727 = ~w873 & ~w8726;
assign w8728 = ~w8718 & w8727;
assign w8729 = ~w8710 & ~w8728;
assign w8730 = pi0662 & ~w525;
assign w8731 = ~w591 & ~w633;
assign w8732 = ~w634 & ~w8731;
assign w8733 = ~w8730 & ~w8732;
assign w8734 = w797 & w37312;
assign w8735 = ~w523 & ~w528;
assign w8736 = ~pi0507 & w8735;
assign w8737 = pi0507 & ~w8735;
assign w8738 = ~w8736 & ~w8737;
assign w8739 = ~pi0662 & ~w8738;
assign w8740 = w526 & w8738;
assign w8741 = ~w8739 & ~w8740;
assign w8742 = (w8741 & ~w797) | (w8741 & w37313) | (~w797 & w37313);
assign w8743 = ~w8734 & ~w8742;
assign w8744 = (w874 & w4379) | (w874 & w37314) | (w4379 & w37314);
assign w8745 = (~w8744 & ~w8743) | (~w8744 & w37315) | (~w8743 & w37315);
assign w8746 = ~w371 & w37316;
assign w8747 = ~w414 & w37317;
assign w8748 = ~w8746 & ~w8747;
assign w8749 = ~w392 & w37318;
assign w8750 = ~w405 & w37319;
assign w8751 = ~w8749 & ~w8750;
assign w8752 = w8748 & w8751;
assign w8753 = w423 & ~w8752;
assign w8754 = w873 & ~w8753;
assign w8755 = (w8754 & ~w8745) | (w8754 & w37320) | (~w8745 & w37320);
assign w8756 = pi2553 & ~w935;
assign w8757 = (w353 & w37321) | (w353 & w37322) | (w37321 & w37322);
assign w8758 = w940 & w37325;
assign w8759 = (w342 & w37326) | (w342 & w37327) | (w37326 & w37327);
assign w8760 = ~w8756 & w37328;
assign w8761 = ~pi0775 & ~w905;
assign w8762 = (~w8761 & w423) | (~w8761 & w37329) | (w423 & w37329);
assign w8763 = ~w8760 & w8762;
assign w8764 = pi2264 & w1314;
assign w8765 = ~w414 & w37330;
assign w8766 = ~w8764 & ~w8765;
assign w8767 = pi2273 & w1316;
assign w8768 = pi1979 & w1309;
assign w8769 = ~w8767 & ~w8768;
assign w8770 = w8766 & w8769;
assign w8771 = w424 & ~w8770;
assign w8772 = ~w873 & ~w8771;
assign w8773 = ~w8763 & w8772;
assign w8774 = ~w8755 & ~w8773;
assign w8775 = ~w424 & w6446;
assign w8776 = w876 & ~w8775;
assign w8777 = (w8776 & w5969) | (w8776 & w37331) | (w5969 & w37331);
assign w8778 = w937 & w6460;
assign w8779 = (pi2645 & w934) | (pi2645 & w37332) | (w934 & w37332);
assign w8780 = ~w8779 & w37333;
assign w8781 = w905 & ~w8780;
assign w8782 = pi0774 & ~w905;
assign w8783 = (~w8782 & w423) | (~w8782 & w37334) | (w423 & w37334);
assign w8784 = ~w8781 & w8783;
assign w8785 = w424 & w6439;
assign w8786 = ~w873 & ~w8785;
assign w8787 = ~w8784 & w8786;
assign w8788 = w948 & w6413;
assign w8789 = ~w8787 & ~w8788;
assign w8790 = ~w8777 & w8789;
assign w8791 = w2905 & w937;
assign w8792 = (pi2797 & w934) | (pi2797 & w37335) | (w934 & w37335);
assign w8793 = ~w8792 & w37336;
assign w8794 = w905 & w8793;
assign w8795 = ~pi0773 & ~w905;
assign w8796 = (~w8795 & w423) | (~w8795 & w37337) | (w423 & w37337);
assign w8797 = ~w8794 & w8796;
assign w8798 = w424 & ~w2856;
assign w8799 = ~w873 & ~w8798;
assign w8800 = ~w8797 & w8799;
assign w8801 = w874 & w40134;
assign w8802 = (~w8801 & w2415) | (~w8801 & w37338) | (w2415 & w37338);
assign w8803 = w423 & ~w2863;
assign w8804 = w873 & ~w8803;
assign w8805 = (w8804 & w8802) | (w8804 & w37339) | (w8802 & w37339);
assign w8806 = ~w8800 & ~w8805;
assign w8807 = ~w424 & ~w4423;
assign w8808 = w876 & ~w8807;
assign w8809 = (w8808 & w4408) | (w8808 & w37340) | (w4408 & w37340);
assign w8810 = w937 & w4431;
assign w8811 = (pi2644 & w934) | (pi2644 & w37341) | (w934 & w37341);
assign w8812 = ~w8811 & w37342;
assign w8813 = w905 & w8812;
assign w8814 = ~pi0861 & ~w905;
assign w8815 = (~w8814 & w423) | (~w8814 & w37343) | (w423 & w37343);
assign w8816 = ~w8813 & w8815;
assign w8817 = w424 & ~w4416;
assign w8818 = ~w873 & ~w8817;
assign w8819 = ~w8816 & w8818;
assign w8820 = w948 & ~w3195;
assign w8821 = ~w8819 & ~w8820;
assign w8822 = ~w8809 & w8821;
assign w8823 = w6556 & w40111;
assign w8824 = ~w6592 & ~w8823;
assign w8825 = (w874 & w6176) | (w874 & w37344) | (w6176 & w37344);
assign w8826 = (~w8825 & ~w8824) | (~w8825 & w37345) | (~w8824 & w37345);
assign w8827 = w423 & w6538;
assign w8828 = w873 & ~w8827;
assign w8829 = (w8828 & w8826) | (w8828 & w37346) | (w8826 & w37346);
assign w8830 = ~pi0862 & ~w905;
assign w8831 = (pi2796 & w934) | (pi2796 & w37347) | (w934 & w37347);
assign w8832 = (w342 & w37350) | (w342 & w37351) | (w37350 & w37351);
assign w8833 = ~w8831 & w37352;
assign w8834 = ~w8830 & ~w8833;
assign w8835 = ~w424 & ~w8834;
assign w8836 = w424 & w6531;
assign w8837 = ~w873 & ~w8836;
assign w8838 = ~w8835 & w8837;
assign w8839 = ~w8829 & ~w8838;
assign w8840 = ~w424 & w3878;
assign w8841 = w876 & ~w8840;
assign w8842 = (w8841 & w3831) | (w8841 & w37353) | (w3831 & w37353);
assign w8843 = w937 & w3886;
assign w8844 = (pi2794 & w934) | (pi2794 & w37354) | (w934 & w37354);
assign w8845 = ~w8844 & w37355;
assign w8846 = w905 & ~w8845;
assign w8847 = pi0845 & ~w905;
assign w8848 = (~w8847 & w423) | (~w8847 & w37356) | (w423 & w37356);
assign w8849 = ~w8846 & w8848;
assign w8850 = w424 & w3871;
assign w8851 = ~w873 & ~w8850;
assign w8852 = ~w8849 & w8851;
assign w8853 = w948 & w4141;
assign w8854 = ~w8852 & ~w8853;
assign w8855 = ~w8842 & w8854;
assign w8856 = ~w424 & w4826;
assign w8857 = w876 & ~w8856;
assign w8858 = (w8857 & ~w4812) | (w8857 & w37357) | (~w4812 & w37357);
assign w8859 = w937 & w5065;
assign w8860 = (pi2788 & w934) | (pi2788 & w37358) | (w934 & w37358);
assign w8861 = ~w8860 & w37359;
assign w8862 = w905 & ~w8861;
assign w8863 = pi0781 & ~w905;
assign w8864 = (~w8863 & w423) | (~w8863 & w37360) | (w423 & w37360);
assign w8865 = ~w8862 & w8864;
assign w8866 = w424 & w4819;
assign w8867 = ~w873 & ~w8866;
assign w8868 = ~w8865 & w8867;
assign w8869 = w948 & w5053;
assign w8870 = ~w8868 & ~w8869;
assign w8871 = ~w8858 & w8870;
assign w8872 = (w424 & w5414) | (w424 & w37361) | (w5414 & w37361);
assign w8873 = ~w424 & w5650;
assign w8874 = w876 & ~w8873;
assign w8875 = ~w8872 & w8874;
assign w8876 = w5920 & w937;
assign w8877 = (pi2953 & w934) | (pi2953 & w37362) | (w934 & w37362);
assign w8878 = ~w8877 & w37363;
assign w8879 = w905 & ~w8878;
assign w8880 = pi0780 & ~w905;
assign w8881 = (~w8880 & w423) | (~w8880 & w37364) | (w423 & w37364);
assign w8882 = ~w8879 & w8881;
assign w8883 = w424 & w5643;
assign w8884 = ~w873 & ~w8883;
assign w8885 = ~w8882 & w8884;
assign w8886 = w948 & w5635;
assign w8887 = ~w8885 & ~w8886;
assign w8888 = ~w8875 & w8887;
assign w8889 = w2958 & ~w8558;
assign w8890 = w2941 & w3732;
assign w8891 = ~pi0749 & w2899;
assign w8892 = ~w354 & ~w8567;
assign w8893 = w8585 & ~w8892;
assign w8894 = (w2417 & w8892) | (w2417 & w37365) | (w8892 & w37365);
assign w8895 = ~w3774 & w37366;
assign w8896 = w2236 & w37367;
assign w8897 = (~w8573 & ~w359) | (~w8573 & w37369) | (~w359 & w37369);
assign w8898 = ~w2899 & w8897;
assign w8899 = w8572 & w40102;
assign w8900 = (pi1039 & w2907) | (pi1039 & w37370) | (w2907 & w37370);
assign w8901 = ~w8899 & ~w8900;
assign w8902 = w8898 & w8901;
assign w8903 = ~w8895 & w8902;
assign w8904 = ~w8894 & w8903;
assign w8905 = ~w8891 & ~w8904;
assign w8906 = w2961 & w8905;
assign w8907 = ~w8890 & ~w8906;
assign w8908 = (w8907 & w3465) | (w8907 & w37371) | (w3465 & w37371);
assign w8909 = ~w8889 & w8908;
assign w8910 = ~w2397 & ~w8909;
assign w8911 = w3813 & w37372;
assign w8912 = (w2397 & ~w2961) | (w2397 & w37373) | (~w2961 & w37373);
assign w8913 = ~w3775 & w8893;
assign w8914 = w2958 & w8913;
assign w8915 = w3433 & ~w3711;
assign w8916 = ~w8914 & ~w8915;
assign w8917 = w8912 & w8916;
assign w8918 = ~w8911 & w8917;
assign w8919 = ~w8910 & ~w8918;
assign w8920 = w2958 & ~w8602;
assign w8921 = ~w4480 & w37374;
assign w8922 = (~w354 & ~w8608) | (~w354 & w37375) | (~w8608 & w37375);
assign w8923 = w8619 & ~w8922;
assign w8924 = w2236 & w37376;
assign w8925 = (~w8924 & w8923) | (~w8924 & w37377) | (w8923 & w37377);
assign w8926 = (w2365 & ~w8925) | (w2365 & w37378) | (~w8925 & w37378);
assign w8927 = pi1012 & ~w2908;
assign w8928 = (w342 & w37381) | (w342 & w37382) | (w37381 & w37382);
assign w8929 = ~w8927 & w8928;
assign w8930 = (~w2899 & w8926) | (~w2899 & w37383) | (w8926 & w37383);
assign w8931 = pi0778 & w2899;
assign w8932 = w2961 & w37384;
assign w8933 = (~w2397 & ~w2941) | (~w2397 & w37385) | (~w2941 & w37385);
assign w8934 = ~w8932 & w8933;
assign w8935 = (w8934 & ~w4502) | (w8934 & w37386) | (~w4502 & w37386);
assign w8936 = ~w8920 & w8935;
assign w8937 = w1308 & ~w2387;
assign w8938 = w2425 & w4749;
assign w8939 = ~w2958 & ~w8938;
assign w8940 = ~w8937 & w8939;
assign w8941 = ~w4481 & w8923;
assign w8942 = (w2397 & ~w2958) | (w2397 & w37387) | (~w2958 & w37387);
assign w8943 = ~w8940 & w8942;
assign w8944 = (~w8943 & ~w4464) | (~w8943 & w37388) | (~w4464 & w37388);
assign w8945 = ~w8936 & w8944;
assign w8946 = w2941 & ~w5670;
assign w8947 = ~w5949 & w37389;
assign w8948 = (~w354 & ~w8670) | (~w354 & w37390) | (~w8670 & w37390);
assign w8949 = w8648 & ~w8948;
assign w8950 = w2236 & w37391;
assign w8951 = (~w8950 & w8949) | (~w8950 & w37392) | (w8949 & w37392);
assign w8952 = (w2365 & ~w8951) | (w2365 & w37393) | (~w8951 & w37393);
assign w8953 = pi1034 & ~w2908;
assign w8954 = (w342 & w37396) | (w342 & w37397) | (w37396 & w37397);
assign w8955 = ~w8953 & w8954;
assign w8956 = (~w2899 & w8952) | (~w2899 & w37398) | (w8952 & w37398);
assign w8957 = pi0777 & w2899;
assign w8958 = w2961 & w37399;
assign w8959 = ~w8946 & ~w8958;
assign w8960 = (w8959 & w5397) | (w8959 & w37400) | (w5397 & w37400);
assign w8961 = ~w2397 & ~w8960;
assign w8962 = ~w2826 & ~w5429;
assign w8963 = ~w5423 & ~w8962;
assign w8964 = w2961 & ~w5635;
assign w8965 = w3433 & ~w5914;
assign w8966 = ~w5950 & w8949;
assign w8967 = w2958 & w8966;
assign w8968 = ~w8965 & ~w8967;
assign w8969 = ~w8964 & w8968;
assign w8970 = (w8969 & ~w8963) | (w8969 & w37401) | (~w8963 & w37401);
assign w8971 = w3782 & ~w8665;
assign w8972 = (~w8971 & w8970) | (~w8971 & w37402) | (w8970 & w37402);
assign w8973 = ~w8961 & w8972;
assign w8974 = w2941 & w4846;
assign w8975 = w2236 & w37403;
assign w8976 = ~w5359 & w37404;
assign w8977 = (w2365 & w8976) | (w2365 & w37405) | (w8976 & w37405);
assign w8978 = ~w354 & ~w8707;
assign w8979 = w8725 & ~w8978;
assign w8980 = (w2417 & w8978) | (w2417 & w37406) | (w8978 & w37406);
assign w8981 = ~w2899 & ~w8713;
assign w8982 = w8712 & w40102;
assign w8983 = (pi1033 & w2907) | (pi1033 & w37407) | (w2907 & w37407);
assign w8984 = ~w8983 & w37408;
assign w8985 = ~w8980 & w8984;
assign w8986 = ~w8977 & w8985;
assign w8987 = ~pi0776 & w2899;
assign w8988 = w2961 & w37409;
assign w8989 = ~w8974 & ~w8988;
assign w8990 = (w8989 & ~w5377) | (w8989 & w37410) | (~w5377 & w37410);
assign w8991 = ~w2397 & ~w8990;
assign w8992 = w5340 & w37411;
assign w8993 = (w2397 & ~w2961) | (w2397 & w37412) | (~w2961 & w37412);
assign w8994 = ~w5360 & w8979;
assign w8995 = w2958 & w8994;
assign w8996 = w3433 & ~w5320;
assign w8997 = ~w8995 & ~w8996;
assign w8998 = w8993 & w8997;
assign w8999 = ~w8992 & w8998;
assign w9000 = w3782 & ~w8697;
assign w9001 = ~w8999 & ~w9000;
assign w9002 = ~w8991 & w9001;
assign w9003 = ~w2826 & ~w3843;
assign w9004 = ~w3838 & ~w9003;
assign w9005 = w2961 & ~w4141;
assign w9006 = w3433 & ~w4380;
assign w9007 = ~w354 & ~w8752;
assign w9008 = w8770 & ~w9007;
assign w9009 = ~w3911 & w9008;
assign w9010 = w2958 & w9009;
assign w9011 = ~w9006 & ~w9010;
assign w9012 = ~w9005 & w9011;
assign w9013 = (w9012 & ~w9004) | (w9012 & w37413) | (~w9004 & w37413);
assign w9014 = w2397 & ~w9013;
assign w9015 = w3433 & w3934;
assign w9016 = w2236 & w37414;
assign w9017 = (~w2377 & w9007) | (~w2377 & w37415) | (w9007 & w37415);
assign w9018 = (w2365 & w9017) | (w2365 & w37416) | (w9017 & w37416);
assign w9019 = w2363 & w3911;
assign w9020 = ~w2899 & ~w8758;
assign w9021 = w8757 & w40102;
assign w9022 = (~w9021 & w2908) | (~w9021 & w37417) | (w2908 & w37417);
assign w9023 = w9020 & w9022;
assign w9024 = ~w9019 & w9023;
assign w9025 = ~w9018 & w9024;
assign w9026 = ~pi0775 & w2899;
assign w9027 = w2961 & w37418;
assign w9028 = (~w2397 & ~w2941) | (~w2397 & w37419) | (~w2941 & w37419);
assign w9029 = ~w9027 & w9028;
assign w9030 = (w9029 & w8743) | (w9029 & w37420) | (w8743 & w37420);
assign w9031 = ~w9015 & w9030;
assign w9032 = ~w9014 & ~w9031;
assign w9033 = ~w1770 & w6980;
assign w9034 = ~w2227 & w37421;
assign w9035 = ~w2227 & w37422;
assign w9036 = w1770 & ~w7004;
assign w9037 = ~pi2016 & w7004;
assign w9038 = ~w9036 & ~w9037;
assign w9039 = w6687 & w37424;
assign w9040 = (~w9039 & ~w2227) | (~w9039 & w37425) | (~w2227 & w37425);
assign w9041 = ~w9035 & w9040;
assign w9042 = ~w9034 & w9041;
assign w9043 = (w7076 & w37426) | (w7076 & w37427) | (w37426 & w37427);
assign w9044 = (pi0976 & ~w1743) | (pi0976 & w37428) | (~w1743 & w37428);
assign w9045 = ~w1757 & w6988;
assign w9046 = pi1245 & w1040;
assign w9047 = ~w9045 & ~w9046;
assign w9048 = pi1147 & w1037;
assign w9049 = pi1329 & w1043;
assign w9050 = ~w9048 & ~w9049;
assign w9051 = w9047 & w9050;
assign w9052 = pi1044 & ~pi1119;
assign w9053 = w1045 & ~w9052;
assign w9054 = w1766 & w9053;
assign w9055 = pi1161 & w1382;
assign w9056 = pi1133 & w1409;
assign w9057 = pi1273 & w1414;
assign w9058 = ~w9056 & ~w9057;
assign w9059 = ~w9055 & w9058;
assign w9060 = ~w9054 & w9059;
assign w9061 = w9060 & w37429;
assign w9062 = w6984 & ~w9061;
assign w9063 = ~w9043 & ~w9062;
assign w9064 = w9042 & w9063;
assign w9065 = ~w9033 & w9064;
assign w9066 = (pi0408 & ~w342) | (pi0408 & w37430) | (~w342 & w37430);
assign w9067 = w342 & w37431;
assign w9068 = ~w9066 & ~w9067;
assign w9069 = ~w6674 & w9068;
assign w9070 = ~pi3460 & w6674;
assign w9071 = ~w6685 & w37432;
assign w9072 = ~w9069 & w9071;
assign w9073 = pi0749 & w889;
assign w9074 = ~w8572 & ~w9073;
assign w9075 = ~w350 & w37433;
assign w9076 = ~w9072 & ~w9075;
assign w9077 = (w9076 & w9065) | (w9076 & w37434) | (w9065 & w37434);
assign w9078 = ~w1693 & w6980;
assign w9079 = pi1156 & w1382;
assign w9080 = pi1324 & w1043;
assign w9081 = pi1268 & w1414;
assign w9082 = ~w9080 & ~w9081;
assign w9083 = pi1226 & w1046;
assign w9084 = pi1296 & w1678;
assign w9085 = ~w9083 & ~w9084;
assign w9086 = w9082 & w9085;
assign w9087 = ~w9079 & w9086;
assign w9088 = (pi0976 & w1673) | (pi0976 & w37435) | (w1673 & w37435);
assign w9089 = pi1114 & w1416;
assign w9090 = pi1198 & w1385;
assign w9091 = ~w9089 & ~w9090;
assign w9092 = pi1240 & w1040;
assign w9093 = pi1282 & w1390;
assign w9094 = ~w9092 & ~w9093;
assign w9095 = w9091 & w9094;
assign w9096 = pi1184 & w1411;
assign w9097 = pi1254 & w1661;
assign w9098 = ~w9096 & ~w9097;
assign w9099 = pi1142 & w1037;
assign w9100 = pi1170 & w1388;
assign w9101 = ~w9099 & ~w9100;
assign w9102 = w9098 & w9101;
assign w9103 = w9095 & w9102;
assign w9104 = ~w9088 & w9103;
assign w9105 = w9087 & w9104;
assign w9106 = ~w2227 & w37436;
assign w9107 = ~pi3437 & ~pi3460;
assign w9108 = ~w7054 & ~w9107;
assign w9109 = ~w2227 & w37437;
assign w9110 = w1693 & ~w7004;
assign w9111 = ~pi2015 & w7004;
assign w9112 = ~w9110 & ~w9111;
assign w9113 = w6687 & w37439;
assign w9114 = (~w9113 & ~w2227) | (~w9113 & w37440) | (~w2227 & w37440);
assign w9115 = ~w9109 & w9114;
assign w9116 = ~w9106 & w9115;
assign w9117 = ~pi3400 & ~pi3403;
assign w9118 = ~w7078 & ~w9117;
assign w9119 = (w7076 & w37441) | (w7076 & w37442) | (w37441 & w37442);
assign w9120 = ~w2227 & w37443;
assign w9121 = ~w9119 & ~w9120;
assign w9122 = w9116 & w9121;
assign w9123 = ~w9078 & w9122;
assign w9124 = (pi0413 & ~w342) | (pi0413 & w37444) | (~w342 & w37444);
assign w9125 = w342 & w37445;
assign w9126 = ~w9124 & ~w9125;
assign w9127 = ~w6674 & w9126;
assign w9128 = ~pi3437 & w6674;
assign w9129 = ~w6685 & w37446;
assign w9130 = ~w9127 & w9129;
assign w9131 = pi0778 & w889;
assign w9132 = ~w8623 & ~w9131;
assign w9133 = ~w350 & w37447;
assign w9134 = ~w9130 & ~w9133;
assign w9135 = (w9134 & w9123) | (w9134 & w37448) | (w9123 & w37448);
assign w9136 = ~w1957 & w6980;
assign w9137 = ~w2227 & w37449;
assign w9138 = ~pi3433 & ~w7054;
assign w9139 = ~w7055 & ~w9138;
assign w9140 = ~w2227 & w37450;
assign w9141 = w1957 & ~w7004;
assign w9142 = ~pi2014 & w7004;
assign w9143 = ~w9141 & ~w9142;
assign w9144 = w6687 & w37452;
assign w9145 = w347 & w37453;
assign w9146 = ~pi1048 & ~pi1597;
assign w9147 = ~pi3269 & w9146;
assign w9148 = ~pi1330 & ~pi2019;
assign w9149 = ~pi2474 & w9148;
assign w9150 = w9147 & w9149;
assign w9151 = w9145 & ~w9150;
assign w9152 = ~w9144 & ~w9151;
assign w9153 = (w9152 & ~w2227) | (w9152 & w37454) | (~w2227 & w37454);
assign w9154 = ~w9140 & w9153;
assign w9155 = ~w9137 & w9154;
assign w9156 = ~pi3402 & ~w7078;
assign w9157 = ~w7079 & ~w9156;
assign w9158 = (w7076 & w37455) | (w7076 & w37456) | (w37455 & w37456);
assign w9159 = (pi0976 & ~w1936) | (pi0976 & w37457) | (~w1936 & w37457);
assign w9160 = pi1281 & w1390;
assign w9161 = pi1197 & w1385;
assign w9162 = pi1141 & w1037;
assign w9163 = ~w9161 & ~w9162;
assign w9164 = ~w9160 & w9163;
assign w9165 = pi1239 & w1040;
assign w9166 = pi1169 & w1388;
assign w9167 = ~w9165 & ~w9166;
assign w9168 = pi1295 & w1678;
assign w9169 = pi1267 & w1414;
assign w9170 = ~w9168 & ~w9169;
assign w9171 = w9167 & w9170;
assign w9172 = pi1155 & w1382;
assign w9173 = pi1225 & w1046;
assign w9174 = pi1113 & w1416;
assign w9175 = ~w9173 & ~w9174;
assign w9176 = ~w9172 & w9175;
assign w9177 = w9171 & w9176;
assign w9178 = w9164 & w9177;
assign w9179 = ~w9159 & w9178;
assign w9180 = ~w2227 & w37458;
assign w9181 = ~w9158 & ~w9180;
assign w9182 = w9155 & w9181;
assign w9183 = ~w9136 & w9182;
assign w9184 = (pi0412 & ~w342) | (pi0412 & w37459) | (~w342 & w37459);
assign w9185 = w342 & w37460;
assign w9186 = ~w9184 & ~w9185;
assign w9187 = ~w6674 & w9186;
assign w9188 = ~pi3433 & w6674;
assign w9189 = ~w6685 & w37461;
assign w9190 = ~w9187 & w9189;
assign w9191 = pi0777 & w889;
assign w9192 = ~w8633 & ~w9191;
assign w9193 = ~w350 & w37462;
assign w9194 = ~w9190 & ~w9193;
assign w9195 = (w9194 & w9183) | (w9194 & w37463) | (w9183 & w37463);
assign w9196 = ~w2025 & w6980;
assign w9197 = ~w2227 & w37464;
assign w9198 = (~pi3457 & ~w7054) | (~pi3457 & w37465) | (~w7054 & w37465);
assign w9199 = ~w7056 & ~w9198;
assign w9200 = ~w2227 & w37466;
assign w9201 = w2025 & ~w7004;
assign w9202 = ~pi2013 & w7004;
assign w9203 = ~w9201 & ~w9202;
assign w9204 = w6687 & w37468;
assign w9205 = ~pi1049 & ~pi2018;
assign w9206 = ~pi2777 & w9205;
assign w9207 = w9147 & w9206;
assign w9208 = w9145 & ~w9207;
assign w9209 = ~w9204 & ~w9208;
assign w9210 = (w9209 & ~w2227) | (w9209 & w37469) | (~w2227 & w37469);
assign w9211 = ~w9200 & w9210;
assign w9212 = ~w9197 & w9211;
assign w9213 = (~pi3404 & ~w7078) | (~pi3404 & w37470) | (~w7078 & w37470);
assign w9214 = ~w7080 & ~w9213;
assign w9215 = (w7076 & w37471) | (w7076 & w37472) | (w37471 & w37472);
assign w9216 = pi1182 & w1411;
assign w9217 = pi1126 & w1409;
assign w9218 = ~w9216 & ~w9217;
assign w9219 = pi1322 & w1043;
assign w9220 = pi1196 & w1385;
assign w9221 = ~w9219 & ~w9220;
assign w9222 = pi1308 & w1659;
assign w9223 = pi1140 & w1037;
assign w9224 = ~w9222 & ~w9223;
assign w9225 = w9221 & w9224;
assign w9226 = w9218 & w9225;
assign w9227 = (w1024 & ~w2006) | (w1024 & w37473) | (~w2006 & w37473);
assign w9228 = w1045 & ~w2014;
assign w9229 = pi1294 & w1678;
assign w9230 = pi1280 & w1390;
assign w9231 = pi1238 & w1040;
assign w9232 = ~w9230 & ~w9231;
assign w9233 = ~w9229 & w9232;
assign w9234 = ~w9228 & w9233;
assign w9235 = ~w9227 & w9234;
assign w9236 = w9226 & w9235;
assign w9237 = ~w2227 & w37474;
assign w9238 = ~w9215 & ~w9237;
assign w9239 = w9212 & w9238;
assign w9240 = ~w9196 & w9239;
assign w9241 = (pi0411 & ~w342) | (pi0411 & w37475) | (~w342 & w37475);
assign w9242 = w342 & w37476;
assign w9243 = ~w9241 & ~w9242;
assign w9244 = ~w6674 & w9243;
assign w9245 = ~pi3457 & w6674;
assign w9246 = ~w6685 & w37477;
assign w9247 = ~w9244 & w9246;
assign w9248 = pi0776 & w889;
assign w9249 = ~w8712 & ~w9248;
assign w9250 = ~w350 & w37478;
assign w9251 = ~w9247 & ~w9250;
assign w9252 = (w9251 & w9240) | (w9251 & w37479) | (w9240 & w37479);
assign w9253 = ~w1918 & w6980;
assign w9254 = pi1153 & w1382;
assign w9255 = pi1139 & w1037;
assign w9256 = pi1181 & w1411;
assign w9257 = ~w9255 & ~w9256;
assign w9258 = pi1279 & w1390;
assign w9259 = pi1251 & w1661;
assign w9260 = ~w9258 & ~w9259;
assign w9261 = w9257 & w9260;
assign w9262 = ~w9254 & w9261;
assign w9263 = w1045 & ~w1907;
assign w9264 = pi1237 & w1040;
assign w9265 = pi1209 & w1687;
assign w9266 = pi1307 & w1659;
assign w9267 = ~w9265 & ~w9266;
assign w9268 = ~w9264 & w9267;
assign w9269 = pi1125 & w1409;
assign w9270 = pi1321 & w1043;
assign w9271 = ~w9269 & ~w9270;
assign w9272 = pi1195 & w1385;
assign w9273 = pi1293 & w1678;
assign w9274 = ~w9272 & ~w9273;
assign w9275 = w9271 & w9274;
assign w9276 = w9268 & w9275;
assign w9277 = ~w9263 & w9276;
assign w9278 = w9262 & w9277;
assign w9279 = ~w2227 & w37480;
assign w9280 = w1918 & ~w7004;
assign w9281 = ~pi2012 & w7004;
assign w9282 = ~w9280 & ~w9281;
assign w9283 = w2227 & w37481;
assign w9284 = ~pi3456 & ~w7056;
assign w9285 = ~w7057 & ~w9284;
assign w9286 = ~pi2018 & ~pi2019;
assign w9287 = ~pi1048 & ~pi2017;
assign w9288 = w9286 & w9287;
assign w9289 = w9145 & ~w9288;
assign w9290 = w6687 & w37483;
assign w9291 = ~w9289 & ~w9290;
assign w9292 = (w9291 & w2227) | (w9291 & w37484) | (w2227 & w37484);
assign w9293 = ~w9283 & w9292;
assign w9294 = ~w9279 & w9293;
assign w9295 = ~pi3414 & ~w7080;
assign w9296 = ~w7081 & ~w9295;
assign w9297 = (w7076 & w37485) | (w7076 & w37486) | (w37485 & w37486);
assign w9298 = ~w2227 & w37487;
assign w9299 = ~w9297 & ~w9298;
assign w9300 = w9294 & w9299;
assign w9301 = ~w9253 & w9300;
assign w9302 = (pi0410 & ~w342) | (pi0410 & w37488) | (~w342 & w37488);
assign w9303 = w342 & w37489;
assign w9304 = ~w9302 & ~w9303;
assign w9305 = ~w6674 & w9304;
assign w9306 = ~pi3456 & w6674;
assign w9307 = ~w6685 & w37490;
assign w9308 = ~w9305 & w9307;
assign w9309 = pi0775 & w889;
assign w9310 = ~w8757 & ~w9309;
assign w9311 = ~w350 & w37491;
assign w9312 = ~w9308 & ~w9311;
assign w9313 = (w9312 & w9301) | (w9312 & w37492) | (w9301 & w37492);
assign w9314 = ~w2134 & w6980;
assign w9315 = pi0976 & w2116;
assign w9316 = (w1045 & ~w2121) | (w1045 & w37493) | (~w2121 & w37493);
assign w9317 = pi1110 & w1416;
assign w9318 = pi1292 & w1678;
assign w9319 = ~w9317 & ~w9318;
assign w9320 = pi1236 & w1040;
assign w9321 = pi1138 & w1037;
assign w9322 = pi1194 & w1385;
assign w9323 = ~w9321 & ~w9322;
assign w9324 = ~w9320 & w9323;
assign w9325 = w9324 & w37494;
assign w9326 = ~w9315 & w9325;
assign w9327 = ~w2227 & w37495;
assign w9328 = w2134 & ~w7004;
assign w9329 = ~pi2011 & w7004;
assign w9330 = ~w9328 & ~w9329;
assign w9331 = w2227 & w37496;
assign w9332 = (~pi3434 & ~w7056) | (~pi3434 & w37497) | (~w7056 & w37497);
assign w9333 = ~w7058 & ~w9332;
assign w9334 = ~pi1049 & ~pi1330;
assign w9335 = ~pi1598 & ~pi3269;
assign w9336 = w9334 & w9335;
assign w9337 = w9145 & ~w9336;
assign w9338 = w6687 & w37499;
assign w9339 = ~w9337 & ~w9338;
assign w9340 = (w9339 & w2227) | (w9339 & w37500) | (w2227 & w37500);
assign w9341 = ~w9331 & w9340;
assign w9342 = ~w9327 & w9341;
assign w9343 = (~pi3405 & ~w7080) | (~pi3405 & w37501) | (~w7080 & w37501);
assign w9344 = ~w7082 & ~w9343;
assign w9345 = (w7076 & w37502) | (w7076 & w37503) | (w37502 & w37503);
assign w9346 = ~w2227 & w37504;
assign w9347 = ~w9345 & ~w9346;
assign w9348 = w9342 & w9347;
assign w9349 = ~w9314 & w9348;
assign w9350 = (pi0409 & ~w342) | (pi0409 & w37505) | (~w342 & w37505);
assign w9351 = w342 & w37506;
assign w9352 = ~w9350 & ~w9351;
assign w9353 = ~w6674 & w9352;
assign w9354 = ~pi3434 & w6674;
assign w9355 = ~w6685 & w37507;
assign w9356 = ~w9353 & w9355;
assign w9357 = pi0774 & w889;
assign w9358 = ~w6460 & ~w9357;
assign w9359 = ~w350 & w37508;
assign w9360 = ~w9356 & ~w9359;
assign w9361 = (w9360 & w9349) | (w9360 & w37509) | (w9349 & w37509);
assign w9362 = ~w1808 & w6980;
assign w9363 = ~w1783 & w37510;
assign w9364 = w1045 & ~w1800;
assign w9365 = pi1179 & w1411;
assign w9366 = ~w1787 & w6988;
assign w9367 = ~w9365 & ~w9366;
assign w9368 = pi1319 & w1043;
assign w9369 = pi1123 & w1409;
assign w9370 = ~w9368 & ~w9369;
assign w9371 = pi1235 & w1040;
assign w9372 = pi1137 & w1037;
assign w9373 = ~w9371 & ~w9372;
assign w9374 = w9370 & w9373;
assign w9375 = w9367 & w9374;
assign w9376 = w9375 & w37511;
assign w9377 = w6984 & ~w9376;
assign w9378 = (~pi3455 & ~w7056) | (~pi3455 & w37512) | (~w7056 & w37512);
assign w9379 = ~w7059 & ~w9378;
assign w9380 = ~w2227 & w37513;
assign w9381 = w1808 & ~w7004;
assign w9382 = ~pi2374 & w7004;
assign w9383 = ~w9381 & ~w9382;
assign w9384 = w6687 & w37515;
assign w9385 = (~w9384 & ~w2227) | (~w9384 & w37516) | (~w2227 & w37516);
assign w9386 = ~w9380 & w9385;
assign w9387 = ~w9377 & w9386;
assign w9388 = (~pi3413 & ~w7080) | (~pi3413 & w37517) | (~w7080 & w37517);
assign w9389 = ~w7083 & ~w9388;
assign w9390 = (w7076 & w37518) | (w7076 & w37519) | (w37518 & w37519);
assign w9391 = ~w2227 & w37520;
assign w9392 = ~w9390 & ~w9391;
assign w9393 = w9387 & w9392;
assign w9394 = ~w9362 & w9393;
assign w9395 = (pi0426 & ~w342) | (pi0426 & w37521) | (~w342 & w37521);
assign w9396 = w342 & w37522;
assign w9397 = ~w9395 & ~w9396;
assign w9398 = ~w6674 & w9397;
assign w9399 = ~pi3455 & w6674;
assign w9400 = ~w6685 & w37523;
assign w9401 = ~w9398 & w9400;
assign w9402 = pi0773 & w889;
assign w9403 = ~w2905 & ~w9402;
assign w9404 = ~w350 & w37524;
assign w9405 = ~w9401 & ~w9404;
assign w9406 = (w9405 & w9394) | (w9405 & w37525) | (w9394 & w37525);
assign w9407 = ~w1731 & w6980;
assign w9408 = pi0976 & ~w1706;
assign w9409 = pi1234 & w1040;
assign w9410 = pi1136 & w1037;
assign w9411 = pi1108 & w1416;
assign w9412 = ~w9410 & ~w9411;
assign w9413 = ~w9409 & w9412;
assign w9414 = pi1220 & w1046;
assign w9415 = pi1290 & w1678;
assign w9416 = ~w9414 & ~w9415;
assign w9417 = pi1192 & w1385;
assign w9418 = pi1122 & w1409;
assign w9419 = ~w9417 & ~w9418;
assign w9420 = pi1276 & w1390;
assign w9421 = pi1043 & w1045;
assign w9422 = ~w1716 & w9421;
assign w9423 = ~w9420 & ~w9422;
assign w9424 = w9419 & w9423;
assign w9425 = w9416 & w9424;
assign w9426 = w9413 & w9425;
assign w9427 = ~w9408 & w9426;
assign w9428 = ~w2227 & w37526;
assign w9429 = ~pi3454 & ~w7059;
assign w9430 = ~w7060 & ~w9429;
assign w9431 = ~w2227 & w37527;
assign w9432 = w1731 & ~w7004;
assign w9433 = ~pi2010 & w7004;
assign w9434 = ~w9432 & ~w9433;
assign w9435 = w6687 & w37529;
assign w9436 = (~w9435 & ~w2227) | (~w9435 & w37530) | (~w2227 & w37530);
assign w9437 = ~w9431 & w9436;
assign w9438 = ~w9428 & w9437;
assign w9439 = ~pi3406 & ~w7083;
assign w9440 = ~w7084 & ~w9439;
assign w9441 = (w7076 & w37531) | (w7076 & w37532) | (w37531 & w37532);
assign w9442 = ~w2227 & w37533;
assign w9443 = ~w9441 & ~w9442;
assign w9444 = w9438 & w9443;
assign w9445 = ~w9407 & w9444;
assign w9446 = (pi0425 & ~w342) | (pi0425 & w37534) | (~w342 & w37534);
assign w9447 = w342 & w37535;
assign w9448 = ~w9446 & ~w9447;
assign w9449 = ~w6674 & w9448;
assign w9450 = ~pi3454 & w6674;
assign w9451 = ~w6685 & w37536;
assign w9452 = ~w9449 & w9451;
assign w9453 = pi0861 & w889;
assign w9454 = ~w4431 & ~w9453;
assign w9455 = ~w350 & w37537;
assign w9456 = ~w9452 & ~w9455;
assign w9457 = (w9456 & w9445) | (w9456 & w37538) | (w9445 & w37538);
assign w9458 = ~w2167 & w6980;
assign w9459 = pi1149 & w1382;
assign w9460 = pi1205 & w1687;
assign w9461 = pi1135 & w1037;
assign w9462 = ~w9460 & ~w9461;
assign w9463 = pi1317 & w1043;
assign w9464 = pi1107 & w1416;
assign w9465 = ~w9463 & ~w9464;
assign w9466 = w9462 & w9465;
assign w9467 = ~w9459 & w9466;
assign w9468 = pi1303 & w1659;
assign w9469 = pi1163 & w1388;
assign w9470 = pi1219 & w1046;
assign w9471 = ~w9469 & ~w9470;
assign w9472 = ~w9468 & w9471;
assign w9473 = pi1233 & w1040;
assign w9474 = pi1275 & w1390;
assign w9475 = ~w9473 & ~w9474;
assign w9476 = pi1247 & w1661;
assign w9477 = pi1121 & w1409;
assign w9478 = ~w9476 & ~w9477;
assign w9479 = w9475 & w9478;
assign w9480 = pi1289 & w1678;
assign w9481 = pi1261 & w1414;
assign w9482 = ~w9480 & ~w9481;
assign w9483 = pi1191 & w1385;
assign w9484 = pi1177 & w1411;
assign w9485 = ~w9483 & ~w9484;
assign w9486 = w9482 & w9485;
assign w9487 = w9479 & w9486;
assign w9488 = w9472 & w9487;
assign w9489 = w9467 & w9488;
assign w9490 = ~w2227 & w37539;
assign w9491 = (~pi3453 & ~w7059) | (~pi3453 & w37540) | (~w7059 & w37540);
assign w9492 = ~w7061 & ~w9491;
assign w9493 = ~w2227 & w37541;
assign w9494 = w2167 & ~w7004;
assign w9495 = ~pi2373 & w7004;
assign w9496 = ~w9494 & ~w9495;
assign w9497 = w6687 & w37543;
assign w9498 = (~w9497 & ~w2227) | (~w9497 & w37544) | (~w2227 & w37544);
assign w9499 = ~w9493 & w9498;
assign w9500 = ~w9490 & w9499;
assign w9501 = (~pi3411 & ~w7083) | (~pi3411 & w37545) | (~w7083 & w37545);
assign w9502 = ~w7085 & ~w9501;
assign w9503 = (w7076 & w37546) | (w7076 & w37547) | (w37546 & w37547);
assign w9504 = ~w2227 & w37548;
assign w9505 = ~w9503 & ~w9504;
assign w9506 = w9500 & w9505;
assign w9507 = ~w9458 & w9506;
assign w9508 = (pi0406 & ~w342) | (pi0406 & w37549) | (~w342 & w37549);
assign w9509 = w342 & w37550;
assign w9510 = ~w9508 & ~w9509;
assign w9511 = ~w6674 & w9510;
assign w9512 = ~pi3453 & w6674;
assign w9513 = ~w6685 & w37551;
assign w9514 = ~w9511 & w9513;
assign w9515 = pi0862 & w889;
assign w9516 = ~w6566 & ~w9515;
assign w9517 = ~w350 & w37552;
assign w9518 = ~w9514 & ~w9517;
assign w9519 = (w9518 & w9507) | (w9518 & w37553) | (w9507 & w37553);
assign w9520 = ~w2060 & w6980;
assign w9521 = pi0976 & ~w2038;
assign w9522 = w1045 & ~w2049;
assign w9523 = pi1288 & w1678;
assign w9524 = pi1274 & w1390;
assign w9525 = ~w9523 & ~w9524;
assign w9526 = pi1232 & w1040;
assign w9527 = pi1120 & w1409;
assign w9528 = ~w9526 & ~w9527;
assign w9529 = pi1134 & w1037;
assign w9530 = pi1190 & w1385;
assign w9531 = ~w9529 & ~w9530;
assign w9532 = w9528 & w9531;
assign w9533 = w9525 & w9532;
assign w9534 = ~w9522 & w9533;
assign w9535 = ~w9521 & w9534;
assign w9536 = ~w2227 & w37554;
assign w9537 = (~pi3432 & ~w7059) | (~pi3432 & w37555) | (~w7059 & w37555);
assign w9538 = ~w7062 & ~w9537;
assign w9539 = ~w2227 & w37556;
assign w9540 = w2060 & ~w7004;
assign w9541 = ~pi2392 & w7004;
assign w9542 = ~w9540 & ~w9541;
assign w9543 = w6687 & w37558;
assign w9544 = (~w9543 & ~w2227) | (~w9543 & w37559) | (~w2227 & w37559);
assign w9545 = ~w9539 & w9544;
assign w9546 = ~w9536 & w9545;
assign w9547 = (~pi3420 & ~w7083) | (~pi3420 & w37560) | (~w7083 & w37560);
assign w9548 = ~w7086 & ~w9547;
assign w9549 = (w7076 & w37561) | (w7076 & w37562) | (w37561 & w37562);
assign w9550 = ~w2227 & w37563;
assign w9551 = ~w9549 & ~w9550;
assign w9552 = w9546 & w9551;
assign w9553 = ~w9520 & w9552;
assign w9554 = (pi0424 & ~w342) | (pi0424 & w37564) | (~w342 & w37564);
assign w9555 = w342 & w37565;
assign w9556 = ~w9554 & ~w9555;
assign w9557 = ~w6674 & w9556;
assign w9558 = ~pi3432 & w6674;
assign w9559 = ~w6685 & w37566;
assign w9560 = ~w9557 & w9559;
assign w9561 = pi0845 & w889;
assign w9562 = ~w3886 & ~w9561;
assign w9563 = ~w350 & w37567;
assign w9564 = ~w9560 & ~w9563;
assign w9565 = (w9564 & w9553) | (w9564 & w37568) | (w9553 & w37568);
assign w9566 = ~w1845 & w6980;
assign w9567 = pi1146 & w1037;
assign w9568 = pi1188 & w1411;
assign w9569 = ~w9567 & ~w9568;
assign w9570 = pi1244 & w1040;
assign w9571 = pi1272 & w1414;
assign w9572 = ~w9570 & ~w9571;
assign w9573 = ~pi1044 & w1045;
assign w9574 = ~w1825 & w9573;
assign w9575 = pi1132 & w1409;
assign w9576 = ~w9574 & ~w9575;
assign w9577 = w9572 & w9576;
assign w9578 = w9569 & w9577;
assign w9579 = w1024 & ~w1837;
assign w9580 = pi1328 & w1043;
assign w9581 = pi1118 & w1416;
assign w9582 = ~w9580 & ~w9581;
assign w9583 = pi1286 & w1390;
assign w9584 = ~w1818 & w6988;
assign w9585 = ~w9583 & ~w9584;
assign w9586 = w9582 & w9585;
assign w9587 = ~w9579 & w9586;
assign w9588 = w9578 & w9587;
assign w9589 = ~w2227 & w37569;
assign w9590 = (~pi3459 & ~w7059) | (~pi3459 & w37570) | (~w7059 & w37570);
assign w9591 = ~w7063 & ~w9590;
assign w9592 = ~w2227 & w37571;
assign w9593 = w1845 & ~w7004;
assign w9594 = ~pi2378 & w7004;
assign w9595 = ~w9593 & ~w9594;
assign w9596 = w6687 & w37573;
assign w9597 = (~w9596 & ~w2227) | (~w9596 & w37574) | (~w2227 & w37574);
assign w9598 = ~w9592 & w9597;
assign w9599 = ~w9589 & w9598;
assign w9600 = (~pi3401 & ~w7083) | (~pi3401 & w37575) | (~w7083 & w37575);
assign w9601 = ~w7087 & ~w9600;
assign w9602 = (w7076 & w37576) | (w7076 & w37577) | (w37576 & w37577);
assign w9603 = ~w2227 & w37578;
assign w9604 = ~w9602 & ~w9603;
assign w9605 = w9599 & w9604;
assign w9606 = ~w9566 & w9605;
assign w9607 = (pi0423 & ~w342) | (pi0423 & w37579) | (~w342 & w37579);
assign w9608 = w342 & w37580;
assign w9609 = ~w9607 & ~w9608;
assign w9610 = ~w6674 & w9609;
assign w9611 = ~pi3459 & w6674;
assign w9612 = ~w6685 & w37581;
assign w9613 = ~w9610 & w9612;
assign w9614 = pi0781 & w889;
assign w9615 = ~w5065 & ~w9614;
assign w9616 = ~w350 & w37582;
assign w9617 = ~w9613 & ~w9616;
assign w9618 = (w9617 & w9606) | (w9617 & w37583) | (w9606 & w37583);
assign w9619 = ~w1879 & w6980;
assign w9620 = ~w2227 & w37584;
assign w9621 = ~pi3478 & ~w7063;
assign w9622 = ~w7064 & ~w9621;
assign w9623 = ~w2227 & w37585;
assign w9624 = w1879 & ~w7004;
assign w9625 = ~pi2377 & w7004;
assign w9626 = ~w9624 & ~w9625;
assign w9627 = pi0816 & w7068;
assign w9628 = (~w9627 & ~w2227) | (~w9627 & w37587) | (~w2227 & w37587);
assign w9629 = ~w9623 & w9628;
assign w9630 = ~w9620 & w9629;
assign w9631 = ~pi3422 & ~w7087;
assign w9632 = ~w7088 & ~w9631;
assign w9633 = (w7076 & w37588) | (w7076 & w37589) | (w37588 & w37589);
assign w9634 = pi1201 & w1385;
assign w9635 = pi1243 & w1040;
assign w9636 = ~w9634 & ~w9635;
assign w9637 = pi1257 & w1661;
assign w9638 = pi1313 & w1659;
assign w9639 = ~w9637 & ~w9638;
assign w9640 = w9636 & w9639;
assign w9641 = pi1159 & w1382;
assign w9642 = pi1327 & w1043;
assign w9643 = pi1299 & w1678;
assign w9644 = ~w9642 & ~w9643;
assign w9645 = ~w9641 & w9644;
assign w9646 = w9640 & w9645;
assign w9647 = pi1271 & w1414;
assign w9648 = pi1131 & w1409;
assign w9649 = ~w9647 & ~w9648;
assign w9650 = pi1285 & w1390;
assign w9651 = pi1117 & w1416;
assign w9652 = ~w9650 & ~w9651;
assign w9653 = w9649 & w9652;
assign w9654 = pi1215 & w1687;
assign w9655 = ~w1859 & w9573;
assign w9656 = ~w9654 & ~w9655;
assign w9657 = pi1187 & w1411;
assign w9658 = pi1145 & w1037;
assign w9659 = ~w9657 & ~w9658;
assign w9660 = w9656 & w9659;
assign w9661 = w9653 & w9660;
assign w9662 = w9646 & w9661;
assign w9663 = ~w2227 & w37590;
assign w9664 = ~w9633 & ~w9663;
assign w9665 = w9630 & w9664;
assign w9666 = ~w9619 & w9665;
assign w9667 = (pi0422 & ~w342) | (pi0422 & w37591) | (~w342 & w37591);
assign w9668 = w342 & w37592;
assign w9669 = ~w9667 & ~w9668;
assign w9670 = ~w6674 & w9669;
assign w9671 = ~pi3478 & w6674;
assign w9672 = ~w6685 & w37593;
assign w9673 = ~w9670 & w9672;
assign w9674 = pi0780 & w889;
assign w9675 = ~w5920 & ~w9674;
assign w9676 = ~w350 & w37594;
assign w9677 = ~w9673 & ~w9676;
assign w9678 = (w9677 & w9666) | (w9677 & w37595) | (w9666 & w37595);
assign w9679 = ~pi0434 & w938;
assign w9680 = pi0393 & ~w7234;
assign w9681 = (~w938 & ~w7234) | (~w938 & w37596) | (~w7234 & w37596);
assign w9682 = ~w9680 & w9681;
assign w9683 = ~w9679 & ~w9682;
assign w9684 = (w353 & w37597) | (w353 & w37598) | (w37597 & w37598);
assign w9685 = pi0390 & ~w7234;
assign w9686 = (~w938 & ~w7234) | (~w938 & w37599) | (~w7234 & w37599);
assign w9687 = ~w9685 & w9686;
assign w9688 = ~w9684 & ~w9687;
assign w9689 = (w353 & w37600) | (w353 & w37601) | (w37600 & w37601);
assign w9690 = pi0389 & ~w7234;
assign w9691 = (~w938 & ~w7234) | (~w938 & w37602) | (~w7234 & w37602);
assign w9692 = ~w9690 & w9691;
assign w9693 = ~w9689 & ~w9692;
assign w9694 = (w353 & w37603) | (w353 & w37604) | (w37603 & w37604);
assign w9695 = pi0388 & ~w7234;
assign w9696 = (~w938 & ~w7234) | (~w938 & w37605) | (~w7234 & w37605);
assign w9697 = ~w9695 & w9696;
assign w9698 = ~w9694 & ~w9697;
assign w9699 = (w353 & w37606) | (w353 & w37607) | (w37606 & w37607);
assign w9700 = pi0387 & ~w7234;
assign w9701 = (~w938 & ~w7234) | (~w938 & w37608) | (~w7234 & w37608);
assign w9702 = ~w9700 & w9701;
assign w9703 = ~w9699 & ~w9702;
assign w9704 = (w353 & w37609) | (w353 & w37610) | (w37609 & w37610);
assign w9705 = pi0386 & ~w7234;
assign w9706 = (~w938 & ~w7234) | (~w938 & w37611) | (~w7234 & w37611);
assign w9707 = ~w9705 & w9706;
assign w9708 = ~w9704 & ~w9707;
assign w9709 = (w353 & w37612) | (w353 & w37613) | (w37612 & w37613);
assign w9710 = pi0385 & ~w7234;
assign w9711 = (~w938 & ~w7234) | (~w938 & w37614) | (~w7234 & w37614);
assign w9712 = ~w9710 & w9711;
assign w9713 = ~w9709 & ~w9712;
assign w9714 = (w353 & w37615) | (w353 & w37616) | (w37615 & w37616);
assign w9715 = pi0384 & ~w7234;
assign w9716 = (~w938 & ~w7234) | (~w938 & w37617) | (~w7234 & w37617);
assign w9717 = ~w9715 & w9716;
assign w9718 = ~w9714 & ~w9717;
assign w9719 = (w353 & w37618) | (w353 & w37619) | (w37618 & w37619);
assign w9720 = pi0383 & ~w7234;
assign w9721 = (~w938 & ~w7234) | (~w938 & w37620) | (~w7234 & w37620);
assign w9722 = ~w9720 & w9721;
assign w9723 = ~w9719 & ~w9722;
assign w9724 = (w353 & w37621) | (w353 & w37622) | (w37621 & w37622);
assign w9725 = pi0382 & ~w7234;
assign w9726 = (~w938 & ~w7234) | (~w938 & w37623) | (~w7234 & w37623);
assign w9727 = ~w9725 & w9726;
assign w9728 = ~w9724 & ~w9727;
assign w9729 = (w353 & w37624) | (w353 & w37625) | (w37624 & w37625);
assign w9730 = pi0392 & ~w7234;
assign w9731 = (~w938 & ~w7234) | (~w938 & w37626) | (~w7234 & w37626);
assign w9732 = ~w9730 & w9731;
assign w9733 = ~w9729 & ~w9732;
assign w9734 = (w353 & w37627) | (w353 & w37628) | (w37627 & w37628);
assign w9735 = pi0391 & ~w7234;
assign w9736 = (~w938 & ~w7234) | (~w938 & w37629) | (~w7234 & w37629);
assign w9737 = ~w9735 & w9736;
assign w9738 = ~w9734 & ~w9737;
assign w9739 = (w353 & w37630) | (w353 & w37631) | (w37630 & w37631);
assign w9740 = pi0381 & ~w7234;
assign w9741 = (~w938 & ~w7234) | (~w938 & w37632) | (~w7234 & w37632);
assign w9742 = ~w9740 & w9741;
assign w9743 = ~w9739 & ~w9742;
assign w9744 = (w353 & w37633) | (w353 & w37634) | (w37633 & w37634);
assign w9745 = pi0378 & ~w7234;
assign w9746 = (~w938 & ~w7234) | (~w938 & w37635) | (~w7234 & w37635);
assign w9747 = ~w9745 & w9746;
assign w9748 = ~w9744 & ~w9747;
assign w9749 = (w353 & w37636) | (w353 & w37637) | (w37636 & w37637);
assign w9750 = pi0377 & ~w7234;
assign w9751 = (~w938 & ~w7234) | (~w938 & w37638) | (~w7234 & w37638);
assign w9752 = ~w9750 & w9751;
assign w9753 = ~w9749 & ~w9752;
assign w9754 = (w353 & w37639) | (w353 & w37640) | (w37639 & w37640);
assign w9755 = pi0376 & ~w7234;
assign w9756 = (~w938 & ~w7234) | (~w938 & w37641) | (~w7234 & w37641);
assign w9757 = ~w9755 & w9756;
assign w9758 = ~w9754 & ~w9757;
assign w9759 = (w353 & w37642) | (w353 & w37643) | (w37642 & w37643);
assign w9760 = pi0375 & ~w7234;
assign w9761 = (~w938 & ~w7234) | (~w938 & w37644) | (~w7234 & w37644);
assign w9762 = ~w9760 & w9761;
assign w9763 = ~w9759 & ~w9762;
assign w9764 = (w353 & w37645) | (w353 & w37646) | (w37645 & w37646);
assign w9765 = pi0374 & ~w7234;
assign w9766 = (~w938 & ~w7234) | (~w938 & w37647) | (~w7234 & w37647);
assign w9767 = ~w9765 & w9766;
assign w9768 = ~w9764 & ~w9767;
assign w9769 = (w353 & w37648) | (w353 & w37649) | (w37648 & w37649);
assign w9770 = pi0373 & ~w7234;
assign w9771 = (~w938 & ~w7234) | (~w938 & w37650) | (~w7234 & w37650);
assign w9772 = ~w9770 & w9771;
assign w9773 = ~w9769 & ~w9772;
assign w9774 = (w353 & w37651) | (w353 & w37652) | (w37651 & w37652);
assign w9775 = pi0372 & ~w7234;
assign w9776 = (~w938 & ~w7234) | (~w938 & w37653) | (~w7234 & w37653);
assign w9777 = ~w9775 & w9776;
assign w9778 = ~w9774 & ~w9777;
assign w9779 = (w353 & w37654) | (w353 & w37655) | (w37654 & w37655);
assign w9780 = pi0371 & ~w7234;
assign w9781 = (~w938 & ~w7234) | (~w938 & w37656) | (~w7234 & w37656);
assign w9782 = ~w9780 & w9781;
assign w9783 = ~w9779 & ~w9782;
assign w9784 = (w353 & w37657) | (w353 & w37658) | (w37657 & w37658);
assign w9785 = pi0369 & ~w7234;
assign w9786 = (~w938 & ~w7234) | (~w938 & w37659) | (~w7234 & w37659);
assign w9787 = ~w9785 & w9786;
assign w9788 = ~w9784 & ~w9787;
assign w9789 = (w353 & w37660) | (w353 & w37661) | (w37660 & w37661);
assign w9790 = pi0380 & ~w7234;
assign w9791 = (~w938 & ~w7234) | (~w938 & w37662) | (~w7234 & w37662);
assign w9792 = ~w9790 & w9791;
assign w9793 = ~w9789 & ~w9792;
assign w9794 = (w353 & w37663) | (w353 & w37664) | (w37663 & w37664);
assign w9795 = pi0379 & ~w7234;
assign w9796 = (~w938 & ~w7234) | (~w938 & w37665) | (~w7234 & w37665);
assign w9797 = ~w9795 & w9796;
assign w9798 = ~w9794 & ~w9797;
assign w9799 = ~w6683 & w9065;
assign w9800 = w342 & w37666;
assign w9801 = ~w9799 & ~w9800;
assign w9802 = ~w6683 & w9123;
assign w9803 = w342 & w37667;
assign w9804 = ~w9802 & ~w9803;
assign w9805 = ~w6683 & w9183;
assign w9806 = w342 & w37668;
assign w9807 = ~w9805 & ~w9806;
assign w9808 = ~w6683 & w9240;
assign w9809 = w342 & w37669;
assign w9810 = ~w9808 & ~w9809;
assign w9811 = ~w6683 & w9301;
assign w9812 = w342 & w37670;
assign w9813 = ~w9811 & ~w9812;
assign w9814 = pi3114 & ~w2214;
assign w9815 = (w2211 & w37671) | (w2211 & w37672) | (w37671 & w37672);
assign w9816 = ~pi3118 & ~w9815;
assign w9817 = ~w9814 & ~w9816;
assign w9818 = pi3118 & ~w9815;
assign w9819 = ~w9814 & ~w9818;
assign w9820 = pi2763 & pi2951;
assign w9821 = ~pi2763 & pi2952;
assign w9822 = ~w9820 & ~w9821;
assign w9823 = ~pi3209 & ~w9822;
assign w9824 = pi3208 & ~w9822;
assign w9825 = pi3405 & w9822;
assign w9826 = ~w9824 & ~w9825;
assign w9827 = pi3235 & ~w9822;
assign w9828 = pi3413 & w9822;
assign w9829 = ~w9827 & ~w9828;
assign w9830 = pi3234 & ~w9822;
assign w9831 = pi3406 & w9822;
assign w9832 = ~w9830 & ~w9831;
assign w9833 = pi3207 & ~w9822;
assign w9834 = pi3411 & w9822;
assign w9835 = ~w9833 & ~w9834;
assign w9836 = pi3206 & ~w9822;
assign w9837 = pi3420 & w9822;
assign w9838 = ~w9836 & ~w9837;
assign w9839 = pi3231 & ~w9822;
assign w9840 = pi3401 & w9822;
assign w9841 = ~w9839 & ~w9840;
assign w9842 = pi3230 & ~w9822;
assign w9843 = pi3422 & w9822;
assign w9844 = ~w9842 & ~w9843;
assign w9845 = pi3229 & ~w9822;
assign w9846 = pi3421 & w9822;
assign w9847 = ~w9845 & ~w9846;
assign w9848 = pi3228 & ~w9822;
assign w9849 = pi3430 & w9822;
assign w9850 = ~w9848 & ~w9849;
assign w9851 = (w2211 & w37673) | (w2211 & w37674) | (w37673 & w37674);
assign w9852 = (pi3121 & ~w341) | (pi3121 & w37675) | (~w341 & w37675);
assign w9853 = ~w9851 & w9852;
assign w9854 = ~pi0939 & pi1930;
assign w9855 = ~pi2492 & w9854;
assign w9856 = pi3195 & w9821;
assign w9857 = (~w2214 & ~w2174) | (~w2214 & w37676) | (~w2174 & w37676);
assign w9858 = ~w9857 & w37677;
assign w9859 = pi2763 & w40135;
assign w9860 = ~w9858 & w9859;
assign w9861 = ~w9856 & ~w9860;
assign w9862 = pi3124 & w9821;
assign w9863 = (~w9112 & w9857) | (~w9112 & w37679) | (w9857 & w37679);
assign w9864 = (pi2763 & w9857) | (pi2763 & w37681) | (w9857 & w37681);
assign w9865 = ~w9863 & w9864;
assign w9866 = ~w9862 & ~w9865;
assign w9867 = pi3194 & w9821;
assign w9868 = (~w9143 & w9857) | (~w9143 & w37682) | (w9857 & w37682);
assign w9869 = (pi2763 & w9857) | (pi2763 & w37684) | (w9857 & w37684);
assign w9870 = ~w9868 & w9869;
assign w9871 = ~w9867 & ~w9870;
assign w9872 = pi3139 & w9821;
assign w9873 = (~w9203 & w9857) | (~w9203 & w37685) | (w9857 & w37685);
assign w9874 = (pi2763 & w9857) | (pi2763 & w37687) | (w9857 & w37687);
assign w9875 = ~w9873 & w9874;
assign w9876 = ~w9872 & ~w9875;
assign w9877 = pi3135 & w9821;
assign w9878 = (~w9282 & w9857) | (~w9282 & w37688) | (w9857 & w37688);
assign w9879 = (pi2763 & w9857) | (pi2763 & w37690) | (w9857 & w37690);
assign w9880 = ~w9878 & w9879;
assign w9881 = ~w9877 & ~w9880;
assign w9882 = pi3187 & w9821;
assign w9883 = (~w9330 & w9857) | (~w9330 & w37691) | (w9857 & w37691);
assign w9884 = (pi2763 & w9857) | (pi2763 & w37693) | (w9857 & w37693);
assign w9885 = ~w9883 & w9884;
assign w9886 = ~w9882 & ~w9885;
assign w9887 = pi3193 & w9821;
assign w9888 = ~w9857 & w37694;
assign w9889 = pi2763 & w40136;
assign w9890 = ~w9888 & w9889;
assign w9891 = ~w9887 & ~w9890;
assign w9892 = pi3192 & w9821;
assign w9893 = ~w9857 & w37696;
assign w9894 = pi2763 & w40137;
assign w9895 = ~w9893 & w9894;
assign w9896 = ~w9892 & ~w9895;
assign w9897 = pi3117 & w9821;
assign w9898 = ~w9857 & w37698;
assign w9899 = pi2763 & w40138;
assign w9900 = ~w9898 & w9899;
assign w9901 = ~w9897 & ~w9900;
assign w9902 = pi3116 & w9821;
assign w9903 = (~w9542 & w9857) | (~w9542 & w37700) | (w9857 & w37700);
assign w9904 = (pi2763 & w9857) | (pi2763 & w37702) | (w9857 & w37702);
assign w9905 = ~w9903 & w9904;
assign w9906 = ~w9902 & ~w9905;
assign w9907 = pi3198 & w9821;
assign w9908 = (~w9595 & w9857) | (~w9595 & w37703) | (w9857 & w37703);
assign w9909 = (pi2763 & w9857) | (pi2763 & w37705) | (w9857 & w37705);
assign w9910 = ~w9908 & w9909;
assign w9911 = ~w9907 & ~w9910;
assign w9912 = pi3115 & w9821;
assign w9913 = (~w9626 & w9857) | (~w9626 & w37706) | (w9857 & w37706);
assign w9914 = (pi2763 & w9857) | (pi2763 & w37708) | (w9857 & w37708);
assign w9915 = ~w9913 & w9914;
assign w9916 = ~w9912 & ~w9915;
assign w9917 = pi3197 & w9821;
assign w9918 = (~w7007 & w9857) | (~w7007 & w37709) | (w9857 & w37709);
assign w9919 = (pi2763 & w9857) | (pi2763 & w37711) | (w9857 & w37711);
assign w9920 = ~w9918 & w9919;
assign w9921 = ~w9917 & ~w9920;
assign w9922 = pi3196 & w9821;
assign w9923 = (~w7117 & w9857) | (~w7117 & w37712) | (w9857 & w37712);
assign w9924 = ~w9857 & w37713;
assign w9925 = pi2763 & ~w9924;
assign w9926 = ~w9923 & w9925;
assign w9927 = ~w9922 & ~w9926;
assign w9928 = ~w7004 & ~w9820;
assign w9929 = ~w370 & ~w9928;
assign w9930 = ~pi3509 & ~pi3517;
assign w9931 = pi3508 & w9930;
assign w9932 = ~w8220 & w9931;
assign w9933 = pi3509 & pi3517;
assign w9934 = ~pi3508 & w9933;
assign w9935 = ~w1143 & w9934;
assign w9936 = ~w9932 & ~w9935;
assign w9937 = ~pi3509 & pi3517;
assign w9938 = ~pi3508 & w9937;
assign w9939 = ~w8157 & w9938;
assign w9940 = pi3509 & ~pi3517;
assign w9941 = pi3508 & w9940;
assign w9942 = ~w8172 & w9941;
assign w9943 = ~w9939 & ~w9942;
assign w9944 = pi3508 & w9937;
assign w9945 = ~w8203 & w9944;
assign w9946 = pi3508 & w9933;
assign w9947 = ~w8195 & w9946;
assign w9948 = ~w9945 & ~w9947;
assign w9949 = w9943 & w9948;
assign w9950 = pi3509 & w8215;
assign w9951 = ~pi3508 & ~pi3517;
assign w9952 = (w9951 & ~w8224) | (w9951 & w37714) | (~w8224 & w37714);
assign w9953 = ~w9950 & w9952;
assign w9954 = w9949 & w37715;
assign w9955 = ~pi1974 & ~pi1975;
assign w9956 = ~pi1972 & ~pi1973;
assign w9957 = w9955 & w9956;
assign w9958 = pi2758 & pi3065;
assign w9959 = pi2142 & w9958;
assign w9960 = ~pi0143 & ~pi3065;
assign w9961 = ~w9959 & ~w9960;
assign w9962 = pi1974 & pi1975;
assign w9963 = ~pi3065 & w9962;
assign w9964 = ~pi1972 & pi1973;
assign w9965 = ~w9963 & w9964;
assign w9966 = (w9954 & w37717) | (w9954 & w37718) | (w37717 & w37718);
assign w9967 = ~w9956 & w37719;
assign w9968 = (pi1974 & w9967) | (pi1974 & w37720) | (w9967 & w37720);
assign w9969 = ~w9959 & ~w9968;
assign w9970 = ~w7982 & w9931;
assign w9971 = ~w9935 & ~w9970;
assign w9972 = ~w7958 & w9944;
assign w9973 = ~w7927 & w9941;
assign w9974 = ~w9972 & ~w9973;
assign w9975 = ~w7942 & w9938;
assign w9976 = ~w7950 & w9946;
assign w9977 = ~w9975 & ~w9976;
assign w9978 = w9974 & w9977;
assign w9979 = pi3509 & w7974;
assign w9980 = (w9951 & ~w7969) | (w9951 & w37714) | (~w7969 & w37714);
assign w9981 = ~w9979 & w9980;
assign w9982 = w9978 & w37721;
assign w9983 = w9969 & ~w9982;
assign w9984 = ~w9966 & w9983;
assign w9985 = w9966 & ~w9983;
assign w9986 = ~w9984 & ~w9985;
assign w9987 = pi1972 & ~pi1973;
assign w9988 = ~w9959 & ~w9987;
assign w9989 = ~pi1972 & w9955;
assign w9990 = ~w9959 & ~w9989;
assign w9991 = ~pi3510 & ~pi3511;
assign w9992 = ~pi3520 & ~pi3521;
assign w9993 = w9991 & w9992;
assign w9994 = ~pi2982 & ~w9993;
assign w9995 = w9990 & w9994;
assign w9996 = ~pi1794 & w9995;
assign w9997 = w9990 & ~w9994;
assign w9998 = pi0242 & pi0979;
assign w9999 = ~pi3516 & pi3518;
assign w10000 = pi0244 & ~pi0979;
assign w10001 = w9999 & ~w10000;
assign w10002 = ~w9998 & w10001;
assign w10003 = ~pi3516 & ~pi3518;
assign w10004 = ~w7965 & w10003;
assign w10005 = pi3516 & ~pi3518;
assign w10006 = ~w7978 & w10005;
assign w10007 = ~w10004 & ~w10006;
assign w10008 = ~w10002 & w10007;
assign w10009 = w9997 & ~w10008;
assign w10010 = ~w10009 & w37722;
assign w10011 = (w9988 & w10009) | (w9988 & w37723) | (w10009 & w37723);
assign w10012 = ~w10010 & ~w10011;
assign w10013 = ~w9986 & w10012;
assign w10014 = ~w1449 & w9931;
assign w10015 = ~w9935 & ~w10014;
assign w10016 = ~w1509 & w9938;
assign w10017 = ~w1548 & w9944;
assign w10018 = ~w10016 & ~w10017;
assign w10019 = ~w1517 & w9941;
assign w10020 = ~w1540 & w9946;
assign w10021 = ~w10019 & ~w10020;
assign w10022 = w10018 & w10021;
assign w10023 = pi3509 & w1432;
assign w10024 = (w9951 & ~w1441) | (w9951 & w37714) | (~w1441 & w37714);
assign w10025 = ~w10023 & w10024;
assign w10026 = w10022 & w37724;
assign w10027 = w9969 & ~w10026;
assign w10028 = ~w9966 & w10027;
assign w10029 = w9966 & ~w10027;
assign w10030 = ~w10028 & ~w10029;
assign w10031 = ~pi1795 & w9995;
assign w10032 = pi0243 & pi0979;
assign w10033 = pi0245 & ~pi0979;
assign w10034 = w9999 & ~w10033;
assign w10035 = ~w10032 & w10034;
assign w10036 = ~w1436 & w10005;
assign w10037 = ~w1445 & w10003;
assign w10038 = ~w10036 & ~w10037;
assign w10039 = ~w10035 & w10038;
assign w10040 = w9997 & ~w10039;
assign w10041 = (w9987 & w10040) | (w9987 & w37725) | (w10040 & w37725);
assign w10042 = ~w10040 & w37726;
assign w10043 = ~w10041 & ~w10042;
assign w10044 = w10030 & w10043;
assign w10045 = ~w9954 & w9969;
assign w10046 = ~w9966 & w10045;
assign w10047 = w9966 & ~w10045;
assign w10048 = ~w10046 & ~w10047;
assign w10049 = ~w9993 & w37727;
assign w10050 = ~w8211 & w10003;
assign w10051 = ~w9994 & ~w10050;
assign w10052 = pi0230 & pi0979;
assign w10053 = pi0231 & ~pi0979;
assign w10054 = w9999 & ~w10053;
assign w10055 = ~w10052 & w10054;
assign w10056 = ~w8228 & w10005;
assign w10057 = ~w10055 & ~w10056;
assign w10058 = w10051 & w10057;
assign w10059 = (w9988 & w10058) | (w9988 & w37729) | (w10058 & w37729);
assign w10060 = ~w10058 & w37730;
assign w10061 = ~w10059 & ~w10060;
assign w10062 = ~w10048 & ~w10061;
assign w10063 = ~w1191 & w9944;
assign w10064 = ~w9935 & ~w10063;
assign w10065 = ~w1147 & w9941;
assign w10066 = ~w1136 & w9931;
assign w10067 = ~w10065 & ~w10066;
assign w10068 = ~w1187 & w9946;
assign w10069 = ~w1161 & w9938;
assign w10070 = ~w10068 & ~w10069;
assign w10071 = w10067 & w10070;
assign w10072 = pi3509 & w1123;
assign w10073 = (w9951 & ~w1119) | (w9951 & w37714) | (~w1119 & w37714);
assign w10074 = ~w10072 & w10073;
assign w10075 = w10071 & w37731;
assign w10076 = w9969 & ~w10075;
assign w10077 = ~w9966 & w10076;
assign w10078 = w9966 & ~w10076;
assign w10079 = ~w10077 & ~w10078;
assign w10080 = ~pi1796 & w9995;
assign w10081 = pi0273 & pi0979;
assign w10082 = pi0275 & ~pi0979;
assign w10083 = w9999 & ~w10082;
assign w10084 = ~w10081 & w10083;
assign w10085 = ~w1132 & w10003;
assign w10086 = ~w1128 & w10005;
assign w10087 = ~w10085 & ~w10086;
assign w10088 = ~w10084 & w10087;
assign w10089 = w9997 & ~w10088;
assign w10090 = ~w10089 & w37732;
assign w10091 = (w9988 & w10089) | (w9988 & w37733) | (w10089 & w37733);
assign w10092 = ~w10090 & ~w10091;
assign w10093 = w10079 & ~w10092;
assign w10094 = ~w10062 & w10093;
assign w10095 = ~w10044 & ~w10094;
assign w10096 = (~w10013 & w10094) | (~w10013 & w37734) | (w10094 & w37734);
assign w10097 = w9986 & ~w10012;
assign w10098 = ~w10096 & ~w10097;
assign w10099 = ~w9955 & w9956;
assign w10100 = ~w10048 & w37735;
assign w10101 = ~w10048 & w37736;
assign w10102 = (w10101 & w10096) | (w10101 & w37737) | (w10096 & w37737);
assign w10103 = ~w10030 & ~w10043;
assign w10104 = ~w10079 & w10092;
assign w10105 = ~w10103 & ~w10104;
assign w10106 = ~w10013 & w10105;
assign w10107 = w10105 & w37738;
assign w10108 = pi0828 & w10107;
assign w10109 = ~w10102 & ~w10108;
assign w10110 = ~w3060 & w9941;
assign w10111 = ~w9935 & ~w10110;
assign w10112 = ~w3108 & w9946;
assign w10113 = ~w3075 & w9938;
assign w10114 = ~w10112 & ~w10113;
assign w10115 = ~w3083 & w9931;
assign w10116 = ~w3112 & w9944;
assign w10117 = ~w10115 & ~w10116;
assign w10118 = w10114 & w10117;
assign w10119 = pi3509 & w3101;
assign w10120 = (w9951 & ~w3092) | (w9951 & w37714) | (~w3092 & w37714);
assign w10121 = ~w10119 & w10120;
assign w10122 = w10118 & w37739;
assign w10123 = w9969 & ~w10122;
assign w10124 = ~w9966 & w10123;
assign w10125 = w9966 & ~w10123;
assign w10126 = ~w10124 & ~w10125;
assign w10127 = ~pi2195 & w9995;
assign w10128 = pi0325 & pi0979;
assign w10129 = pi0326 & ~pi0979;
assign w10130 = w9999 & ~w10129;
assign w10131 = ~w10128 & w10130;
assign w10132 = ~w3088 & w10003;
assign w10133 = ~w3097 & w10005;
assign w10134 = ~w10132 & ~w10133;
assign w10135 = ~w10131 & w10134;
assign w10136 = w9997 & ~w10135;
assign w10137 = ~w10136 & w37740;
assign w10138 = (w9988 & w10136) | (w9988 & w37741) | (w10136 & w37741);
assign w10139 = ~w10137 & ~w10138;
assign w10140 = w10126 & ~w10139;
assign w10141 = ~w6304 & w9946;
assign w10142 = ~w9944 & ~w10141;
assign w10143 = ~pi3509 & w6308;
assign w10144 = ~w10142 & ~w10143;
assign w10145 = w6316 & w9933;
assign w10146 = (~pi3508 & ~w6330) | (~pi3508 & w37742) | (~w6330 & w37742);
assign w10147 = ~w10145 & w10146;
assign w10148 = ~w6270 & w9930;
assign w10149 = ~w6320 & w9940;
assign w10150 = ~w10148 & ~w10149;
assign w10151 = ~w10147 & w10150;
assign w10152 = ~w10144 & w10151;
assign w10153 = ~pi3509 & ~w6279;
assign w10154 = (w9951 & w6288) | (w9951 & w37743) | (w6288 & w37743);
assign w10155 = ~w10153 & w10154;
assign w10156 = w9969 & ~w10155;
assign w10157 = ~w10152 & w10156;
assign w10158 = ~w9966 & w10157;
assign w10159 = w9966 & ~w10157;
assign w10160 = ~w10158 & ~w10159;
assign w10161 = ~pi2197 & w9995;
assign w10162 = pi0338 & pi0979;
assign w10163 = pi0340 & ~pi0979;
assign w10164 = w9999 & ~w10163;
assign w10165 = ~w10162 & w10164;
assign w10166 = ~w6275 & w10003;
assign w10167 = ~w6284 & w10005;
assign w10168 = ~w10166 & ~w10167;
assign w10169 = ~w10165 & w10168;
assign w10170 = w9997 & ~w10169;
assign w10171 = (w9987 & w10170) | (w9987 & w37744) | (w10170 & w37744);
assign w10172 = ~w10170 & w37745;
assign w10173 = ~w10171 & ~w10172;
assign w10174 = ~w10160 & ~w10173;
assign w10175 = pi0348 & ~pi0979;
assign w10176 = pi0346 & pi0979;
assign w10177 = w9999 & ~w10176;
assign w10178 = ~w10175 & w10177;
assign w10179 = ~w4298 & w10003;
assign w10180 = ~w4302 & w10005;
assign w10181 = ~w10179 & ~w10180;
assign w10182 = (w9990 & ~w10181) | (w9990 & w37746) | (~w10181 & w37746);
assign w10183 = ~w9987 & w10182;
assign w10184 = (~w9995 & w10182) | (~w9995 & w37747) | (w10182 & w37747);
assign w10185 = ~w10183 & w10184;
assign w10186 = ~w9959 & w9994;
assign w10187 = ~pi2079 & ~w9987;
assign w10188 = pi2079 & w9987;
assign w10189 = ~w10187 & ~w10188;
assign w10190 = w10186 & w10189;
assign w10191 = ~w10185 & ~w10190;
assign w10192 = ~w4323 & w9946;
assign w10193 = ~w4331 & w9944;
assign w10194 = ~w10192 & ~w10193;
assign w10195 = ~w4339 & w9938;
assign w10196 = ~w4366 & w9934;
assign w10197 = ~w10195 & ~w10196;
assign w10198 = ~w4357 & w9941;
assign w10199 = ~w4293 & w9931;
assign w10200 = ~w10198 & ~w10199;
assign w10201 = w10197 & w10200;
assign w10202 = ~pi3509 & w4311;
assign w10203 = (w9951 & ~w4307) | (w9951 & w37743) | (~w4307 & w37743);
assign w10204 = ~w10202 & w10203;
assign w10205 = w10201 & w37748;
assign w10206 = w9969 & ~w10205;
assign w10207 = ~w9966 & w10206;
assign w10208 = w9966 & ~w10206;
assign w10209 = ~w10207 & ~w10208;
assign w10210 = ~w10191 & ~w10209;
assign w10211 = (~pi3508 & ~w5119) | (~pi3508 & w37749) | (~w5119 & w37749);
assign w10212 = ~w5179 & w9930;
assign w10213 = ~w10211 & ~w10212;
assign w10214 = w5123 & w9937;
assign w10215 = ~w10213 & ~w10214;
assign w10216 = ~w5204 & w9946;
assign w10217 = ~w9944 & ~w10216;
assign w10218 = ~pi3509 & w5200;
assign w10219 = ~w5129 & w9940;
assign w10220 = (~w10219 & w10217) | (~w10219 & w37750) | (w10217 & w37750);
assign w10221 = ~w10215 & w10220;
assign w10222 = ~pi3509 & ~w5175;
assign w10223 = (w9951 & w5188) | (w9951 & w37743) | (w5188 & w37743);
assign w10224 = ~w10222 & w10223;
assign w10225 = w9969 & ~w10224;
assign w10226 = ~w10221 & w10225;
assign w10227 = ~w9966 & w10226;
assign w10228 = w9966 & ~w10226;
assign w10229 = ~w10227 & ~w10228;
assign w10230 = ~pi2199 & w9995;
assign w10231 = pi0347 & pi0979;
assign w10232 = pi0349 & ~pi0979;
assign w10233 = w9999 & ~w10232;
assign w10234 = ~w10231 & w10233;
assign w10235 = ~w5192 & w10005;
assign w10236 = ~w5183 & w10003;
assign w10237 = ~w10235 & ~w10236;
assign w10238 = ~w10234 & w10237;
assign w10239 = w9997 & ~w10238;
assign w10240 = (w9987 & w10239) | (w9987 & w37751) | (w10239 & w37751);
assign w10241 = ~w10239 & w37752;
assign w10242 = ~w10240 & ~w10241;
assign w10243 = ~w10229 & ~w10242;
assign w10244 = ~w5767 & w9946;
assign w10245 = ~w5703 & w9941;
assign w10246 = ~w10244 & ~w10245;
assign w10247 = ~w5718 & w9938;
assign w10248 = ~w5783 & w9931;
assign w10249 = ~w10247 & ~w10248;
assign w10250 = ~w5758 & w9944;
assign w10251 = ~w5695 & w9934;
assign w10252 = ~w10250 & ~w10251;
assign w10253 = w10249 & w10252;
assign w10254 = pi3509 & w5796;
assign w10255 = (w9951 & ~w5792) | (w9951 & w37714) | (~w5792 & w37714);
assign w10256 = ~w10254 & w10255;
assign w10257 = w10253 & w37753;
assign w10258 = w9969 & ~w10257;
assign w10259 = ~w9966 & w10258;
assign w10260 = w9966 & ~w10258;
assign w10261 = ~w10259 & ~w10260;
assign w10262 = ~w9993 & w37754;
assign w10263 = ~w5778 & w10003;
assign w10264 = ~w9994 & ~w10263;
assign w10265 = pi0401 & pi0979;
assign w10266 = pi0402 & ~pi0979;
assign w10267 = w9999 & ~w10266;
assign w10268 = ~w10265 & w10267;
assign w10269 = ~w5787 & w10005;
assign w10270 = ~w10268 & ~w10269;
assign w10271 = w10264 & w10270;
assign w10272 = (w9988 & w10271) | (w9988 & w37755) | (w10271 & w37755);
assign w10273 = ~w9987 & ~w9989;
assign w10274 = ~w9959 & ~w10273;
assign w10275 = ~w10271 & w37756;
assign w10276 = ~w10272 & ~w10275;
assign w10277 = ~w10261 & ~w10276;
assign w10278 = (pi3516 & w4734) | (pi3516 & w37757) | (w4734 & w37757);
assign w10279 = ~pi0437 & ~pi0979;
assign w10280 = ~pi0436 & pi0979;
assign w10281 = pi3518 & ~w10280;
assign w10282 = ~w10279 & w10281;
assign w10283 = w4716 & w10003;
assign w10284 = w9990 & ~w10283;
assign w10285 = w10284 & w37758;
assign w10286 = ~w9987 & w10285;
assign w10287 = (~w9995 & w10285) | (~w9995 & w37747) | (w10285 & w37747);
assign w10288 = ~w10286 & w10287;
assign w10289 = ~pi2083 & ~w9987;
assign w10290 = pi2083 & w9987;
assign w10291 = ~w10289 & ~w10290;
assign w10292 = w10186 & w10291;
assign w10293 = ~w10288 & ~w10292;
assign w10294 = ~w4661 & w9946;
assign w10295 = ~w4721 & w9931;
assign w10296 = ~w10294 & ~w10295;
assign w10297 = ~w4695 & w9938;
assign w10298 = ~w4685 & w9941;
assign w10299 = ~w10297 & ~w10298;
assign w10300 = ~w4689 & w9934;
assign w10301 = ~w4657 & w9944;
assign w10302 = ~w10300 & ~w10301;
assign w10303 = w10299 & w10302;
assign w10304 = pi3509 & w4725;
assign w10305 = (w9951 & ~w4730) | (w9951 & w37714) | (~w4730 & w37714);
assign w10306 = ~w10304 & w10305;
assign w10307 = w10303 & w37759;
assign w10308 = w9969 & ~w10307;
assign w10309 = ~w9966 & w10308;
assign w10310 = w9966 & ~w10308;
assign w10311 = ~w10309 & ~w10310;
assign w10312 = w10293 & w10311;
assign w10313 = ~pi3509 & w3613;
assign w10314 = (~pi3508 & ~w3627) | (~pi3508 & w37760) | (~w3627 & w37760);
assign w10315 = ~w10313 & w10314;
assign w10316 = (~w9951 & w3588) | (~w9951 & w37761) | (w3588 & w37761);
assign w10317 = ~w3576 & w9946;
assign w10318 = ~w3580 & w9944;
assign w10319 = ~w3631 & w9940;
assign w10320 = ~w10318 & ~w10319;
assign w10321 = w10320 & w37762;
assign w10322 = ~w10315 & w10321;
assign w10323 = pi3509 & ~w3602;
assign w10324 = (w9951 & w3597) | (w9951 & w37714) | (w3597 & w37714);
assign w10325 = ~w10323 & w10324;
assign w10326 = w9969 & ~w10325;
assign w10327 = ~w10322 & w10326;
assign w10328 = ~w9966 & w10327;
assign w10329 = w9966 & ~w10327;
assign w10330 = ~w10328 & ~w10329;
assign w10331 = ~w9993 & w37763;
assign w10332 = ~w3593 & w10003;
assign w10333 = ~w9994 & ~w10332;
assign w10334 = pi0463 & pi0979;
assign w10335 = pi0464 & ~pi0979;
assign w10336 = w9999 & ~w10335;
assign w10337 = ~w10334 & w10336;
assign w10338 = ~w3606 & w10005;
assign w10339 = ~w10337 & ~w10338;
assign w10340 = w10333 & w10339;
assign w10341 = (w9988 & w10340) | (w9988 & w37764) | (w10340 & w37764);
assign w10342 = ~w10340 & w37765;
assign w10343 = ~w10341 & ~w10342;
assign w10344 = w10330 & w10343;
assign w10345 = ~w10293 & ~w10311;
assign w10346 = pi1973 & w9955;
assign w10347 = pi0196 & ~pi1974;
assign w10348 = pi1975 & ~w10347;
assign w10349 = ~w9956 & ~w10348;
assign w10350 = ~w10346 & w10349;
assign w10351 = (w9954 & w37766) | (w9954 & w37767) | (w37766 & w37767);
assign w10352 = ~w10345 & ~w10351;
assign w10353 = ~w10330 & ~w10343;
assign w10354 = (~w10353 & w10352) | (~w10353 & w37768) | (w10352 & w37768);
assign w10355 = (w10354 & w37770) | (w10354 & w37771) | (w37770 & w37771);
assign w10356 = w10229 & w10242;
assign w10357 = w10261 & w10276;
assign w10358 = ~w10174 & w10357;
assign w10359 = ~w10356 & ~w10358;
assign w10360 = (~w10210 & w10355) | (~w10210 & w37772) | (w10355 & w37772);
assign w10361 = w3335 & w9933;
assign w10362 = (~pi3508 & ~w3350) | (~pi3508 & w37742) | (~w3350 & w37742);
assign w10363 = ~w10361 & w10362;
assign w10364 = ~w3396 & w9946;
assign w10365 = ~w3387 & w9944;
assign w10366 = ~w10364 & ~w10365;
assign w10367 = ~w3367 & w9930;
assign w10368 = ~w3354 & w9940;
assign w10369 = ~w10367 & ~w10368;
assign w10370 = w10366 & w10369;
assign w10371 = ~w10363 & w10370;
assign w10372 = ~pi3509 & ~w3371;
assign w10373 = (w9951 & w3376) | (w9951 & w37743) | (w3376 & w37743);
assign w10374 = ~w10372 & w10373;
assign w10375 = w9969 & ~w10374;
assign w10376 = ~w10371 & w10375;
assign w10377 = ~w9966 & w10376;
assign w10378 = w9966 & ~w10376;
assign w10379 = ~w10377 & ~w10378;
assign w10380 = ~w9993 & w37773;
assign w10381 = ~w3362 & w10003;
assign w10382 = ~w9994 & ~w10381;
assign w10383 = pi0339 & ~pi0979;
assign w10384 = pi0337 & pi0979;
assign w10385 = w9999 & ~w10384;
assign w10386 = ~w10383 & w10385;
assign w10387 = ~w3380 & w10005;
assign w10388 = ~w10386 & ~w10387;
assign w10389 = w10382 & w10388;
assign w10390 = (w9988 & w10389) | (w9988 & w37774) | (w10389 & w37774);
assign w10391 = ~w10389 & w37775;
assign w10392 = ~w10390 & ~w10391;
assign w10393 = w10379 & w10392;
assign w10394 = w10160 & w10173;
assign w10395 = w10191 & w10209;
assign w10396 = ~w10243 & w10395;
assign w10397 = ~w10394 & ~w10396;
assign w10398 = ~w10396 & w37776;
assign w10399 = ~w10126 & w10139;
assign w10400 = ~w10379 & ~w10392;
assign w10401 = ~w10399 & ~w10400;
assign w10402 = (w10360 & w37778) | (w10360 & w37779) | (w37778 & w37779);
assign w10403 = ~w10140 & ~w10402;
assign w10404 = ~w9993 & w37780;
assign w10405 = ~pi0302 & w9999;
assign w10406 = pi2916 & w10005;
assign w10407 = ~w10405 & ~w10406;
assign w10408 = ~pi0979 & ~w10407;
assign w10409 = ~pi0301 & w9999;
assign w10410 = pi2144 & w10005;
assign w10411 = ~w10409 & ~w10410;
assign w10412 = pi0979 & ~w10411;
assign w10413 = ~w4068 & w10003;
assign w10414 = ~w9994 & ~w10413;
assign w10415 = ~w10412 & w10414;
assign w10416 = (~w10404 & ~w10415) | (~w10404 & w37781) | (~w10415 & w37781);
assign w10417 = w9987 & ~w10416;
assign w10418 = (~w9959 & ~w10416) | (~w9959 & w10274) | (~w10416 & w10274);
assign w10419 = ~w10417 & w10418;
assign w10420 = ~w4023 & w9938;
assign w10421 = ~w9935 & ~w10420;
assign w10422 = ~w4042 & w9941;
assign w10423 = ~w4075 & w9944;
assign w10424 = ~w10422 & ~w10423;
assign w10425 = ~w4083 & w9946;
assign w10426 = ~w4064 & w9931;
assign w10427 = ~w10425 & ~w10426;
assign w10428 = w10424 & w10427;
assign w10429 = w10421 & w10428;
assign w10430 = ~pi2931 & pi3509;
assign w10431 = ~pi2939 & ~pi3509;
assign w10432 = ~pi0979 & ~w10431;
assign w10433 = ~w10430 & w10432;
assign w10434 = ~pi2161 & pi3509;
assign w10435 = ~pi2177 & ~pi3509;
assign w10436 = pi0979 & ~w10435;
assign w10437 = ~w10434 & w10436;
assign w10438 = ~w10433 & ~w10437;
assign w10439 = w9951 & ~w10438;
assign w10440 = (w9969 & ~w10429) | (w9969 & w37782) | (~w10429 & w37782);
assign w10441 = ~w9966 & w10440;
assign w10442 = w9966 & ~w10440;
assign w10443 = ~w10441 & ~w10442;
assign w10444 = w10419 & ~w10443;
assign w10445 = ~w6091 & w9944;
assign w10446 = ~w9935 & ~w10445;
assign w10447 = ~w6060 & w9938;
assign w10448 = ~w6111 & w9931;
assign w10449 = ~w10447 & ~w10448;
assign w10450 = ~w6087 & w9946;
assign w10451 = ~w6056 & w9941;
assign w10452 = ~w10450 & ~w10451;
assign w10453 = w10449 & w10452;
assign w10454 = pi3509 & w6119;
assign w10455 = (w9951 & ~w6102) | (w9951 & w37714) | (~w6102 & w37714);
assign w10456 = ~w10454 & w10455;
assign w10457 = w10453 & w37783;
assign w10458 = w9969 & ~w10457;
assign w10459 = ~w9966 & w10458;
assign w10460 = w9966 & ~w10458;
assign w10461 = ~w10459 & ~w10460;
assign w10462 = ~pi2086 & w9995;
assign w10463 = pi0322 & ~pi0979;
assign w10464 = pi0321 & pi0979;
assign w10465 = w9999 & ~w10464;
assign w10466 = ~w10463 & w10465;
assign w10467 = ~w6106 & w10005;
assign w10468 = ~w6115 & w10003;
assign w10469 = ~w10467 & ~w10468;
assign w10470 = ~w10466 & w10469;
assign w10471 = w9997 & ~w10470;
assign w10472 = ~w10471 & w37784;
assign w10473 = (w9988 & w10471) | (w9988 & w37785) | (w10471 & w37785);
assign w10474 = ~w10472 & ~w10473;
assign w10475 = ~w10461 & w10474;
assign w10476 = ~w10444 & ~w10475;
assign w10477 = ~w5566 & w9931;
assign w10478 = ~w9935 & ~w10477;
assign w10479 = ~w5605 & w9941;
assign w10480 = ~w5613 & w9946;
assign w10481 = ~w10479 & ~w10480;
assign w10482 = ~w5590 & w9938;
assign w10483 = ~w5617 & w9944;
assign w10484 = ~w10482 & ~w10483;
assign w10485 = w10481 & w10484;
assign w10486 = pi3509 & w5570;
assign w10487 = (w9951 & ~w5574) | (w9951 & w37714) | (~w5574 & w37714);
assign w10488 = ~w10486 & w10487;
assign w10489 = w10485 & w37786;
assign w10490 = w9969 & ~w10489;
assign w10491 = ~w9966 & w10490;
assign w10492 = w9966 & ~w10490;
assign w10493 = ~w10491 & ~w10492;
assign w10494 = ~w9993 & w37787;
assign w10495 = ~w5557 & w10003;
assign w10496 = ~w9994 & ~w10495;
assign w10497 = pi0274 & pi0979;
assign w10498 = pi0276 & ~pi0979;
assign w10499 = w9999 & ~w10498;
assign w10500 = ~w10497 & w10499;
assign w10501 = ~w5561 & w10005;
assign w10502 = ~w10500 & ~w10501;
assign w10503 = w10496 & w10502;
assign w10504 = (w9988 & w10503) | (w9988 & w37788) | (w10503 & w37788);
assign w10505 = ~w10503 & w37789;
assign w10506 = ~w10504 & ~w10505;
assign w10507 = w10493 & w10506;
assign w10508 = ~w4962 & w9931;
assign w10509 = ~w9935 & ~w10508;
assign w10510 = ~w4933 & w9944;
assign w10511 = ~w4973 & w9941;
assign w10512 = ~w10510 & ~w10511;
assign w10513 = ~w4977 & w9938;
assign w10514 = ~w4941 & w9946;
assign w10515 = ~w10513 & ~w10514;
assign w10516 = w10512 & w10515;
assign w10517 = ~pi3509 & w4966;
assign w10518 = (w9951 & ~w4953) | (w9951 & w37743) | (~w4953 & w37743);
assign w10519 = ~w10517 & w10518;
assign w10520 = w10516 & w37790;
assign w10521 = w9969 & ~w10520;
assign w10522 = ~w9966 & w10521;
assign w10523 = w9966 & ~w10521;
assign w10524 = ~w10522 & ~w10523;
assign w10525 = ~pi2080 & w9995;
assign w10526 = pi0295 & pi0979;
assign w10527 = pi0296 & ~pi0979;
assign w10528 = w9999 & ~w10527;
assign w10529 = ~w10526 & w10528;
assign w10530 = ~w4958 & w10005;
assign w10531 = ~w4949 & w10003;
assign w10532 = ~w10530 & ~w10531;
assign w10533 = ~w10529 & w10532;
assign w10534 = w9997 & ~w10533;
assign w10535 = ~w10534 & w37791;
assign w10536 = (w9988 & w10534) | (w9988 & w37792) | (w10534 & w37792);
assign w10537 = ~w10535 & ~w10536;
assign w10538 = w10524 & ~w10537;
assign w10539 = ~w10444 & w10538;
assign w10540 = ~w10507 & ~w10539;
assign w10541 = ~w10493 & ~w10506;
assign w10542 = ~w10524 & w10537;
assign w10543 = ~w10541 & ~w10542;
assign w10544 = (w10476 & ~w10540) | (w10476 & w37793) | (~w10540 & w37793);
assign w10545 = ~w10419 & w10443;
assign w10546 = w10461 & ~w10474;
assign w10547 = ~w10541 & w10546;
assign w10548 = ~w10545 & ~w10547;
assign w10549 = w10543 & ~w10548;
assign w10550 = w10540 & ~w10549;
assign w10551 = ~w10102 & w10550;
assign w10552 = (w10551 & w10403) | (w10551 & w37794) | (w10403 & w37794);
assign w10553 = ~w10109 & ~w10552;
assign w10554 = pi3210 & ~w2214;
assign w10555 = ~pi2487 & ~pi3330;
assign w10556 = ~w10554 & ~w10555;
assign w10557 = pi3394 & ~w10554;
assign w10558 = ~w10556 & ~w10557;
assign w10559 = pi1042 & pi1093;
assign w10560 = pi1588 & w10559;
assign w10561 = ~pi1042 & ~pi1093;
assign w10562 = pi1540 & w10561;
assign w10563 = ~w10560 & ~w10562;
assign w10564 = pi1042 & ~pi1093;
assign w10565 = pi1557 & w10564;
assign w10566 = ~pi1042 & pi1093;
assign w10567 = pi1625 & w10566;
assign w10568 = ~w10565 & ~w10567;
assign w10569 = w10563 & w10568;
assign w10570 = pi1041 & ~w10569;
assign w10571 = (~pi1041 & ~w10566) | (~pi1041 & w37796) | (~w10566 & w37796);
assign w10572 = ~pi1521 & w10559;
assign w10573 = ~pi1485 & w10564;
assign w10574 = ~w10572 & ~w10573;
assign w10575 = w10571 & w10574;
assign w10576 = ~w10570 & ~w10575;
assign w10577 = w10558 & w10576;
assign w10578 = (~w10577 & w4748) | (~w10577 & w37797) | (w4748 & w37797);
assign w10579 = w10106 & w10544;
assign w10580 = w10578 & w10579;
assign w10581 = ~w10403 & w10580;
assign w10582 = w10048 & w10061;
assign w10583 = w10048 & w37798;
assign w10584 = (w10106 & w10549) | (w10106 & w37799) | (w10549 & w37799);
assign w10585 = ~w10584 & w37800;
assign w10586 = (w10578 & ~w10585) | (w10578 & w37801) | (~w10585 & w37801);
assign w10587 = ~w10581 & ~w10586;
assign w10588 = w10553 & ~w10587;
assign w10589 = w10107 & w10544;
assign w10590 = (w10589 & w10402) | (w10589 & w37802) | (w10402 & w37802);
assign w10591 = (w10100 & w10584) | (w10100 & w37803) | (w10584 & w37803);
assign w10592 = ~w10590 & ~w10591;
assign w10593 = pi1974 & w9956;
assign w10594 = w9956 & w9962;
assign w10595 = (~w10594 & w10048) | (~w10594 & w37804) | (w10048 & w37804);
assign w10596 = ~w10582 & w10595;
assign w10597 = w10048 & w37805;
assign w10598 = (w10099 & w10596) | (w10099 & w37806) | (w10596 & w37806);
assign w10599 = w10579 & ~w10598;
assign w10600 = ~w10403 & w10599;
assign w10601 = ~w10584 & w37807;
assign w10602 = ~w10598 & ~w10601;
assign w10603 = ~w10600 & ~w10602;
assign w10604 = w10592 & ~w10603;
assign w10605 = pi1975 & w9956;
assign w10606 = w10048 & w37808;
assign w10607 = w10544 & w37809;
assign w10608 = (w10607 & w10402) | (w10607 & w37810) | (w10402 & w37810);
assign w10609 = (w10606 & w10584) | (w10606 & w37811) | (w10584 & w37811);
assign w10610 = ~w10608 & ~w10609;
assign w10611 = ~w10587 & w10610;
assign w10612 = w10604 & w10611;
assign w10613 = (w2211 & w37812) | (w2211 & w37813) | (w37812 & w37813);
assign w10614 = ~pi3426 & ~w10613;
assign w10615 = ~w10613 & w37814;
assign w10616 = (w4748 & w37815) | (w4748 & w37816) | (w37815 & w37816);
assign w10617 = pi0407 & w397;
assign w10618 = w10617 & ~w10616;
assign w10619 = ~w10612 & w37817;
assign w10620 = pi0152 & pi0829;
assign w10621 = ~w10585 & ~w10620;
assign w10622 = w10544 & w37818;
assign w10623 = (w10622 & w10402) | (w10622 & w37819) | (w10402 & w37819);
assign w10624 = ~w10621 & ~w10623;
assign w10625 = w10592 & ~w10624;
assign w10626 = ~pi1041 & w10561;
assign w10627 = w10558 & ~w10626;
assign w10628 = ~pi1481 & w10564;
assign w10629 = ~pi1517 & w10559;
assign w10630 = ~pi1499 & w10566;
assign w10631 = ~w10629 & ~w10630;
assign w10632 = (~pi1041 & ~w10631) | (~pi1041 & w37822) | (~w10631 & w37822);
assign w10633 = (pi1041 & ~w10566) | (pi1041 & w37823) | (~w10566 & w37823);
assign w10634 = pi1417 & w10561;
assign w10635 = pi1553 & w10564;
assign w10636 = pi1585 & w10559;
assign w10637 = ~w10635 & ~w10636;
assign w10638 = w10637 & w37824;
assign w10639 = ~w10632 & ~w10638;
assign w10640 = w10558 & w37825;
assign w10641 = (w5893 & w37826) | (w5893 & w37827) | (w37826 & w37827);
assign w10642 = w10615 & w10641;
assign w10643 = pi0427 & w397;
assign w10644 = ~w10625 & w37828;
assign w10645 = ~pi0427 & w10641;
assign w10646 = pi0427 & ~w10641;
assign w10647 = ~w10645 & ~w10646;
assign w10648 = w397 & ~w10647;
assign w10649 = (w10648 & w10625) | (w10648 & w37829) | (w10625 & w37829);
assign w10650 = ~w10644 & ~w10649;
assign w10651 = ~w10619 & w10650;
assign w10652 = ~w10612 & w37830;
assign w10653 = pi0407 & pi0427;
assign w10654 = ~w10625 & w37831;
assign w10655 = pi0407 & ~w10647;
assign w10656 = (w10655 & w10625) | (w10655 & w37832) | (w10625 & w37832);
assign w10657 = ~w10654 & ~w10656;
assign w10658 = w10652 & ~w10657;
assign w10659 = ~w10651 & ~w10658;
assign w10660 = (w10550 & w10403) | (w10550 & w37833) | (w10403 & w37833);
assign w10661 = w10097 & ~w10103;
assign w10662 = ~w10582 & ~w10661;
assign w10663 = ~w10096 & w10662;
assign w10664 = w10062 & ~w10661;
assign w10665 = ~w10613 & w37835;
assign w10666 = (w10665 & w10661) | (w10665 & w37836) | (w10661 & w37836);
assign w10667 = w10666 & w40139;
assign w10668 = (~pi1041 & ~w10559) | (~pi1041 & w37838) | (~w10559 & w37838);
assign w10669 = ~pi1498 & w10566;
assign w10670 = ~pi1406 & w10564;
assign w10671 = ~w10669 & ~w10670;
assign w10672 = w10668 & w10671;
assign w10673 = (pi1041 & ~w10566) | (pi1041 & w37839) | (~w10566 & w37839);
assign w10674 = ~pi1535 & w10561;
assign w10675 = ~pi1409 & w10564;
assign w10676 = ~pi1584 & w10559;
assign w10677 = ~w10675 & ~w10676;
assign w10678 = w10677 & w37840;
assign w10679 = ~w10672 & ~w10678;
assign w10680 = w10558 & w37841;
assign w10681 = (~w10680 & w5319) | (~w10680 & w37842) | (w5319 & w37842);
assign w10682 = ~w10667 & w10681;
assign w10683 = pi0407 & ~pi0427;
assign w10684 = w385 & w10683;
assign w10685 = ~pi0407 & ~pi0427;
assign w10686 = ~pi0835 & w6668;
assign w10687 = ~w370 & w10558;
assign w10688 = w10558 & w37843;
assign w10689 = (~w10686 & ~w10558) | (~w10686 & w37844) | (~w10558 & w37844);
assign w10690 = ~w370 & w10615;
assign w10691 = ~pi1971 & w9957;
assign w10692 = w10615 & w37845;
assign w10693 = w10689 & ~w10692;
assign w10694 = (~pi1041 & ~w10564) | (~pi1041 & w37847) | (~w10564 & w37847);
assign w10695 = ~pi1626 & w10566;
assign w10696 = ~pi1515 & w10559;
assign w10697 = ~w10695 & ~w10696;
assign w10698 = w10694 & w10697;
assign w10699 = (pi1041 & ~w10564) | (pi1041 & w37848) | (~w10564 & w37848);
assign w10700 = ~pi1583 & w10559;
assign w10701 = ~pi1394 & w10566;
assign w10702 = ~pi1534 & w10561;
assign w10703 = ~w10701 & ~w10702;
assign w10704 = w10703 & w37849;
assign w10705 = ~w10698 & ~w10704;
assign w10706 = w10558 & w37850;
assign w10707 = (~w10706 & w4379) | (~w10706 & w37851) | (w4379 & w37851);
assign w10708 = w10689 & w37852;
assign w10709 = ~w9954 & w10692;
assign w10710 = ~w10708 & ~w10709;
assign w10711 = (w10710 & w10707) | (w10710 & w37853) | (w10707 & w37853);
assign w10712 = ~pi0407 & ~pi0415;
assign w10713 = w10712 & ~w10711;
assign w10714 = ~w10685 & ~w10713;
assign w10715 = ~pi0415 & ~pi0427;
assign w10716 = w10715 & ~w10711;
assign w10717 = pi0414 & ~w10716;
assign w10718 = ~w10714 & w10717;
assign w10719 = w10689 & ~w10690;
assign w10720 = w385 & w10653;
assign w10721 = pi0196 & ~w10720;
assign w10722 = ~pi0196 & ~w10684;
assign w10723 = ~w10721 & ~w10722;
assign w10724 = pi0134 & pi0407;
assign w10725 = ~pi0152 & pi0427;
assign w10726 = pi0152 & ~pi0427;
assign w10727 = ~w10725 & ~w10726;
assign w10728 = w10724 & w10727;
assign w10729 = (w397 & w10727) | (w397 & w37854) | (w10727 & w37854);
assign w10730 = ~w10728 & w10729;
assign w10731 = ~w10723 & ~w10730;
assign w10732 = w10689 & w37855;
assign w10733 = ~w343 & ~w10732;
assign w10734 = ~w10718 & w37856;
assign w10735 = w10682 & w10734;
assign w10736 = ~w10718 & w37857;
assign w10737 = ~w10682 & w10736;
assign w10738 = ~w10735 & ~w10737;
assign w10739 = ~w10659 & ~w10738;
assign w10740 = ~w10718 & w37858;
assign w10741 = ~pi3377 & pi3642;
assign w10742 = (w10741 & ~w342) | (w10741 & w37860) | (~w342 & w37860);
assign w10743 = ~w10740 & w10742;
assign w10744 = ~w10739 & w10743;
assign w10745 = ~w8265 & w37862;
assign w10746 = (~w10745 & w8239) | (~w10745 & w37863) | (w8239 & w37863);
assign w10747 = ~pi2757 & ~pi3633;
assign w10748 = ~pi0714 & ~w10747;
assign w10749 = w10748 & w40209;
assign w10750 = (pi0979 & ~w341) | (pi0979 & w37866) | (~w341 & w37866);
assign w10751 = ~w10613 & w37867;
assign w10752 = w10750 & w10751;
assign w10753 = w10747 & w40209;
assign w10754 = pi0051 & w40140;
assign w10755 = (~w10754 & ~w10751) | (~w10754 & w37868) | (~w10751 & w37868);
assign w10756 = (w10755 & w10746) | (w10755 & w37869) | (w10746 & w37869);
assign w10757 = ~pi0713 & w40209;
assign w10758 = (pi3245 & w7569) | (pi3245 & w37870) | (w7569 & w37870);
assign w10759 = ~w10749 & ~w10753;
assign w10760 = (~pi0039 & ~w40209) | (~pi0039 & w37874) | (~w40209 & w37874);
assign w10761 = w10759 & ~w10760;
assign w10762 = (w10761 & w40176) | (w10761 & w37875) | (w40176 & w37875);
assign w10763 = w10756 & ~w10762;
assign w10764 = ~pi0095 & ~pi0096;
assign w10765 = pi0095 & pi0096;
assign w10766 = ~w10764 & ~w10765;
assign w10767 = ~pi0098 & pi1425;
assign w10768 = pi0098 & ~pi1425;
assign w10769 = ~w10767 & ~w10768;
assign w10770 = ~pi0114 & ~w10769;
assign w10771 = pi0114 & w10769;
assign w10772 = ~w10770 & ~w10771;
assign w10773 = w10766 & ~w10772;
assign w10774 = pi1472 & pi2384;
assign w10775 = ~pi0868 & w10774;
assign w10776 = ~w6056 & w10775;
assign w10777 = pi0868 & w10774;
assign w10778 = ~w3060 & w10777;
assign w10779 = ~w10776 & ~w10778;
assign w10780 = ~pi0096 & pi1469;
assign w10781 = pi0096 & ~pi1469;
assign w10782 = ~w10780 & ~w10781;
assign w10783 = ~pi0074 & ~pi0075;
assign w10784 = pi0096 & ~w10783;
assign w10785 = pi0074 & pi0075;
assign w10786 = ~pi0096 & ~w10785;
assign w10787 = ~w10784 & ~w10786;
assign w10788 = ~w10782 & w10787;
assign w10789 = pi0108 & pi1473;
assign w10790 = ~pi0108 & ~pi1473;
assign w10791 = ~w10789 & ~w10790;
assign w10792 = pi0066 & ~pi0104;
assign w10793 = w10791 & w10792;
assign w10794 = pi0066 & pi0104;
assign w10795 = pi0078 & pi1473;
assign w10796 = ~pi0078 & ~pi1473;
assign w10797 = ~w10795 & ~w10796;
assign w10798 = w10794 & w10797;
assign w10799 = ~pi0066 & ~pi0104;
assign w10800 = ~w10791 & w10799;
assign w10801 = ~w10798 & ~w10800;
assign w10802 = ~w10793 & w10801;
assign w10803 = ~w10788 & w10802;
assign w10804 = w10788 & ~w10802;
assign w10805 = ~w10803 & ~w10804;
assign w10806 = ~w10779 & w10805;
assign w10807 = w10779 & ~w10805;
assign w10808 = ~w10806 & ~w10807;
assign w10809 = ~w10783 & ~w10785;
assign w10810 = ~w10782 & w10809;
assign w10811 = ~w3354 & w10777;
assign w10812 = ~w3060 & w10775;
assign w10813 = ~w10811 & ~w10812;
assign w10814 = ~w10810 & w10813;
assign w10815 = w10810 & ~w10813;
assign w10816 = ~w10814 & ~w10815;
assign w10817 = w10792 & w10797;
assign w10818 = pi0079 & pi1473;
assign w10819 = ~pi0079 & ~pi1473;
assign w10820 = ~w10818 & ~w10819;
assign w10821 = w10794 & w10820;
assign w10822 = ~w10797 & w10799;
assign w10823 = ~w10821 & ~w10822;
assign w10824 = ~w10817 & w10823;
assign w10825 = w10816 & w10824;
assign w10826 = (~w10814 & ~w10816) | (~w10814 & w37876) | (~w10816 & w37876);
assign w10827 = ~w10808 & ~w10826;
assign w10828 = w10808 & w10826;
assign w10829 = ~w10827 & ~w10828;
assign w10830 = pi0076 & pi0097;
assign w10831 = ~pi0076 & ~pi0097;
assign w10832 = ~w10830 & ~w10831;
assign w10833 = ~pi0075 & pi1468;
assign w10834 = pi0075 & ~pi1468;
assign w10835 = ~w10833 & ~w10834;
assign w10836 = ~pi0106 & ~w10835;
assign w10837 = pi0106 & w10835;
assign w10838 = ~w10836 & ~w10837;
assign w10839 = w10832 & ~w10838;
assign w10840 = ~pi0075 & ~w10830;
assign w10841 = pi0075 & ~w10831;
assign w10842 = ~w10840 & ~w10841;
assign w10843 = ~pi0056 & ~w10835;
assign w10844 = pi0056 & w10835;
assign w10845 = ~w10843 & ~w10844;
assign w10846 = w10842 & ~w10845;
assign w10847 = ~w10839 & ~w10846;
assign w10848 = pi0055 & ~pi0066;
assign w10849 = ~pi0055 & pi0066;
assign w10850 = ~w10848 & ~w10849;
assign w10851 = pi0097 & pi1424;
assign w10852 = ~pi0097 & ~pi1424;
assign w10853 = ~w10851 & ~w10852;
assign w10854 = ~pi0079 & w10853;
assign w10855 = pi0079 & ~w10853;
assign w10856 = ~w10854 & ~w10855;
assign w10857 = w10850 & ~w10856;
assign w10858 = ~pi0097 & w10848;
assign w10859 = pi0097 & w10849;
assign w10860 = ~w10858 & ~w10859;
assign w10861 = ~pi0080 & w10853;
assign w10862 = pi0080 & ~w10853;
assign w10863 = ~w10861 & ~w10862;
assign w10864 = ~w10860 & ~w10863;
assign w10865 = ~w10857 & ~w10864;
assign w10866 = ~pi0067 & ~w10782;
assign w10867 = pi0067 & w10782;
assign w10868 = ~w10866 & ~w10867;
assign w10869 = w10809 & ~w10868;
assign w10870 = ~pi0114 & ~w10782;
assign w10871 = pi0114 & w10782;
assign w10872 = ~w10870 & ~w10871;
assign w10873 = w10787 & ~w10872;
assign w10874 = ~w10869 & ~w10873;
assign w10875 = ~w10865 & w10874;
assign w10876 = w10865 & ~w10874;
assign w10877 = ~w10875 & ~w10876;
assign w10878 = ~w10847 & ~w10877;
assign w10879 = w10847 & w10877;
assign w10880 = ~w10878 & ~w10879;
assign w10881 = w10850 & ~w10863;
assign w10882 = ~pi0106 & w10853;
assign w10883 = pi0106 & ~w10853;
assign w10884 = ~w10882 & ~w10883;
assign w10885 = ~w10860 & ~w10884;
assign w10886 = ~w10881 & ~w10885;
assign w10887 = w10809 & ~w10872;
assign w10888 = w10886 & ~w10887;
assign w10889 = ~w10886 & w10887;
assign w10890 = w10832 & ~w10845;
assign w10891 = ~pi0067 & ~w10835;
assign w10892 = pi0067 & w10835;
assign w10893 = ~w10891 & ~w10892;
assign w10894 = w10842 & ~w10893;
assign w10895 = ~w10890 & ~w10894;
assign w10896 = ~w10889 & w10895;
assign w10897 = ~w10888 & ~w10896;
assign w10898 = ~w10880 & ~w10897;
assign w10899 = w10880 & w10897;
assign w10900 = ~w10898 & ~w10899;
assign w10901 = ~w10829 & ~w10900;
assign w10902 = ~w10816 & ~w10824;
assign w10903 = ~w10825 & ~w10902;
assign w10904 = ~w10835 & w10842;
assign w10905 = ~w6320 & w10777;
assign w10906 = ~w3354 & w10775;
assign w10907 = ~w10905 & ~w10906;
assign w10908 = w10904 & ~w10907;
assign w10909 = ~w10904 & w10907;
assign w10910 = ~w10908 & ~w10909;
assign w10911 = w10792 & w10820;
assign w10912 = pi0080 & pi1473;
assign w10913 = ~pi0080 & ~pi1473;
assign w10914 = ~w10912 & ~w10913;
assign w10915 = w10794 & w10914;
assign w10916 = w10799 & ~w10820;
assign w10917 = ~w10915 & ~w10916;
assign w10918 = ~w10911 & w10917;
assign w10919 = w10910 & ~w10918;
assign w10920 = (~w10908 & ~w10910) | (~w10908 & w37877) | (~w10910 & w37877);
assign w10921 = w10903 & w10920;
assign w10922 = ~pi0056 & w10853;
assign w10923 = pi0056 & ~w10853;
assign w10924 = ~w10922 & ~w10923;
assign w10925 = ~w10860 & ~w10924;
assign w10926 = w10850 & ~w10884;
assign w10927 = ~w10925 & ~w10926;
assign w10928 = w10832 & ~w10893;
assign w10929 = ~pi0114 & ~w10835;
assign w10930 = pi0114 & w10835;
assign w10931 = ~w10929 & ~w10930;
assign w10932 = w10842 & ~w10931;
assign w10933 = ~w10928 & ~w10932;
assign w10934 = ~w10927 & ~w10933;
assign w10935 = ~w10888 & ~w10889;
assign w10936 = w10895 & w10935;
assign w10937 = ~w10895 & ~w10935;
assign w10938 = ~w10936 & ~w10937;
assign w10939 = ~w10934 & w10938;
assign w10940 = (~w10921 & ~w10938) | (~w10921 & w37878) | (~w10938 & w37878);
assign w10941 = (~w10940 & w10900) | (~w10940 & w37879) | (w10900 & w37879);
assign w10942 = w10829 & w10900;
assign w10943 = w10827 & w10898;
assign w10944 = ~w10942 & ~w10943;
assign w10945 = ~w10941 & w10944;
assign w10946 = w10944 & w37880;
assign w10947 = (~w10804 & ~w10805) | (~w10804 & w37881) | (~w10805 & w37881);
assign w10948 = ~w6056 & w10777;
assign w10949 = ~w4042 & w10775;
assign w10950 = ~w10948 & ~w10949;
assign w10951 = w10766 & ~w10769;
assign w10952 = pi0107 & pi1473;
assign w10953 = ~pi0107 & ~pi1473;
assign w10954 = ~w10952 & ~w10953;
assign w10955 = w10792 & w10954;
assign w10956 = w10791 & w10794;
assign w10957 = w10799 & ~w10954;
assign w10958 = ~w10956 & ~w10957;
assign w10959 = w10958 & w37882;
assign w10960 = (w10951 & ~w10958) | (w10951 & w37883) | (~w10958 & w37883);
assign w10961 = ~w10959 & ~w10960;
assign w10962 = ~w10950 & w10961;
assign w10963 = w10950 & ~w10961;
assign w10964 = ~w10962 & ~w10963;
assign w10965 = w10947 & ~w10964;
assign w10966 = ~w10947 & w10964;
assign w10967 = ~w10965 & ~w10966;
assign w10968 = ~w10827 & ~w10898;
assign w10969 = ~w10865 & ~w10874;
assign w10970 = (~w10969 & w10877) | (~w10969 & w37884) | (w10877 & w37884);
assign w10971 = ~w10856 & ~w10860;
assign w10972 = ~pi0078 & w10853;
assign w10973 = pi0078 & ~w10853;
assign w10974 = ~w10972 & ~w10973;
assign w10975 = w10850 & ~w10974;
assign w10976 = ~w10971 & ~w10975;
assign w10977 = ~w10838 & w10842;
assign w10978 = ~pi0080 & ~w10835;
assign w10979 = pi0080 & w10835;
assign w10980 = ~w10978 & ~w10979;
assign w10981 = w10832 & ~w10980;
assign w10982 = ~w10977 & ~w10981;
assign w10983 = w10787 & ~w10868;
assign w10984 = ~pi0056 & ~w10782;
assign w10985 = pi0056 & w10782;
assign w10986 = ~w10984 & ~w10985;
assign w10987 = w10809 & ~w10986;
assign w10988 = ~w10983 & ~w10987;
assign w10989 = ~w10982 & w10988;
assign w10990 = w10982 & ~w10988;
assign w10991 = ~w10989 & ~w10990;
assign w10992 = ~w10976 & ~w10991;
assign w10993 = w10976 & w10991;
assign w10994 = ~w10992 & ~w10993;
assign w10995 = w10970 & ~w10994;
assign w10996 = ~w10970 & w10994;
assign w10997 = ~w10995 & ~w10996;
assign w10998 = w10968 & ~w10997;
assign w10999 = ~w10968 & w10997;
assign w11000 = ~w10998 & ~w10999;
assign w11001 = w10967 & ~w11000;
assign w11002 = ~w10967 & w11000;
assign w11003 = ~w11001 & ~w11002;
assign w11004 = ~w10946 & ~w11003;
assign w11005 = (w10773 & w11003) | (w10773 & w37885) | (w11003 & w37885);
assign w11006 = w10967 & ~w10998;
assign w11007 = ~w10994 & w37886;
assign w11008 = ~w10999 & ~w11007;
assign w11009 = ~w11006 & w11008;
assign w11010 = ~w10982 & ~w10988;
assign w11011 = (~w11010 & w10991) | (~w11010 & w37887) | (w10991 & w37887);
assign w11012 = w10842 & ~w10980;
assign w11013 = ~pi0079 & ~w10835;
assign w11014 = pi0079 & w10835;
assign w11015 = ~w11013 & ~w11014;
assign w11016 = w10832 & ~w11015;
assign w11017 = ~w11012 & ~w11016;
assign w11018 = ~w10860 & ~w10974;
assign w11019 = ~pi0108 & w10853;
assign w11020 = pi0108 & ~w10853;
assign w11021 = ~w11019 & ~w11020;
assign w11022 = w10850 & ~w11021;
assign w11023 = ~w11018 & ~w11022;
assign w11024 = w10787 & ~w10986;
assign w11025 = ~pi0106 & ~w10782;
assign w11026 = pi0106 & w10782;
assign w11027 = ~w11025 & ~w11026;
assign w11028 = w10809 & ~w11027;
assign w11029 = ~w11024 & ~w11028;
assign w11030 = ~w11023 & w11029;
assign w11031 = w11023 & ~w11029;
assign w11032 = ~w11030 & ~w11031;
assign w11033 = ~w11017 & ~w11032;
assign w11034 = w11017 & w11032;
assign w11035 = ~w11033 & ~w11034;
assign w11036 = w11011 & ~w11035;
assign w11037 = ~w11011 & w11035;
assign w11038 = ~w11036 & ~w11037;
assign w11039 = ~w4973 & w10775;
assign w11040 = ~w4042 & w10777;
assign w11041 = ~w11039 & ~w11040;
assign w11042 = pi0098 & w10764;
assign w11043 = ~pi0098 & w10765;
assign w11044 = ~w11042 & ~w11043;
assign w11045 = ~w10769 & ~w11044;
assign w11046 = pi0105 & pi1473;
assign w11047 = ~pi0105 & ~pi1473;
assign w11048 = ~w11046 & ~w11047;
assign w11049 = w10792 & w11048;
assign w11050 = w10799 & ~w11048;
assign w11051 = w10794 & w10954;
assign w11052 = ~w11050 & ~w11051;
assign w11053 = ~w11049 & w11052;
assign w11054 = ~w11045 & w11053;
assign w11055 = w11045 & ~w11053;
assign w11056 = ~w11054 & ~w11055;
assign w11057 = w11041 & w11056;
assign w11058 = ~w11041 & ~w11056;
assign w11059 = ~w11057 & ~w11058;
assign w11060 = (~w10960 & ~w10961) | (~w10960 & w37888) | (~w10961 & w37888);
assign w11061 = w11059 & w11060;
assign w11062 = ~w11059 & ~w11060;
assign w11063 = ~w11061 & ~w11062;
assign w11064 = ~w11038 & ~w11063;
assign w11065 = w11038 & w11063;
assign w11066 = ~w11064 & ~w11065;
assign w11067 = ~w10772 & ~w11044;
assign w11068 = ~pi0067 & ~w10769;
assign w11069 = pi0067 & w10769;
assign w11070 = ~w11068 & ~w11069;
assign w11071 = w10766 & ~w11070;
assign w11072 = ~w11067 & ~w11071;
assign w11073 = (~w10965 & w10994) | (~w10965 & w37889) | (w10994 & w37889);
assign w11074 = ~w11072 & w11073;
assign w11075 = w11072 & ~w11073;
assign w11076 = ~w11074 & ~w11075;
assign w11077 = w11066 & ~w11076;
assign w11078 = ~w11066 & w11076;
assign w11079 = ~w11077 & ~w11078;
assign w11080 = ~w11009 & w11079;
assign w11081 = w11009 & ~w11079;
assign w11082 = ~w11080 & ~w11081;
assign w11083 = ~w11005 & w11082;
assign w11084 = ~w10910 & w10918;
assign w11085 = ~w10919 & ~w11084;
assign w11086 = w10832 & ~w10835;
assign w11087 = ~w6320 & w10775;
assign w11088 = ~w4357 & w10777;
assign w11089 = ~w11087 & ~w11088;
assign w11090 = w11086 & ~w11089;
assign w11091 = ~w11086 & w11089;
assign w11092 = ~w11090 & ~w11091;
assign w11093 = w10792 & w10914;
assign w11094 = pi0106 & pi1473;
assign w11095 = ~pi0106 & ~pi1473;
assign w11096 = ~w11094 & ~w11095;
assign w11097 = w10794 & w11096;
assign w11098 = w10799 & ~w10914;
assign w11099 = ~w11097 & ~w11098;
assign w11100 = ~w11093 & w11099;
assign w11101 = w11092 & ~w11100;
assign w11102 = (~w11090 & ~w11092) | (~w11090 & w37890) | (~w11092 & w37890);
assign w11103 = ~w11085 & w11102;
assign w11104 = w10850 & ~w10924;
assign w11105 = ~pi0067 & w10853;
assign w11106 = pi0067 & ~w10853;
assign w11107 = ~w11105 & ~w11106;
assign w11108 = ~w10860 & ~w11107;
assign w11109 = ~w11104 & ~w11108;
assign w11110 = w10832 & ~w10931;
assign w11111 = ~w11109 & w11110;
assign w11112 = w10927 & w10933;
assign w11113 = ~w10934 & ~w11112;
assign w11114 = ~w11111 & ~w11113;
assign w11115 = ~w11103 & ~w11114;
assign w11116 = w10934 & ~w10938;
assign w11117 = ~w10903 & ~w10920;
assign w11118 = (~w11117 & w10938) | (~w11117 & w37891) | (w10938 & w37891);
assign w11119 = w10940 & ~w11118;
assign w11120 = w10938 & w37892;
assign w11121 = ~w11119 & ~w11120;
assign w11122 = (w11115 & w11119) | (w11115 & w37893) | (w11119 & w37893);
assign w11123 = ~w10901 & ~w10942;
assign w11124 = ~w10940 & ~w11116;
assign w11125 = ~w11115 & ~w11117;
assign w11126 = w11124 & w11125;
assign w11127 = w11123 & w37894;
assign w11128 = w11115 & w11121;
assign w11129 = ~w11124 & w11125;
assign w11130 = ~w11123 & ~w11129;
assign w11131 = ~w11128 & w11130;
assign w11132 = ~w11127 & ~w11131;
assign w11133 = ~w11115 & w11117;
assign w11134 = ~w11116 & w11133;
assign w11135 = ~w11123 & ~w11134;
assign w11136 = ~w11123 & w37895;
assign w11137 = ~w10940 & w11123;
assign w11138 = ~w11136 & ~w11137;
assign w11139 = ~w11132 & ~w11138;
assign w11140 = w11085 & ~w11102;
assign w11141 = ~w11103 & ~w11140;
assign w11142 = w11111 & w11113;
assign w11143 = ~w11114 & ~w11142;
assign w11144 = ~w11141 & ~w11143;
assign w11145 = w11109 & ~w11110;
assign w11146 = ~w11111 & ~w11145;
assign w11147 = w10853 & ~w10860;
assign w11148 = ~w5129 & w10777;
assign w11149 = ~w4357 & w10775;
assign w11150 = ~w11148 & ~w11149;
assign w11151 = w11147 & ~w11150;
assign w11152 = ~w11147 & w11150;
assign w11153 = ~w11151 & ~w11152;
assign w11154 = w10792 & w11096;
assign w11155 = pi0056 & pi1473;
assign w11156 = ~pi0056 & ~pi1473;
assign w11157 = w10794 & ~w11156;
assign w11158 = ~w11155 & w11157;
assign w11159 = w10799 & ~w11096;
assign w11160 = ~w11158 & ~w11159;
assign w11161 = ~w11154 & w11160;
assign w11162 = w11153 & ~w11161;
assign w11163 = (~w11151 & ~w11153) | (~w11151 & w37896) | (~w11153 & w37896);
assign w11164 = ~w11092 & w11100;
assign w11165 = ~w11101 & ~w11164;
assign w11166 = w11163 & ~w11165;
assign w11167 = w11146 & ~w11166;
assign w11168 = ~w11144 & ~w11167;
assign w11169 = w11141 & w11143;
assign w11170 = w11103 & w11114;
assign w11171 = ~w11169 & ~w11170;
assign w11172 = ~w11168 & w11171;
assign w11173 = ~w10939 & ~w11116;
assign w11174 = ~w10921 & ~w11117;
assign w11175 = ~w11115 & w11174;
assign w11176 = w11115 & ~w11174;
assign w11177 = ~w11175 & ~w11176;
assign w11178 = w11173 & ~w11177;
assign w11179 = ~w11173 & w11177;
assign w11180 = ~w11178 & ~w11179;
assign w11181 = ~w11172 & ~w11180;
assign w11182 = w10850 & ~w11107;
assign w11183 = ~pi0114 & w10853;
assign w11184 = pi0114 & ~w10853;
assign w11185 = ~w11183 & ~w11184;
assign w11186 = ~w10860 & ~w11185;
assign w11187 = ~w11182 & ~w11186;
assign w11188 = ~w11153 & w11161;
assign w11189 = ~w11162 & ~w11188;
assign w11190 = ~w5703 & w10777;
assign w11191 = ~w5129 & w10775;
assign w11192 = ~w11190 & ~w11191;
assign w11193 = w10850 & w10853;
assign w11194 = w11192 & ~w11193;
assign w11195 = ~w11192 & w11193;
assign w11196 = pi0067 & pi1473;
assign w11197 = ~pi0067 & ~pi1473;
assign w11198 = w10794 & ~w11197;
assign w11199 = ~w11196 & w11198;
assign w11200 = ~pi0066 & pi1473;
assign w11201 = pi0066 & ~pi1473;
assign w11202 = ~w11200 & ~w11201;
assign w11203 = ~pi0056 & ~w11202;
assign w11204 = (~pi0104 & ~w11202) | (~pi0104 & w37897) | (~w11202 & w37897);
assign w11205 = ~w11203 & w11204;
assign w11206 = ~w11199 & ~w11205;
assign w11207 = ~w11195 & w11206;
assign w11208 = ~w11194 & ~w11207;
assign w11209 = w11189 & w11208;
assign w11210 = w11189 & w37898;
assign w11211 = ~w11189 & ~w11208;
assign w11212 = ~w11209 & ~w11211;
assign w11213 = w11187 & ~w11212;
assign w11214 = ~w11187 & w11212;
assign w11215 = ~w11213 & ~w11214;
assign w11216 = ~pi0104 & pi0114;
assign w11217 = (w11216 & w4685) | (w11216 & w37899) | (w4685 & w37899);
assign w11218 = ~pi0868 & w11217;
assign w11219 = ~w3631 & w10774;
assign w11220 = pi0868 & w11216;
assign w11221 = ~w11219 & w11220;
assign w11222 = (~pi0104 & w11202) | (~pi0104 & w11216) | (w11202 & w11216);
assign w11223 = ~w11221 & w11222;
assign w11224 = ~w11218 & w11223;
assign w11225 = pi0114 & w10794;
assign w11226 = pi0067 & w11202;
assign w11227 = (~pi0104 & w11202) | (~pi0104 & w37900) | (w11202 & w37900);
assign w11228 = ~w11226 & w11227;
assign w11229 = ~w11225 & ~w11228;
assign w11230 = ~w5703 & w10775;
assign w11231 = ~w4685 & w10777;
assign w11232 = ~w11230 & ~w11231;
assign w11233 = ~w11229 & w11232;
assign w11234 = w11229 & ~w11232;
assign w11235 = ~w11233 & ~w11234;
assign w11236 = w11224 & ~w11235;
assign w11237 = ~pi0114 & pi1473;
assign w11238 = w10794 & w11237;
assign w11239 = (~w11238 & w11229) | (~w11238 & w37901) | (w11229 & w37901);
assign w11240 = ~w11236 & w11239;
assign w11241 = pi0114 & w10850;
assign w11242 = ~w11192 & w11241;
assign w11243 = w11192 & ~w11241;
assign w11244 = ~w11242 & ~w11243;
assign w11245 = ~w11206 & w11244;
assign w11246 = w11206 & ~w11244;
assign w11247 = ~w11245 & ~w11246;
assign w11248 = w11240 & w11247;
assign w11249 = w10850 & ~w11185;
assign w11250 = ~w11247 & ~w11249;
assign w11251 = ~w11248 & ~w11250;
assign w11252 = w11215 & w11251;
assign w11253 = (~w11210 & ~w11215) | (~w11210 & w37902) | (~w11215 & w37902);
assign w11254 = w11146 & ~w11163;
assign w11255 = ~w11146 & w11163;
assign w11256 = ~w11254 & ~w11255;
assign w11257 = (~w11187 & w11189) | (~w11187 & w37903) | (w11189 & w37903);
assign w11258 = ~w11165 & ~w11257;
assign w11259 = w11165 & ~w11187;
assign w11260 = ~w11211 & w11259;
assign w11261 = ~w11258 & ~w11260;
assign w11262 = w11256 & ~w11261;
assign w11263 = ~w11256 & w11261;
assign w11264 = ~w11262 & ~w11263;
assign w11265 = ~w11253 & ~w11264;
assign w11266 = ~w11144 & ~w11169;
assign w11267 = ~w11254 & w11258;
assign w11268 = w11254 & w11260;
assign w11269 = w11255 & ~w11260;
assign w11270 = ~w11268 & ~w11269;
assign w11271 = ~w11267 & w11270;
assign w11272 = w11266 & ~w11271;
assign w11273 = ~w11266 & w11271;
assign w11274 = ~w11272 & ~w11273;
assign w11275 = w11265 & ~w11274;
assign w11276 = ~w11266 & w11268;
assign w11277 = ~w11167 & w11266;
assign w11278 = w11271 & w11277;
assign w11279 = ~w11276 & ~w11278;
assign w11280 = w11172 & w11180;
assign w11281 = w11279 & ~w11280;
assign w11282 = ~w11275 & w11281;
assign w11283 = ~w11181 & ~w11282;
assign w11284 = ~w10938 & w37904;
assign w11285 = w11123 & ~w11284;
assign w11286 = ~w11135 & ~w11285;
assign w11287 = ~w11132 & ~w11286;
assign w11288 = w11283 & ~w11287;
assign w11289 = ~w11139 & ~w11288;
assign w11290 = w10946 & w11003;
assign w11291 = ~w11082 & w11290;
assign w11292 = (~w11083 & w11289) | (~w11083 & w37905) | (w11289 & w37905);
assign w11293 = ~w10773 & ~w10945;
assign w11294 = ~w11004 & ~w11293;
assign w11295 = ~w11003 & w11293;
assign w11296 = (~w11295 & w11288) | (~w11295 & w37906) | (w11288 & w37906);
assign w11297 = ~w11294 & ~w11296;
assign w11298 = ~w11292 & ~w11297;
assign w11299 = (~w11073 & w11038) | (~w11073 & w37907) | (w11038 & w37907);
assign w11300 = w11036 & w11061;
assign w11301 = ~w11065 & ~w11300;
assign w11302 = ~w11299 & w11301;
assign w11303 = ~pi0098 & ~pi0103;
assign w11304 = pi0098 & pi0103;
assign w11305 = ~w11303 & ~w11304;
assign w11306 = ~pi0102 & pi1470;
assign w11307 = pi0102 & ~pi1470;
assign w11308 = ~w11306 & ~w11307;
assign w11309 = ~pi0114 & w11308;
assign w11310 = pi0114 & ~w11308;
assign w11311 = ~w11309 & ~w11310;
assign w11312 = w11305 & w11311;
assign w11313 = ~w11044 & ~w11070;
assign w11314 = ~pi0056 & ~w10769;
assign w11315 = pi0056 & w10769;
assign w11316 = ~w11314 & ~w11315;
assign w11317 = w10766 & ~w11316;
assign w11318 = ~w11313 & ~w11317;
assign w11319 = w11312 & ~w11318;
assign w11320 = ~w11312 & w11318;
assign w11321 = ~w11319 & ~w11320;
assign w11322 = ~w11036 & ~w11061;
assign w11323 = (~w11054 & ~w11056) | (~w11054 & w37908) | (~w11056 & w37908);
assign w11324 = ~w5605 & w10775;
assign w11325 = ~w4973 & w10777;
assign w11326 = ~w11324 & ~w11325;
assign w11327 = w11305 & ~w11308;
assign w11328 = pi0113 & ~pi1473;
assign w11329 = ~pi0113 & pi1473;
assign w11330 = ~w11328 & ~w11329;
assign w11331 = w10799 & w11330;
assign w11332 = w10792 & ~w11330;
assign w11333 = w10794 & w11048;
assign w11334 = ~w11332 & ~w11333;
assign w11335 = (w11327 & ~w11334) | (w11327 & w37909) | (~w11334 & w37909);
assign w11336 = w11334 & w37910;
assign w11337 = ~w11335 & ~w11336;
assign w11338 = w11326 & ~w11337;
assign w11339 = ~w11326 & w11337;
assign w11340 = ~w11338 & ~w11339;
assign w11341 = ~w11323 & ~w11340;
assign w11342 = w11323 & w11340;
assign w11343 = ~w11341 & ~w11342;
assign w11344 = ~w11023 & ~w11029;
assign w11345 = (~w11344 & w11032) | (~w11344 & w37911) | (w11032 & w37911);
assign w11346 = w10842 & ~w11015;
assign w11347 = ~pi0078 & ~w10835;
assign w11348 = pi0078 & w10835;
assign w11349 = ~w11347 & ~w11348;
assign w11350 = w10832 & ~w11349;
assign w11351 = ~w11346 & ~w11350;
assign w11352 = w10787 & ~w11027;
assign w11353 = ~pi0080 & ~w10782;
assign w11354 = pi0080 & w10782;
assign w11355 = ~w11353 & ~w11354;
assign w11356 = w10809 & ~w11355;
assign w11357 = ~w11352 & ~w11356;
assign w11358 = ~w10860 & ~w11021;
assign w11359 = ~pi0107 & w10853;
assign w11360 = pi0107 & ~w10853;
assign w11361 = ~w11359 & ~w11360;
assign w11362 = w10850 & ~w11361;
assign w11363 = ~w11358 & ~w11362;
assign w11364 = w11357 & w11363;
assign w11365 = ~w11357 & ~w11363;
assign w11366 = ~w11364 & ~w11365;
assign w11367 = w11351 & ~w11366;
assign w11368 = ~w11351 & w11366;
assign w11369 = ~w11367 & ~w11368;
assign w11370 = w11345 & ~w11369;
assign w11371 = ~w11345 & w11369;
assign w11372 = ~w11370 & ~w11371;
assign w11373 = w11343 & w11372;
assign w11374 = ~w11343 & ~w11372;
assign w11375 = ~w11373 & ~w11374;
assign w11376 = ~w11322 & w11375;
assign w11377 = w11322 & ~w11375;
assign w11378 = ~w11376 & ~w11377;
assign w11379 = w11321 & ~w11378;
assign w11380 = ~w11321 & w11378;
assign w11381 = ~w11379 & ~w11380;
assign w11382 = w11302 & w11381;
assign w11383 = ~w11302 & ~w11381;
assign w11384 = ~w11382 & ~w11383;
assign w11385 = w11005 & ~w11079;
assign w11386 = ~w11066 & w11073;
assign w11387 = w11066 & ~w11073;
assign w11388 = ~w11386 & ~w11387;
assign w11389 = ~w11072 & ~w11388;
assign w11390 = (~w11009 & w11388) | (~w11009 & w37912) | (w11388 & w37912);
assign w11391 = ~w11385 & w11390;
assign w11392 = ~w11388 & w11495;
assign w11393 = w11005 & w11392;
assign w11394 = w11072 & w11388;
assign w11395 = ~w11005 & w11394;
assign w11396 = ~w11393 & ~w11395;
assign w11397 = ~w11391 & w11396;
assign w11398 = w11384 & ~w11397;
assign w11399 = ~w11384 & w11397;
assign w11400 = ~w11398 & ~w11399;
assign w11401 = w11298 & ~w11400;
assign w11402 = pi0102 & w11303;
assign w11403 = ~pi0102 & w11304;
assign w11404 = ~w11402 & ~w11403;
assign w11405 = w11311 & ~w11404;
assign w11406 = ~pi0067 & w11308;
assign w11407 = pi0067 & ~w11308;
assign w11408 = ~w11406 & ~w11407;
assign w11409 = w11305 & w11408;
assign w11410 = ~w11405 & ~w11409;
assign w11411 = ~w11044 & ~w11316;
assign w11412 = ~pi0106 & ~w10769;
assign w11413 = pi0106 & w10769;
assign w11414 = ~w11412 & ~w11413;
assign w11415 = w10766 & ~w11414;
assign w11416 = ~w11411 & ~w11415;
assign w11417 = ~w11410 & ~w11416;
assign w11418 = w11410 & w11416;
assign w11419 = ~w11417 & ~w11418;
assign w11420 = w11319 & w11419;
assign w11421 = ~w11319 & ~w11419;
assign w11422 = ~w11420 & ~w11421;
assign w11423 = ~w11369 & w37913;
assign w11424 = (~w11423 & ~w11372) | (~w11423 & w37914) | (~w11372 & w37914);
assign w11425 = (w11424 & ~w11375) | (w11424 & w37915) | (~w11375 & w37915);
assign w11426 = w10787 & ~w11355;
assign w11427 = ~pi0079 & ~w10782;
assign w11428 = pi0079 & w10782;
assign w11429 = ~w11427 & ~w11428;
assign w11430 = w10809 & ~w11429;
assign w11431 = ~w11426 & ~w11430;
assign w11432 = w10842 & ~w11349;
assign w11433 = ~pi0108 & ~w10835;
assign w11434 = pi0108 & w10835;
assign w11435 = ~w11433 & ~w11434;
assign w11436 = w10832 & ~w11435;
assign w11437 = ~w11432 & ~w11436;
assign w11438 = ~w10860 & ~w11361;
assign w11439 = ~pi0105 & w10853;
assign w11440 = pi0105 & ~w10853;
assign w11441 = ~w11439 & ~w11440;
assign w11442 = w10850 & ~w11441;
assign w11443 = ~w11438 & ~w11442;
assign w11444 = ~w11437 & w11443;
assign w11445 = w11437 & ~w11443;
assign w11446 = ~w11444 & ~w11445;
assign w11447 = ~w11431 & ~w11446;
assign w11448 = w11431 & w11446;
assign w11449 = ~w11447 & ~w11448;
assign w11450 = ~w11351 & ~w11364;
assign w11451 = ~w11365 & ~w11450;
assign w11452 = ~w11449 & w11451;
assign w11453 = w11449 & ~w11451;
assign w11454 = ~w11452 & ~w11453;
assign w11455 = (~w11341 & w11369) | (~w11341 & w37916) | (w11369 & w37916);
assign w11456 = pi0112 & pi1473;
assign w11457 = ~pi0112 & ~pi1473;
assign w11458 = ~w11456 & ~w11457;
assign w11459 = w10792 & w11458;
assign w11460 = w10799 & ~w11458;
assign w11461 = w10794 & ~w11330;
assign w11462 = ~w11460 & ~w11461;
assign w11463 = ~w11459 & w11462;
assign w11464 = (pi1470 & ~w11304) | (pi1470 & w12571) | (~w11304 & w12571);
assign w11465 = (~pi1470 & ~w11303) | (~pi1470 & w12569) | (~w11303 & w12569);
assign w11466 = ~w11464 & ~w11465;
assign w11467 = ~w5605 & w10777;
assign w11468 = ~w1147 & w10775;
assign w11469 = ~w11467 & ~w11468;
assign w11470 = w11466 & ~w11469;
assign w11471 = ~w11466 & w11469;
assign w11472 = ~w11470 & ~w11471;
assign w11473 = ~w11463 & w11472;
assign w11474 = w11463 & ~w11472;
assign w11475 = ~w11473 & ~w11474;
assign w11476 = w11326 & ~w11335;
assign w11477 = ~w11336 & ~w11476;
assign w11478 = ~w11475 & ~w11477;
assign w11479 = w11475 & w11477;
assign w11480 = ~w11478 & ~w11479;
assign w11481 = ~w11455 & w11480;
assign w11482 = w11455 & ~w11480;
assign w11483 = ~w11481 & ~w11482;
assign w11484 = w11454 & ~w11483;
assign w11485 = ~w11454 & w11483;
assign w11486 = ~w11484 & ~w11485;
assign w11487 = ~w11425 & ~w11486;
assign w11488 = w11425 & w11486;
assign w11489 = ~w11487 & ~w11488;
assign w11490 = w11422 & ~w11489;
assign w11491 = ~w11422 & w11489;
assign w11492 = ~w11490 & ~w11491;
assign w11493 = w11301 & w37917;
assign w11494 = ~w11492 & ~w11493;
assign w11495 = w11009 & ~w11072;
assign w11496 = ~w11389 & ~w11495;
assign w11497 = ~w11382 & w11496;
assign w11498 = ~w11383 & ~w11497;
assign w11499 = (~w11378 & w11389) | (~w11378 & w37918) | (w11389 & w37918);
assign w11500 = w11493 & w11499;
assign w11501 = w11492 & w11500;
assign w11502 = (~w11501 & ~w11498) | (~w11501 & w37919) | (~w11498 & w37919);
assign w11503 = ~w11384 & w11393;
assign w11504 = w11384 & w11496;
assign w11505 = w11397 & w11504;
assign w11506 = ~w11503 & ~w11505;
assign w11507 = w11502 & w11506;
assign w11508 = ~w11401 & w11507;
assign w11509 = ~w11378 & w37920;
assign w11510 = ~w11492 & w11509;
assign w11511 = ~w11489 & w37921;
assign w11512 = ~w11488 & ~w11493;
assign w11513 = ~w11422 & ~w11487;
assign w11514 = ~w11512 & w11513;
assign w11515 = ~w11511 & ~w11514;
assign w11516 = ~w11510 & w11515;
assign w11517 = w11319 & w11417;
assign w11518 = ~w11487 & w11517;
assign w11519 = (~w11417 & ~w11419) | (~w11417 & w37922) | (~w11419 & w37922);
assign w11520 = ~w11319 & w11418;
assign w11521 = (~w11520 & ~w11487) | (~w11520 & w37923) | (~w11487 & w37923);
assign w11522 = ~w11518 & w11521;
assign w11523 = w11454 & ~w11482;
assign w11524 = ~w11449 & w37924;
assign w11525 = ~w11481 & ~w11524;
assign w11526 = ~w11523 & w11525;
assign w11527 = ~w11437 & ~w11443;
assign w11528 = (~w11527 & w11446) | (~w11527 & w37925) | (w11446 & w37925);
assign w11529 = ~w10860 & ~w11441;
assign w11530 = ~pi0113 & w10853;
assign w11531 = pi0113 & ~w10853;
assign w11532 = ~w11530 & ~w11531;
assign w11533 = w10850 & ~w11532;
assign w11534 = ~w11529 & ~w11533;
assign w11535 = w10842 & ~w11435;
assign w11536 = ~pi0107 & ~w10835;
assign w11537 = pi0107 & w10835;
assign w11538 = ~w11536 & ~w11537;
assign w11539 = w10832 & ~w11538;
assign w11540 = ~w11535 & ~w11539;
assign w11541 = w10787 & ~w11429;
assign w11542 = ~pi0078 & ~w10782;
assign w11543 = pi0078 & w10782;
assign w11544 = ~w11542 & ~w11543;
assign w11545 = w10809 & ~w11544;
assign w11546 = ~w11541 & ~w11545;
assign w11547 = ~w11540 & w11546;
assign w11548 = w11540 & ~w11546;
assign w11549 = ~w11547 & ~w11548;
assign w11550 = ~w11534 & ~w11549;
assign w11551 = w11534 & w11549;
assign w11552 = ~w11550 & ~w11551;
assign w11553 = w11528 & ~w11552;
assign w11554 = ~w11528 & w11552;
assign w11555 = ~w11553 & ~w11554;
assign w11556 = pi0101 & pi0102;
assign w11557 = ~pi0101 & ~pi0102;
assign w11558 = ~w11556 & ~w11557;
assign w11559 = ~pi0100 & pi1418;
assign w11560 = pi0100 & ~pi1418;
assign w11561 = ~w11559 & ~w11560;
assign w11562 = w11558 & ~w11561;
assign w11563 = ~w1517 & w10775;
assign w11564 = ~w1147 & w10777;
assign w11565 = ~w11563 & ~w11564;
assign w11566 = ~w11562 & w11565;
assign w11567 = w11562 & ~w11565;
assign w11568 = ~w11566 & ~w11567;
assign w11569 = pi0111 & pi1473;
assign w11570 = ~pi0111 & ~pi1473;
assign w11571 = ~w11569 & ~w11570;
assign w11572 = w10792 & w11571;
assign w11573 = w10799 & ~w11571;
assign w11574 = w10794 & w11458;
assign w11575 = ~w11573 & ~w11574;
assign w11576 = ~w11572 & w11575;
assign w11577 = w11568 & w11576;
assign w11578 = ~w11568 & ~w11576;
assign w11579 = ~w11577 & ~w11578;
assign w11580 = w11463 & ~w11470;
assign w11581 = ~w11471 & ~w11580;
assign w11582 = w11579 & ~w11581;
assign w11583 = ~w11579 & w11581;
assign w11584 = ~w11582 & ~w11583;
assign w11585 = ~w11478 & ~w11584;
assign w11586 = ~w11452 & w11585;
assign w11587 = (~w11478 & w11449) | (~w11478 & w37926) | (w11449 & w37926);
assign w11588 = w11584 & ~w11587;
assign w11589 = ~w11586 & ~w11588;
assign w11590 = w11555 & ~w11589;
assign w11591 = ~w11555 & w11589;
assign w11592 = ~w11590 & ~w11591;
assign w11593 = ~w11526 & ~w11592;
assign w11594 = w11526 & w11592;
assign w11595 = ~w11593 & ~w11594;
assign w11596 = ~pi0114 & ~w11561;
assign w11597 = pi0114 & w11561;
assign w11598 = ~w11596 & ~w11597;
assign w11599 = w11558 & ~w11598;
assign w11600 = ~w11404 & w11408;
assign w11601 = ~pi0056 & w11308;
assign w11602 = pi0056 & ~w11308;
assign w11603 = ~w11601 & ~w11602;
assign w11604 = w11305 & w11603;
assign w11605 = ~w11600 & ~w11604;
assign w11606 = ~w11044 & ~w11414;
assign w11607 = ~pi0080 & ~w10769;
assign w11608 = pi0080 & w10769;
assign w11609 = ~w11607 & ~w11608;
assign w11610 = w10766 & ~w11609;
assign w11611 = ~w11606 & ~w11610;
assign w11612 = ~w11605 & w11611;
assign w11613 = w11605 & ~w11611;
assign w11614 = ~w11612 & ~w11613;
assign w11615 = ~w11599 & ~w11614;
assign w11616 = w11599 & w11614;
assign w11617 = ~w11615 & ~w11616;
assign w11618 = w11595 & ~w11617;
assign w11619 = ~w11595 & w11617;
assign w11620 = ~w11618 & ~w11619;
assign w11621 = ~w11522 & w11620;
assign w11622 = w11522 & ~w11620;
assign w11623 = ~w11621 & ~w11622;
assign w11624 = ~w11516 & ~w11623;
assign w11625 = w11516 & w11623;
assign w11626 = ~w11624 & ~w11625;
assign w11627 = (~w11321 & ~w11301) | (~w11321 & w37927) | (~w11301 & w37927);
assign w11628 = w11492 & ~w11627;
assign w11629 = (~w11499 & w11492) | (~w11499 & w37928) | (w11492 & w37928);
assign w11630 = ~w11628 & w11629;
assign w11631 = w11378 & w11492;
assign w11632 = w11497 & w11631;
assign w11633 = ~w11510 & ~w11632;
assign w11634 = ~w11630 & w11633;
assign w11635 = w11626 & w11634;
assign w11636 = ~w11508 & w11635;
assign w11637 = ~w11540 & ~w11546;
assign w11638 = (~w11637 & w11549) | (~w11637 & w37929) | (w11549 & w37929);
assign w11639 = ~w10860 & ~w11532;
assign w11640 = ~pi0112 & w10853;
assign w11641 = pi0112 & ~w10853;
assign w11642 = ~w11640 & ~w11641;
assign w11643 = w10850 & ~w11642;
assign w11644 = ~w11639 & ~w11643;
assign w11645 = ~pi0105 & ~w10835;
assign w11646 = pi0105 & w10835;
assign w11647 = ~w11645 & ~w11646;
assign w11648 = w10832 & ~w11647;
assign w11649 = w10842 & ~w11538;
assign w11650 = ~w11648 & ~w11649;
assign w11651 = ~pi0108 & ~w10782;
assign w11652 = pi0108 & w10782;
assign w11653 = ~w11651 & ~w11652;
assign w11654 = w10809 & ~w11653;
assign w11655 = w10787 & ~w11544;
assign w11656 = ~w11654 & ~w11655;
assign w11657 = ~w11650 & w11656;
assign w11658 = w11650 & ~w11656;
assign w11659 = ~w11657 & ~w11658;
assign w11660 = ~w11644 & ~w11659;
assign w11661 = w11644 & w11659;
assign w11662 = ~w11660 & ~w11661;
assign w11663 = w11638 & ~w11662;
assign w11664 = ~w11638 & w11662;
assign w11665 = ~w11663 & ~w11664;
assign w11666 = (~w11566 & ~w11568) | (~w11566 & w37930) | (~w11568 & w37930);
assign w11667 = ~w7927 & w10775;
assign w11668 = ~w1517 & w10777;
assign w11669 = ~w11667 & ~w11668;
assign w11670 = ~pi0100 & ~w11556;
assign w11671 = pi0100 & ~w11557;
assign w11672 = ~w11670 & ~w11671;
assign w11673 = ~w11561 & w11672;
assign w11674 = pi0110 & pi1473;
assign w11675 = ~pi0110 & ~pi1473;
assign w11676 = ~w11674 & ~w11675;
assign w11677 = w10792 & w11676;
assign w11678 = w10794 & w11571;
assign w11679 = w10799 & ~w11676;
assign w11680 = ~w11678 & ~w11679;
assign w11681 = ~w11677 & w11680;
assign w11682 = ~w11673 & w11681;
assign w11683 = w11673 & ~w11681;
assign w11684 = ~w11682 & ~w11683;
assign w11685 = ~w11669 & w11684;
assign w11686 = w11669 & ~w11684;
assign w11687 = ~w11685 & ~w11686;
assign w11688 = ~w11666 & ~w11687;
assign w11689 = w11666 & w11687;
assign w11690 = ~w11688 & ~w11689;
assign w11691 = ~w11665 & ~w11690;
assign w11692 = w11665 & w11690;
assign w11693 = ~w11691 & ~w11692;
assign w11694 = w11528 & w11584;
assign w11695 = ~w11582 & ~w11587;
assign w11696 = ~w11694 & ~w11695;
assign w11697 = ~w11528 & ~w11584;
assign w11698 = ~w11694 & ~w11697;
assign w11699 = ~w11555 & ~w11587;
assign w11700 = ~w11698 & w11699;
assign w11701 = ~w11696 & ~w11700;
assign w11702 = w11555 & ~w11586;
assign w11703 = (w11582 & w11552) | (w11582 & w37931) | (w11552 & w37931);
assign w11704 = ~w11702 & w11703;
assign w11705 = (w11693 & w11701) | (w11693 & w37932) | (w11701 & w37932);
assign w11706 = ~w11582 & ~w11693;
assign w11707 = w11582 & w11693;
assign w11708 = w11552 & w11587;
assign w11709 = ~w11695 & ~w11697;
assign w11710 = ~w11708 & w11709;
assign w11711 = ~w11707 & w11710;
assign w11712 = ~w11706 & w11711;
assign w11713 = ~w11705 & ~w11712;
assign w11714 = ~w11693 & ~w11704;
assign w11715 = ~w11701 & w11714;
assign w11716 = ~w11555 & w11698;
assign w11717 = ~w11589 & w11716;
assign w11718 = w11555 & w11698;
assign w11719 = w11589 & w11718;
assign w11720 = ~w11717 & ~w11719;
assign w11721 = w11715 & w11720;
assign w11722 = w11713 & ~w11721;
assign w11723 = w11417 & ~w11617;
assign w11724 = ~pi0067 & ~w11561;
assign w11725 = pi0067 & w11561;
assign w11726 = ~w11724 & ~w11725;
assign w11727 = w11558 & ~w11726;
assign w11728 = ~w11598 & w11672;
assign w11729 = ~w11727 & ~w11728;
assign w11730 = ~w11404 & w11603;
assign w11731 = ~pi0106 & w11308;
assign w11732 = pi0106 & ~w11308;
assign w11733 = ~w11731 & ~w11732;
assign w11734 = w11305 & w11733;
assign w11735 = ~w11730 & ~w11734;
assign w11736 = ~pi0079 & ~w10769;
assign w11737 = pi0079 & w10769;
assign w11738 = ~w11736 & ~w11737;
assign w11739 = w10766 & ~w11738;
assign w11740 = ~w11044 & ~w11609;
assign w11741 = ~w11739 & ~w11740;
assign w11742 = ~w11735 & w11741;
assign w11743 = w11735 & ~w11741;
assign w11744 = ~w11742 & ~w11743;
assign w11745 = ~w11729 & w11744;
assign w11746 = w11729 & ~w11744;
assign w11747 = ~w11745 & ~w11746;
assign w11748 = w11605 & w11611;
assign w11749 = (~w11748 & w11614) | (~w11748 & w37933) | (w11614 & w37933);
assign w11750 = ~w11747 & w11749;
assign w11751 = w11747 & ~w11749;
assign w11752 = ~w11750 & ~w11751;
assign w11753 = ~w11723 & ~w11752;
assign w11754 = w11723 & w11752;
assign w11755 = ~w11753 & ~w11754;
assign w11756 = (w11755 & ~w11713) | (w11755 & w37934) | (~w11713 & w37934);
assign w11757 = w11713 & w37935;
assign w11758 = ~w11756 & ~w11757;
assign w11759 = w11422 & ~w11487;
assign w11760 = ~w11593 & ~w11759;
assign w11761 = (~w11594 & w11758) | (~w11594 & w37936) | (w11758 & w37936);
assign w11762 = ~w11417 & w11617;
assign w11763 = ~w11723 & ~w11762;
assign w11764 = ~w11420 & ~w11763;
assign w11765 = (~w11764 & w11592) | (~w11764 & w37937) | (w11592 & w37937);
assign w11766 = ~w11758 & w11765;
assign w11767 = ~w11593 & w11757;
assign w11768 = (w11755 & w11592) | (w11755 & w37938) | (w11592 & w37938);
assign w11769 = (w11768 & ~w11713) | (w11768 & w37939) | (~w11713 & w37939);
assign w11770 = w11420 & ~w11617;
assign w11771 = ~w11487 & w37940;
assign w11772 = (~w11770 & w11487) | (~w11770 & w37941) | (w11487 & w37941);
assign w11773 = ~w11769 & w11772;
assign w11774 = ~w11767 & w11773;
assign w11775 = ~w11766 & ~w11774;
assign w11776 = ~w11761 & w11775;
assign w11777 = ~w11624 & ~w11776;
assign w11778 = ~w11650 & ~w11656;
assign w11779 = (~w11778 & w11659) | (~w11778 & w37942) | (w11659 & w37942);
assign w11780 = ~w10860 & ~w11642;
assign w11781 = ~pi0111 & w10853;
assign w11782 = pi0111 & ~w10853;
assign w11783 = ~w11781 & ~w11782;
assign w11784 = w10850 & ~w11783;
assign w11785 = ~w11780 & ~w11784;
assign w11786 = ~pi0113 & ~w10835;
assign w11787 = pi0113 & w10835;
assign w11788 = ~w11786 & ~w11787;
assign w11789 = w10832 & ~w11788;
assign w11790 = w10842 & ~w11647;
assign w11791 = ~w11789 & ~w11790;
assign w11792 = ~pi0107 & ~w10782;
assign w11793 = pi0107 & w10782;
assign w11794 = ~w11792 & ~w11793;
assign w11795 = w10809 & ~w11794;
assign w11796 = w10787 & ~w11653;
assign w11797 = ~w11795 & ~w11796;
assign w11798 = ~w11791 & w11797;
assign w11799 = w11791 & ~w11797;
assign w11800 = ~w11798 & ~w11799;
assign w11801 = ~w11785 & ~w11800;
assign w11802 = w11785 & w11800;
assign w11803 = ~w11801 & ~w11802;
assign w11804 = w11779 & ~w11803;
assign w11805 = ~w8172 & w10775;
assign w11806 = ~w7927 & w10777;
assign w11807 = ~w11805 & ~w11806;
assign w11808 = pi0099 & pi0100;
assign w11809 = ~pi0099 & ~pi0100;
assign w11810 = ~w11808 & ~w11809;
assign w11811 = ~pi0077 & pi1471;
assign w11812 = pi0077 & ~pi1471;
assign w11813 = ~w11811 & ~w11812;
assign w11814 = w11810 & ~w11813;
assign w11815 = pi0109 & pi1473;
assign w11816 = ~pi0109 & ~pi1473;
assign w11817 = ~w11815 & ~w11816;
assign w11818 = w10792 & w11817;
assign w11819 = w10794 & w11676;
assign w11820 = w10799 & ~w11817;
assign w11821 = ~w11819 & ~w11820;
assign w11822 = (w11814 & ~w11821) | (w11814 & w37943) | (~w11821 & w37943);
assign w11823 = w11821 & w37944;
assign w11824 = ~w11822 & ~w11823;
assign w11825 = ~w11807 & w11824;
assign w11826 = w11807 & ~w11824;
assign w11827 = ~w11825 & ~w11826;
assign w11828 = (~w11683 & ~w11684) | (~w11683 & w37945) | (~w11684 & w37945);
assign w11829 = ~w11827 & w11828;
assign w11830 = (~w11829 & w11803) | (~w11829 & w37946) | (w11803 & w37946);
assign w11831 = (~w11822 & ~w11824) | (~w11822 & w37947) | (~w11824 & w37947);
assign w11832 = ~w8172 & w10777;
assign w11833 = ~pi0077 & ~w11808;
assign w11834 = pi0077 & ~w11809;
assign w11835 = ~w11833 & ~w11834;
assign w11836 = ~w11813 & w11835;
assign w11837 = (~pi0104 & ~w11202) | (~pi0104 & w37948) | (~w11202 & w37948);
assign w11838 = ~pi0081 & ~w11202;
assign w11839 = w11837 & ~w11838;
assign w11840 = w10794 & w11817;
assign w11841 = ~w11839 & ~w11840;
assign w11842 = w11836 & ~w11841;
assign w11843 = ~w11836 & w11841;
assign w11844 = ~w11842 & ~w11843;
assign w11845 = w11832 & w11844;
assign w11846 = ~w11832 & ~w11844;
assign w11847 = ~w11845 & ~w11846;
assign w11848 = w11831 & ~w11847;
assign w11849 = ~w11831 & w11847;
assign w11850 = ~w11848 & ~w11849;
assign w11851 = ~w11791 & ~w11797;
assign w11852 = (~w11851 & w11800) | (~w11851 & w37949) | (w11800 & w37949);
assign w11853 = ~pi0112 & ~w10835;
assign w11854 = pi0112 & w10835;
assign w11855 = ~w11853 & ~w11854;
assign w11856 = w10832 & ~w11855;
assign w11857 = w10842 & ~w11788;
assign w11858 = ~w11856 & ~w11857;
assign w11859 = ~pi0105 & ~w10782;
assign w11860 = pi0105 & w10782;
assign w11861 = ~w11859 & ~w11860;
assign w11862 = w10809 & ~w11861;
assign w11863 = w10787 & ~w11794;
assign w11864 = ~w11862 & ~w11863;
assign w11865 = ~w10860 & ~w11783;
assign w11866 = ~pi0110 & w10853;
assign w11867 = pi0110 & ~w10853;
assign w11868 = ~w11866 & ~w11867;
assign w11869 = w10850 & ~w11868;
assign w11870 = ~w11865 & ~w11869;
assign w11871 = ~w11864 & w11870;
assign w11872 = w11864 & ~w11870;
assign w11873 = ~w11871 & ~w11872;
assign w11874 = ~w11858 & ~w11873;
assign w11875 = w11858 & w11873;
assign w11876 = ~w11874 & ~w11875;
assign w11877 = w11852 & ~w11876;
assign w11878 = ~w11852 & w11876;
assign w11879 = ~w11877 & ~w11878;
assign w11880 = w11850 & w11879;
assign w11881 = ~w11850 & ~w11879;
assign w11882 = ~w11880 & ~w11881;
assign w11883 = ~w11830 & w11882;
assign w11884 = w11830 & ~w11882;
assign w11885 = ~w11883 & ~w11884;
assign w11886 = ~w11663 & ~w11688;
assign w11887 = ~w11779 & w11803;
assign w11888 = ~w11804 & ~w11887;
assign w11889 = w11827 & ~w11828;
assign w11890 = ~w11829 & ~w11889;
assign w11891 = ~w11888 & ~w11890;
assign w11892 = ~w11886 & ~w11891;
assign w11893 = w11888 & w11890;
assign w11894 = ~w11803 & w37950;
assign w11895 = (~w11894 & ~w11888) | (~w11894 & w37951) | (~w11888 & w37951);
assign w11896 = ~w11892 & w11895;
assign w11897 = w11885 & ~w11896;
assign w11898 = ~w11885 & w11896;
assign w11899 = ~w11897 & ~w11898;
assign w11900 = ~pi0078 & ~w10769;
assign w11901 = pi0078 & w10769;
assign w11902 = ~w11900 & ~w11901;
assign w11903 = w10766 & ~w11902;
assign w11904 = ~w11044 & ~w11738;
assign w11905 = ~w11903 & ~w11904;
assign w11906 = ~w11404 & w11733;
assign w11907 = ~pi0080 & w11308;
assign w11908 = pi0080 & ~w11308;
assign w11909 = ~w11907 & ~w11908;
assign w11910 = w11305 & w11909;
assign w11911 = ~w11906 & ~w11910;
assign w11912 = ~pi0056 & ~w11561;
assign w11913 = pi0056 & w11561;
assign w11914 = ~w11912 & ~w11913;
assign w11915 = w11558 & ~w11914;
assign w11916 = w11672 & ~w11726;
assign w11917 = ~w11915 & ~w11916;
assign w11918 = ~w11911 & w11917;
assign w11919 = w11911 & ~w11917;
assign w11920 = ~w11918 & ~w11919;
assign w11921 = w11905 & ~w11920;
assign w11922 = ~w11905 & w11920;
assign w11923 = ~w11921 & ~w11922;
assign w11924 = w11735 & w11741;
assign w11925 = (~w11924 & w11744) | (~w11924 & w37952) | (w11744 & w37952);
assign w11926 = ~w11923 & w11925;
assign w11927 = ~pi0114 & ~w11813;
assign w11928 = pi0114 & w11813;
assign w11929 = ~w11927 & ~w11928;
assign w11930 = ~pi0868 & ~pi1789;
assign w11931 = ~w11929 & w37953;
assign w11932 = (~w11930 & w11929) | (~w11930 & w37954) | (w11929 & w37954);
assign w11933 = ~w11931 & ~w11932;
assign w11934 = w11923 & ~w11925;
assign w11935 = (w11933 & ~w11923) | (w11933 & w37955) | (~w11923 & w37955);
assign w11936 = ~w11926 & ~w11935;
assign w11937 = w11911 & w11917;
assign w11938 = (~w11937 & w11920) | (~w11937 & w37956) | (w11920 & w37956);
assign w11939 = ~pi0108 & ~w10769;
assign w11940 = pi0108 & w10769;
assign w11941 = ~w11939 & ~w11940;
assign w11942 = w10766 & ~w11941;
assign w11943 = ~w11044 & ~w11902;
assign w11944 = ~w11942 & ~w11943;
assign w11945 = ~pi0106 & ~w11561;
assign w11946 = pi0106 & w11561;
assign w11947 = ~w11945 & ~w11946;
assign w11948 = w11558 & ~w11947;
assign w11949 = w11672 & ~w11914;
assign w11950 = ~w11948 & ~w11949;
assign w11951 = ~w11404 & w11909;
assign w11952 = ~pi0079 & w11308;
assign w11953 = pi0079 & ~w11308;
assign w11954 = ~w11952 & ~w11953;
assign w11955 = w11305 & w11954;
assign w11956 = ~w11951 & ~w11955;
assign w11957 = ~w11950 & w11956;
assign w11958 = w11950 & ~w11956;
assign w11959 = ~w11957 & ~w11958;
assign w11960 = w11944 & ~w11959;
assign w11961 = ~w11944 & w11959;
assign w11962 = ~w11960 & ~w11961;
assign w11963 = ~w11938 & w11962;
assign w11964 = w11938 & ~w11962;
assign w11965 = ~w11963 & ~w11964;
assign w11966 = pi0868 & ~pi1789;
assign w11967 = (~w11966 & w11929) | (~w11966 & w37957) | (w11929 & w37957);
assign w11968 = ~pi0067 & ~w11813;
assign w11969 = pi0067 & w11813;
assign w11970 = ~w11968 & ~w11969;
assign w11971 = w11810 & ~w11970;
assign w11972 = w11835 & ~w11929;
assign w11973 = ~w11971 & ~w11972;
assign w11974 = ~w3613 & w10775;
assign w11975 = ~w11973 & w11974;
assign w11976 = w11973 & ~w11974;
assign w11977 = ~w11975 & ~w11976;
assign w11978 = w11967 & ~w11977;
assign w11979 = ~w11967 & w11977;
assign w11980 = ~w11978 & ~w11979;
assign w11981 = w11965 & ~w11980;
assign w11982 = ~w11965 & w11980;
assign w11983 = ~w11981 & ~w11982;
assign w11984 = ~w11936 & ~w11983;
assign w11985 = w11936 & w11983;
assign w11986 = ~w11984 & ~w11985;
assign w11987 = ~w11899 & ~w11986;
assign w11988 = w11899 & w11986;
assign w11989 = ~w11987 & ~w11988;
assign w11990 = ~w11926 & ~w11934;
assign w11991 = w11933 & ~w11990;
assign w11992 = ~w11933 & w11990;
assign w11993 = ~w11991 & ~w11992;
assign w11994 = ~w11750 & w11993;
assign w11995 = (~w11582 & w11552) | (~w11582 & w37958) | (w11552 & w37958);
assign w11996 = (~w11995 & w11665) | (~w11995 & w37959) | (w11665 & w37959);
assign w11997 = w11663 & w11688;
assign w11998 = ~w11692 & ~w11997;
assign w11999 = ~w11996 & w11998;
assign w12000 = ~w11891 & ~w11893;
assign w12001 = w11886 & ~w12000;
assign w12002 = ~w11886 & w12000;
assign w12003 = ~w12001 & ~w12002;
assign w12004 = ~w11999 & w12003;
assign w12005 = (~w11994 & ~w12003) | (~w11994 & w37960) | (~w12003 & w37960);
assign w12006 = ~w11989 & w12005;
assign w12007 = w12003 & w37961;
assign w12008 = ~w12005 & ~w12007;
assign w12009 = w11989 & w12008;
assign w12010 = ~w12006 & ~w12009;
assign w12011 = w11750 & ~w11993;
assign w12012 = ~w11994 & ~w12011;
assign w12013 = w11999 & ~w12003;
assign w12014 = ~w12004 & ~w12013;
assign w12015 = ~w12012 & ~w12014;
assign w12016 = (~w11753 & ~w11715) | (~w11753 & w37962) | (~w11715 & w37962);
assign w12017 = ~w11552 & w37963;
assign w12018 = ~w11588 & ~w12017;
assign w12019 = ~w11702 & w12018;
assign w12020 = ~w11753 & w12019;
assign w12021 = (~w12020 & ~w11713) | (~w12020 & w37964) | (~w11713 & w37964);
assign w12022 = ~w12015 & w12021;
assign w12023 = w12012 & w12014;
assign w12024 = ~w12022 & ~w12023;
assign w12025 = ~w12010 & w12024;
assign w12026 = ~w11752 & ~w12019;
assign w12027 = ~w11755 & ~w12026;
assign w12028 = (w12027 & ~w11713) | (w12027 & w37965) | (~w11713 & w37965);
assign w12029 = (~w12028 & w11758) | (~w12028 & w37966) | (w11758 & w37966);
assign w12030 = ~w12015 & ~w12023;
assign w12031 = w12021 & ~w12030;
assign w12032 = ~w12021 & w12030;
assign w12033 = ~w12031 & ~w12032;
assign w12034 = ~w12029 & w12033;
assign w12035 = ~w12025 & ~w12034;
assign w12036 = w11777 & w12035;
assign w12037 = ~w11636 & w12036;
assign w12038 = (~w12011 & w12003) | (~w12011 & w37967) | (w12003 & w37967);
assign w12039 = ~w11999 & ~w12038;
assign w12040 = (w12039 & w12021) | (w12039 & w37968) | (w12021 & w37968);
assign w12041 = w11994 & w12003;
assign w12042 = (w11999 & ~w12003) | (w11999 & w37960) | (~w12003 & w37960);
assign w12043 = ~w12003 & w12011;
assign w12044 = w12042 & ~w12043;
assign w12045 = w12021 & w12044;
assign w12046 = w12038 & w12042;
assign w12047 = ~w11989 & ~w12046;
assign w12048 = w12047 & w37969;
assign w12049 = w12038 & ~w12042;
assign w12050 = w12021 & w12049;
assign w12051 = ~w12041 & ~w12043;
assign w12052 = ~w12014 & ~w12051;
assign w12053 = w11989 & ~w12052;
assign w12054 = ~w12050 & w12053;
assign w12055 = ~w12048 & ~w12054;
assign w12056 = ~w11994 & ~w12014;
assign w12057 = ~w12021 & w12056;
assign w12058 = w12010 & w12057;
assign w12059 = w11989 & ~w12011;
assign w12060 = ~w11989 & ~w11994;
assign w12061 = ~w12004 & ~w12021;
assign w12062 = ~w12060 & w12061;
assign w12063 = ~w12059 & w12062;
assign w12064 = ~w12058 & ~w12063;
assign w12065 = w12064 & w37970;
assign w12066 = ~w11592 & w37971;
assign w12067 = w11758 & ~w12066;
assign w12068 = w11420 & ~w11526;
assign w12069 = w11592 & w12068;
assign w12070 = w11420 & w11526;
assign w12071 = ~w11592 & w12070;
assign w12072 = ~w12069 & ~w12071;
assign w12073 = w11713 & w40078;
assign w12074 = w11755 & w12072;
assign w12075 = (~w11771 & w11722) | (~w11771 & w37972) | (w11722 & w37972);
assign w12076 = ~w12073 & w12075;
assign w12077 = ~w12067 & w12076;
assign w12078 = (~w11763 & ~w11592) | (~w11763 & w37973) | (~w11592 & w37973);
assign w12079 = ~w11759 & w12078;
assign w12080 = w12072 & w12079;
assign w12081 = w11758 & ~w12080;
assign w12082 = w11595 & w11763;
assign w12083 = (~w11770 & w11526) | (~w11770 & w37974) | (w11526 & w37974);
assign w12084 = w11765 & w12083;
assign w12085 = (w12084 & w12082) | (w12084 & w37975) | (w12082 & w37975);
assign w12086 = ~w11758 & ~w12085;
assign w12087 = ~w12081 & ~w12086;
assign w12088 = ~w12077 & ~w12087;
assign w12089 = w12029 & ~w12033;
assign w12090 = w12088 & ~w12089;
assign w12091 = w12035 & ~w12090;
assign w12092 = ~w12065 & ~w12091;
assign w12093 = ~w12037 & w12092;
assign w12094 = w11848 & w11877;
assign w12095 = ~w11880 & ~w12094;
assign w12096 = ~w11883 & w12095;
assign w12097 = (~w11842 & ~w11844) | (~w11842 & w37976) | (~w11844 & w37976);
assign w12098 = ~pi0077 & ~pi1647;
assign w12099 = ~pi1424 & w12098;
assign w12100 = pi0081 & pi1640;
assign w12101 = pi0081 & ~pi1640;
assign w12102 = w10794 & w12101;
assign w12103 = (w11201 & w12102) | (w11201 & w37977) | (w12102 & w37977);
assign w12104 = ~pi0066 & pi0104;
assign w12105 = w11202 & w37978;
assign w12106 = ~w12103 & ~w12105;
assign w12107 = (~w12100 & ~w11202) | (~w12100 & w37979) | (~w11202 & w37979);
assign w12108 = ~w11837 & w12100;
assign w12109 = w12106 & w12108;
assign w12110 = ~w12107 & ~w12109;
assign w12111 = (w12106 & w12109) | (w12106 & w37981) | (w12109 & w37981);
assign w12112 = ~w12099 & w12111;
assign w12113 = w12099 & ~w12111;
assign w12114 = ~w12112 & ~w12113;
assign w12115 = w12097 & ~w12114;
assign w12116 = ~w12097 & w12114;
assign w12117 = ~w12115 & ~w12116;
assign w12118 = ~w11848 & ~w11877;
assign w12119 = ~w11864 & ~w11870;
assign w12120 = (~w12119 & w11873) | (~w12119 & w37982) | (w11873 & w37982);
assign w12121 = ~pi0111 & ~w10835;
assign w12122 = pi0111 & w10835;
assign w12123 = ~w12121 & ~w12122;
assign w12124 = w10832 & ~w12123;
assign w12125 = w10842 & ~w11855;
assign w12126 = ~w12124 & ~w12125;
assign w12127 = ~pi0113 & ~w10782;
assign w12128 = pi0113 & w10782;
assign w12129 = ~w12127 & ~w12128;
assign w12130 = w10809 & ~w12129;
assign w12131 = w10787 & ~w11861;
assign w12132 = ~w12130 & ~w12131;
assign w12133 = ~w10860 & ~w11868;
assign w12134 = ~pi0109 & w10853;
assign w12135 = pi0109 & ~w10853;
assign w12136 = ~w12134 & ~w12135;
assign w12137 = w10850 & ~w12136;
assign w12138 = ~w12133 & ~w12137;
assign w12139 = ~w12132 & ~w12138;
assign w12140 = w12132 & w12138;
assign w12141 = ~w12139 & ~w12140;
assign w12142 = w12126 & ~w12141;
assign w12143 = ~w12126 & w12141;
assign w12144 = ~w12142 & ~w12143;
assign w12145 = w12120 & ~w12144;
assign w12146 = ~w12120 & w12144;
assign w12147 = ~w12145 & ~w12146;
assign w12148 = ~w12118 & w12147;
assign w12149 = w12118 & ~w12147;
assign w12150 = ~w12148 & ~w12149;
assign w12151 = w12117 & w12150;
assign w12152 = ~w12117 & ~w12150;
assign w12153 = ~w12151 & ~w12152;
assign w12154 = ~w12096 & w12153;
assign w12155 = ~w11931 & ~w11980;
assign w12156 = ~w11963 & ~w12155;
assign w12157 = w11950 & w11956;
assign w12158 = (~w12157 & w11959) | (~w12157 & w37983) | (w11959 & w37983);
assign w12159 = ~pi0107 & ~w10769;
assign w12160 = pi0107 & w10769;
assign w12161 = ~w12159 & ~w12160;
assign w12162 = w10766 & ~w12161;
assign w12163 = ~w11044 & ~w11941;
assign w12164 = ~w12162 & ~w12163;
assign w12165 = ~w11404 & w11954;
assign w12166 = ~pi0078 & w11308;
assign w12167 = pi0078 & ~w11308;
assign w12168 = ~w12166 & ~w12167;
assign w12169 = w11305 & w12168;
assign w12170 = ~w12165 & ~w12169;
assign w12171 = ~pi0080 & ~w11561;
assign w12172 = pi0080 & w11561;
assign w12173 = ~w12171 & ~w12172;
assign w12174 = w11558 & ~w12173;
assign w12175 = w11672 & ~w11947;
assign w12176 = ~w12174 & ~w12175;
assign w12177 = ~w12170 & w12176;
assign w12178 = w12170 & ~w12176;
assign w12179 = ~w12177 & ~w12178;
assign w12180 = ~w12164 & ~w12179;
assign w12181 = w12164 & w12179;
assign w12182 = ~w12180 & ~w12181;
assign w12183 = ~w12158 & ~w12182;
assign w12184 = w12158 & w12182;
assign w12185 = ~w12183 & ~w12184;
assign w12186 = ~w11966 & ~w11974;
assign w12187 = ~w11973 & ~w12186;
assign w12188 = ~pi0056 & ~w11813;
assign w12189 = pi0056 & w11813;
assign w12190 = ~w12188 & ~w12189;
assign w12191 = w11810 & ~w12190;
assign w12192 = w11835 & ~w11970;
assign w12193 = ~w12191 & ~w12192;
assign w12194 = ~pi0114 & pi1424;
assign w12195 = pi0114 & ~pi1473;
assign w12196 = w12098 & ~w12195;
assign w12197 = ~w12194 & w12196;
assign w12198 = ~w3613 & w10777;
assign w12199 = ~w4695 & w10775;
assign w12200 = ~w12198 & ~w12199;
assign w12201 = ~w12197 & w12200;
assign w12202 = w12197 & ~w12200;
assign w12203 = ~w12201 & ~w12202;
assign w12204 = w12193 & ~w12203;
assign w12205 = ~w12193 & w12203;
assign w12206 = ~w12204 & ~w12205;
assign w12207 = ~w12187 & ~w12206;
assign w12208 = w12187 & w12206;
assign w12209 = ~w12207 & ~w12208;
assign w12210 = w12185 & w12209;
assign w12211 = ~w12185 & ~w12209;
assign w12212 = ~w12210 & ~w12211;
assign w12213 = w11963 & ~w11980;
assign w12214 = w11931 & w11977;
assign w12215 = (~w12214 & w12213) | (~w12214 & w37984) | (w12213 & w37984);
assign w12216 = ~w11964 & ~w12215;
assign w12217 = w11964 & w12155;
assign w12218 = ~w11963 & w11980;
assign w12219 = ~w11935 & w12218;
assign w12220 = ~w12217 & ~w12219;
assign w12221 = ~w12216 & w12220;
assign w12222 = w12212 & ~w12221;
assign w12223 = (w12156 & w12221) | (w12156 & w37985) | (w12221 & w37985);
assign w12224 = ~w12212 & w12221;
assign w12225 = (~w12156 & ~w12221) | (~w12156 & w37986) | (~w12221 & w37986);
assign w12226 = ~w12223 & ~w12225;
assign w12227 = ~w12154 & ~w12226;
assign w12228 = ~w12156 & ~w12211;
assign w12229 = ~w12182 & w37987;
assign w12230 = (~w12229 & ~w12185) | (~w12229 & w37988) | (~w12185 & w37988);
assign w12231 = ~w12228 & w12230;
assign w12232 = (~w12207 & w12182) | (~w12207 & w37989) | (w12182 & w37989);
assign w12233 = ~w12170 & ~w12176;
assign w12234 = (~w12233 & w12179) | (~w12233 & w37990) | (w12179 & w37990);
assign w12235 = ~pi0108 & w11308;
assign w12236 = pi0108 & ~w11308;
assign w12237 = ~w12235 & ~w12236;
assign w12238 = w11305 & w12237;
assign w12239 = ~w11404 & w12168;
assign w12240 = ~w12238 & ~w12239;
assign w12241 = ~pi0105 & ~w10769;
assign w12242 = pi0105 & w10769;
assign w12243 = ~w12241 & ~w12242;
assign w12244 = w10766 & ~w12243;
assign w12245 = ~w11044 & ~w12161;
assign w12246 = ~w12244 & ~w12245;
assign w12247 = ~pi0079 & ~w11561;
assign w12248 = pi0079 & w11561;
assign w12249 = ~w12247 & ~w12248;
assign w12250 = w11558 & ~w12249;
assign w12251 = w11672 & ~w12173;
assign w12252 = ~w12250 & ~w12251;
assign w12253 = w12246 & w12252;
assign w12254 = ~w12246 & ~w12252;
assign w12255 = ~w12253 & ~w12254;
assign w12256 = w12240 & ~w12255;
assign w12257 = ~w12240 & w12255;
assign w12258 = ~w12256 & ~w12257;
assign w12259 = w12234 & ~w12258;
assign w12260 = ~w12234 & w12258;
assign w12261 = ~w12259 & ~w12260;
assign w12262 = ~w12232 & w12261;
assign w12263 = w12232 & ~w12261;
assign w12264 = ~w12262 & ~w12263;
assign w12265 = ~pi0106 & ~w11813;
assign w12266 = pi0106 & w11813;
assign w12267 = ~w12265 & ~w12266;
assign w12268 = w11810 & ~w12267;
assign w12269 = w11835 & ~w12190;
assign w12270 = ~w12268 & ~w12269;
assign w12271 = ~w5718 & w10775;
assign w12272 = ~w4695 & w10777;
assign w12273 = ~w12271 & ~w12272;
assign w12274 = ~pi0067 & ~pi1424;
assign w12275 = ~w11196 & ~w12274;
assign w12276 = w12098 & ~w12275;
assign w12277 = ~w12273 & w12276;
assign w12278 = w12273 & ~w12276;
assign w12279 = ~w12277 & ~w12278;
assign w12280 = w12270 & w12279;
assign w12281 = ~w12270 & ~w12279;
assign w12282 = ~w12280 & ~w12281;
assign w12283 = (~w12201 & ~w12193) | (~w12201 & w37991) | (~w12193 & w37991);
assign w12284 = w12282 & ~w12283;
assign w12285 = ~w12282 & w12283;
assign w12286 = ~w12284 & ~w12285;
assign w12287 = w12264 & ~w12286;
assign w12288 = ~w12264 & w12286;
assign w12289 = ~w12287 & ~w12288;
assign w12290 = ~w12231 & ~w12289;
assign w12291 = w12231 & w12289;
assign w12292 = ~w12290 & ~w12291;
assign w12293 = ~w12144 & w37992;
assign w12294 = ~w12148 & ~w12293;
assign w12295 = (~w12115 & w12144) | (~w12115 & w37993) | (w12144 & w37993);
assign w12296 = ~pi0081 & w10853;
assign w12297 = pi0081 & ~w10853;
assign w12298 = ~w12296 & ~w12297;
assign w12299 = w10850 & ~w12298;
assign w12300 = ~w10860 & ~w12136;
assign w12301 = ~w12299 & ~w12300;
assign w12302 = ~pi0112 & ~w10782;
assign w12303 = pi0112 & w10782;
assign w12304 = ~w12302 & ~w12303;
assign w12305 = w10809 & ~w12304;
assign w12306 = w10787 & ~w12129;
assign w12307 = ~w12305 & ~w12306;
assign w12308 = ~pi0110 & ~w10835;
assign w12309 = pi0110 & w10835;
assign w12310 = ~w12308 & ~w12309;
assign w12311 = w10832 & ~w12310;
assign w12312 = w10842 & ~w12123;
assign w12313 = ~w12311 & ~w12312;
assign w12314 = ~w12307 & w12313;
assign w12315 = w12307 & ~w12313;
assign w12316 = ~w12314 & ~w12315;
assign w12317 = ~w12301 & ~w12316;
assign w12318 = w12301 & w12316;
assign w12319 = ~w12317 & ~w12318;
assign w12320 = ~w12126 & ~w12140;
assign w12321 = ~w12139 & ~w12320;
assign w12322 = w12099 & w12102;
assign w12323 = (~w12322 & w12109) | (~w12322 & w37995) | (w12109 & w37995);
assign w12324 = (w12323 & w12320) | (w12323 & w40049) | (w12320 & w40049);
assign w12325 = ~w12320 & w37996;
assign w12326 = ~w12324 & ~w12325;
assign w12327 = w12319 & ~w12326;
assign w12328 = ~w12319 & w12326;
assign w12329 = ~w12327 & ~w12328;
assign w12330 = ~w12295 & w12329;
assign w12331 = w12295 & ~w12329;
assign w12332 = ~w12330 & ~w12331;
assign w12333 = (w12332 & w12151) | (w12332 & w40050) | (w12151 & w40050);
assign w12334 = ~w12151 & w40051;
assign w12335 = ~w12333 & ~w12334;
assign w12336 = w12292 & w12335;
assign w12337 = ~w12292 & ~w12335;
assign w12338 = ~w12336 & ~w12337;
assign w12339 = ~w12227 & w12338;
assign w12340 = w12290 & w12333;
assign w12341 = ~w12336 & ~w12340;
assign w12342 = ~w12339 & w12341;
assign w12343 = w12099 & ~w12106;
assign w12344 = ~w12110 & ~w12343;
assign w12345 = ~w12319 & w37997;
assign w12346 = w12319 & ~w12321;
assign w12347 = (~w12323 & w12319) | (~w12323 & w37998) | (w12319 & w37998);
assign w12348 = ~w12346 & w12347;
assign w12349 = ~w12345 & ~w12348;
assign w12350 = ~w12330 & w12349;
assign w12351 = ~w12307 & ~w12313;
assign w12352 = (~w12351 & w12316) | (~w12351 & w37999) | (w12316 & w37999);
assign w12353 = ~pi1640 & ~w10848;
assign w12354 = pi0097 & ~w10848;
assign w12355 = (pi1424 & w10848) | (pi1424 & w38000) | (w10848 & w38000);
assign w12356 = ~w12353 & w12355;
assign w12357 = pi0097 & pi1640;
assign w12358 = ~w10849 & ~w12357;
assign w12359 = (pi0081 & w12358) | (pi0081 & w38001) | (w12358 & w38001);
assign w12360 = ~w12356 & w12359;
assign w12361 = ~w12296 & ~w12360;
assign w12362 = ~pi1424 & ~pi1640;
assign w12363 = w10850 & ~w12362;
assign w12364 = ~w10858 & ~w12354;
assign w12365 = ~w12363 & w12364;
assign w12366 = w10851 & w12358;
assign w12367 = ~w12365 & ~w12366;
assign w12368 = ~w12361 & w12367;
assign w12369 = ~pi0109 & ~w10835;
assign w12370 = pi0109 & w10835;
assign w12371 = ~w12369 & ~w12370;
assign w12372 = w10832 & ~w12371;
assign w12373 = w10842 & ~w12310;
assign w12374 = ~w12372 & ~w12373;
assign w12375 = ~pi0111 & ~w10782;
assign w12376 = pi0111 & w10782;
assign w12377 = ~w12375 & ~w12376;
assign w12378 = w10809 & ~w12377;
assign w12379 = w10787 & ~w12304;
assign w12380 = ~w12378 & ~w12379;
assign w12381 = ~w12374 & ~w12380;
assign w12382 = w12374 & w12380;
assign w12383 = ~w12381 & ~w12382;
assign w12384 = ~w12368 & w12383;
assign w12385 = w12368 & ~w12383;
assign w12386 = ~w12384 & ~w12385;
assign w12387 = w12352 & w12386;
assign w12388 = ~w12352 & ~w12386;
assign w12389 = ~w12387 & ~w12388;
assign w12390 = ~w12319 & w38002;
assign w12391 = w11201 & w12322;
assign w12392 = (w12391 & w12319) | (w12391 & w38003) | (w12319 & w38003);
assign w12393 = ~w12390 & ~w12392;
assign w12394 = w12389 & ~w12393;
assign w12395 = ~w12389 & w12393;
assign w12396 = ~w12394 & ~w12395;
assign w12397 = ~w12350 & ~w12396;
assign w12398 = w12350 & w12396;
assign w12399 = ~w12397 & ~w12398;
assign w12400 = (w12399 & w12290) | (w12399 & w40052) | (w12290 & w40052);
assign w12401 = ~w12290 & w40053;
assign w12402 = ~w12400 & ~w12401;
assign w12403 = ~w11044 & ~w12243;
assign w12404 = ~pi0113 & ~w10769;
assign w12405 = pi0113 & w10769;
assign w12406 = ~w12404 & ~w12405;
assign w12407 = w10766 & ~w12406;
assign w12408 = ~w12403 & ~w12407;
assign w12409 = ~w11404 & w12237;
assign w12410 = ~pi0107 & w11308;
assign w12411 = pi0107 & ~w11308;
assign w12412 = w11305 & ~w12411;
assign w12413 = ~w12410 & w12412;
assign w12414 = ~w12409 & ~w12413;
assign w12415 = w11672 & ~w12249;
assign w12416 = ~pi0078 & ~w11561;
assign w12417 = pi0078 & w11561;
assign w12418 = ~w12416 & ~w12417;
assign w12419 = w11558 & ~w12418;
assign w12420 = ~w12415 & ~w12419;
assign w12421 = ~w12414 & w12420;
assign w12422 = w12414 & ~w12420;
assign w12423 = ~w12421 & ~w12422;
assign w12424 = ~w12408 & ~w12423;
assign w12425 = w12408 & w12423;
assign w12426 = ~w12424 & ~w12425;
assign w12427 = ~w12240 & ~w12253;
assign w12428 = ~w12254 & ~w12427;
assign w12429 = (~w12277 & w12270) | (~w12277 & w38004) | (w12270 & w38004);
assign w12430 = ~w12427 & w40054;
assign w12431 = ~w12426 & w12430;
assign w12432 = ~pi0080 & ~w11813;
assign w12433 = pi0080 & w11813;
assign w12434 = ~w12432 & ~w12433;
assign w12435 = w11810 & ~w12434;
assign w12436 = w11835 & ~w12267;
assign w12437 = ~w12435 & ~w12436;
assign w12438 = ~w5718 & w10777;
assign w12439 = ~w5123 & w10775;
assign w12440 = ~w12438 & ~w12439;
assign w12441 = ~pi0056 & ~pi1424;
assign w12442 = ~w11155 & ~w12441;
assign w12443 = w12098 & ~w12442;
assign w12444 = ~w12440 & w12443;
assign w12445 = w12440 & ~w12443;
assign w12446 = ~w12444 & ~w12445;
assign w12447 = ~w12437 & w12446;
assign w12448 = w12437 & ~w12446;
assign w12449 = ~w12447 & ~w12448;
assign w12450 = w12429 & ~w12449;
assign w12451 = ~w12429 & w12449;
assign w12452 = ~w12450 & ~w12451;
assign w12453 = ~w12431 & ~w12452;
assign w12454 = ~w12426 & w40055;
assign w12455 = ~w12453 & ~w12454;
assign w12456 = ~w12427 & w38005;
assign w12457 = ~w12426 & w12456;
assign w12458 = w12426 & ~w12428;
assign w12459 = ~w12457 & ~w12458;
assign w12460 = w12455 & ~w12459;
assign w12461 = ~w12455 & w12459;
assign w12462 = ~w12460 & ~w12461;
assign w12463 = ~w12207 & ~w12284;
assign w12464 = ~w12183 & w12463;
assign w12465 = ~w12261 & w12464;
assign w12466 = ~w12285 & ~w12465;
assign w12467 = ~w12262 & ~w12466;
assign w12468 = (~w12284 & w12258) | (~w12284 & w38006) | (w12258 & w38006);
assign w12469 = (~w12259 & ~w12261) | (~w12259 & w38007) | (~w12261 & w38007);
assign w12470 = ~w12468 & ~w12469;
assign w12471 = (w12259 & w12465) | (w12259 & w38008) | (w12465 & w38008);
assign w12472 = (~w12471 & w12467) | (~w12471 & w38009) | (w12467 & w38009);
assign w12473 = w12462 & w12472;
assign w12474 = ~w12462 & ~w12472;
assign w12475 = ~w12473 & ~w12474;
assign w12476 = w12402 & ~w12475;
assign w12477 = ~w12402 & w12475;
assign w12478 = ~w12476 & ~w12477;
assign w12479 = w12342 & w12478;
assign w12480 = w12227 & ~w12338;
assign w12481 = ~w12339 & ~w12480;
assign w12482 = w12096 & ~w12153;
assign w12483 = ~w12154 & ~w12482;
assign w12484 = w11935 & ~w11983;
assign w12485 = ~w11985 & ~w12484;
assign w12486 = ~w11897 & w12485;
assign w12487 = ~w12222 & ~w12224;
assign w12488 = ~w12486 & w12487;
assign w12489 = w12486 & ~w12487;
assign w12490 = ~w12488 & ~w12489;
assign w12491 = w12483 & w12490;
assign w12492 = w12154 & w12226;
assign w12493 = ~w12488 & ~w12492;
assign w12494 = ~w12491 & w12493;
assign w12495 = ~w12481 & w12494;
assign w12496 = (~w12005 & w11899) | (~w12005 & w38010) | (w11899 & w38010);
assign w12497 = w11897 & ~w12485;
assign w12498 = ~w11988 & ~w12497;
assign w12499 = ~w12496 & w12498;
assign w12500 = ~w12483 & ~w12490;
assign w12501 = ~w12491 & ~w12500;
assign w12502 = w12499 & ~w12501;
assign w12503 = ~w12495 & ~w12502;
assign w12504 = ~w12479 & w12503;
assign w12505 = (w12504 & w12037) | (w12504 & w38011) | (w12037 & w38011);
assign w12506 = w11835 & ~w12434;
assign w12507 = ~pi0079 & w11813;
assign w12508 = pi0079 & ~w11813;
assign w12509 = w11810 & ~w12508;
assign w12510 = ~w12507 & w12509;
assign w12511 = ~w12506 & ~w12510;
assign w12512 = ~pi0106 & ~pi1424;
assign w12513 = ~w11094 & ~w12512;
assign w12514 = w12098 & ~w12513;
assign w12515 = ~w12511 & w12514;
assign w12516 = ~w5123 & w10777;
assign w12517 = ~w4339 & w10775;
assign w12518 = ~w12516 & ~w12517;
assign w12519 = w12511 & ~w12514;
assign w12520 = ~w12515 & ~w12519;
assign w12521 = ~w12518 & w12520;
assign w12522 = (~w12515 & ~w12520) | (~w12515 & w38012) | (~w12520 & w38012);
assign w12523 = ~w6330 & w10775;
assign w12524 = ~w4339 & w10777;
assign w12525 = ~w12523 & ~w12524;
assign w12526 = ~pi0079 & w11835;
assign w12527 = ~pi0078 & w11810;
assign w12528 = ~w12526 & ~w12527;
assign w12529 = (~w11813 & w12526) | (~w11813 & w38013) | (w12526 & w38013);
assign w12530 = pi1471 & w11808;
assign w12531 = ~pi1471 & w11809;
assign w12532 = ~w12530 & ~w12531;
assign w12533 = w11813 & w12532;
assign w12534 = w12528 & w12533;
assign w12535 = (~w12525 & w12534) | (~w12525 & w38014) | (w12534 & w38014);
assign w12536 = ~w12534 & w38015;
assign w12537 = ~w12535 & ~w12536;
assign w12538 = ~pi0080 & ~pi1424;
assign w12539 = ~w10912 & ~w12538;
assign w12540 = w12098 & ~w12539;
assign w12541 = ~w12537 & w12540;
assign w12542 = w12537 & ~w12540;
assign w12543 = ~w12541 & ~w12542;
assign w12544 = w12522 & w12543;
assign w12545 = ~w12522 & ~w12543;
assign w12546 = ~w12544 & ~w12545;
assign w12547 = ~w12414 & ~w12420;
assign w12548 = (~w12547 & w12423) | (~w12547 & w38016) | (w12423 & w38016);
assign w12549 = w11672 & ~w12418;
assign w12550 = pi0108 & ~w11561;
assign w12551 = ~pi0108 & w11561;
assign w12552 = w11558 & ~w12551;
assign w12553 = ~w12550 & w12552;
assign w12554 = ~w12549 & ~w12553;
assign w12555 = ~w11044 & ~w12406;
assign w12556 = ~pi0112 & ~w10769;
assign w12557 = pi0112 & w10769;
assign w12558 = ~w12556 & ~w12557;
assign w12559 = w10766 & ~w12558;
assign w12560 = ~w12555 & ~w12559;
assign w12561 = ~pi0098 & pi0102;
assign w12562 = ~w11304 & ~w12561;
assign w12563 = pi0102 & pi0103;
assign w12564 = ~pi0107 & ~w12563;
assign w12565 = ~w12562 & w12564;
assign w12566 = ~pi0105 & w11305;
assign w12567 = ~w12565 & ~w12566;
assign w12568 = w11308 & ~w12567;
assign w12569 = ~pi0102 & ~pi1470;
assign w12570 = ~w11303 & w12569;
assign w12571 = pi0102 & pi1470;
assign w12572 = ~w11304 & w12571;
assign w12573 = ~w12570 & ~w12572;
assign w12574 = w12567 & w12573;
assign w12575 = ~w12568 & ~w12574;
assign w12576 = ~w12560 & w12575;
assign w12577 = w12560 & ~w12575;
assign w12578 = ~w12576 & ~w12577;
assign w12579 = ~w12554 & w12578;
assign w12580 = w12554 & ~w12578;
assign w12581 = ~w12579 & ~w12580;
assign w12582 = w12548 & ~w12581;
assign w12583 = w12518 & ~w12520;
assign w12584 = ~w12521 & ~w12583;
assign w12585 = ~w12444 & ~w12447;
assign w12586 = ~w12584 & w12585;
assign w12587 = ~w12582 & ~w12586;
assign w12588 = ~w11044 & ~w12558;
assign w12589 = ~pi0111 & ~w10769;
assign w12590 = pi0111 & w10769;
assign w12591 = ~w12589 & ~w12590;
assign w12592 = w10766 & ~w12591;
assign w12593 = ~w12588 & ~w12592;
assign w12594 = ~pi0105 & ~w12563;
assign w12595 = ~w12562 & w12594;
assign w12596 = ~pi0113 & w11305;
assign w12597 = ~w12595 & ~w12596;
assign w12598 = w11308 & ~w12597;
assign w12599 = w12573 & w12597;
assign w12600 = ~w12598 & ~w12599;
assign w12601 = ~w12593 & w12600;
assign w12602 = w12593 & ~w12600;
assign w12603 = ~w12601 & ~w12602;
assign w12604 = ~pi0108 & w11672;
assign w12605 = ~pi0107 & w11558;
assign w12606 = ~w12604 & ~w12605;
assign w12607 = (~w11561 & w12604) | (~w11561 & w38017) | (w12604 & w38017);
assign w12608 = ~w11558 & ~w11672;
assign w12609 = (w11561 & w11672) | (w11561 & w38018) | (w11672 & w38018);
assign w12610 = w12606 & w12609;
assign w12611 = ~w12607 & ~w12610;
assign w12612 = w12603 & ~w12611;
assign w12613 = ~w12603 & w12611;
assign w12614 = ~w12612 & ~w12613;
assign w12615 = (~w12576 & ~w12578) | (~w12576 & w38019) | (~w12578 & w38019);
assign w12616 = ~w12614 & w12615;
assign w12617 = w12614 & ~w12615;
assign w12618 = ~w12616 & ~w12617;
assign w12619 = w12587 & ~w12618;
assign w12620 = ~w12587 & w12618;
assign w12621 = ~w12619 & ~w12620;
assign w12622 = ~w12546 & w12621;
assign w12623 = w12546 & ~w12621;
assign w12624 = ~w12622 & ~w12623;
assign w12625 = (~w12450 & w12426) | (~w12450 & w38020) | (w12426 & w38020);
assign w12626 = ~w12548 & w12581;
assign w12627 = ~w12582 & ~w12626;
assign w12628 = w12584 & ~w12585;
assign w12629 = ~w12586 & ~w12628;
assign w12630 = w12627 & w12629;
assign w12631 = ~w12627 & ~w12629;
assign w12632 = ~w12630 & ~w12631;
assign w12633 = ~w12625 & w12632;
assign w12634 = w12582 & w12586;
assign w12635 = ~w12630 & ~w12634;
assign w12636 = ~w12633 & w12635;
assign w12637 = ~w12624 & ~w12636;
assign w12638 = w12624 & w12636;
assign w12639 = ~w12637 & ~w12638;
assign w12640 = pi0081 & w10835;
assign w12641 = ~pi0081 & ~w10835;
assign w12642 = ~w12640 & ~w12641;
assign w12643 = w10832 & ~w12642;
assign w12644 = w10842 & ~w12371;
assign w12645 = ~w12643 & ~w12644;
assign w12646 = ~w10853 & ~w12100;
assign w12647 = w10853 & w12100;
assign w12648 = ~w12646 & ~w12647;
assign w12649 = ~w12365 & w12648;
assign w12650 = ~pi0110 & ~w10782;
assign w12651 = pi0110 & w10782;
assign w12652 = ~w12650 & ~w12651;
assign w12653 = w10809 & ~w12652;
assign w12654 = w10787 & ~w12377;
assign w12655 = ~w12653 & ~w12654;
assign w12656 = ~w12649 & w12655;
assign w12657 = w12649 & ~w12655;
assign w12658 = ~w12656 & ~w12657;
assign w12659 = w12645 & ~w12658;
assign w12660 = ~w12645 & w12658;
assign w12661 = ~w12659 & ~w12660;
assign w12662 = w12368 & ~w12382;
assign w12663 = ~w12381 & ~w12662;
assign w12664 = ~w12661 & w12663;
assign w12665 = ~w12661 & w38021;
assign w12666 = w12387 & w12665;
assign w12667 = w12386 & w38022;
assign w12668 = w12661 & ~w12663;
assign w12669 = ~w12667 & w12668;
assign w12670 = ~w12666 & ~w12669;
assign w12671 = w10787 & ~w12652;
assign w12672 = ~pi0109 & ~w10782;
assign w12673 = pi0109 & w10782;
assign w12674 = ~w12672 & ~w12673;
assign w12675 = w10809 & ~w12674;
assign w12676 = ~w12671 & ~w12675;
assign w12677 = ~pi1468 & ~pi1640;
assign w12678 = ~w10831 & ~w12677;
assign w12679 = w10840 & ~w12678;
assign w12680 = (~w10830 & ~w12678) | (~w10830 & w38023) | (~w12678 & w38023);
assign w12681 = pi0075 & ~w12680;
assign w12682 = ~w12679 & ~w12681;
assign w12683 = ~w10835 & ~w12100;
assign w12684 = ~w12640 & ~w12683;
assign w12685 = pi1468 & ~w10830;
assign w12686 = (pi0081 & w10831) | (pi0081 & w38024) | (w10831 & w38024);
assign w12687 = ~w12685 & w12686;
assign w12688 = ~w12684 & ~w12687;
assign w12689 = w12682 & w12688;
assign w12690 = ~w12676 & w12689;
assign w12691 = w12676 & ~w12689;
assign w12692 = ~w12690 & ~w12691;
assign w12693 = w12645 & ~w12655;
assign w12694 = ~w12645 & w12649;
assign w12695 = ~w12656 & ~w12694;
assign w12696 = ~w12693 & w12695;
assign w12697 = w12692 & ~w12696;
assign w12698 = ~w12692 & w12696;
assign w12699 = ~w12697 & ~w12698;
assign w12700 = ~w12670 & w12699;
assign w12701 = w12670 & ~w12699;
assign w12702 = ~w12700 & ~w12701;
assign w12703 = ~w12639 & w12702;
assign w12704 = w12639 & ~w12702;
assign w12705 = ~w12703 & ~w12704;
assign w12706 = ~w12664 & ~w12668;
assign w12707 = ~w12387 & w12706;
assign w12708 = w12387 & ~w12706;
assign w12709 = ~w12707 & ~w12708;
assign w12710 = (~w12390 & ~w12389) | (~w12390 & w38025) | (~w12389 & w38025);
assign w12711 = w12709 & ~w12710;
assign w12712 = ~w12706 & w38026;
assign w12713 = (~w12712 & ~w12709) | (~w12712 & w38027) | (~w12709 & w38027);
assign w12714 = w12625 & ~w12632;
assign w12715 = ~w12633 & ~w12714;
assign w12716 = w12459 & ~w12468;
assign w12717 = ~w12455 & ~w12716;
assign w12718 = ~w12459 & w12468;
assign w12719 = ~w12717 & ~w12718;
assign w12720 = w12715 & w12719;
assign w12721 = (w12713 & ~w12715) | (w12713 & w38028) | (~w12715 & w38028);
assign w12722 = w12705 & ~w12721;
assign w12723 = ~w12705 & w12721;
assign w12724 = ~w12722 & ~w12723;
assign w12725 = ~w12709 & w12710;
assign w12726 = ~w12711 & ~w12725;
assign w12727 = ~w12715 & ~w12719;
assign w12728 = ~w12720 & ~w12727;
assign w12729 = ~w12726 & ~w12728;
assign w12730 = w12462 & ~w12470;
assign w12731 = ~w12459 & ~w12468;
assign w12732 = w12455 & ~w12731;
assign w12733 = ~w12717 & ~w12732;
assign w12734 = ~w12467 & ~w12733;
assign w12735 = ~w12730 & w12734;
assign w12736 = ~w12397 & w12726;
assign w12737 = ~w12735 & w12736;
assign w12738 = ~w12728 & w12737;
assign w12739 = ~w12397 & ~w12726;
assign w12740 = ~w12735 & w12739;
assign w12741 = w12728 & w12740;
assign w12742 = ~w12738 & ~w12741;
assign w12743 = ~w12729 & w12742;
assign w12744 = w12719 & ~w12725;
assign w12745 = w12713 & ~w12744;
assign w12746 = w12715 & ~w12745;
assign w12747 = w12742 & w12746;
assign w12748 = ~w12743 & ~w12747;
assign w12749 = ~w12724 & w12748;
assign w12750 = ~w12397 & ~w12735;
assign w12751 = w12726 & w12728;
assign w12752 = ~w12729 & ~w12751;
assign w12753 = ~w12750 & ~w12752;
assign w12754 = w12397 & w12735;
assign w12755 = ~w12400 & ~w12754;
assign w12756 = (~w12755 & w12753) | (~w12755 & w38029) | (w12753 & w38029);
assign w12757 = ~w12401 & w12475;
assign w12758 = w12397 & ~w12752;
assign w12759 = (w12757 & w12758) | (w12757 & w38030) | (w12758 & w38030);
assign w12760 = ~w12756 & ~w12759;
assign w12761 = ~w12749 & ~w12760;
assign w12762 = w12544 & w12616;
assign w12763 = (~w12619 & ~w12621) | (~w12619 & w38031) | (~w12621 & w38031);
assign w12764 = ~w12762 & ~w12763;
assign w12765 = ~w12544 & ~w12616;
assign w12766 = ~w11044 & ~w12591;
assign w12767 = ~pi0110 & ~w10769;
assign w12768 = pi0110 & w10769;
assign w12769 = ~w12767 & ~w12768;
assign w12770 = w10766 & ~w12769;
assign w12771 = ~w12766 & ~w12770;
assign w12772 = ~pi0113 & ~w12563;
assign w12773 = ~w12562 & w12772;
assign w12774 = ~pi0112 & w11305;
assign w12775 = ~w12773 & ~w12774;
assign w12776 = w11308 & ~w12775;
assign w12777 = w12573 & w12775;
assign w12778 = ~w12776 & ~w12777;
assign w12779 = w12771 & ~w12778;
assign w12780 = ~w12771 & w12778;
assign w12781 = ~w12779 & ~w12780;
assign w12782 = ~pi0107 & w11672;
assign w12783 = ~pi0105 & w11558;
assign w12784 = ~w12782 & ~w12783;
assign w12785 = (~w11561 & w12782) | (~w11561 & w38032) | (w12782 & w38032);
assign w12786 = w12609 & w12784;
assign w12787 = ~w12785 & ~w12786;
assign w12788 = w12781 & w12787;
assign w12789 = ~w12781 & ~w12787;
assign w12790 = ~w12788 & ~w12789;
assign w12791 = (~w12601 & ~w12603) | (~w12601 & w38033) | (~w12603 & w38033);
assign w12792 = w12790 & w12791;
assign w12793 = ~w12790 & ~w12791;
assign w12794 = ~w12792 & ~w12793;
assign w12795 = ~w12536 & w12540;
assign w12796 = ~w12535 & ~w12795;
assign w12797 = pi0078 & w11835;
assign w12798 = pi0108 & w11810;
assign w12799 = (w11813 & w12797) | (w11813 & w38034) | (w12797 & w38034);
assign w12800 = ~pi0108 & w11814;
assign w12801 = w11835 & w38035;
assign w12802 = ~w12800 & ~w12801;
assign w12803 = ~w12799 & w12802;
assign w12804 = ~w6330 & w10777;
assign w12805 = ~w3350 & w10775;
assign w12806 = ~w12804 & ~w12805;
assign w12807 = ~pi0079 & ~pi1424;
assign w12808 = ~w10818 & ~w12807;
assign w12809 = w12098 & ~w12808;
assign w12810 = ~w12806 & w12809;
assign w12811 = w12806 & ~w12809;
assign w12812 = ~w12810 & ~w12811;
assign w12813 = ~w12803 & w12812;
assign w12814 = w12803 & ~w12812;
assign w12815 = ~w12813 & ~w12814;
assign w12816 = w12796 & ~w12815;
assign w12817 = ~w12796 & w12815;
assign w12818 = ~w12816 & ~w12817;
assign w12819 = w12794 & ~w12818;
assign w12820 = ~w12794 & w12818;
assign w12821 = ~w12819 & ~w12820;
assign w12822 = ~w12765 & ~w12821;
assign w12823 = w12765 & w12821;
assign w12824 = ~w12822 & ~w12823;
assign w12825 = ~w12764 & w12824;
assign w12826 = ~w12665 & w12699;
assign w12827 = w12645 & ~w12657;
assign w12828 = ~w12656 & ~w12827;
assign w12829 = w12826 & w12828;
assign w12830 = w12699 & ~w12828;
assign w12831 = w12665 & w12830;
assign w12832 = ~w12829 & ~w12831;
assign w12833 = ~pi0081 & ~w10782;
assign w12834 = pi0081 & w10782;
assign w12835 = ~w12833 & ~w12834;
assign w12836 = w10809 & ~w12835;
assign w12837 = w10787 & ~w12674;
assign w12838 = ~w12836 & ~w12837;
assign w12839 = w10835 & w12100;
assign w12840 = ~w12683 & ~w12839;
assign w12841 = w12682 & ~w12840;
assign w12842 = w12649 & w12841;
assign w12843 = w12838 & w12842;
assign w12844 = ~w12649 & ~w12841;
assign w12845 = ~w12838 & w12844;
assign w12846 = w12838 & ~w12844;
assign w12847 = ~w12842 & ~w12846;
assign w12848 = (~w12843 & ~w12847) | (~w12843 & w38036) | (~w12847 & w38036);
assign w12849 = w12649 & ~w12691;
assign w12850 = ~w12690 & ~w12849;
assign w12851 = w12848 & ~w12850;
assign w12852 = ~w12848 & w12850;
assign w12853 = ~w12851 & ~w12852;
assign w12854 = w12832 & w12853;
assign w12855 = ~w12832 & ~w12853;
assign w12856 = ~w12854 & ~w12855;
assign w12857 = w12828 & w12848;
assign w12858 = (w12857 & w12826) | (w12857 & w38037) | (w12826 & w38037);
assign w12859 = ~w12656 & ~w12850;
assign w12860 = ~w12848 & w12859;
assign w12861 = w12699 & w38038;
assign w12862 = (~w12860 & ~w12861) | (~w12860 & w38039) | (~w12861 & w38039);
assign w12863 = ~w12858 & w12862;
assign w12864 = w12856 & w12863;
assign w12865 = ~w12825 & ~w12864;
assign w12866 = w12851 & ~w12861;
assign w12867 = w12852 & w12861;
assign w12868 = ~w12866 & ~w12867;
assign w12869 = pi1469 & ~pi1640;
assign w12870 = ~w10785 & ~w12869;
assign w12871 = w10784 & ~w12870;
assign w12872 = ~pi1469 & ~pi1640;
assign w12873 = ~w10783 & ~w12872;
assign w12874 = w10786 & ~w12873;
assign w12875 = ~w12871 & ~w12874;
assign w12876 = (~w12101 & ~w10782) | (~w12101 & w38040) | (~w10782 & w38040);
assign w12877 = pi1469 & w10785;
assign w12878 = ~pi1469 & w10783;
assign w12879 = ~w12877 & ~w12878;
assign w12880 = ~w12876 & w12879;
assign w12881 = ~w12833 & ~w12880;
assign w12882 = w12875 & ~w12881;
assign w12883 = (w12882 & w12846) | (w12882 & w38041) | (w12846 & w38041);
assign w12884 = ~w12846 & w38042;
assign w12885 = ~w12883 & ~w12884;
assign w12886 = w12868 & w12885;
assign w12887 = ~w12868 & ~w12885;
assign w12888 = ~w12886 & ~w12887;
assign w12889 = ~w12793 & ~w12817;
assign w12890 = w12821 & w12889;
assign w12891 = ~w12822 & ~w12890;
assign w12892 = ~w3350 & w10777;
assign w12893 = ~w3075 & w10775;
assign w12894 = ~w12892 & ~w12893;
assign w12895 = ~pi0078 & ~pi1424;
assign w12896 = ~w10795 & ~w12895;
assign w12897 = w12098 & ~w12896;
assign w12898 = w12894 & ~w12897;
assign w12899 = ~w12894 & w12897;
assign w12900 = ~w12898 & ~w12899;
assign w12901 = ~pi0108 & w11835;
assign w12902 = ~pi0107 & w11810;
assign w12903 = ~w12901 & ~w12902;
assign w12904 = (~w11813 & w12901) | (~w11813 & w38043) | (w12901 & w38043);
assign w12905 = w12533 & w12903;
assign w12906 = ~w12904 & ~w12905;
assign w12907 = w12900 & w12906;
assign w12908 = ~w12900 & ~w12906;
assign w12909 = ~w12907 & ~w12908;
assign w12910 = (~w12810 & w12803) | (~w12810 & w38044) | (w12803 & w38044);
assign w12911 = w12909 & w12910;
assign w12912 = ~w12909 & ~w12910;
assign w12913 = ~w12911 & ~w12912;
assign w12914 = ~w12792 & ~w12816;
assign w12915 = ~w11044 & ~w12769;
assign w12916 = ~pi0109 & ~w10769;
assign w12917 = pi0109 & w10769;
assign w12918 = ~w12916 & ~w12917;
assign w12919 = w10766 & ~w12918;
assign w12920 = ~w12915 & ~w12919;
assign w12921 = pi0113 & ~w11561;
assign w12922 = ~pi0113 & w11561;
assign w12923 = w11558 & ~w12922;
assign w12924 = ~w12921 & w12923;
assign w12925 = ~pi0105 & w11561;
assign w12926 = pi0105 & ~w11561;
assign w12927 = w11672 & ~w12926;
assign w12928 = ~w12925 & w12927;
assign w12929 = ~w12924 & ~w12928;
assign w12930 = ~pi0112 & ~w12563;
assign w12931 = ~w12562 & w12930;
assign w12932 = ~pi0111 & w11305;
assign w12933 = ~w12931 & ~w12932;
assign w12934 = w11308 & ~w12933;
assign w12935 = w12573 & w12933;
assign w12936 = ~w12934 & ~w12935;
assign w12937 = w12929 & ~w12936;
assign w12938 = ~w12929 & w12936;
assign w12939 = ~w12937 & ~w12938;
assign w12940 = w12920 & w12939;
assign w12941 = ~w12920 & ~w12939;
assign w12942 = ~w12940 & ~w12941;
assign w12943 = (~w12779 & ~w12781) | (~w12779 & w38045) | (~w12781 & w38045);
assign w12944 = w12942 & ~w12943;
assign w12945 = ~w12942 & w12943;
assign w12946 = ~w12944 & ~w12945;
assign w12947 = w12914 & ~w12946;
assign w12948 = ~w12914 & w12946;
assign w12949 = ~w12947 & ~w12948;
assign w12950 = w12913 & ~w12949;
assign w12951 = ~w12913 & w12949;
assign w12952 = ~w12950 & ~w12951;
assign w12953 = ~w12891 & ~w12952;
assign w12954 = w12891 & w12952;
assign w12955 = ~w12953 & ~w12954;
assign w12956 = ~w12888 & w12955;
assign w12957 = w12888 & ~w12955;
assign w12958 = ~w12956 & ~w12957;
assign w12959 = ~w12865 & w12958;
assign w12960 = w12865 & ~w12958;
assign w12961 = ~w12959 & ~w12960;
assign w12962 = ~w12666 & ~w12826;
assign w12963 = ~w12700 & ~w12962;
assign w12964 = ~w12637 & w38046;
assign w12965 = ~w12825 & w12964;
assign w12966 = (~w12856 & w12637) | (~w12856 & w38047) | (w12637 & w38047);
assign w12967 = w12764 & ~w12824;
assign w12968 = w12864 & ~w12967;
assign w12969 = ~w12825 & ~w12967;
assign w12970 = ~w12968 & ~w12969;
assign w12971 = ~w12966 & w12970;
assign w12972 = ~w12965 & ~w12971;
assign w12973 = w12961 & w12972;
assign w12974 = w12637 & w12963;
assign w12975 = ~w12704 & ~w12974;
assign w12976 = ~w12722 & w12975;
assign w12977 = ~w12964 & ~w12966;
assign w12978 = w12969 & ~w12977;
assign w12979 = ~w12969 & w12977;
assign w12980 = ~w12978 & ~w12979;
assign w12981 = ~w12976 & ~w12980;
assign w12982 = ~w12973 & ~w12981;
assign w12983 = w12724 & ~w12748;
assign w12984 = (~w12882 & w12846) | (~w12882 & w38048) | (w12846 & w38048);
assign w12985 = (~w12882 & ~w12844) | (~w12882 & w38049) | (~w12844 & w38049);
assign w12986 = ~w12843 & ~w12985;
assign w12987 = ~w12849 & w38050;
assign w12988 = ~w12986 & w12987;
assign w12989 = ~w12984 & ~w12988;
assign w12990 = (w12989 & w12861) | (w12989 & w38051) | (w12861 & w38051);
assign w12991 = (w12990 & ~w12868) | (w12990 & w38052) | (~w12868 & w38052);
assign w12992 = w12953 & w12991;
assign w12993 = ~w12956 & ~w12992;
assign w12994 = ~w12959 & w12993;
assign w12995 = w10782 & w12100;
assign w12996 = ~w10782 & ~w12100;
assign w12997 = ~w12995 & ~w12996;
assign w12998 = w12875 & ~w12997;
assign w12999 = (w12998 & w12988) | (w12998 & w38053) | (w12988 & w38053);
assign w13000 = ~w12988 & w38054;
assign w13001 = ~w12999 & ~w13000;
assign w13002 = ~w12953 & ~w12991;
assign w13003 = ~w12911 & w12947;
assign w13004 = w12942 & w38055;
assign w13005 = ~w12913 & ~w13004;
assign w13006 = ~w12948 & w13005;
assign w13007 = ~w13003 & ~w13006;
assign w13008 = ~w12911 & ~w12944;
assign w13009 = ~w11044 & ~w12918;
assign w13010 = ~pi0081 & w10769;
assign w13011 = pi0081 & ~w10769;
assign w13012 = w10766 & ~w13011;
assign w13013 = ~w13010 & w13012;
assign w13014 = ~w13009 & ~w13013;
assign w13015 = ~pi0111 & ~w12563;
assign w13016 = ~w12562 & w13015;
assign w13017 = ~pi0110 & w11305;
assign w13018 = ~w13016 & ~w13017;
assign w13019 = w11308 & ~w13018;
assign w13020 = w12573 & w13018;
assign w13021 = ~w13019 & ~w13020;
assign w13022 = w13014 & ~w13021;
assign w13023 = ~w13014 & w13021;
assign w13024 = ~w13022 & ~w13023;
assign w13025 = ~pi0113 & w11672;
assign w13026 = ~pi0112 & w11558;
assign w13027 = ~w13025 & ~w13026;
assign w13028 = (~w11561 & w13025) | (~w11561 & w38056) | (w13025 & w38056);
assign w13029 = w12609 & w13027;
assign w13030 = ~w13028 & ~w13029;
assign w13031 = w13024 & w13030;
assign w13032 = ~w13024 & ~w13030;
assign w13033 = ~w13031 & ~w13032;
assign w13034 = (~w12937 & ~w12939) | (~w12937 & w38057) | (~w12939 & w38057);
assign w13035 = w13033 & ~w13034;
assign w13036 = ~w13033 & w13034;
assign w13037 = ~w13035 & ~w13036;
assign w13038 = ~w13008 & w13037;
assign w13039 = w13008 & ~w13037;
assign w13040 = ~w13038 & ~w13039;
assign w13041 = ~w6060 & w10775;
assign w13042 = ~w3075 & w10777;
assign w13043 = ~w13041 & ~w13042;
assign w13044 = ~pi0108 & ~pi1424;
assign w13045 = ~w10789 & ~w13044;
assign w13046 = w12098 & ~w13045;
assign w13047 = ~w13043 & w13046;
assign w13048 = w13043 & ~w13046;
assign w13049 = ~w13047 & ~w13048;
assign w13050 = ~pi0107 & w11835;
assign w13051 = ~pi0105 & w11810;
assign w13052 = ~w13050 & ~w13051;
assign w13053 = (~w11813 & w13050) | (~w11813 & w38058) | (w13050 & w38058);
assign w13054 = w12533 & w13052;
assign w13055 = ~w13053 & ~w13054;
assign w13056 = w13049 & ~w13055;
assign w13057 = ~w13049 & w13055;
assign w13058 = ~w13056 & ~w13057;
assign w13059 = (~w12898 & ~w12906) | (~w12898 & w38059) | (~w12906 & w38059);
assign w13060 = ~w13058 & ~w13059;
assign w13061 = w13058 & w13059;
assign w13062 = ~w13060 & ~w13061;
assign w13063 = w13040 & w13062;
assign w13064 = ~w13040 & ~w13062;
assign w13065 = ~w13063 & ~w13064;
assign w13066 = w13007 & w13065;
assign w13067 = ~w13007 & ~w13065;
assign w13068 = ~w13066 & ~w13067;
assign w13069 = ~w13002 & w13068;
assign w13070 = w13002 & ~w13068;
assign w13071 = ~w13069 & ~w13070;
assign w13072 = w13001 & w13071;
assign w13073 = ~w13001 & ~w13071;
assign w13074 = ~w13072 & ~w13073;
assign w13075 = ~w12994 & w13074;
assign w13076 = ~w13001 & ~w13069;
assign w13077 = ~w13070 & ~w13076;
assign w13078 = ~w12944 & w38060;
assign w13079 = w13033 & w38061;
assign w13080 = (~w13078 & w13038) | (~w13078 & w38062) | (w13038 & w38062);
assign w13081 = ~w13063 & ~w13080;
assign w13082 = ~w13035 & ~w13060;
assign w13083 = w10769 & w12100;
assign w13084 = ~w10769 & ~w12100;
assign w13085 = ~w13083 & ~w13084;
assign w13086 = ~pi0098 & w10764;
assign w13087 = pi0098 & w10765;
assign w13088 = ~w13086 & ~w13087;
assign w13089 = pi0096 & pi1425;
assign w13090 = ~w10764 & ~w13089;
assign w13091 = ~pi0095 & pi1425;
assign w13092 = pi0081 & ~w13091;
assign w13093 = ~w13090 & w13092;
assign w13094 = w13088 & ~w13093;
assign w13095 = ~w13085 & w13094;
assign w13096 = ~w11044 & w12101;
assign w13097 = ~w13093 & w13096;
assign w13098 = ~w13095 & ~w13097;
assign w13099 = pi0110 & w12573;
assign w13100 = ~pi0110 & w11308;
assign w13101 = ~w11404 & ~w13100;
assign w13102 = ~w13099 & w13101;
assign w13103 = ~pi0109 & w11308;
assign w13104 = pi0109 & ~w11308;
assign w13105 = w11305 & ~w13104;
assign w13106 = ~w13103 & w13105;
assign w13107 = ~w13102 & ~w13106;
assign w13108 = w13098 & w13107;
assign w13109 = ~w13098 & ~w13107;
assign w13110 = ~w13108 & ~w13109;
assign w13111 = ~pi0111 & ~w11561;
assign w13112 = pi0111 & w11561;
assign w13113 = ~w13111 & ~w13112;
assign w13114 = w11558 & ~w13113;
assign w13115 = ~pi0112 & w11561;
assign w13116 = pi0112 & ~w11561;
assign w13117 = w11672 & ~w13116;
assign w13118 = ~w13115 & w13117;
assign w13119 = ~w13114 & ~w13118;
assign w13120 = w13110 & w13119;
assign w13121 = ~w13110 & ~w13119;
assign w13122 = ~w13120 & ~w13121;
assign w13123 = (~w13022 & ~w13024) | (~w13022 & w38063) | (~w13024 & w38063);
assign w13124 = w13122 & ~w13123;
assign w13125 = ~w13122 & w13123;
assign w13126 = ~w13124 & ~w13125;
assign w13127 = (~w13047 & w13055) | (~w13047 & w38064) | (w13055 & w38064);
assign w13128 = ~w6060 & w10777;
assign w13129 = ~w4023 & w10775;
assign w13130 = ~w13128 & ~w13129;
assign w13131 = pi0113 & ~w11813;
assign w13132 = ~pi0113 & w11813;
assign w13133 = w11810 & ~w13132;
assign w13134 = ~w13131 & w13133;
assign w13135 = ~pi0105 & w11813;
assign w13136 = pi0105 & ~w11813;
assign w13137 = w11835 & ~w13136;
assign w13138 = ~w13135 & w13137;
assign w13139 = ~w13134 & ~w13138;
assign w13140 = ~w13130 & w13139;
assign w13141 = w13130 & ~w13139;
assign w13142 = ~w13140 & ~w13141;
assign w13143 = ~pi0107 & ~pi1424;
assign w13144 = ~w10952 & ~w13143;
assign w13145 = w12098 & ~w13144;
assign w13146 = ~w13142 & ~w13145;
assign w13147 = w13142 & w13145;
assign w13148 = ~w13146 & ~w13147;
assign w13149 = w13127 & w13148;
assign w13150 = ~w13127 & ~w13148;
assign w13151 = ~w13149 & ~w13150;
assign w13152 = ~w13126 & ~w13151;
assign w13153 = w13126 & w13151;
assign w13154 = ~w13152 & ~w13153;
assign w13155 = w13082 & ~w13154;
assign w13156 = ~w13082 & w13154;
assign w13157 = ~w13155 & ~w13156;
assign w13158 = w13081 & ~w13157;
assign w13159 = ~w13081 & w13157;
assign w13160 = ~w13158 & ~w13159;
assign w13161 = w13065 & w38065;
assign w13162 = (w12999 & ~w13065) | (w12999 & w38066) | (~w13065 & w38066);
assign w13163 = ~w13161 & ~w13162;
assign w13164 = w13160 & w13163;
assign w13165 = ~w13160 & ~w13163;
assign w13166 = ~w13164 & ~w13165;
assign w13167 = (~w12999 & ~w13065) | (~w12999 & w38067) | (~w13065 & w38067);
assign w13168 = ~w12110 & ~w12998;
assign w13169 = w12844 & w13168;
assign w13170 = ~w12844 & w38068;
assign w13171 = ~w12881 & w38069;
assign w13172 = ~w12842 & w13171;
assign w13173 = ~w13170 & w13172;
assign w13174 = ~w13169 & ~w13173;
assign w13175 = ~w13167 & w13174;
assign w13176 = ~w13160 & w13175;
assign w13177 = w13160 & ~w13175;
assign w13178 = ~w13176 & ~w13177;
assign w13179 = (w13178 & w13077) | (w13178 & w38070) | (w13077 & w38070);
assign w13180 = ~w13075 & ~w13179;
assign w13181 = ~w12983 & w13180;
assign w13182 = w12982 & w13181;
assign w13183 = w13181 & w38071;
assign w13184 = w12481 & ~w12494;
assign w13185 = ~w12495 & ~w13184;
assign w13186 = ~w12342 & ~w12478;
assign w13187 = ~w12499 & w12501;
assign w13188 = ~w13186 & ~w13187;
assign w13189 = w13185 & w13188;
assign w13190 = ~w12479 & ~w12495;
assign w13191 = ~w13186 & ~w13190;
assign w13192 = ~w13189 & ~w13191;
assign w13193 = ~w5590 & w10775;
assign w13194 = ~w4977 & w10777;
assign w13195 = ~w13193 & ~w13194;
assign w13196 = ~pi0113 & pi1424;
assign w13197 = ~w11328 & w12098;
assign w13198 = ~w13196 & w13197;
assign w13199 = ~w13195 & w13198;
assign w13200 = w13195 & ~w13198;
assign w13201 = ~pi0112 & w11835;
assign w13202 = ~pi0111 & w11810;
assign w13203 = ~w13201 & ~w13202;
assign w13204 = (~w11813 & w13201) | (~w11813 & w38072) | (w13201 & w38072);
assign w13205 = w12533 & w13203;
assign w13206 = ~w13204 & ~w13205;
assign w13207 = (~w13200 & w13205) | (~w13200 & w38073) | (w13205 & w38073);
assign w13208 = ~w13199 & ~w13207;
assign w13209 = ~w5590 & w10777;
assign w13210 = ~w1161 & w10775;
assign w13211 = ~w13209 & ~w13210;
assign w13212 = ~pi0112 & ~pi1424;
assign w13213 = ~w11456 & ~w13212;
assign w13214 = w12098 & ~w13213;
assign w13215 = w13211 & ~w13214;
assign w13216 = ~w13211 & w13214;
assign w13217 = ~w13215 & ~w13216;
assign w13218 = ~pi0111 & w11835;
assign w13219 = ~pi0110 & w11810;
assign w13220 = ~w13218 & ~w13219;
assign w13221 = (~w11813 & w13218) | (~w11813 & w38074) | (w13218 & w38074);
assign w13222 = w12533 & w13220;
assign w13223 = ~w13221 & ~w13222;
assign w13224 = w13217 & ~w13223;
assign w13225 = ~w13217 & w13223;
assign w13226 = ~w13224 & ~w13225;
assign w13227 = w13208 & ~w13226;
assign w13228 = ~pi0102 & w11303;
assign w13229 = pi0102 & w11304;
assign w13230 = ~w13228 & ~w13229;
assign w13231 = ~w11308 & w12100;
assign w13232 = w11308 & ~w12100;
assign w13233 = ~w13231 & ~w13232;
assign w13234 = w13230 & w13233;
assign w13235 = ~pi0109 & ~w11561;
assign w13236 = pi0109 & w11561;
assign w13237 = ~w13235 & ~w13236;
assign w13238 = w11672 & ~w13237;
assign w13239 = ~pi0081 & w11561;
assign w13240 = pi0081 & ~w11561;
assign w13241 = w11558 & ~w13240;
assign w13242 = ~w13239 & w13241;
assign w13243 = ~w13238 & ~w13242;
assign w13244 = ~w13234 & w13243;
assign w13245 = w13234 & ~w13243;
assign w13246 = ~w13244 & ~w13245;
assign w13247 = ~w13085 & w13088;
assign w13248 = pi0103 & pi1470;
assign w13249 = ~w11303 & ~w13248;
assign w13250 = ~pi0098 & pi1470;
assign w13251 = pi0081 & ~w13250;
assign w13252 = ~w13249 & w13251;
assign w13253 = w13230 & ~w13252;
assign w13254 = w13233 & w13253;
assign w13255 = ~w11404 & w12101;
assign w13256 = ~w13252 & w13255;
assign w13257 = ~w13254 & ~w13256;
assign w13258 = w11558 & ~w13237;
assign w13259 = ~pi0110 & ~w11561;
assign w13260 = pi0110 & w11561;
assign w13261 = ~w13259 & ~w13260;
assign w13262 = w11672 & ~w13261;
assign w13263 = ~w13258 & ~w13262;
assign w13264 = w13257 & w13263;
assign w13265 = w13247 & ~w13264;
assign w13266 = ~w13257 & ~w13263;
assign w13267 = ~w13247 & ~w13266;
assign w13268 = ~w13265 & ~w13267;
assign w13269 = w13246 & ~w13268;
assign w13270 = ~w13246 & w13268;
assign w13271 = ~w13269 & ~w13270;
assign w13272 = (~w13266 & w13246) | (~w13266 & w13267) | (w13246 & w13267);
assign w13273 = (~w13227 & ~w13271) | (~w13227 & w38075) | (~w13271 & w38075);
assign w13274 = ~pi0109 & ~w11813;
assign w13275 = pi0109 & w11813;
assign w13276 = ~w13274 & ~w13275;
assign w13277 = w11810 & ~w13276;
assign w13278 = ~pi0110 & w11813;
assign w13279 = pi0110 & ~w11813;
assign w13280 = w11835 & ~w13279;
assign w13281 = ~w13278 & w13280;
assign w13282 = ~w13277 & ~w13281;
assign w13283 = ~w1509 & w10775;
assign w13284 = ~w1161 & w10777;
assign w13285 = ~w13283 & ~w13284;
assign w13286 = ~pi0111 & ~pi1424;
assign w13287 = ~w11569 & ~w13286;
assign w13288 = w12098 & ~w13287;
assign w13289 = w13285 & ~w13288;
assign w13290 = ~w13285 & w13288;
assign w13291 = ~w13289 & ~w13290;
assign w13292 = ~w13282 & w13291;
assign w13293 = w13282 & ~w13291;
assign w13294 = ~w13292 & ~w13293;
assign w13295 = (~w13215 & w13222) | (~w13215 & w38076) | (w13222 & w38076);
assign w13296 = ~w13216 & ~w13295;
assign w13297 = ~w13294 & w13296;
assign w13298 = w13294 & ~w13296;
assign w13299 = ~w13297 & ~w13298;
assign w13300 = ~w13234 & ~w13247;
assign w13301 = w13243 & ~w13300;
assign w13302 = pi1418 & ~w11556;
assign w13303 = (pi0081 & w11557) | (pi0081 & w38077) | (w11557 & w38077);
assign w13304 = ~w13302 & w13303;
assign w13305 = ~w11561 & w12100;
assign w13306 = ~w13239 & ~w13305;
assign w13307 = ~pi1418 & ~pi1640;
assign w13308 = ~w11557 & ~w13307;
assign w13309 = w11670 & ~w13308;
assign w13310 = pi1418 & ~pi1640;
assign w13311 = ~w11556 & ~w13310;
assign w13312 = w11671 & ~w13311;
assign w13313 = ~w13309 & ~w13312;
assign w13314 = w13306 & w13313;
assign w13315 = ~w13304 & w13314;
assign w13316 = w13234 & w13247;
assign w13317 = w13315 & ~w13316;
assign w13318 = ~w13301 & w13317;
assign w13319 = (~w13315 & w13301) | (~w13315 & w38078) | (w13301 & w38078);
assign w13320 = ~w13318 & ~w13319;
assign w13321 = ~w13299 & w13320;
assign w13322 = w13299 & ~w13320;
assign w13323 = ~w13321 & ~w13322;
assign w13324 = ~w13273 & w13323;
assign w13325 = w13273 & ~w13323;
assign w13326 = ~w13324 & ~w13325;
assign w13327 = w13271 & w38079;
assign w13328 = ~w13199 & ~w13200;
assign w13329 = ~w13206 & w13328;
assign w13330 = w13206 & ~w13328;
assign w13331 = ~w13329 & ~w13330;
assign w13332 = ~w4977 & w10775;
assign w13333 = ~w4023 & w10777;
assign w13334 = ~w13332 & ~w13333;
assign w13335 = ~pi0112 & w11810;
assign w13336 = ~pi0077 & pi0099;
assign w13337 = ~w11809 & ~w13336;
assign w13338 = ~pi0077 & ~pi0100;
assign w13339 = ~pi0113 & ~w13338;
assign w13340 = ~w13337 & w13339;
assign w13341 = ~w13335 & ~w13340;
assign w13342 = ~w11813 & ~w13341;
assign w13343 = w12533 & w13341;
assign w13344 = ~w13342 & ~w13343;
assign w13345 = ~w13334 & ~w13344;
assign w13346 = w13334 & w13344;
assign w13347 = ~pi0105 & ~pi1424;
assign w13348 = ~w11046 & ~w13347;
assign w13349 = w12098 & ~w13348;
assign w13350 = (w13349 & ~w13344) | (w13349 & w38080) | (~w13344 & w38080);
assign w13351 = ~w13345 & ~w13350;
assign w13352 = ~w13331 & w13351;
assign w13353 = ~w13264 & ~w13266;
assign w13354 = w11672 & ~w13113;
assign w13355 = w11558 & ~w13261;
assign w13356 = ~w13354 & ~w13355;
assign w13357 = ~pi0081 & w11305;
assign w13358 = ~pi0109 & ~w12563;
assign w13359 = ~w12562 & w13358;
assign w13360 = ~w13357 & ~w13359;
assign w13361 = w11308 & ~w13360;
assign w13362 = w12573 & w13360;
assign w13363 = ~w13361 & ~w13362;
assign w13364 = ~w13356 & w13363;
assign w13365 = ~w13247 & ~w13364;
assign w13366 = ~w13353 & ~w13365;
assign w13367 = w13356 & ~w13363;
assign w13368 = w13247 & w13367;
assign w13369 = w13353 & ~w13368;
assign w13370 = ~w13366 & ~w13369;
assign w13371 = ~w13352 & ~w13370;
assign w13372 = ~w13271 & ~w13371;
assign w13373 = ~w13208 & w13226;
assign w13374 = ~w13227 & ~w13373;
assign w13375 = ~w13372 & ~w13374;
assign w13376 = ~w13327 & w13375;
assign w13377 = w13271 & w13371;
assign w13378 = ~w13227 & w13377;
assign w13379 = ~w13376 & ~w13378;
assign w13380 = w13326 & w13379;
assign w13381 = w13379 & w38081;
assign w13382 = ~w13300 & ~w13317;
assign w13383 = ~w13318 & ~w13382;
assign w13384 = w13297 & w13383;
assign w13385 = ~w13322 & ~w13384;
assign w13386 = ~w13324 & w13385;
assign w13387 = (~w13289 & ~w13282) | (~w13289 & w38082) | (~w13282 & w38082);
assign w13388 = w11835 & ~w13276;
assign w13389 = ~pi0081 & w11813;
assign w13390 = pi0081 & ~w11813;
assign w13391 = w11810 & ~w13390;
assign w13392 = ~w13389 & w13391;
assign w13393 = ~w13388 & ~w13392;
assign w13394 = ~w7942 & w10775;
assign w13395 = ~w1509 & w10777;
assign w13396 = ~w13394 & ~w13395;
assign w13397 = ~pi0110 & ~pi1424;
assign w13398 = ~w11674 & ~w13397;
assign w13399 = w12098 & ~w13398;
assign w13400 = w13396 & ~w13399;
assign w13401 = ~w13396 & w13399;
assign w13402 = ~w13400 & ~w13401;
assign w13403 = ~w13393 & w13402;
assign w13404 = w13393 & ~w13402;
assign w13405 = ~w13403 & ~w13404;
assign w13406 = ~w13387 & ~w13405;
assign w13407 = w13387 & w13405;
assign w13408 = ~w13406 & ~w13407;
assign w13409 = w11561 & ~w12100;
assign w13410 = ~w13305 & ~w13409;
assign w13411 = ~w12608 & w13410;
assign w13412 = ~w13318 & w13411;
assign w13413 = w13318 & ~w13411;
assign w13414 = ~w13412 & ~w13413;
assign w13415 = ~w13297 & w13414;
assign w13416 = ~w13317 & w38083;
assign w13417 = (~w13411 & w13317) | (~w13411 & w13567) | (w13317 & w13567);
assign w13418 = ~w13416 & ~w13417;
assign w13419 = w13297 & ~w13418;
assign w13420 = (w13408 & w13415) | (w13408 & w38084) | (w13415 & w38084);
assign w13421 = ~w13415 & w38085;
assign w13422 = ~w13420 & ~w13421;
assign w13423 = w13386 & ~w13422;
assign w13424 = ~w13386 & w13422;
assign w13425 = ~w13423 & ~w13424;
assign w13426 = ~w13381 & ~w13425;
assign w13427 = ~w13326 & ~w13379;
assign w13428 = (~w13108 & ~w13110) | (~w13108 & w38086) | (~w13110 & w38086);
assign w13429 = ~w13364 & ~w13367;
assign w13430 = w13247 & ~w13429;
assign w13431 = ~w13247 & w13429;
assign w13432 = ~w13430 & ~w13431;
assign w13433 = ~w13428 & w13432;
assign w13434 = w13130 & w13139;
assign w13435 = (~w13434 & w13142) | (~w13434 & w38087) | (w13142 & w38087);
assign w13436 = ~w13345 & ~w13346;
assign w13437 = ~w13349 & w13436;
assign w13438 = w13349 & ~w13436;
assign w13439 = ~w13437 & ~w13438;
assign w13440 = ~w13435 & w13439;
assign w13441 = ~w13433 & ~w13440;
assign w13442 = w13331 & ~w13351;
assign w13443 = ~w13352 & ~w13442;
assign w13444 = ~w13247 & w13364;
assign w13445 = ~w13368 & ~w13444;
assign w13446 = w13353 & ~w13445;
assign w13447 = ~w13353 & w13445;
assign w13448 = ~w13446 & ~w13447;
assign w13449 = ~w13443 & ~w13448;
assign w13450 = ~w13441 & ~w13449;
assign w13451 = w13443 & w13448;
assign w13452 = w13352 & w13370;
assign w13453 = ~w13451 & ~w13452;
assign w13454 = ~w13450 & w13453;
assign w13455 = ~w13372 & ~w13377;
assign w13456 = w13374 & ~w13455;
assign w13457 = ~w13374 & w13455;
assign w13458 = ~w13456 & ~w13457;
assign w13459 = ~w13454 & ~w13458;
assign w13460 = ~w13458 & w38088;
assign w13461 = w13427 & ~w13460;
assign w13462 = w13426 & ~w13461;
assign w13463 = ~w13380 & ~w13427;
assign w13464 = w13460 & ~w13463;
assign w13465 = w13425 & ~w13427;
assign w13466 = w13464 & w13465;
assign w13467 = ~w13462 & ~w13466;
assign w13468 = w13428 & ~w13432;
assign w13469 = ~w13433 & ~w13468;
assign w13470 = ~w13124 & ~w13149;
assign w13471 = w13435 & ~w13439;
assign w13472 = ~w13440 & ~w13471;
assign w13473 = w13470 & ~w13472;
assign w13474 = w13469 & ~w13473;
assign w13475 = ~w13470 & w13472;
assign w13476 = w13433 & w13440;
assign w13477 = ~w13475 & ~w13476;
assign w13478 = ~w13474 & w13477;
assign w13479 = ~w13449 & ~w13451;
assign w13480 = w13441 & ~w13479;
assign w13481 = ~w13441 & w13479;
assign w13482 = ~w13480 & ~w13481;
assign w13483 = ~w13169 & w13482;
assign w13484 = ~w13478 & w13483;
assign w13485 = w13459 & w13484;
assign w13486 = w13463 & ~w13485;
assign w13487 = w13454 & w13458;
assign w13488 = ~w13484 & w13487;
assign w13489 = ~w13464 & ~w13488;
assign w13490 = ~w13486 & w13489;
assign w13491 = w13467 & ~w13490;
assign w13492 = w13159 & ~w13169;
assign w13493 = ~w13158 & ~w13492;
assign w13494 = ~w13175 & ~w13493;
assign w13495 = ~w13082 & ~w13152;
assign w13496 = w13124 & w13149;
assign w13497 = ~w13153 & ~w13496;
assign w13498 = ~w13495 & w13497;
assign w13499 = ~w13473 & ~w13475;
assign w13500 = w13469 & ~w13499;
assign w13501 = ~w13469 & w13499;
assign w13502 = ~w13500 & ~w13501;
assign w13503 = ~w13498 & ~w13502;
assign w13504 = w13498 & w13502;
assign w13505 = ~w13503 & ~w13504;
assign w13506 = ~w13492 & w13505;
assign w13507 = w13492 & ~w13505;
assign w13508 = ~w13506 & ~w13507;
assign w13509 = ~w13494 & w13508;
assign w13510 = ~w13478 & ~w13482;
assign w13511 = w13478 & w13482;
assign w13512 = ~w13510 & ~w13511;
assign w13513 = w13503 & w13512;
assign w13514 = ~w13503 & ~w13512;
assign w13515 = ~w13513 & ~w13514;
assign w13516 = w13492 & ~w13515;
assign w13517 = ~w13504 & w13512;
assign w13518 = w13504 & ~w13512;
assign w13519 = ~w13492 & ~w13518;
assign w13520 = ~w13517 & w13519;
assign w13521 = ~w13516 & ~w13520;
assign w13522 = w13509 & ~w13521;
assign w13523 = ~w13169 & ~w13498;
assign w13524 = ~w13502 & w13523;
assign w13525 = (~w13510 & w13524) | (~w13510 & w38089) | (w13524 & w38089);
assign w13526 = ~w13459 & ~w13487;
assign w13527 = ~w13478 & w13526;
assign w13528 = w13478 & ~w13526;
assign w13529 = ~w13527 & ~w13528;
assign w13530 = w13525 & ~w13529;
assign w13531 = ~w13525 & w13529;
assign w13532 = ~w13530 & ~w13531;
assign w13533 = ~w13502 & w38090;
assign w13534 = ~w13515 & ~w13533;
assign w13535 = w13517 & ~w13524;
assign w13536 = ~w13492 & ~w13535;
assign w13537 = ~w13534 & ~w13536;
assign w13538 = w13532 & ~w13537;
assign w13539 = ~w13522 & w13538;
assign w13540 = w13491 & w13539;
assign w13541 = ~pi1471 & ~pi1640;
assign w13542 = ~w11809 & ~w13541;
assign w13543 = (~w11808 & ~w13542) | (~w11808 & w38091) | (~w13542 & w38091);
assign w13544 = pi0077 & ~w13543;
assign w13545 = pi0081 & ~w12532;
assign w13546 = ~w11813 & w12100;
assign w13547 = w11833 & ~w13542;
assign w13548 = ~w13389 & ~w13547;
assign w13549 = ~w13546 & w13548;
assign w13550 = w13549 & w38092;
assign w13551 = ~w8157 & w10775;
assign w13552 = ~w7942 & w10777;
assign w13553 = ~w13551 & ~w13552;
assign w13554 = ~pi0109 & ~pi1424;
assign w13555 = ~w11815 & ~w13554;
assign w13556 = w12098 & ~w13555;
assign w13557 = ~w13553 & w13556;
assign w13558 = w13553 & ~w13556;
assign w13559 = ~w13557 & ~w13558;
assign w13560 = ~w13550 & w13559;
assign w13561 = w13550 & ~w13559;
assign w13562 = ~w13560 & ~w13561;
assign w13563 = (~w13400 & ~w13393) | (~w13400 & w38093) | (~w13393 & w38093);
assign w13564 = w13562 & ~w13563;
assign w13565 = w13316 & w13411;
assign w13566 = (w13565 & ~w13562) | (w13565 & w38094) | (~w13562 & w38094);
assign w13567 = w13300 & ~w13411;
assign w13568 = ~pi0081 & pi1424;
assign w13569 = pi0081 & ~pi1473;
assign w13570 = w12098 & ~w13569;
assign w13571 = ~w13568 & w13570;
assign w13572 = ~w11810 & ~w11835;
assign w13573 = w11813 & ~w12100;
assign w13574 = ~w13546 & ~w13573;
assign w13575 = ~w13572 & w13574;
assign w13576 = ~w8157 & w10777;
assign w13577 = ~w3627 & w10775;
assign w13578 = ~w13576 & ~w13577;
assign w13579 = ~w13575 & w13578;
assign w13580 = w13575 & ~w13578;
assign w13581 = ~w13579 & ~w13580;
assign w13582 = w13571 & w13581;
assign w13583 = ~w13571 & ~w13581;
assign w13584 = ~w13582 & ~w13583;
assign w13585 = (~w13558 & w13550) | (~w13558 & w38095) | (w13550 & w38095);
assign w13586 = w13584 & w13585;
assign w13587 = (w13567 & ~w13584) | (w13567 & w38096) | (~w13584 & w38096);
assign w13588 = ~w13565 & ~w13567;
assign w13589 = w13564 & w13588;
assign w13590 = ~w13584 & ~w13585;
assign w13591 = ~w13586 & ~w13590;
assign w13592 = ~w13591 & w38097;
assign w13593 = ~w13566 & ~w13592;
assign w13594 = ~w13584 & w38098;
assign w13595 = (w13565 & w13584) | (w13565 & w38099) | (w13584 & w38099);
assign w13596 = ~w13594 & ~w13595;
assign w13597 = (~w13580 & ~w13581) | (~w13580 & w38100) | (~w13581 & w38100);
assign w13598 = pi0868 & ~w3627;
assign w13599 = ~pi0868 & ~w4689;
assign w13600 = ~w13598 & ~w13599;
assign w13601 = w10774 & ~w13600;
assign w13602 = w13570 & w38101;
assign w13603 = w12098 & w12362;
assign w13604 = ~w13602 & ~w13603;
assign w13605 = w13575 & ~w13604;
assign w13606 = ~w13575 & w13604;
assign w13607 = ~w13605 & ~w13606;
assign w13608 = ~w13601 & w13607;
assign w13609 = w13601 & ~w13607;
assign w13610 = ~w13608 & ~w13609;
assign w13611 = w13597 & w13610;
assign w13612 = ~w13597 & ~w13610;
assign w13613 = ~w13611 & ~w13612;
assign w13614 = w13596 & ~w13613;
assign w13615 = ~w13596 & w13613;
assign w13616 = ~w13614 & ~w13615;
assign w13617 = w13593 & ~w13616;
assign w13618 = w13610 & w38102;
assign w13619 = ~w13595 & ~w13612;
assign w13620 = (~w13594 & ~w13619) | (~w13594 & w38103) | (~w13619 & w38103);
assign w13621 = ~w5695 & w10775;
assign w13622 = ~w4689 & w10777;
assign w13623 = ~w13621 & ~w13622;
assign w13624 = w13601 & ~w13605;
assign w13625 = (w13623 & w13624) | (w13623 & w38104) | (w13624 & w38104);
assign w13626 = ~w13624 & w38105;
assign w13627 = ~w13625 & ~w13626;
assign w13628 = w13565 & w13627;
assign w13629 = ~w13565 & ~w13627;
assign w13630 = ~w13628 & ~w13629;
assign w13631 = ~w13618 & w13630;
assign w13632 = w13618 & ~w13630;
assign w13633 = ~w13631 & ~w13632;
assign w13634 = w13620 & ~w13633;
assign w13635 = ~w13620 & w13633;
assign w13636 = ~w13634 & ~w13635;
assign w13637 = w13617 & w13636;
assign w13638 = ~w13169 & ~w13566;
assign w13639 = ~w13592 & w13638;
assign w13640 = ~w13616 & w13639;
assign w13641 = ~w13636 & ~w13640;
assign w13642 = ~w13637 & ~w13641;
assign w13643 = ~w13562 & w13563;
assign w13644 = ~w13564 & ~w13643;
assign w13645 = ~w13405 & w38106;
assign w13646 = w13416 & ~w13645;
assign w13647 = w13406 & w13588;
assign w13648 = ~w13646 & ~w13647;
assign w13649 = ~w13644 & w13648;
assign w13650 = (w13565 & w13405) | (w13565 & w38107) | (w13405 & w38107);
assign w13651 = (~w13650 & ~w13648) | (~w13650 & w38108) | (~w13648 & w38108);
assign w13652 = w13562 & w38109;
assign w13653 = ~w13651 & ~w13652;
assign w13654 = ~w13566 & ~w13589;
assign w13655 = w13591 & ~w13654;
assign w13656 = ~w13591 & w13654;
assign w13657 = ~w13655 & ~w13656;
assign w13658 = ~w13653 & ~w13657;
assign w13659 = ~w13169 & w13658;
assign w13660 = ~w13593 & w13616;
assign w13661 = (~w13660 & ~w13636) | (~w13660 & w13681) | (~w13636 & w13681);
assign w13662 = ~w13659 & ~w13661;
assign w13663 = ~w13642 & ~w13662;
assign w13664 = w13644 & ~w13648;
assign w13665 = ~w13649 & ~w13664;
assign w13666 = ~w13297 & ~w13412;
assign w13667 = ~w13408 & w13666;
assign w13668 = w13418 & ~w13667;
assign w13669 = ~w13297 & ~w13383;
assign w13670 = w13408 & ~w13669;
assign w13671 = ~w13416 & ~w13567;
assign w13672 = ~w13405 & w38110;
assign w13673 = ~w13671 & w13672;
assign w13674 = ~w13670 & ~w13673;
assign w13675 = ~w13668 & w13674;
assign w13676 = ~w13665 & ~w13675;
assign w13677 = ~w13169 & w13676;
assign w13678 = w13653 & w13657;
assign w13679 = ~w13659 & ~w13678;
assign w13680 = ~w13677 & ~w13679;
assign w13681 = ~w13617 & ~w13660;
assign w13682 = ~w13659 & ~w13681;
assign w13683 = w13659 & w13681;
assign w13684 = ~w13682 & ~w13683;
assign w13685 = w13680 & w13684;
assign w13686 = ~w13663 & w13685;
assign w13687 = w13642 & w13682;
assign w13688 = (w13623 & w13575) | (w13623 & w38111) | (w13575 & w38111);
assign w13689 = ~w13605 & ~w13688;
assign w13690 = (w13600 & w13575) | (w13600 & w38112) | (w13575 & w38112);
assign w13691 = ~w13623 & ~w13690;
assign w13692 = ~w13567 & ~w13691;
assign w13693 = w13689 & ~w13692;
assign w13694 = ~w5695 & w10777;
assign w13695 = ~w5119 & w10775;
assign w13696 = ~w13694 & ~w13695;
assign w13697 = (w13696 & ~w13316) | (w13696 & w38113) | (~w13316 & w38113);
assign w13698 = w13316 & w38114;
assign w13699 = ~w13697 & ~w13698;
assign w13700 = w13693 & w13699;
assign w13701 = ~w13693 & ~w13699;
assign w13702 = ~w13700 & ~w13701;
assign w13703 = (~w13567 & ~w13610) | (~w13567 & w38115) | (~w13610 & w38115);
assign w13704 = ~w13630 & w13703;
assign w13705 = w13565 & ~w13688;
assign w13706 = ~w13691 & w13705;
assign w13707 = ~w13588 & ~w13689;
assign w13708 = ~w13627 & w13707;
assign w13709 = ~w13706 & ~w13708;
assign w13710 = (~w13702 & w13704) | (~w13702 & w38116) | (w13704 & w38116);
assign w13711 = ~w13704 & w38117;
assign w13712 = ~w13710 & ~w13711;
assign w13713 = w13634 & ~w13640;
assign w13714 = w13635 & w13640;
assign w13715 = ~w13713 & ~w13714;
assign w13716 = w13712 & ~w13715;
assign w13717 = ~w13712 & w13715;
assign w13718 = ~w13716 & ~w13717;
assign w13719 = ~w13687 & w13718;
assign w13720 = ~w13686 & w13719;
assign w13721 = ~w13169 & w13422;
assign w13722 = ~w13386 & w13721;
assign w13723 = w13665 & w13675;
assign w13724 = ~w13676 & ~w13723;
assign w13725 = ~w13722 & ~w13724;
assign w13726 = ~w13423 & w13725;
assign w13727 = w13424 & w13724;
assign w13728 = ~w13725 & ~w13727;
assign w13729 = w13381 & ~w13728;
assign w13730 = ~w13726 & ~w13729;
assign w13731 = ~w13658 & ~w13678;
assign w13732 = ~w13722 & w13723;
assign w13733 = w13424 & w13677;
assign w13734 = ~w13732 & ~w13733;
assign w13735 = w13731 & ~w13734;
assign w13736 = ~w13731 & w13734;
assign w13737 = ~w13735 & ~w13736;
assign w13738 = w13730 & w13737;
assign w13739 = w13731 & w13732;
assign w13740 = w13677 & ~w13731;
assign w13741 = ~w13739 & ~w13740;
assign w13742 = ~w13738 & w13741;
assign w13743 = ~w13680 & ~w13684;
assign w13744 = ~w13663 & ~w13743;
assign w13745 = (w13744 & w13738) | (w13744 & w38118) | (w13738 & w38118);
assign w13746 = w13633 & w38119;
assign w13747 = ~w13634 & ~w13746;
assign w13748 = ~w13640 & ~w13747;
assign w13749 = ~w13718 & ~w13748;
assign w13750 = (~w13749 & w13745) | (~w13749 & w38120) | (w13745 & w38120);
assign w13751 = w13539 & w38121;
assign w13752 = ~w13192 & w13751;
assign w13753 = w13183 & w13752;
assign w13754 = ~w12505 & w13753;
assign w13755 = w13494 & ~w13508;
assign w13756 = ~w13521 & ~w13755;
assign w13757 = w13179 & w13756;
assign w13758 = w13540 & ~w13757;
assign w13759 = ~w13483 & ~w13526;
assign w13760 = w13529 & w38122;
assign w13761 = w13463 & w13487;
assign w13762 = ~w13464 & ~w13761;
assign w13763 = ~w13484 & ~w13762;
assign w13764 = ~w13760 & ~w13763;
assign w13765 = w13491 & ~w13764;
assign w13766 = w13426 & w13728;
assign w13767 = ~w13426 & ~w13460;
assign w13768 = ~w13465 & w13767;
assign w13769 = ~w13766 & ~w13768;
assign w13770 = w13737 & w13769;
assign w13771 = w13720 & w13770;
assign w13772 = ~w13765 & w13771;
assign w13773 = (w13772 & ~w13540) | (w13772 & w38123) | (~w13540 & w38123);
assign w13774 = ~w12961 & ~w12972;
assign w13775 = w12976 & w12980;
assign w13776 = ~w13774 & ~w13775;
assign w13777 = ~w12973 & ~w13075;
assign w13778 = ~w13776 & w13777;
assign w13779 = w12994 & ~w13074;
assign w13780 = ~w13077 & ~w13166;
assign w13781 = w13756 & ~w13780;
assign w13782 = ~w13779 & w13781;
assign w13783 = w13772 & w13782;
assign w13784 = ~w13778 & w13783;
assign w13785 = ~w13773 & ~w13784;
assign w13786 = ~w13784 & w38124;
assign w13787 = ~w12715 & w12745;
assign w13788 = (w13787 & ~w12742) | (w13787 & w38125) | (~w12742 & w38125);
assign w13789 = ~w12713 & w12719;
assign w13790 = (w13789 & w12735) | (w13789 & w38126) | (w12735 & w38126);
assign w13791 = (~w12712 & w12717) | (~w12712 & w38127) | (w12717 & w38127);
assign w13792 = w12725 & w13791;
assign w13793 = ~w12735 & w38128;
assign w13794 = ~w13790 & ~w13793;
assign w13795 = (w13794 & ~w12742) | (w13794 & w38129) | (~w12742 & w38129);
assign w13796 = ~w13788 & w13795;
assign w13797 = ~w12705 & ~w13796;
assign w13798 = w12755 & ~w12757;
assign w13799 = ~w12753 & w40056;
assign w13800 = w12705 & w13794;
assign w13801 = ~w12747 & w13800;
assign w13802 = ~w13788 & w13801;
assign w13803 = ~w13799 & ~w13802;
assign w13804 = ~w13797 & w13803;
assign w13805 = ~w12761 & ~w13804;
assign w13806 = w13182 & w13805;
assign w13807 = w13751 & w13806;
assign w13808 = ~w13169 & w13711;
assign w13809 = ~w13710 & ~w13808;
assign w13810 = ~w13746 & ~w13809;
assign w13811 = ~w13688 & ~w13696;
assign w13812 = (w13696 & w13575) | (w13696 & w38130) | (w13575 & w38130);
assign w13813 = w13567 & ~w13812;
assign w13814 = (~w13605 & w13813) | (~w13605 & w38131) | (w13813 & w38131);
assign w13815 = w13701 & w13814;
assign w13816 = (~w13565 & w13701) | (~w13565 & w38132) | (w13701 & w38132);
assign w13817 = ~w13815 & ~w13816;
assign w13818 = ~w5119 & w10777;
assign w13819 = ~w4366 & w10775;
assign w13820 = ~w13818 & ~w13819;
assign w13821 = (w13820 & ~w13316) | (w13820 & w38133) | (~w13316 & w38133);
assign w13822 = w13316 & w38134;
assign w13823 = ~w13821 & ~w13822;
assign w13824 = w13814 & w13823;
assign w13825 = ~w13814 & ~w13823;
assign w13826 = ~w13824 & ~w13825;
assign w13827 = ~w13817 & w13826;
assign w13828 = w13817 & ~w13826;
assign w13829 = ~w13827 & ~w13828;
assign w13830 = ~w13808 & ~w13829;
assign w13831 = w13808 & w13829;
assign w13832 = ~w13830 & ~w13831;
assign w13833 = w13810 & w13832;
assign w13834 = ~w13810 & ~w13832;
assign w13835 = ~w13833 & ~w13834;
assign w13836 = pi0868 & ~w13835;
assign w13837 = ~w13807 & w38135;
assign w13838 = ~w13754 & w13837;
assign w13839 = pi0868 & w13835;
assign w13840 = (~w13839 & w13807) | (~w13839 & w38136) | (w13807 & w38136);
assign w13841 = w13752 & w38137;
assign w13842 = ~w12505 & w13841;
assign w13843 = ~w13840 & ~w13842;
assign w13844 = ~w13838 & w13843;
assign w13845 = w13540 & ~w13804;
assign w13846 = w13183 & w13845;
assign w13847 = ~w13785 & ~w13846;
assign w13848 = w13687 & ~w13718;
assign w13849 = ~pi0868 & ~w13848;
assign w13850 = (w13849 & w13745) | (w13849 & w38138) | (w13745 & w38138);
assign w13851 = ~w13847 & w13850;
assign w13852 = ~w13192 & w13540;
assign w13853 = w13183 & w13852;
assign w13854 = w13852 & w38139;
assign w13855 = ~w12505 & w13854;
assign w13856 = ~w13851 & ~w13855;
assign w13857 = w13769 & w38140;
assign w13858 = ~w13765 & w13857;
assign w13859 = (w13858 & ~w13540) | (w13858 & w38141) | (~w13540 & w38141);
assign w13860 = w13782 & w13858;
assign w13861 = ~w13778 & w13860;
assign w13862 = ~w13859 & ~w13861;
assign w13863 = ~w13686 & ~w13745;
assign w13864 = ~w13861 & w38142;
assign w13865 = w13539 & w38143;
assign w13866 = w13806 & w13865;
assign w13867 = (~w13718 & w13866) | (~w13718 & w38144) | (w13866 & w38144);
assign w13868 = ~w13192 & w13865;
assign w13869 = w13183 & w13868;
assign w13870 = w13868 & w38145;
assign w13871 = ~w12505 & w13870;
assign w13872 = ~w13867 & ~w13871;
assign w13873 = ~w13856 & w13872;
assign w13874 = ~w13844 & ~w13873;
assign w13875 = w10752 & ~w13874;
assign w13876 = ~w10763 & ~w13875;
assign w13877 = (~w13743 & w13738) | (~w13743 & w38146) | (w13738 & w38146);
assign w13878 = w13852 & w38147;
assign w13879 = ~w12505 & w13878;
assign w13880 = ~w13804 & w38148;
assign w13881 = w13183 & w13880;
assign w13882 = ~w13765 & w13770;
assign w13883 = (w13882 & ~w13540) | (w13882 & w38149) | (~w13540 & w38149);
assign w13884 = w13782 & w13882;
assign w13885 = ~w13778 & w13884;
assign w13886 = ~w13885 & w38150;
assign w13887 = ~w13881 & ~w13886;
assign w13888 = ~w13663 & ~w13687;
assign w13889 = ~w13685 & ~w13888;
assign w13890 = w13887 & w13889;
assign w13891 = ~w13879 & w13890;
assign w13892 = pi0868 & ~w13719;
assign w13893 = ~w13892 & w40142;
assign w13894 = ~w13862 & ~w13892;
assign w13895 = (~w13893 & ~w13894) | (~w13893 & w38152) | (~w13894 & w38152);
assign w13896 = w13852 & w40057;
assign w13897 = ~w12505 & w13896;
assign w13898 = ~w13895 & ~w13897;
assign w13899 = ~w13891 & w13898;
assign w13900 = ~w12505 & w13869;
assign w13901 = pi0868 & w13719;
assign w13902 = ~w13866 & w38153;
assign w13903 = ~w13900 & w13902;
assign w13904 = pi0868 & ~w13718;
assign w13905 = w13687 & w13904;
assign w13906 = (~w13905 & w13861) | (~w13905 & w38154) | (w13861 & w38154);
assign w13907 = ~w13846 & w13906;
assign w13908 = (w13904 & w13745) | (w13904 & w38156) | (w13745 & w38156);
assign w13909 = ~w13907 & w13908;
assign w13910 = w13852 & w38157;
assign w13911 = ~w12505 & w13910;
assign w13912 = ~w13909 & ~w13911;
assign w13913 = ~w13903 & w13912;
assign w13914 = ~w13899 & w38158;
assign w13915 = pi3245 & ~w7537;
assign w13916 = ~w13915 & w40143;
assign w13917 = (~pi0040 & ~w40209) | (~pi0040 & w38161) | (~w40209 & w38161);
assign w13918 = w10759 & ~w13917;
assign w13919 = (w13918 & w13916) | (w13918 & w38162) | (w13916 & w38162);
assign w13920 = w10756 & ~w13919;
assign w13921 = ~w13914 & ~w13920;
assign w13922 = (~pi0979 & ~w341) | (~pi0979 & w38163) | (~w341 & w38163);
assign w13923 = w10751 & w13922;
assign w13924 = ~w13874 & w13923;
assign w13925 = w10747 & w40144;
assign w13926 = pi0053 & w40145;
assign w13927 = (~w13926 & ~w10751) | (~w13926 & w38166) | (~w10751 & w38166);
assign w13928 = ~pi0714 & w40144;
assign w13929 = ~w10747 & w40146;
assign w13930 = (w13927 & w10746) | (w13927 & w38167) | (w10746 & w38167);
assign w13931 = ~pi0713 & w40144;
assign w13932 = (w5319 & w38168) | (w5319 & w38169) | (w38168 & w38169);
assign w13933 = ~w13925 & ~w13928;
assign w13934 = (~pi0041 & ~w40144) | (~pi0041 & w38170) | (~w40144 & w38170);
assign w13935 = w13933 & ~w13934;
assign w13936 = ~w13932 & w13935;
assign w13937 = w13930 & ~w13936;
assign w13938 = ~w13924 & ~w13937;
assign w13939 = ~w13899 & w38171;
assign w13940 = (~pi0042 & ~w40144) | (~pi0042 & w38172) | (~w40144 & w38172);
assign w13941 = w13933 & ~w13940;
assign w13942 = (w13941 & w13916) | (w13941 & w38173) | (w13916 & w38173);
assign w13943 = w13930 & ~w13942;
assign w13944 = ~w13939 & ~w13943;
assign w13945 = ~w370 & w10614;
assign w13946 = w10614 & w38174;
assign w13947 = pi0043 & ~w13946;
assign w13948 = w13874 & w13946;
assign w13949 = ~w13947 & ~w13948;
assign w13950 = (w13946 & w13899) | (w13946 & w38175) | (w13899 & w38175);
assign w13951 = pi0044 & ~w13946;
assign w13952 = ~w13950 & ~w13951;
assign w13953 = ~pi1798 & ~pi2340;
assign w13954 = pi1798 & ~pi2329;
assign w13955 = pi1713 & ~w13954;
assign w13956 = ~w13953 & w13955;
assign w13957 = pi2354 & w6760;
assign w13958 = pi2364 & w6758;
assign w13959 = ~w13957 & ~w13958;
assign w13960 = ~w13956 & w13959;
assign w13961 = pi0134 & ~w13960;
assign w13962 = ~pi1798 & ~pi2519;
assign w13963 = pi1798 & ~pi2335;
assign w13964 = pi1713 & ~w13963;
assign w13965 = ~w13962 & w13964;
assign w13966 = pi2358 & w6760;
assign w13967 = pi2471 & w6758;
assign w13968 = ~w13966 & ~w13967;
assign w13969 = ~w13965 & w13968;
assign w13970 = ~pi0152 & w13969;
assign w13971 = pi0152 & ~w13969;
assign w13972 = ~w13970 & ~w13971;
assign w13973 = ~w13961 & ~w13972;
assign w13974 = ~pi1798 & ~pi2338;
assign w13975 = pi1798 & ~pi1990;
assign w13976 = pi1713 & ~w13975;
assign w13977 = ~w13974 & w13976;
assign w13978 = pi2001 & w6760;
assign w13979 = pi2362 & w6758;
assign w13980 = ~w13978 & ~w13979;
assign w13981 = ~w13977 & w13980;
assign w13982 = ~pi1798 & ~pi2406;
assign w13983 = pi1798 & ~pi2328;
assign w13984 = pi1713 & ~w13983;
assign w13985 = ~w13982 & w13984;
assign w13986 = pi2353 & w6760;
assign w13987 = pi2407 & w6758;
assign w13988 = ~w13986 & ~w13987;
assign w13989 = ~w13985 & w13988;
assign w13990 = w13981 & ~w13989;
assign w13991 = (w13990 & ~w13972) | (w13990 & w38176) | (~w13972 & w38176);
assign w13992 = ~w13973 & w13991;
assign w13993 = pi0196 & ~w13969;
assign w13994 = ~w13960 & ~w13993;
assign w13995 = ~w13981 & w13989;
assign w13996 = ~pi0196 & w13969;
assign w13997 = w13995 & ~w13996;
assign w13998 = w13994 & w13997;
assign w13999 = ~w13992 & ~w13998;
assign w14000 = w10689 & w38177;
assign w14001 = ~w343 & ~w14000;
assign w14002 = w13960 & ~w13969;
assign w14003 = (w10707 & w38178) | (w10707 & w38179) | (w38178 & w38179);
assign w14004 = w13960 & w13969;
assign w14005 = w14004 & ~w10711;
assign w14006 = ~w14003 & ~w14005;
assign w14007 = (~w13960 & ~w10689) | (~w13960 & w38180) | (~w10689 & w38180);
assign w14008 = w13969 & w14007;
assign w14009 = (w13995 & ~w14006) | (w13995 & w38181) | (~w14006 & w38181);
assign w14010 = w14001 & ~w14009;
assign w14011 = ~w10682 & w14010;
assign w14012 = ~w13969 & w14007;
assign w14013 = (w13995 & ~w14006) | (w13995 & w38182) | (~w14006 & w38182);
assign w14014 = w14001 & ~w14013;
assign w14015 = w10682 & w14014;
assign w14016 = (w10741 & ~w342) | (w10741 & w38184) | (~w342 & w38184);
assign w14017 = ~w14015 & w14016;
assign w14018 = ~w14011 & w14017;
assign w14019 = (w13990 & ~w10689) | (w13990 & w38185) | (~w10689 & w38185);
assign w14020 = ~w13960 & w14019;
assign w14021 = ~w10625 & w38186;
assign w14022 = ~w10641 & w13969;
assign w14023 = w10641 & ~w13969;
assign w14024 = ~w14022 & ~w14023;
assign w14025 = w14019 & w40147;
assign w14026 = ~w14021 & w14025;
assign w14027 = (~w14026 & ~w10652) | (~w14026 & w38188) | (~w10652 & w38188);
assign w14028 = ~w13960 & w13969;
assign w14029 = ~w10625 & w38189;
assign w14030 = ~w13960 & ~w14024;
assign w14031 = (~w14030 & w10625) | (~w14030 & w38190) | (w10625 & w38190);
assign w14032 = ~w14029 & ~w14031;
assign w14033 = (w14016 & ~w10652) | (w14016 & w38191) | (~w10652 & w38191);
assign w14034 = ~w14027 & w14033;
assign w14035 = ~w14018 & ~w14034;
assign w14036 = (pi3245 & w7504) | (pi3245 & w38192) | (w7504 & w38192);
assign w14037 = (~pi0046 & ~w40209) | (~pi0046 & w38196) | (~w40209 & w38196);
assign w14038 = w10759 & ~w14037;
assign w14039 = (w14038 & w40159) | (w14038 & w38197) | (w40159 & w38197);
assign w14040 = w10756 & ~w14039;
assign w14041 = (~w10752 & w14039) | (~w10752 & w38198) | (w14039 & w38198);
assign w14042 = w13539 & w38199;
assign w14043 = ~w13192 & w14042;
assign w14044 = w13183 & w14043;
assign w14045 = ~w12505 & w14044;
assign w14046 = ~w13885 & w38200;
assign w14047 = w13806 & w14042;
assign w14048 = ~w13685 & ~w13743;
assign w14049 = ~pi0868 & ~w14048;
assign w14050 = ~w14047 & w38201;
assign w14051 = ~w14045 & w14050;
assign w14052 = ~pi0868 & w14048;
assign w14053 = (~w14052 & w14047) | (~w14052 & w38202) | (w14047 & w38202);
assign w14054 = w14043 & w38203;
assign w14055 = ~w12505 & w14054;
assign w14056 = ~w14053 & ~w14055;
assign w14057 = ~w14051 & w14056;
assign w14058 = ~w13685 & w13887;
assign w14059 = ~w13879 & w14058;
assign w14060 = pi0868 & w13888;
assign w14061 = ~w14059 & w14060;
assign w14062 = ~w14057 & ~w14061;
assign w14063 = (~w14040 & ~w13891) | (~w14040 & w38204) | (~w13891 & w38204);
assign w14064 = w14062 & w14063;
assign w14065 = ~w14041 & ~w14064;
assign w14066 = (w4748 & w38205) | (w4748 & w38206) | (w38205 & w38206);
assign w14067 = (~pi0047 & ~w40144) | (~pi0047 & w38207) | (~w40144 & w38207);
assign w14068 = w13933 & ~w14067;
assign w14069 = ~w14066 & w14068;
assign w14070 = w13930 & ~w14069;
assign w14071 = (~w13923 & w14069) | (~w13923 & w38208) | (w14069 & w38208);
assign w14072 = (~w14070 & ~w13891) | (~w14070 & w38209) | (~w13891 & w38209);
assign w14073 = w14062 & w14072;
assign w14074 = ~w14071 & ~w14073;
assign w14075 = pi0048 & ~w13946;
assign w14076 = (w13946 & ~w13891) | (w13946 & w38210) | (~w13891 & w38210);
assign w14077 = w14062 & w14076;
assign w14078 = ~w14075 & ~w14077;
assign w14079 = pi0868 & w14048;
assign w14080 = ~w14047 & w38211;
assign w14081 = ~w14045 & w14080;
assign w14082 = pi0868 & ~w14048;
assign w14083 = (~w14082 & w14047) | (~w14082 & w38212) | (w14047 & w38212);
assign w14084 = w14043 & w40058;
assign w14085 = ~w12505 & w14084;
assign w14086 = ~w14083 & ~w14085;
assign w14087 = ~w14081 & w14086;
assign w14088 = w13539 & w38213;
assign w14089 = ~w13192 & w14088;
assign w14090 = w13183 & w14089;
assign w14091 = ~w12505 & w14090;
assign w14092 = w13806 & w14088;
assign w14093 = ~w13765 & w13769;
assign w14094 = ~w13778 & w13782;
assign w14095 = ~w13778 & w38214;
assign w14096 = (w14093 & ~w13540) | (w14093 & w38215) | (~w13540 & w38215);
assign w14097 = w13730 & ~w14096;
assign w14098 = ~w14095 & w14097;
assign w14099 = ~w14092 & ~w14098;
assign w14100 = ~pi0868 & w13737;
assign w14101 = ~w14092 & w38216;
assign w14102 = ~w14091 & w14101;
assign w14103 = ~pi0868 & ~w13737;
assign w14104 = (w14103 & w14092) | (w14103 & w38217) | (w14092 & w38217);
assign w14105 = w14089 & w38218;
assign w14106 = ~w12505 & w14105;
assign w14107 = ~w14104 & ~w14106;
assign w14108 = ~w14102 & w14107;
assign w14109 = ~w14087 & w38219;
assign w14110 = pi3245 & ~w7473;
assign w14111 = (~pi0049 & ~w40209) | (~pi0049 & w38223) | (~w40209 & w38223);
assign w14112 = w10759 & ~w14111;
assign w14113 = (w14112 & w40171) | (w14112 & w38224) | (w40171 & w38224);
assign w14114 = w10756 & ~w14113;
assign w14115 = ~w14109 & ~w14114;
assign w14116 = ~w14087 & w38225;
assign w14117 = (w3710 & w38226) | (w3710 & w38227) | (w38226 & w38227);
assign w14118 = (~pi0050 & ~w40144) | (~pi0050 & w38228) | (~w40144 & w38228);
assign w14119 = w13933 & ~w14118;
assign w14120 = ~w14117 & w14119;
assign w14121 = w13930 & ~w14120;
assign w14122 = ~w14116 & ~w14121;
assign w14123 = ~w6316 & w10775;
assign w14124 = ~w4366 & w10777;
assign w14125 = ~w14123 & ~w14124;
assign w14126 = ~w13812 & ~w13820;
assign w14127 = ~w13567 & ~w14126;
assign w14128 = (~w13820 & ~w13575) | (~w13820 & w38229) | (~w13575 & w38229);
assign w14129 = ~w13606 & ~w14128;
assign w14130 = (w13565 & w14127) | (w13565 & w38230) | (w14127 & w38230);
assign w14131 = ~w14125 & w14130;
assign w14132 = ~w14127 & w38231;
assign w14133 = ~w14130 & ~w14132;
assign w14134 = w13826 & w38232;
assign w14135 = ~w14131 & ~w14134;
assign w14136 = w14125 & ~w14132;
assign w14137 = (~w14125 & w13826) | (~w14125 & w38233) | (w13826 & w38233);
assign w14138 = ~w14136 & ~w14137;
assign w14139 = w14135 & ~w14138;
assign w14140 = ~w13827 & w14139;
assign w14141 = w13827 & ~w14139;
assign w14142 = ~w14140 & ~w14141;
assign w14143 = ~w13817 & w38234;
assign w14144 = ~w13828 & ~w14143;
assign w14145 = ~w13808 & ~w14144;
assign w14146 = ~w14142 & w14145;
assign w14147 = ~w13833 & ~w14146;
assign w14148 = w13719 & w14147;
assign w14149 = ~w13686 & w14148;
assign w14150 = w13770 & w14149;
assign w14151 = ~w13765 & w14150;
assign w14152 = (w14151 & ~w13540) | (w14151 & w38235) | (~w13540 & w38235);
assign w14153 = w13782 & w14151;
assign w14154 = ~w13778 & w14153;
assign w14155 = ~w14152 & ~w14154;
assign w14156 = ~w14137 & w38236;
assign w14157 = ~w6316 & w10777;
assign w14158 = ~w3335 & w10775;
assign w14159 = ~w14157 & ~w14158;
assign w14160 = ~w14125 & ~w14129;
assign w14161 = w13565 & ~w14160;
assign w14162 = w13588 & w14160;
assign w14163 = (w14125 & w13575) | (w14125 & w38237) | (w13575 & w38237);
assign w14164 = ~w13605 & ~w14163;
assign w14165 = w13567 & w14164;
assign w14166 = ~w14162 & ~w14165;
assign w14167 = (w14159 & ~w14166) | (w14159 & w38238) | (~w14166 & w38238);
assign w14168 = w14166 & w38239;
assign w14169 = ~w14167 & ~w14168;
assign w14170 = ~w14130 & w14166;
assign w14171 = (~w14161 & ~w14170) | (~w14161 & w38240) | (~w14170 & w38240);
assign w14172 = w14169 & ~w14171;
assign w14173 = ~w14156 & w14172;
assign w14174 = ~w14169 & w14171;
assign w14175 = ~w13169 & w14174;
assign w14176 = w14138 & w14175;
assign w14177 = ~w14173 & ~w14176;
assign w14178 = ~w3335 & w10777;
assign w14179 = ~w1143 & w10775;
assign w14180 = ~w14178 & ~w14179;
assign w14181 = ~w13588 & w14180;
assign w14182 = w13588 & ~w14180;
assign w14183 = ~w14181 & ~w14182;
assign w14184 = (~w14159 & ~w13575) | (~w14159 & w38241) | (~w13575 & w38241);
assign w14185 = ~w13606 & ~w14184;
assign w14186 = w14183 & ~w14185;
assign w14187 = ~w14183 & w14185;
assign w14188 = ~w14186 & ~w14187;
assign w14189 = ~w14159 & ~w14163;
assign w14190 = ~w14185 & ~w14189;
assign w14191 = ~w13567 & ~w14190;
assign w14192 = ~w14188 & w14191;
assign w14193 = w14188 & ~w14191;
assign w14194 = ~w14192 & ~w14193;
assign w14195 = w13567 & ~w14185;
assign w14196 = w13565 & w14160;
assign w14197 = ~w14159 & ~w14164;
assign w14198 = ~w14196 & ~w14197;
assign w14199 = (~w14195 & w14167) | (~w14195 & w38242) | (w14167 & w38242);
assign w14200 = w14194 & ~w14199;
assign w14201 = ~w14194 & w14199;
assign w14202 = ~w14200 & ~w14201;
assign w14203 = w14177 & ~w14202;
assign w14204 = ~w14177 & w14202;
assign w14205 = ~w14203 & ~w14204;
assign w14206 = ~w13827 & w14156;
assign w14207 = ~w14135 & ~w14143;
assign w14208 = ~w14206 & ~w14207;
assign w14209 = ~w14156 & ~w14207;
assign w14210 = ~w14172 & ~w14174;
assign w14211 = (w14210 & w14209) | (w14210 & w38243) | (w14209 & w38243);
assign w14212 = ~w14209 & w38244;
assign w14213 = ~w14211 & ~w14212;
assign w14214 = ~w14208 & w14213;
assign w14215 = ~w14205 & ~w14214;
assign w14216 = (~w14173 & ~w14202) | (~w14173 & w38245) | (~w14202 & w38245);
assign w14217 = ~w14203 & w14216;
assign w14218 = ~w14215 & ~w14217;
assign w14219 = (~w14218 & w14154) | (~w14218 & w38246) | (w14154 & w38246);
assign w14220 = ~w13846 & w14219;
assign w14221 = ~w13745 & w14149;
assign w14222 = ~w14139 & w14144;
assign w14223 = (~w14222 & ~w14142) | (~w14222 & w38247) | (~w14142 & w38247);
assign w14224 = ~w13749 & ~w13834;
assign w14225 = (w14147 & w13749) | (w14147 & w38248) | (w13749 & w38248);
assign w14226 = w14223 & ~w14225;
assign w14227 = ~w14225 & w38249;
assign w14228 = ~w14221 & w14227;
assign w14229 = (w14215 & w14221) | (w14215 & w38250) | (w14221 & w38250);
assign w14230 = ~w14217 & ~w14229;
assign w14231 = ~w14220 & w14230;
assign w14232 = w13852 & w38251;
assign w14233 = ~w12505 & w14232;
assign w14234 = ~w14231 & ~w14233;
assign w14235 = w14174 & w38252;
assign w14236 = (~w14180 & ~w13575) | (~w14180 & w38253) | (~w13575 & w38253);
assign w14237 = ~w13606 & ~w14236;
assign w14238 = ~w13565 & ~w14237;
assign w14239 = (w14180 & ~w13316) | (w14180 & w38254) | (~w13316 & w38254);
assign w14240 = w14185 & w14239;
assign w14241 = ~w14238 & ~w14240;
assign w14242 = ~w14235 & ~w14241;
assign w14243 = (~w14237 & ~w13588) | (~w14237 & w38255) | (~w13588 & w38255);
assign w14244 = w14235 & ~w14243;
assign w14245 = (w14199 & ~w14174) | (w14199 & w38256) | (~w14174 & w38256);
assign w14246 = w14188 & ~w14245;
assign w14247 = ~w14244 & w14246;
assign w14248 = ~w14242 & w14247;
assign w14249 = w14192 & ~w14235;
assign w14250 = ~w14191 & w14241;
assign w14251 = w14191 & ~w14241;
assign w14252 = ~w14250 & ~w14251;
assign w14253 = w14188 & w14252;
assign w14254 = w14245 & ~w14253;
assign w14255 = ~w14249 & ~w14254;
assign w14256 = ~w1143 & w10774;
assign w14257 = w13588 & ~w14188;
assign w14258 = (w14183 & w38258) | (w14183 & w38259) | (w38258 & w38259);
assign w14259 = ~w14257 & w38260;
assign w14260 = (w14256 & w14257) | (w14256 & w38261) | (w14257 & w38261);
assign w14261 = ~w14259 & ~w14260;
assign w14262 = (w14261 & w14248) | (w14261 & w38262) | (w14248 & w38262);
assign w14263 = ~w14248 & w38263;
assign w14264 = ~w14262 & ~w14263;
assign w14265 = pi0868 & w14264;
assign w14266 = w14234 & w14265;
assign w14267 = pi0868 & ~w14264;
assign w14268 = ~w14234 & w14267;
assign w14269 = ~w14266 & ~w14268;
assign w14270 = w13540 & w14228;
assign w14271 = ~w13192 & w14270;
assign w14272 = w13183 & w14271;
assign w14273 = ~w12505 & w14272;
assign w14274 = ~w14154 & w38264;
assign w14275 = w13806 & w14270;
assign w14276 = ~pi0868 & w14215;
assign w14277 = ~w14275 & w38265;
assign w14278 = ~w14273 & w14277;
assign w14279 = ~w13846 & ~w14155;
assign w14280 = ~pi0868 & w14205;
assign w14281 = ~w14221 & w38266;
assign w14282 = ~w14279 & w14281;
assign w14283 = w13852 & w38267;
assign w14284 = ~w12505 & w14283;
assign w14285 = ~w14282 & ~w14284;
assign w14286 = ~w14278 & w14285;
assign w14287 = (w10752 & ~w14280) | (w10752 & w38268) | (~w14280 & w38268);
assign w14288 = w14286 & w14287;
assign w14289 = w14269 & w14288;
assign w14290 = (pi3245 & w7699) | (pi3245 & w38269) | (w7699 & w38269);
assign w14291 = (~pi0051 & ~w40209) | (~pi0051 & w38273) | (~w40209 & w38273);
assign w14292 = w10759 & ~w14291;
assign w14293 = (w14292 & w40174) | (w14292 & w38274) | (w40174 & w38274);
assign w14294 = w10756 & ~w14293;
assign w14295 = ~w14289 & ~w14294;
assign w14296 = ~w14221 & w14226;
assign w14297 = w13852 & w38275;
assign w14298 = ~w12505 & w14297;
assign w14299 = ~w14154 & w38276;
assign w14300 = ~w13804 & w38277;
assign w14301 = w13183 & w14300;
assign w14302 = ~w14299 & ~w14301;
assign w14303 = w14213 & w14302;
assign w14304 = ~w14298 & w14303;
assign w14305 = ~w14275 & w38278;
assign w14306 = ~w14273 & w14305;
assign w14307 = ~w14304 & w14306;
assign w14308 = pi0868 & w14215;
assign w14309 = ~w14275 & w38279;
assign w14310 = ~w14273 & w14309;
assign w14311 = pi0868 & w14205;
assign w14312 = w14214 & w14311;
assign w14313 = (~w14312 & w14154) | (~w14312 & w38280) | (w14154 & w38280);
assign w14314 = ~w13846 & w14313;
assign w14315 = (~w14214 & w14221) | (~w14214 & w38281) | (w14221 & w38281);
assign w14316 = w14311 & ~w14315;
assign w14317 = ~w14314 & w14316;
assign w14318 = w13852 & w38282;
assign w14319 = ~w12505 & w14318;
assign w14320 = ~w14317 & ~w14319;
assign w14321 = ~w14310 & w14320;
assign w14322 = ~w14307 & w14321;
assign w14323 = w10752 & w14322;
assign w14324 = (pi3245 & w7667) | (pi3245 & w38283) | (w7667 & w38283);
assign w14325 = ~w14324 & w40151;
assign w14326 = (~pi0052 & ~w40209) | (~pi0052 & w38286) | (~w40209 & w38286);
assign w14327 = w10759 & ~w14326;
assign w14328 = (w14327 & w14325) | (w14327 & w38287) | (w14325 & w38287);
assign w14329 = w10756 & ~w14328;
assign w14330 = ~w14323 & ~w14329;
assign w14331 = (w3194 & w38288) | (w3194 & w38289) | (w38288 & w38289);
assign w14332 = (pi0053 & ~w40144) | (pi0053 & w38290) | (~w40144 & w38290);
assign w14333 = ~w13928 & ~w14332;
assign w14334 = (w14333 & w14331) | (w14333 & w38291) | (w14331 & w38291);
assign w14335 = ~pi0053 & w40145;
assign w14336 = (~w14335 & ~w10751) | (~w14335 & w38292) | (~w10751 & w38292);
assign w14337 = (w14336 & ~w10746) | (w14336 & w38293) | (~w10746 & w38293);
assign w14338 = ~w14334 & w14337;
assign w14339 = (~w14338 & ~w14280) | (~w14338 & w38294) | (~w14280 & w38294);
assign w14340 = w14286 & w14339;
assign w14341 = w14269 & w14340;
assign w14342 = (~w13923 & w14334) | (~w13923 & w38295) | (w14334 & w38295);
assign w14343 = ~w14341 & ~w14342;
assign w14344 = w13923 & w14322;
assign w14345 = (~pi0054 & ~w40144) | (~pi0054 & w38296) | (~w40144 & w38296);
assign w14346 = w13933 & ~w14345;
assign w14347 = (w14346 & w14325) | (w14346 & w38297) | (w14325 & w38297);
assign w14348 = w13930 & ~w14347;
assign w14349 = ~w14344 & ~w14348;
assign w14350 = pi0425 & ~w923;
assign w14351 = (w921 & w38298) | (w921 & w38299) | (w38298 & w38299);
assign w14352 = ~w14350 & ~w14351;
assign w14353 = pi0406 & ~w923;
assign w14354 = (w921 & w38300) | (w921 & w38301) | (w38300 & w38301);
assign w14355 = ~w14353 & ~w14354;
assign w14356 = ~w14352 & ~w14355;
assign w14357 = ~pi0416 & w374;
assign w14358 = w374 & w38302;
assign w14359 = ~pi0419 & w14358;
assign w14360 = w14358 & w38303;
assign w14361 = ~w923 & w14360;
assign w14362 = (w921 & w38304) | (w921 & w38305) | (w38304 & w38305);
assign w14363 = ~w14361 & ~w14362;
assign w14364 = ~w14356 & ~w14363;
assign w14365 = ~pi0426 & ~pi0715;
assign w14366 = ~pi0405 & ~pi0422;
assign w14367 = ~pi0423 & ~pi0424;
assign w14368 = w14366 & w14367;
assign w14369 = ~pi0421 & ~w14368;
assign w14370 = ~pi0416 & w2241;
assign w14371 = w374 & ~w14370;
assign w14372 = ~w2237 & ~w2355;
assign w14373 = ~w14371 & w14372;
assign w14374 = (w14369 & ~w14372) | (w14369 & w38306) | (~w14372 & w38306);
assign w14375 = ~pi3426 & w14374;
assign w14376 = pi0410 & pi0426;
assign w14377 = pi0709 & w14376;
assign w14378 = pi0426 & ~pi0710;
assign w14379 = ~pi0410 & ~w14365;
assign w14380 = ~w14378 & w14379;
assign w14381 = ~w14377 & ~w14380;
assign w14382 = ~pi0410 & ~pi2020;
assign w14383 = ~pi0426 & ~w14382;
assign w14384 = pi0426 & pi2140;
assign w14385 = ~w14383 & ~w14384;
assign w14386 = (w14381 & w10613) | (w14381 & w38307) | (w10613 & w38307);
assign w14387 = ~pi0409 & pi0426;
assign w14388 = ~pi0714 & w14387;
assign w14389 = pi0409 & pi0410;
assign w14390 = ~pi0426 & w14389;
assign w14391 = w14389 & w38308;
assign w14392 = ~w14388 & ~w14391;
assign w14393 = ~w14387 & ~w14390;
assign w14394 = (w10747 & w14390) | (w10747 & w38309) | (w14390 & w38309);
assign w14395 = ~pi0409 & ~pi0713;
assign w14396 = w14376 & w14395;
assign w14397 = ~w14394 & ~w14396;
assign w14398 = w14392 & w14397;
assign w14399 = (w14398 & w14386) | (w14398 & w38310) | (w14386 & w38310);
assign w14400 = pi0409 & ~w923;
assign w14401 = ~w14399 & w38313;
assign w14402 = w10048 & w38314;
assign w14403 = ~w10096 & w38315;
assign w14404 = (w14403 & w10660) | (w14403 & w38316) | (w10660 & w38316);
assign w14405 = ~w10553 & ~w14404;
assign w14406 = ~w10664 & w40139;
assign w14407 = ~w14405 & ~w14406;
assign w14408 = ~w14405 & w38317;
assign w14409 = (w14401 & w10552) | (w14401 & w38318) | (w10552 & w38318);
assign w14410 = ~w14404 & w14409;
assign w14411 = ~w10261 & w38319;
assign w14412 = (w14411 & w10354) | (w14411 & w38320) | (w10354 & w38320);
assign w14413 = (~w10605 & w10354) | (~w10605 & w38321) | (w10354 & w38321);
assign w14414 = ~w10357 & ~w14413;
assign w14415 = (w10354 & w38322) | (w10354 & w38323) | (w38322 & w38323);
assign w14416 = ~w10593 & ~w14415;
assign w14417 = ~w14414 & w14416;
assign w14418 = (w10594 & ~w10261) | (w10594 & w38324) | (~w10261 & w38324);
assign w14419 = ~w10277 & ~w14418;
assign w14420 = (~w14412 & w14417) | (~w14412 & w38325) | (w14417 & w38325);
assign w14421 = w14410 & ~w14420;
assign w14422 = ~w14399 & w38326;
assign w14423 = ~w8199 & w9951;
assign w14424 = w9949 & w38327;
assign w14425 = ~pi3504 & pi3514;
assign w14426 = ~w14424 & w14425;
assign w14427 = pi3504 & ~pi3514;
assign w14428 = w3567 & w4670;
assign w14429 = w14428 & w18917;
assign w14430 = w14429 & w38329;
assign w14431 = ~w14430 & w38330;
assign w14432 = ~pi2486 & ~w14427;
assign w14433 = w1182 & ~w14432;
assign w14434 = ~pi3521 & w14432;
assign w14435 = ~w14434 & w40152;
assign w14436 = ~w14431 & w14435;
assign w14437 = (w14427 & ~w14429) | (w14427 & w38332) | (~w14429 & w38332);
assign w14438 = ~w3392 & ~w14432;
assign w14439 = ~w14437 & w14438;
assign w14440 = ~w14427 & w38333;
assign w14441 = (~w14440 & ~w14437) | (~w14440 & w38334) | (~w14437 & w38334);
assign w14442 = ~w14439 & w14441;
assign w14443 = ~w6295 & ~w14432;
assign w14444 = (w14429 & w38336) | (w14429 & w38337) | (w38336 & w38337);
assign w14445 = w6295 & w40153;
assign w14446 = pi3511 & w14432;
assign w14447 = ~w14445 & ~w14446;
assign w14448 = ~w14444 & w14447;
assign w14449 = pi3504 & pi3514;
assign w14450 = ~pi2021 & ~w14449;
assign w14451 = (w14450 & ~w14447) | (w14450 & w38338) | (~w14447 & w38338);
assign w14452 = ~w14442 & w14451;
assign w14453 = w14436 & w14452;
assign w14454 = w14452 & w38339;
assign w14455 = w14426 & w14454;
assign w14456 = (w14427 & ~w14428) | (w14427 & w38340) | (~w14428 & w38340);
assign w14457 = w5209 & w14456;
assign w14458 = ~w5209 & ~w14432;
assign w14459 = ~w14427 & w38341;
assign w14460 = (~w14459 & w14456) | (~w14459 & w38342) | (w14456 & w38342);
assign w14461 = ~w14457 & w14460;
assign w14462 = ~w3567 & w14427;
assign w14463 = ~w4670 & w14462;
assign w14464 = w4670 & ~w14432;
assign w14465 = ~w14462 & w14464;
assign w14466 = ~w14427 & w38343;
assign w14467 = ~w14465 & ~w14466;
assign w14468 = ~w14463 & w14467;
assign w14469 = ~w14461 & ~w14468;
assign w14470 = ~w4327 & ~w14432;
assign w14471 = (w14470 & w14429) | (w14470 & w38344) | (w14429 & w38344);
assign w14472 = pi3520 & w14432;
assign w14473 = (~w14472 & w14429) | (~w14472 & w38346) | (w14429 & w38346);
assign w14474 = ~w14471 & w14473;
assign w14475 = ~w5763 & ~w14428;
assign w14476 = w14456 & ~w14475;
assign w14477 = pi2486 & ~w14427;
assign w14478 = ~w5763 & w14477;
assign w14479 = ~w14427 & w38347;
assign w14480 = ~w14478 & ~w14479;
assign w14481 = ~w14476 & w14480;
assign w14482 = ~w14476 & w38348;
assign w14483 = ~w14474 & w14482;
assign w14484 = w14469 & w14483;
assign w14485 = w3567 & ~w14432;
assign w14486 = ~w14427 & w38349;
assign w14487 = ~w14485 & ~w14486;
assign w14488 = w14484 & w14487;
assign w14489 = w14467 & w38350;
assign w14490 = ~w14461 & w14489;
assign w14491 = w14483 & w14490;
assign w14492 = ~w14487 & w14491;
assign w14493 = ~w14488 & ~w14492;
assign w14494 = w14455 & ~w14493;
assign w14495 = w14452 & w38351;
assign w14496 = pi0152 & pi0196;
assign w14497 = ~pi3518 & w14496;
assign w14498 = w14427 & w14497;
assign w14499 = (~w14498 & w14424) | (~w14498 & w38352) | (w14424 & w38352);
assign w14500 = w14495 & ~w14499;
assign w14501 = w14495 & w38353;
assign w14502 = (w14450 & w14476) | (w14450 & w38354) | (w14476 & w38354);
assign w14503 = w14474 & w14502;
assign w14504 = w14461 & w14489;
assign w14505 = w14503 & w14504;
assign w14506 = w14495 & w38355;
assign w14507 = w14474 & w14481;
assign w14508 = w14504 & w14507;
assign w14509 = w14495 & w38357;
assign w14510 = ~pi2021 & pi3518;
assign w14511 = ~w14424 & w38358;
assign w14512 = w14436 & w14511;
assign w14513 = w14483 & w14504;
assign w14514 = (w14487 & ~w14447) | (w14487 & w38359) | (~w14447 & w38359);
assign w14515 = (~w14442 & ~w14513) | (~w14442 & w38360) | (~w14513 & w38360);
assign w14516 = w14512 & ~w14515;
assign w14517 = ~w14509 & ~w14516;
assign w14518 = ~w14506 & w14517;
assign w14519 = w14490 & w14507;
assign w14520 = w14495 & w14519;
assign w14521 = (w14450 & w14485) | (w14450 & w38361) | (w14485 & w38361);
assign w14522 = w14521 & ~w14499;
assign w14523 = w14495 & w38362;
assign w14524 = w14461 & ~w14468;
assign w14525 = w14442 & w14448;
assign w14526 = ~w14436 & w14525;
assign w14527 = w14525 & w38363;
assign w14528 = w14527 & w38364;
assign w14529 = ~w14523 & ~w14528;
assign w14530 = w14483 & w14524;
assign w14531 = w14490 & w14503;
assign w14532 = ~w14530 & ~w14531;
assign w14533 = w14501 & ~w14532;
assign w14534 = w14450 & w14469;
assign w14535 = w14507 & w14534;
assign w14536 = w14500 & w14535;
assign w14537 = ~w14533 & ~w14536;
assign w14538 = w14529 & w14537;
assign w14539 = w14538 & w38365;
assign w14540 = ~w14448 & ~w14474;
assign w14541 = ~w14442 & ~w14540;
assign w14542 = w14512 & w14541;
assign w14543 = w14450 & ~w14507;
assign w14544 = w14524 & ~w14543;
assign w14545 = w14500 & w14544;
assign w14546 = ~w14542 & ~w14545;
assign w14547 = w14495 & w38366;
assign w14548 = w14503 & w14524;
assign w14549 = w14495 & w38367;
assign w14550 = w14450 & ~w14499;
assign w14551 = ~w14499 & w38368;
assign w14552 = w14436 & w14551;
assign w14553 = ~w14452 & w14552;
assign w14554 = ~w14549 & ~w14553;
assign w14555 = ~w14547 & w14554;
assign w14556 = w14546 & w14555;
assign w14557 = w14452 & w38369;
assign w14558 = w14557 & w38370;
assign w14559 = ~w14485 & w38371;
assign w14560 = w14469 & w14503;
assign w14561 = w14495 & w38372;
assign w14562 = ~w14499 & w14561;
assign w14563 = ~w14558 & ~w14562;
assign w14564 = w14495 & w38373;
assign w14565 = w14550 & w14564;
assign w14566 = ~w14474 & w14502;
assign w14567 = w14469 & w14566;
assign w14568 = w14559 & ~w14567;
assign w14569 = ~w14468 & w14566;
assign w14570 = ~w14568 & w14569;
assign w14571 = w14455 & w14570;
assign w14572 = w14559 & w14560;
assign w14573 = w14500 & w14572;
assign w14574 = ~w14571 & ~w14573;
assign w14575 = ~w14565 & w14574;
assign w14576 = w14563 & w14575;
assign w14577 = w14452 & w38374;
assign w14578 = w14511 & w14577;
assign w14579 = ~pi3518 & w14474;
assign w14580 = pi3518 & ~w14474;
assign w14581 = ~w14579 & ~w14580;
assign w14582 = ~w14482 & ~w14507;
assign w14583 = ~w14581 & ~w14582;
assign w14584 = (~pi3518 & w14449) | (~pi3518 & w38375) | (w14449 & w38375);
assign w14585 = w14450 & ~w14524;
assign w14586 = (~w14585 & w14583) | (~w14585 & w38376) | (w14583 & w38376);
assign w14587 = w14578 & w14586;
assign w14588 = w14531 & w14551;
assign w14589 = w14557 & w14588;
assign w14590 = ~w14587 & ~w14589;
assign w14591 = w14557 & w38377;
assign w14592 = w14490 & w14566;
assign w14593 = w14577 & w38378;
assign w14594 = ~w14591 & ~w14593;
assign w14595 = w14590 & w14594;
assign w14596 = w14576 & w14595;
assign w14597 = w14576 & w38379;
assign w14598 = w14454 & w38380;
assign w14599 = w14426 & w14598;
assign w14600 = w14504 & w14566;
assign w14601 = w14454 & w14600;
assign w14602 = w14454 & w38381;
assign w14603 = ~w14559 & w14602;
assign w14604 = ~w14599 & ~w14603;
assign w14605 = w14597 & w14604;
assign w14606 = w14597 & w38382;
assign w14607 = ~w4079 & w9951;
assign w14608 = w10428 & w38383;
assign w14609 = w14559 & ~w14608;
assign w14610 = w14525 & w38384;
assign w14611 = w14535 & w14610;
assign w14612 = w14488 & w14495;
assign w14613 = w14495 & w38385;
assign w14614 = ~w14611 & ~w14613;
assign w14615 = (~w14612 & w14614) | (~w14612 & w38386) | (w14614 & w38386);
assign w14616 = ~w14611 & w14615;
assign w14617 = (w14609 & ~w14615) | (w14609 & w38387) | (~w14615 & w38387);
assign w14618 = ~w3116 & w9951;
assign w14619 = w10118 & w38388;
assign w14620 = w14559 & ~w14619;
assign w14621 = ~w6095 & w9951;
assign w14622 = w10453 & w38389;
assign w14623 = w14521 & ~w14622;
assign w14624 = ~w14620 & ~w14623;
assign w14625 = w14519 & w14610;
assign w14626 = w14491 & w14495;
assign w14627 = ~w14625 & ~w14626;
assign w14628 = ~w14624 & ~w14627;
assign w14629 = w14505 & w14610;
assign w14630 = w14495 & w14600;
assign w14631 = ~w14629 & ~w14630;
assign w14632 = ~w5621 & w9951;
assign w14633 = w10485 & w38390;
assign w14634 = w14559 & ~w14633;
assign w14635 = ~w1195 & w9951;
assign w14636 = w10071 & w38391;
assign w14637 = w14521 & ~w14636;
assign w14638 = ~w14634 & ~w14637;
assign w14639 = ~w14631 & ~w14638;
assign w14640 = ~w14424 & w14559;
assign w14641 = w14495 & w14513;
assign w14642 = w14508 & w14610;
assign w14643 = ~w14641 & ~w14642;
assign w14644 = w14640 & ~w14643;
assign w14645 = ~w14639 & ~w14644;
assign w14646 = ~w14628 & w14645;
assign w14647 = ~w1544 & w9951;
assign w14648 = w10022 & w38392;
assign w14649 = w14559 & ~w14648;
assign w14650 = ~w7954 & w9951;
assign w14651 = w9978 & w38393;
assign w14652 = w14521 & ~w14651;
assign w14653 = ~w14649 & ~w14652;
assign w14654 = w14524 & w14566;
assign w14655 = w14495 & w14654;
assign w14656 = w14450 & w14610;
assign w14657 = w14610 & w38394;
assign w14658 = ~w14655 & ~w14657;
assign w14659 = ~w14653 & ~w14658;
assign w14660 = w5213 & w9951;
assign w14661 = ~w10221 & ~w14660;
assign w14662 = ~w10221 & w38395;
assign w14663 = ~w4318 & w9951;
assign w14664 = w10201 & w38396;
assign w14665 = w14521 & ~w14664;
assign w14666 = ~w14662 & ~w14665;
assign w14667 = w14495 & w14592;
assign w14668 = w14610 & w38397;
assign w14669 = ~w14667 & ~w14668;
assign w14670 = ~w14666 & ~w14669;
assign w14671 = w6300 & w9951;
assign w14672 = ~w10152 & ~w14671;
assign w14673 = ~w10152 & w38398;
assign w14674 = w3400 & w9951;
assign w14675 = (~w14674 & ~w10370) | (~w14674 & w38399) | (~w10370 & w38399);
assign w14676 = ~w14559 & w14675;
assign w14677 = ~w14673 & ~w14676;
assign w14678 = w14560 & w14610;
assign w14679 = w14495 & w14567;
assign w14680 = ~w14678 & ~w14679;
assign w14681 = ~w14677 & ~w14680;
assign w14682 = pi3516 & ~w5767;
assign w14683 = ~w4666 & w9951;
assign w14684 = w10303 & w38400;
assign w14685 = w14559 & ~w14684;
assign w14686 = ~w5771 & w9951;
assign w14687 = w10253 & w38401;
assign w14688 = w14521 & ~w14687;
assign w14689 = ~w14685 & ~w14688;
assign w14690 = w14526 & w14586;
assign w14691 = w14586 & w38402;
assign w14692 = ~w14682 & ~w14691;
assign w14693 = ~w14681 & w14692;
assign w14694 = w14693 & w38403;
assign w14695 = w14646 & w14694;
assign w14696 = ~w4937 & w9951;
assign w14697 = w10516 & w38404;
assign w14698 = w14450 & ~w14697;
assign w14699 = ~w14614 & w14698;
assign w14700 = w14495 & w38405;
assign w14701 = w3572 & w9951;
assign w14702 = (~w14701 & ~w10321) | (~w14701 & w38406) | (~w10321 & w38406);
assign w14703 = w14450 & w14702;
assign w14704 = w14504 & w14583;
assign w14705 = w14704 & w38407;
assign w14706 = ~w14700 & ~w14705;
assign w14707 = ~w14699 & w14706;
assign w14708 = ~w14487 & ~w14707;
assign w14709 = w14559 & ~w14499;
assign w14710 = w14502 & ~w14581;
assign w14711 = ~w14581 & w38408;
assign w14712 = w14453 & w14711;
assign w14713 = w14452 & w38409;
assign w14714 = w14583 & w14713;
assign w14715 = ~w14712 & ~w14714;
assign w14716 = w14709 & ~w14715;
assign w14717 = w14454 & w38410;
assign w14718 = w14495 & w38411;
assign w14719 = ~w14717 & ~w14718;
assign w14720 = w14550 & ~w14719;
assign w14721 = w14610 & w38412;
assign w14722 = w14454 & w38413;
assign w14723 = ~w14721 & ~w14722;
assign w14724 = ~w14720 & w14723;
assign w14725 = ~w14716 & w14724;
assign w14726 = ~w14708 & w14725;
assign w14727 = w14695 & w14726;
assign w14728 = ~w14617 & w14727;
assign w14729 = (~pi0709 & ~w14728) | (~pi0709 & w38414) | (~w14728 & w38414);
assign w14730 = w14422 & w14729;
assign w14731 = pi0342 & ~pi0343;
assign w14732 = (w5893 & w38415) | (w5893 & w38416) | (w38415 & w38416);
assign w14733 = ~pi0341 & ~pi0342;
assign w14734 = ~pi0343 & w14733;
assign w14735 = ~pi0341 & pi0342;
assign w14736 = (w921 & w38417) | (w921 & w38418) | (w38417 & w38418);
assign w14737 = ~pi0426 & w14400;
assign w14738 = ~w14736 & w40154;
assign w14739 = ~w5703 & ~w14738;
assign w14740 = w14374 & w38422;
assign w14741 = ~w1143 & ~w14376;
assign w14742 = w1143 & w14376;
assign w14743 = ~w14741 & ~w14742;
assign w14744 = w14394 & w14743;
assign w14745 = (~pi0343 & ~w14740) | (~pi0343 & w38423) | (~w14740 & w38423);
assign w14746 = ~w14739 & w14745;
assign w14747 = (w921 & w38424) | (w921 & w38425) | (w38424 & w38425);
assign w14748 = w14387 & ~w923;
assign w14749 = ~w14747 & w40155;
assign w14750 = ~w5695 & ~w14749;
assign w14751 = (w921 & w38428) | (w921 & w38429) | (w38428 & w38429);
assign w14752 = ~w14751 & w40156;
assign w14753 = ~w5718 & ~w14752;
assign w14754 = ~w14750 & ~w14753;
assign w14755 = w14746 & w14754;
assign w14756 = (~w14734 & w14755) | (~w14734 & w38433) | (w14755 & w38433);
assign w14757 = ~w14732 & ~w14756;
assign w14758 = ~w14399 & w38434;
assign w14759 = ~w14653 & w14712;
assign w14760 = w14534 & w14583;
assign w14761 = w14453 & w14760;
assign w14762 = w14521 & ~w14697;
assign w14763 = ~w14609 & ~w14762;
assign w14764 = w14760 & w38435;
assign w14765 = w14442 & w14512;
assign w14766 = pi3516 & ~w5758;
assign w14767 = (~w14766 & ~w14512) | (~w14766 & w38436) | (~w14512 & w38436);
assign w14768 = ~w14764 & w14767;
assign w14769 = w14768 & w38437;
assign w14770 = w14450 & ~w14636;
assign w14771 = w14564 & w14770;
assign w14772 = w14521 & w14702;
assign w14773 = ~w14643 & w14772;
assign w14774 = w14583 & w38438;
assign w14775 = w14469 & ~w14677;
assign w14776 = w14490 & ~w14666;
assign w14777 = w14504 & w14634;
assign w14778 = ~w14776 & ~w14777;
assign w14779 = (w14710 & ~w14778) | (w14710 & w38439) | (~w14778 & w38439);
assign w14780 = w14640 & w14704;
assign w14781 = ~w14779 & ~w14780;
assign w14782 = (w14453 & ~w14781) | (w14453 & w38440) | (~w14781 & w38440);
assign w14783 = ~w14782 & w38441;
assign w14784 = w14769 & w14783;
assign w14785 = ~w14591 & ~w14599;
assign w14786 = ~w14587 & w14785;
assign w14787 = w14495 & w14530;
assign w14788 = w14527 & w38442;
assign w14789 = ~w14787 & ~w14788;
assign w14790 = w14450 & ~w14789;
assign w14791 = ~w14789 & w38443;
assign w14792 = ~w14553 & ~w14603;
assign w14793 = w14546 & w14792;
assign w14794 = ~w14791 & w14793;
assign w14795 = w14786 & w14794;
assign w14796 = w14784 & w14795;
assign w14797 = w14758 & ~w14796;
assign w14798 = ~w14399 & w38444;
assign w14799 = w13916 & w14798;
assign w14800 = pi0341 & ~pi0342;
assign w14801 = pi0343 & ~w10746;
assign w14802 = ~w10746 & w38445;
assign w14803 = pi0343 & w14733;
assign w14804 = ~pi0343 & w14800;
assign w14805 = ~w14803 & ~w14804;
assign w14806 = ~pi2384 & ~w14374;
assign w14807 = w342 & w38446;
assign w14808 = ~w14806 & ~w14807;
assign w14809 = (w921 & w38447) | (w921 & w38448) | (w38447 & w38448);
assign w14810 = ~pi0409 & ~pi0426;
assign w14811 = w14810 & ~w923;
assign w14812 = (w342 & w38450) | (w342 & w38451) | (w38450 & w38451);
assign w14813 = w14808 & w14812;
assign w14814 = (w14813 & ~w7537) | (w14813 & w38452) | (~w7537 & w38452);
assign w14815 = (w921 & w38453) | (w921 & w38454) | (w38453 & w38454);
assign w14816 = ~w14815 & w40157;
assign w14817 = ~w5783 & ~w14816;
assign w14818 = (w921 & w38457) | (w921 & w38458) | (w38457 & w38458);
assign w14819 = pi0426 & w14400;
assign w14820 = (w14399 & w38459) | (w14399 & w38460) | (w38459 & w38460);
assign w14821 = ~w14818 & ~w14820;
assign w14822 = (~w5758 & w14820) | (~w5758 & w38461) | (w14820 & w38461);
assign w14823 = (w921 & w38462) | (w921 & w38463) | (w38462 & w38463);
assign w14824 = (w14399 & w38464) | (w14399 & w38465) | (w38464 & w38465);
assign w14825 = ~w14823 & ~w14824;
assign w14826 = (~w5767 & w14824) | (~w5767 & w38466) | (w14824 & w38466);
assign w14827 = ~w14822 & ~w14826;
assign w14828 = ~w14817 & w14827;
assign w14829 = ~w14802 & w38467;
assign w14830 = ~w14799 & w14829;
assign w14831 = ~w14797 & w38468;
assign w14832 = ~w14730 & w14831;
assign w14833 = ~w14421 & w14832;
assign w14834 = ~w14408 & w14833;
assign w14835 = w14833 & w38469;
assign w14836 = w14364 & ~w14812;
assign w14837 = ~pi0410 & pi0579;
assign w14838 = pi0410 & pi0597;
assign w14839 = w14810 & ~w14838;
assign w14840 = ~w14837 & w14839;
assign w14841 = w14740 & w14840;
assign w14842 = w14836 & w14841;
assign w14843 = pi0425 & pi0596;
assign w14844 = ~pi0425 & pi0580;
assign w14845 = ~pi0406 & ~w14844;
assign w14846 = ~w14843 & w14845;
assign w14847 = ~w14360 & w14846;
assign w14848 = w14740 & w14847;
assign w14849 = ~w343 & w14848;
assign w14850 = ~pi3344 & w14849;
assign w14851 = ~w14842 & ~w14850;
assign w14852 = ~pi3245 & ~w14851;
assign w14853 = w14852 & w40133;
assign w14854 = w14836 & w38470;
assign w14855 = ~w14849 & ~w14854;
assign w14856 = ~pi3245 & ~pi3344;
assign w14857 = w7537 & ~w14856;
assign w14858 = ~w14855 & w14857;
assign w14859 = w14363 & ~w14848;
assign w14860 = w14859 & w38471;
assign w14861 = w5713 & ~w14352;
assign w14862 = w5722 & w14352;
assign w14863 = ~w14861 & ~w14862;
assign w14864 = w14860 & w14863;
assign w14865 = pi0410 & ~w923;
assign w14866 = (w921 & w38472) | (w921 & w38473) | (w38472 & w38473);
assign w14867 = ~w14865 & ~w14866;
assign w14868 = w5699 & ~w14867;
assign w14869 = w5709 & w14867;
assign w14870 = ~w14841 & w38474;
assign w14871 = w14836 & w14870;
assign w14872 = w14352 & ~w14355;
assign w14873 = w14859 & w38475;
assign w14874 = pi0220 & pi0979;
assign w14875 = pi0222 & ~pi0979;
assign w14876 = ~w14874 & ~w14875;
assign w14877 = w14873 & w14876;
assign w14878 = ~w14871 & ~w14877;
assign w14879 = ~w14864 & w14878;
assign w14880 = ~w14858 & w14879;
assign w14881 = ~w14853 & w14880;
assign w14882 = w14808 & w38476;
assign w14883 = (~pi0055 & w14807) | (~pi0055 & w38477) | (w14807 & w38477);
assign w14884 = ~w14882 & ~w14883;
assign w14885 = (w14884 & w14881) | (w14884 & w38478) | (w14881 & w38478);
assign w14886 = ~w14835 & ~w14885;
assign w14887 = (w14374 & ~w342) | (w14374 & w38479) | (~w342 & w38479);
assign w14888 = (w921 & w38480) | (w921 & w38481) | (w38480 & w38481);
assign w14889 = ~w14887 & ~w14888;
assign w14890 = (~w14870 & ~w13916) | (~w14870 & w38482) | (~w13916 & w38482);
assign w14891 = ~w14887 & w38483;
assign w14892 = ~w14813 & ~w14891;
assign w14893 = (w14892 & w14890) | (w14892 & w38484) | (w14890 & w38484);
assign w14894 = ~w14834 & ~w14893;
assign w14895 = (w13946 & w14087) | (w13946 & w38485) | (w14087 & w38485);
assign w14896 = pi0057 & ~w13946;
assign w14897 = ~w14895 & ~w14896;
assign w14898 = pi0058 & w10759;
assign w14899 = (w10746 & w38486) | (w10746 & w38487) | (w38486 & w38487);
assign w14900 = ~w10752 & ~w14899;
assign w14901 = ~w14091 & w14099;
assign w14902 = w13730 & ~w13766;
assign w14903 = (~pi0868 & ~w13730) | (~pi0868 & w38488) | (~w13730 & w38488);
assign w14904 = pi0868 & ~w13737;
assign w14905 = ~w14903 & ~w14904;
assign w14906 = ~w14901 & w14905;
assign w14907 = ~w12505 & w13853;
assign w14908 = ~w13768 & w14903;
assign w14909 = ~w13765 & w14908;
assign w14910 = (w14909 & w14094) | (w14909 & w38489) | (w14094 & w38489);
assign w14911 = ~w13846 & w14910;
assign w14912 = ~w14907 & w14911;
assign w14913 = ~w14906 & ~w14912;
assign w14914 = (~w14899 & ~w14901) | (~w14899 & w38490) | (~w14901 & w38490);
assign w14915 = w14913 & w14914;
assign w14916 = ~w14900 & ~w14915;
assign w14917 = pi0059 & w13933;
assign w14918 = (w10746 & w38491) | (w10746 & w38492) | (w38491 & w38492);
assign w14919 = ~w13923 & ~w14918;
assign w14920 = (~w14918 & ~w14901) | (~w14918 & w38493) | (~w14901 & w38493);
assign w14921 = w14913 & w14920;
assign w14922 = ~w14919 & ~w14921;
assign w14923 = (w13946 & ~w14280) | (w13946 & w38494) | (~w14280 & w38494);
assign w14924 = w14286 & w14923;
assign w14925 = w14269 & w14924;
assign w14926 = ~pi0060 & ~w13946;
assign w14927 = ~w14925 & ~w14926;
assign w14928 = w13946 & ~w14322;
assign w14929 = pi0061 & ~w13946;
assign w14930 = ~w14928 & ~w14929;
assign w14931 = w13830 & ~w14142;
assign w14932 = w14223 & ~w14931;
assign w14933 = w13833 & ~w14932;
assign w14934 = (~w14933 & w13784) | (~w14933 & w38495) | (w13784 & w38495);
assign w14935 = ~w13846 & w14934;
assign w14936 = (w14224 & w13745) | (w14224 & w38496) | (w13745 & w38496);
assign w14937 = (~w14932 & w14936) | (~w14932 & w14933) | (w14936 & w14933);
assign w14938 = ~w14935 & w14937;
assign w14939 = w13852 & w38497;
assign w14940 = ~w12505 & w14939;
assign w14941 = ~w14938 & ~w14940;
assign w14942 = ~w13833 & w14932;
assign w14943 = (~pi0868 & ~w14932) | (~pi0868 & w38498) | (~w14932 & w38498);
assign w14944 = (~w14943 & w13784) | (~w14943 & w38499) | (w13784 & w38499);
assign w14945 = ~w13846 & w14944;
assign w14946 = (~pi0868 & w14936) | (~pi0868 & w38500) | (w14936 & w38500);
assign w14947 = ~w14945 & w14946;
assign w14948 = w13852 & w38501;
assign w14949 = ~w12505 & w14948;
assign w14950 = ~w14947 & ~w14949;
assign w14951 = w14941 & ~w14950;
assign w14952 = pi0868 & w14213;
assign w14953 = w14302 & w14952;
assign w14954 = ~w14298 & w14953;
assign w14955 = (pi0868 & w14275) | (pi0868 & w38502) | (w14275 & w38502);
assign w14956 = w14271 & w38818;
assign w14957 = ~w12505 & w14956;
assign w14958 = ~w14955 & ~w14957;
assign w14959 = ~w14954 & w14958;
assign w14960 = (w10752 & ~w14959) | (w10752 & w38503) | (~w14959 & w38503);
assign w14961 = (pi3245 & w7634) | (pi3245 & w38504) | (w7634 & w38504);
assign w14962 = (w6410 & w38507) | (w6410 & w38508) | (w38507 & w38508);
assign w14963 = (~pi0062 & ~w40209) | (~pi0062 & w38509) | (~w40209 & w38509);
assign w14964 = w10759 & ~w14963;
assign w14965 = (w14964 & w14962) | (w14964 & w38510) | (w14962 & w38510);
assign w14966 = w10756 & ~w14965;
assign w14967 = ~w14960 & ~w14966;
assign w14968 = (pi0868 & w13809) | (pi0868 & w38511) | (w13809 & w38511);
assign w14969 = w13835 & ~w14968;
assign w14970 = pi0868 & ~w14932;
assign w14971 = ~w14969 & ~w14970;
assign w14972 = ~w13807 & w38512;
assign w14973 = ~w13754 & w14972;
assign w14974 = ~w14971 & ~w14973;
assign w14975 = ~w13835 & ~w14968;
assign w14976 = ~w13807 & w38513;
assign w14977 = ~w13754 & w14976;
assign w14978 = pi0868 & w14936;
assign w14979 = ~w13847 & w14978;
assign w14980 = w13852 & w38514;
assign w14981 = ~w12505 & w14980;
assign w14982 = ~w14979 & ~w14981;
assign w14983 = ~w14977 & w14982;
assign w14984 = ~w14974 & w14983;
assign w14985 = (w10752 & w14941) | (w10752 & w38515) | (w14941 & w38515);
assign w14986 = ~w14984 & w14985;
assign w14987 = (pi3245 & w7601) | (pi3245 & w38516) | (w7601 & w38516);
assign w14988 = (~pi0063 & ~w40209) | (~pi0063 & w38520) | (~w40209 & w38520);
assign w14989 = w10759 & ~w14988;
assign w14990 = (w14989 & w40168) | (w14989 & w38521) | (w40168 & w38521);
assign w14991 = w10756 & ~w14990;
assign w14992 = ~w14986 & ~w14991;
assign w14993 = (w13923 & ~w14959) | (w13923 & w38522) | (~w14959 & w38522);
assign w14994 = (~pi0064 & ~w40144) | (~pi0064 & w38523) | (~w40144 & w38523);
assign w14995 = w13933 & ~w14994;
assign w14996 = (w14995 & w14962) | (w14995 & w38524) | (w14962 & w38524);
assign w14997 = w13930 & ~w14996;
assign w14998 = ~w14993 & ~w14997;
assign w14999 = (w13923 & w14941) | (w13923 & w38525) | (w14941 & w38525);
assign w15000 = ~w14984 & w14999;
assign w15001 = (w4379 & w38526) | (w4379 & w38527) | (w38526 & w38527);
assign w15002 = (~pi0065 & ~w40144) | (~pi0065 & w38528) | (~w40144 & w38528);
assign w15003 = w13933 & ~w15002;
assign w15004 = ~w15001 & w15003;
assign w15005 = w13930 & ~w15004;
assign w15006 = ~w15000 & ~w15005;
assign w15007 = (~w10099 & w10352) | (~w10099 & w38529) | (w10352 & w38529);
assign w15008 = w10312 & w10593;
assign w15009 = (~w10594 & ~w10311) | (~w10594 & w38530) | (~w10311 & w38530);
assign w15010 = ~w10345 & w15009;
assign w15011 = ~w15008 & ~w15010;
assign w15012 = ~w15007 & w15011;
assign w15013 = w15007 & ~w15011;
assign w15014 = ~w15012 & ~w15013;
assign w15015 = w14410 & w15014;
assign w15016 = w14539 & ~w14716;
assign w15017 = w14597 & w15016;
assign w15018 = w14521 & ~w14608;
assign w15019 = w14559 & ~w14622;
assign w15020 = ~w15018 & ~w15019;
assign w15021 = (~w15020 & ~w14615) | (~w15020 & w38531) | (~w14615 & w38531);
assign w15022 = w14559 & ~w14687;
assign w15023 = ~w10221 & w38532;
assign w15024 = ~w15022 & ~w15023;
assign w15025 = ~w14669 & ~w15024;
assign w15026 = ~w14720 & ~w15025;
assign w15027 = w14521 & ~w14648;
assign w15028 = ~w14636 & w38533;
assign w15029 = ~w15027 & ~w15028;
assign w15030 = ~w14658 & ~w15029;
assign w15031 = ~w14520 & ~w14712;
assign w15032 = (w14709 & ~w15031) | (w14709 & w38534) | (~w15031 & w38534);
assign w15033 = ~w15030 & ~w15032;
assign w15034 = w15026 & w15033;
assign w15035 = w14521 & ~w14619;
assign w15036 = w14559 & w14675;
assign w15037 = ~w15035 & ~w15036;
assign w15038 = ~w14627 & ~w15037;
assign w15039 = w14559 & ~w14697;
assign w15040 = w14521 & ~w14633;
assign w15041 = ~w15039 & ~w15040;
assign w15042 = ~w14631 & ~w15041;
assign w15043 = w14559 & ~w14664;
assign w15044 = ~w10152 & w38535;
assign w15045 = ~w15043 & ~w15044;
assign w15046 = ~w14680 & ~w15045;
assign w15047 = ~w15042 & ~w15046;
assign w15048 = ~w15038 & w15047;
assign w15049 = w14559 & ~w14651;
assign w15050 = ~w14424 & w14521;
assign w15051 = ~w15049 & ~w15050;
assign w15052 = ~w14643 & ~w15051;
assign w15053 = pi3516 & ~w4661;
assign w15054 = w14521 & ~w14684;
assign w15055 = w14559 & w14702;
assign w15056 = ~w15054 & ~w15055;
assign w15057 = w14586 & w38536;
assign w15058 = ~w15053 & ~w15057;
assign w15059 = ~w15052 & w15058;
assign w15060 = w14604 & w15059;
assign w15061 = w15048 & w15060;
assign w15062 = w15061 & w38537;
assign w15063 = w15017 & w15062;
assign w15064 = ~w15063 & w38538;
assign w15065 = (~w14731 & w4748) | (~w14731 & w38539) | (w4748 & w38539);
assign w15066 = (w14745 & w14738) | (w14745 & w38540) | (w14738 & w38540);
assign w15067 = ~w4695 & ~w14752;
assign w15068 = ~w4689 & ~w14749;
assign w15069 = ~w15067 & ~w15068;
assign w15070 = (w14735 & ~w15069) | (w14735 & w38541) | (~w15069 & w38541);
assign w15071 = ~w14734 & ~w15070;
assign w15072 = ~w15065 & ~w15071;
assign w15073 = w14450 & ~w14633;
assign w15074 = w14564 & w15073;
assign w15075 = ~w14591 & ~w14765;
assign w15076 = pi3516 & ~w4657;
assign w15077 = ~w14587 & ~w15076;
assign w15078 = w15077 & w38542;
assign w15079 = w14793 & w15078;
assign w15080 = w14710 & ~w15024;
assign w15081 = (~w15037 & w14583) | (~w15037 & w38543) | (w14583 & w38543);
assign w15082 = ~w15080 & ~w15081;
assign w15083 = w14490 & ~w15082;
assign w15084 = w14583 & w38544;
assign w15085 = ~w14581 & w38545;
assign w15086 = ~w15045 & w15085;
assign w15087 = ~w15084 & ~w15086;
assign w15088 = w14583 & w38546;
assign w15089 = ~w14581 & w38547;
assign w15090 = w15039 & w15089;
assign w15091 = w14711 & ~w15029;
assign w15092 = ~w15090 & ~w15091;
assign w15093 = ~w15088 & w15092;
assign w15094 = w15087 & w15093;
assign w15095 = (w14453 & ~w15094) | (w14453 & w38548) | (~w15094 & w38548);
assign w15096 = w14790 & ~w15056;
assign w15097 = ~w15095 & ~w15096;
assign w15098 = (w14758 & ~w15097) | (w14758 & w38549) | (~w15097 & w38549);
assign w15099 = w14798 & w40159;
assign w15100 = (w14813 & w10746) | (w14813 & w38550) | (w10746 & w38550);
assign w15101 = ~w7504 & w38551;
assign w15102 = (~w4661 & w14824) | (~w4661 & w38552) | (w14824 & w38552);
assign w15103 = ~w15101 & ~w15102;
assign w15104 = (~w4657 & w14820) | (~w4657 & w38553) | (w14820 & w38553);
assign w15105 = ~w4721 & ~w14816;
assign w15106 = ~w15104 & ~w15105;
assign w15107 = w15103 & w15106;
assign w15108 = w15100 & w15107;
assign w15109 = ~w15099 & w15108;
assign w15110 = ~w15098 & w15109;
assign w15111 = ~w15072 & w15110;
assign w15112 = ~w15064 & w15111;
assign w15113 = ~w15015 & w15112;
assign w15114 = ~w14408 & w15113;
assign w15115 = w15113 & w38469;
assign w15116 = ~w7504 & w38554;
assign w15117 = ~w14855 & w15116;
assign w15118 = pi0214 & ~pi0979;
assign w15119 = pi0213 & pi0979;
assign w15120 = ~w15118 & ~w15119;
assign w15121 = w14873 & w15120;
assign w15122 = w4704 & ~w14867;
assign w15123 = w4699 & w14867;
assign w15124 = ~w14841 & w38555;
assign w15125 = w14836 & w15124;
assign w15126 = w4681 & ~w14352;
assign w15127 = w4708 & w14352;
assign w15128 = ~w15126 & ~w15127;
assign w15129 = w14860 & w15128;
assign w15130 = ~w15125 & ~w15129;
assign w15131 = ~w15121 & w15130;
assign w15132 = ~w15117 & w15131;
assign w15133 = ~w14806 & ~w15132;
assign w15134 = (pi0066 & w14807) | (pi0066 & w38557) | (w14807 & w38557);
assign w15135 = ~w14882 & ~w15134;
assign w15136 = (w15135 & w4748) | (w15135 & w38558) | (w4748 & w38558);
assign w15137 = ~w15133 & w15136;
assign w15138 = ~w15115 & ~w15137;
assign w15139 = w14841 & w40159;
assign w15140 = pi0067 & w14889;
assign w15141 = ~w14813 & ~w15140;
assign w15142 = w15141 & w40160;
assign w15143 = ~w15114 & ~w15142;
assign w15144 = ~w13509 & ~w13755;
assign w15145 = (~w13179 & w13778) | (~w13179 & w38560) | (w13778 & w38560);
assign w15146 = ~w13509 & w13521;
assign w15147 = (w15146 & w13806) | (w15146 & w40085) | (w13806 & w40085);
assign w15148 = w13183 & ~w13192;
assign w15149 = w15146 & w15148;
assign w15150 = ~w12505 & w15149;
assign w15151 = ~w15147 & ~w15150;
assign w15152 = (~w13757 & w13778) | (~w13757 & w38562) | (w13778 & w38562);
assign w15153 = pi0868 & ~w13522;
assign w15154 = (w15153 & w13806) | (w15153 & w38563) | (w13806 & w38563);
assign w15155 = w15148 & w15153;
assign w15156 = ~w12505 & w15155;
assign w15157 = ~w15154 & ~w15156;
assign w15158 = w15151 & ~w15157;
assign w15159 = (~w15144 & w13806) | (~w15144 & w38564) | (w13806 & w38564);
assign w15160 = ~w15144 & w15148;
assign w15161 = ~w12505 & w15160;
assign w15162 = ~w15159 & ~w15161;
assign w15163 = ~pi0868 & w15148;
assign w15164 = ~w12505 & w15163;
assign w15165 = (~pi0868 & w13806) | (~pi0868 & w40086) | (w13806 & w40086);
assign w15166 = ~w15164 & ~w15165;
assign w15167 = w15162 & ~w15166;
assign w15168 = ~w15158 & ~w15167;
assign w15169 = w10752 & ~w15168;
assign w15170 = (pi3245 & w7795) | (pi3245 & w38565) | (w7795 & w38565);
assign w15171 = ~w15170 & w40161;
assign w15172 = ~pi0051 & w40140;
assign w15173 = (~w15172 & ~w10751) | (~w15172 & w38569) | (~w10751 & w38569);
assign w15174 = pi0068 & w10759;
assign w15175 = w15173 & ~w15174;
assign w15176 = (w15175 & ~w15171) | (w15175 & w38570) | (~w15171 & w38570);
assign w15177 = ~w15169 & ~w15176;
assign w15178 = w13923 & w15168;
assign w15179 = (w5052 & w38571) | (w5052 & w38572) | (w38571 & w38572);
assign w15180 = ~pi0069 & w13933;
assign w15181 = w13927 & ~w15180;
assign w15182 = ~w15179 & w15181;
assign w15183 = ~w15178 & ~w15182;
assign w15184 = ~w10613 & w38573;
assign w15185 = w10750 & w15184;
assign w15186 = ~w15168 & w15185;
assign w15187 = (pi0070 & ~w15184) | (pi0070 & w38574) | (~w15184 & w38574);
assign w15188 = ~w15186 & ~w15187;
assign w15189 = w13922 & w15184;
assign w15190 = ~w15168 & w15189;
assign w15191 = (pi0071 & ~w15184) | (pi0071 & w38575) | (~w15184 & w38575);
assign w15192 = ~w15190 & ~w15191;
assign w15193 = ~pi1743 & ~pi1866;
assign w15194 = ~pi1897 & w15193;
assign w15195 = ~pi1741 & ~pi1867;
assign w15196 = ~pi0314 & ~pi0330;
assign w15197 = ~pi0073 & ~pi0128;
assign w15198 = ~pi0127 & w15197;
assign w15199 = w15197 & w38576;
assign w15200 = w15196 & w15199;
assign w15201 = w15199 & w38577;
assign w15202 = w15195 & w15201;
assign w15203 = w15201 & w38579;
assign w15204 = (w15203 & w38581) | (w15203 & w38582) | (w38581 & w38582);
assign w15205 = pi1743 & pi1866;
assign w15206 = pi1897 & w15205;
assign w15207 = (w15203 & w38585) | (w15203 & w38586) | (w38585 & w38586);
assign w15208 = ~pi1017 & pi1897;
assign w15209 = pi1714 & w15208;
assign w15210 = ~pi1017 & ~pi1897;
assign w15211 = ~pi1714 & w15210;
assign w15212 = ~w15209 & ~w15211;
assign w15213 = (pi1897 & ~w15199) | (pi1897 & w38587) | (~w15199 & w38587);
assign w15214 = ~pi0368 & w15213;
assign w15215 = pi0368 & ~w15213;
assign w15216 = ~w15214 & ~w15215;
assign w15217 = ~pi1017 & ~w15216;
assign w15218 = ~pi0127 & ~pi1897;
assign w15219 = ~pi0073 & ~pi1017;
assign w15220 = ~w15218 & ~w15219;
assign w15221 = pi0127 & pi1897;
assign w15222 = ~pi0072 & ~w15221;
assign w15223 = ~w15220 & w15222;
assign w15224 = (~pi1017 & w15223) | (~pi1017 & w15210) | (w15223 & w15210);
assign w15225 = pi0128 & w15224;
assign w15226 = pi1017 & pi1897;
assign w15227 = ~w15197 & w15226;
assign w15228 = pi0073 & ~pi1017;
assign w15229 = pi0128 & w15228;
assign w15230 = (pi0072 & w15229) | (pi0072 & w38588) | (w15229 & w38588);
assign w15231 = (pi0127 & w15230) | (pi0127 & w38589) | (w15230 & w38589);
assign w15232 = ~pi1897 & ~w15231;
assign w15233 = w15225 & ~w15232;
assign w15234 = pi1897 & ~w15199;
assign w15235 = (w15234 & ~w15224) | (w15234 & w38591) | (~w15224 & w38591);
assign w15236 = (w15233 & w38592) | (w15233 & w38593) | (w38592 & w38593);
assign w15237 = pi0314 & pi1897;
assign w15238 = ~w15236 & w15237;
assign w15239 = ~pi0314 & ~pi1897;
assign w15240 = (w15233 & w38595) | (w15233 & w38596) | (w38595 & w38596);
assign w15241 = ~w15238 & w38597;
assign w15242 = pi1897 & w15195;
assign w15243 = pi1741 & pi1867;
assign w15244 = ~w15242 & w40162;
assign w15245 = ~pi1017 & pi1742;
assign w15246 = pi1017 & pi1741;
assign w15247 = ~w15245 & ~w15246;
assign w15248 = pi1897 & ~w15247;
assign w15249 = ~pi1897 & w15247;
assign w15250 = w15241 & w38600;
assign w15251 = (pi1897 & ~w15201) | (pi1897 & w38601) | (~w15201 & w38601);
assign w15252 = ~pi1745 & w15251;
assign w15253 = pi1745 & ~w15251;
assign w15254 = ~w15252 & ~w15253;
assign w15255 = w15241 & w38602;
assign w15256 = (w15241 & w38604) | (w15241 & w38605) | (w38604 & w38605);
assign w15257 = pi1714 & pi1744;
assign w15258 = ~pi1714 & ~pi1744;
assign w15259 = (~w15258 & w15203) | (~w15258 & w38606) | (w15203 & w38606);
assign w15260 = pi1744 & w40163;
assign w15261 = ~w15204 & ~w15260;
assign w15262 = (~w15261 & ~w15256) | (~w15261 & w38609) | (~w15256 & w38609);
assign w15263 = ~w15207 & w15262;
assign w15264 = w15201 & w38610;
assign w15265 = ~w15212 & ~w15264;
assign w15266 = (w15265 & ~w15241) | (w15265 & w38611) | (~w15241 & w38611);
assign w15267 = ~pi1714 & ~pi1745;
assign w15268 = ~pi1017 & pi1745;
assign w15269 = pi1714 & w15268;
assign w15270 = ~w15267 & ~w15269;
assign w15271 = ~w15269 & w38612;
assign w15272 = w15254 & ~w15271;
assign w15273 = w15268 & w38580;
assign w15274 = (w15273 & ~w15241) | (w15273 & w38613) | (~w15241 & w38613);
assign w15275 = ~w15272 & ~w15274;
assign w15276 = ~w15266 & w15275;
assign w15277 = w15263 & ~w15276;
assign w15278 = w15193 & w38581;
assign w15279 = (w15203 & w38614) | (w15203 & w38615) | (w38614 & w38615);
assign w15280 = (~w15207 & ~w15256) | (~w15207 & w38616) | (~w15256 & w38616);
assign w15281 = ~w15210 & ~w15268;
assign w15282 = (~w15281 & w15251) | (~w15281 & w38617) | (w15251 & w38617);
assign w15283 = ~pi1742 & ~w15268;
assign w15284 = (w15201 & w38619) | (w15201 & w38620) | (w38619 & w38620);
assign w15285 = ~w15251 & w15284;
assign w15286 = ~w15282 & ~w15285;
assign w15287 = pi1742 & w15226;
assign w15288 = (w15287 & ~w15201) | (w15287 & w38622) | (~w15201 & w38622);
assign w15289 = (w15241 & w38623) | (w15241 & w38624) | (w38623 & w38624);
assign w15290 = w15202 & ~w15245;
assign w15291 = pi1017 & ~pi1867;
assign w15292 = ~w15195 & ~w15291;
assign w15293 = w15201 & ~w15292;
assign w15294 = (~w15249 & w15293) | (~w15249 & w38625) | (w15293 & w38625);
assign w15295 = ~w15290 & w15294;
assign w15296 = (~w15295 & ~w15241) | (~w15295 & w38626) | (~w15241 & w38626);
assign w15297 = ~w15250 & ~w15296;
assign w15298 = ~w15289 & w15297;
assign w15299 = w15280 & ~w15298;
assign w15300 = w15277 & ~w15299;
assign w15301 = ~w15255 & w15289;
assign w15302 = ~w15298 & w38627;
assign w15303 = w15277 & w15302;
assign w15304 = ~w15195 & ~w15243;
assign w15305 = w15241 & ~w15304;
assign w15306 = ~pi1017 & ~pi1741;
assign w15307 = (~w15306 & w15201) | (~w15306 & w38628) | (w15201 & w38628);
assign w15308 = ~pi1741 & w15208;
assign w15309 = ~w15291 & ~w15308;
assign w15310 = ~w15307 & w15309;
assign w15311 = pi1897 & ~w15243;
assign w15312 = ~w15208 & ~w15291;
assign w15313 = ~w15311 & ~w15312;
assign w15314 = ~w15293 & ~w15313;
assign w15315 = (w15314 & w15241) | (w15314 & w38629) | (w15241 & w38629);
assign w15316 = ~w15305 & w15315;
assign w15317 = w15280 & ~w15316;
assign w15318 = pi1017 & w15216;
assign w15319 = (w15233 & w38630) | (w15233 & w38631) | (w38630 & w38631);
assign w15320 = ~w15238 & w38632;
assign w15321 = (~pi1867 & w15238) | (~pi1867 & w38633) | (w15238 & w38633);
assign w15322 = ~pi1017 & ~w15321;
assign w15323 = (~w15318 & ~w15322) | (~w15318 & w38634) | (~w15322 & w38634);
assign w15324 = w15317 & ~w15323;
assign w15325 = w15303 & ~w15324;
assign w15326 = ~w15300 & ~w15325;
assign w15327 = (~w15217 & w15238) | (~w15217 & w38635) | (w15238 & w38635);
assign w15328 = ~w15241 & ~w15327;
assign w15329 = ~w15323 & w15328;
assign w15330 = w15317 & ~w15329;
assign w15331 = w15303 & ~w15330;
assign w15332 = (~pi1017 & ~w15233) | (~pi1017 & w38636) | (~w15233 & w38636);
assign w15333 = ~pi0330 & ~w15233;
assign w15334 = w15332 & ~w15333;
assign w15335 = ~w15234 & w15334;
assign w15336 = pi0072 & pi1017;
assign w15337 = (~w15336 & w15334) | (~w15336 & w38637) | (w15334 & w38637);
assign w15338 = ~w15335 & w15337;
assign w15339 = pi0072 & w15226;
assign w15340 = ~w15198 & w15339;
assign w15341 = ~w15338 & ~w15340;
assign w15342 = w15280 & w15341;
assign w15343 = (w15342 & ~w15303) | (w15342 & w38638) | (~w15303 & w38638);
assign w15344 = (w15223 & w38639) | (w15223 & w38640) | (w38639 & w38640);
assign w15345 = pi0314 & w15210;
assign w15346 = ~w15199 & w38641;
assign w15347 = ~w15345 & w40164;
assign w15348 = ~w15233 & ~w15347;
assign w15349 = ~pi0314 & w15208;
assign w15350 = ~w15236 & ~w15349;
assign w15351 = ~w15348 & w15350;
assign w15352 = ~w15344 & ~w15351;
assign w15353 = w15280 & ~w15352;
assign w15354 = w15303 & w38644;
assign w15355 = ~w15343 & ~w15354;
assign w15356 = w15326 & ~w15355;
assign w15357 = w15241 & w38645;
assign w15358 = pi1017 & w15254;
assign w15359 = (~w15273 & ~w15203) | (~w15273 & w38646) | (~w15203 & w38646);
assign w15360 = ~w15358 & w15359;
assign w15361 = (w15241 & w38647) | (w15241 & w38648) | (w38647 & w38648);
assign w15362 = ~w15357 & w15361;
assign w15363 = w15263 & w15362;
assign w15364 = ~w15300 & ~w15363;
assign w15365 = (w15317 & w15300) | (w15317 & w15432) | (w15300 & w15432);
assign w15366 = ~w15302 & ~w15365;
assign w15367 = w15317 & ~w15328;
assign w15368 = w15280 & ~w15323;
assign w15369 = ~w15367 & ~w15368;
assign w15370 = w15303 & w15369;
assign w15371 = ~w15366 & ~w15370;
assign w15372 = ~w15356 & w15371;
assign w15373 = w15280 & w15301;
assign w15374 = (~w15362 & ~w15373) | (~w15362 & w38649) | (~w15373 & w38649);
assign w15375 = ~w15372 & w15374;
assign w15376 = w15303 & w15317;
assign w15377 = ~w15300 & w38650;
assign w15378 = w15318 & ~w15377;
assign w15379 = w15376 & w15378;
assign w15380 = (w15263 & ~w15378) | (w15263 & w38651) | (~w15378 & w38651);
assign w15381 = w15276 & w15301;
assign w15382 = w15380 & ~w15381;
assign w15383 = ~w15262 & w15280;
assign w15384 = ~w15362 & w15383;
assign w15385 = w15378 & w38652;
assign w15386 = ~w15384 & ~w15385;
assign w15387 = (w15386 & w15375) | (w15386 & w38653) | (w15375 & w38653);
assign w15388 = (~pi3427 & ~w6668) | (~pi3427 & w38654) | (~w6668 & w38654);
assign w15389 = w5320 & ~w15388;
assign w15390 = (w6668 & w38657) | (w6668 & w38658) | (w38657 & w38658);
assign w15391 = pi1017 & pi2555;
assign w15392 = (~w15391 & w15389) | (~w15391 & w38659) | (w15389 & w38659);
assign w15393 = ~w15387 & w15392;
assign w15394 = ~pi1017 & pi2555;
assign w15395 = (~w15394 & w15389) | (~w15394 & w38660) | (w15389 & w38660);
assign w15396 = w15387 & w15395;
assign w15397 = ~w15393 & ~w15396;
assign w15398 = ~w15297 & w15383;
assign w15399 = (pi1017 & w15198) | (pi1017 & w38661) | (w15198 & w38661);
assign w15400 = pi0072 & pi0073;
assign w15401 = w15208 & w15400;
assign w15402 = ~pi0072 & ~pi0128;
assign w15403 = w15210 & w15402;
assign w15404 = ~w15401 & ~w15403;
assign w15405 = ~w15223 & w15404;
assign w15406 = ~w15399 & w15405;
assign w15407 = ~w15231 & w15406;
assign w15408 = (~w15398 & ~w15303) | (~w15398 & w38663) | (~w15303 & w38663);
assign w15409 = w15379 & w15408;
assign w15410 = w15280 & w15328;
assign w15411 = w15300 & ~w15410;
assign w15412 = ~w15303 & ~w15411;
assign w15413 = w15325 & w15355;
assign w15414 = pi0127 & ~pi1017;
assign w15415 = ~w15226 & ~w15414;
assign w15416 = pi0128 & ~w15415;
assign w15417 = ~pi0073 & ~w15414;
assign w15418 = ~w15416 & w15417;
assign w15419 = ~pi0128 & w15218;
assign w15420 = (~pi1017 & w15419) | (~pi1017 & w38664) | (w15419 & w38664);
assign w15421 = ~w15416 & ~w15420;
assign w15422 = pi0073 & ~w15421;
assign w15423 = ~w15418 & ~w15422;
assign w15424 = w15423 & w15280;
assign w15425 = (~w15424 & ~w15303) | (~w15424 & w38665) | (~w15303 & w38665);
assign w15426 = ~w15331 & w15425;
assign w15427 = w15299 & ~w15426;
assign w15428 = ~w15413 & w15427;
assign w15429 = ~w15412 & ~w15428;
assign w15430 = ~w15329 & ~w15398;
assign w15431 = (w15430 & w15377) | (w15430 & w38666) | (w15377 & w38666);
assign w15432 = w15317 & w15363;
assign w15433 = w15277 & w15373;
assign w15434 = w15277 & w38667;
assign w15435 = ~w15432 & ~w15434;
assign w15436 = (w15435 & w15431) | (w15435 & w38668) | (w15431 & w38668);
assign w15437 = (~w15409 & w15429) | (~w15409 & w38669) | (w15429 & w38669);
assign w15438 = w4749 & ~w15388;
assign w15439 = (w6668 & w38672) | (w6668 & w38673) | (w38672 & w38673);
assign w15440 = (~w15391 & w15438) | (~w15391 & w38674) | (w15438 & w38674);
assign w15441 = w15437 & ~w15440;
assign w15442 = (~w15394 & w15438) | (~w15394 & w38675) | (w15438 & w38675);
assign w15443 = ~w15437 & ~w15442;
assign w15444 = ~w15441 & ~w15443;
assign w15445 = ~w10379 & w38676;
assign w15446 = ~w10393 & ~w15445;
assign w15447 = (w10397 & ~w10360) | (w10397 & w38677) | (~w10360 & w38677);
assign w15448 = ~w10605 & ~w15447;
assign w15449 = ~w15446 & w40165;
assign w15450 = ~w10400 & ~w10594;
assign w15451 = w15450 & w40166;
assign w15452 = ~w15449 & ~w15451;
assign w15453 = w14410 & ~w15452;
assign w15454 = w14610 & w38680;
assign w15455 = ~w14599 & ~w15454;
assign w15456 = ~w14599 & w38681;
assign w15457 = ~w14499 & w14657;
assign w15458 = w14495 & w38682;
assign w15459 = ~w14720 & w38683;
assign w15460 = ~w15457 & w15459;
assign w15461 = w14597 & w15460;
assign w15462 = w14597 & w38684;
assign w15463 = w14495 & w38685;
assign w15464 = ~w14487 & w15463;
assign w15465 = w14539 & w38686;
assign w15466 = w15462 & w15465;
assign w15467 = (~w14653 & ~w14615) | (~w14653 & w38687) | (~w14615 & w38687);
assign w15468 = ~w14680 & ~w14763;
assign w15469 = w14526 & w15089;
assign w15470 = pi3516 & ~w3396;
assign w15471 = (~w15470 & ~w15469) | (~w15470 & w38688) | (~w15469 & w38688);
assign w15472 = w14526 & w14711;
assign w15473 = ~w14689 & w15472;
assign w15474 = w14704 & w38689;
assign w15475 = ~w15473 & ~w15474;
assign w15476 = w15471 & w15475;
assign w15477 = ~w15468 & w15476;
assign w15478 = ~w14627 & ~w14638;
assign w15479 = w14454 & w38690;
assign w15480 = ~w14633 & w15479;
assign w15481 = ~w15478 & ~w15480;
assign w15482 = ~w14624 & ~w14669;
assign w15483 = w14521 & w14675;
assign w15484 = ~w14673 & ~w15483;
assign w15485 = w14586 & w38691;
assign w15486 = ~w14522 & ~w14640;
assign w15487 = w14610 & w38692;
assign w15488 = w14495 & w38693;
assign w15489 = ~w15487 & ~w15488;
assign w15490 = ~w15485 & w15489;
assign w15491 = ~w15482 & w15490;
assign w15492 = w15477 & w38694;
assign w15493 = ~w15467 & w15492;
assign w15494 = (~pi0709 & ~w15466) | (~pi0709 & w38695) | (~w15466 & w38695);
assign w15495 = w14422 & w15494;
assign w15496 = (w3412 & w38696) | (w3412 & w38697) | (w38696 & w38697);
assign w15497 = (w14745 & w14749) | (w14745 & w38698) | (w14749 & w38698);
assign w15498 = ~w3350 & ~w14752;
assign w15499 = ~w3354 & ~w14738;
assign w15500 = ~w15498 & ~w15499;
assign w15501 = (w14735 & ~w15500) | (w14735 & w38699) | (~w15500 & w38699);
assign w15502 = ~w14734 & ~w15501;
assign w15503 = ~w15496 & ~w15502;
assign w15504 = w14785 & w38700;
assign w15505 = w14556 & w15504;
assign w15506 = w14792 & w15505;
assign w15507 = ~w14789 & ~w15484;
assign w15508 = ~w14658 & ~w14689;
assign w15509 = ~w14638 & w14714;
assign w15510 = w14710 & w14713;
assign w15511 = ~w14624 & w15510;
assign w15512 = w14577 & w15089;
assign w15513 = ~w14424 & w15512;
assign w15514 = ~w15511 & ~w15513;
assign w15515 = ~w15509 & w15514;
assign w15516 = w15515 & w38701;
assign w15517 = w14709 & w14712;
assign w15518 = w14557 & w38702;
assign w15519 = ~w14565 & ~w15518;
assign w15520 = ~w15517 & w15519;
assign w15521 = ~w14643 & ~w14666;
assign w15522 = ~w14631 & w14772;
assign w15523 = w14760 & w38703;
assign w15524 = w14453 & w15085;
assign w15525 = pi3516 & ~w3387;
assign w15526 = (~w15525 & ~w15524) | (~w15525 & w38704) | (~w15524 & w38704);
assign w15527 = ~w15523 & w15526;
assign w15528 = ~w15522 & w15527;
assign w15529 = ~w15521 & w15528;
assign w15530 = w15520 & w15529;
assign w15531 = w15516 & w15530;
assign w15532 = (w14758 & ~w15531) | (w14758 & w38705) | (~w15531 & w38705);
assign w15533 = w14325 & w14798;
assign w15534 = ~w7667 & w38706;
assign w15535 = (~w3387 & w14820) | (~w3387 & w38707) | (w14820 & w38707);
assign w15536 = ~w15534 & ~w15535;
assign w15537 = (~w3396 & w14824) | (~w3396 & w38708) | (w14824 & w38708);
assign w15538 = ~w3367 & ~w14816;
assign w15539 = ~w15537 & ~w15538;
assign w15540 = w15536 & w15539;
assign w15541 = w15100 & w15540;
assign w15542 = ~w15533 & w15541;
assign w15543 = ~w15532 & w38709;
assign w15544 = ~w15495 & w15543;
assign w15545 = ~w15453 & w15544;
assign w15546 = ~w14408 & w15545;
assign w15547 = w15545 & w38469;
assign w15548 = w14852 & w40134;
assign w15549 = ~w7667 & w38710;
assign w15550 = ~w14855 & w15549;
assign w15551 = w3331 & ~w14352;
assign w15552 = w3327 & w14352;
assign w15553 = ~w15551 & ~w15552;
assign w15554 = w14860 & w15553;
assign w15555 = w3345 & ~w14867;
assign w15556 = w3341 & w14867;
assign w15557 = ~w14841 & w38711;
assign w15558 = w14836 & w15557;
assign w15559 = pi0132 & pi0979;
assign w15560 = pi0133 & ~pi0979;
assign w15561 = ~w15559 & ~w15560;
assign w15562 = w14873 & w15561;
assign w15563 = ~w15558 & ~w15562;
assign w15564 = ~w15554 & w15563;
assign w15565 = ~w15550 & w15564;
assign w15566 = ~w15548 & w15565;
assign w15567 = (~pi0074 & w14807) | (~pi0074 & w38712) | (w14807 & w38712);
assign w15568 = ~w14882 & ~w15567;
assign w15569 = (w15568 & w15566) | (w15568 & w38713) | (w15566 & w38713);
assign w15570 = ~w15547 & ~w15569;
assign w15571 = w10394 & ~w10593;
assign w15572 = (w10594 & ~w10160) | (w10594 & w38715) | (~w10160 & w38715);
assign w15573 = ~w10174 & ~w15572;
assign w15574 = ~w15571 & w15573;
assign w15575 = (w10360 & w38716) | (w10360 & w38717) | (w38716 & w38717);
assign w15576 = w15574 & w40167;
assign w15577 = ~w15575 & ~w15576;
assign w15578 = w14410 & ~w15577;
assign w15579 = (~w15029 & ~w14615) | (~w15029 & w38718) | (~w14615 & w38718);
assign w15580 = (~w15479 & w14627) | (~w15479 & w38719) | (w14627 & w38719);
assign w15581 = w14698 & ~w15580;
assign w15582 = ~w14631 & ~w15051;
assign w15583 = ~w14627 & w15040;
assign w15584 = ~w14680 & ~w15020;
assign w15585 = ~w15583 & ~w15584;
assign w15586 = ~w15582 & w15585;
assign w15587 = ~w14669 & ~w15037;
assign w15588 = ~w14485 & w38720;
assign w15589 = w14586 & w38721;
assign w15590 = ~w15045 & w15589;
assign w15591 = w14704 & w38722;
assign w15592 = pi3516 & ~w6304;
assign w15593 = (~w15592 & ~w15472) | (~w15592 & w38723) | (~w15472 & w38723);
assign w15594 = ~w15591 & w15593;
assign w15595 = ~w15590 & w15594;
assign w15596 = ~w15587 & w15595;
assign w15597 = w15586 & w15596;
assign w15598 = w15597 & w38724;
assign w15599 = w15016 & w15598;
assign w15600 = (~pi0709 & ~w15599) | (~pi0709 & w38725) | (~w15599 & w38725);
assign w15601 = w14422 & w15600;
assign w15602 = ~w14731 & ~w6413;
assign w15603 = (w14745 & w14752) | (w14745 & w38726) | (w14752 & w38726);
assign w15604 = ~w6320 & ~w14738;
assign w15605 = ~w6316 & ~w14749;
assign w15606 = ~w15604 & ~w15605;
assign w15607 = (w14735 & ~w15606) | (w14735 & w38727) | (~w15606 & w38727);
assign w15608 = ~w14734 & ~w15607;
assign w15609 = ~w15602 & ~w15608;
assign w15610 = ~w14789 & w38728;
assign w15611 = ~w14643 & ~w15024;
assign w15612 = ~w14603 & ~w15611;
assign w15613 = w14710 & ~w15020;
assign w15614 = w14583 & ~w15029;
assign w15615 = ~w15613 & ~w15614;
assign w15616 = w14534 & ~w15615;
assign w15617 = w14583 & w38729;
assign w15618 = w15049 & w15089;
assign w15619 = ~w15617 & ~w15618;
assign w15620 = (w14453 & w15616) | (w14453 & w38730) | (w15616 & w38730);
assign w15621 = ~w14424 & w14450;
assign w15622 = w14564 & w15621;
assign w15623 = ~w15620 & ~w15622;
assign w15624 = w15612 & w15623;
assign w15625 = ~w14658 & ~w15056;
assign w15626 = ~w15037 & w15510;
assign w15627 = pi3516 & ~w6308;
assign w15628 = (~w15627 & ~w14712) | (~w15627 & w38731) | (~w14712 & w38731);
assign w15629 = ~w15518 & w15628;
assign w15630 = ~w15626 & w15629;
assign w15631 = ~w15625 & w15630;
assign w15632 = w15624 & w38732;
assign w15633 = (w14758 & ~w15632) | (w14758 & w38733) | (~w15632 & w38733);
assign w15634 = w14798 & w14962;
assign w15635 = ~w7634 & w38734;
assign w15636 = ~w6270 & ~w14816;
assign w15637 = ~w15635 & ~w15636;
assign w15638 = (~w6304 & w14824) | (~w6304 & w38735) | (w14824 & w38735);
assign w15639 = (~w6308 & w14820) | (~w6308 & w38736) | (w14820 & w38736);
assign w15640 = ~w15638 & ~w15639;
assign w15641 = w15637 & w15640;
assign w15642 = w15100 & w15641;
assign w15643 = ~w15634 & w15642;
assign w15644 = ~w15633 & w38737;
assign w15645 = ~w15601 & w15644;
assign w15646 = ~w15578 & w15645;
assign w15647 = ~w14408 & w15646;
assign w15648 = w15646 & w38469;
assign w15649 = ~w7634 & w38738;
assign w15650 = ~w14855 & w15649;
assign w15651 = pi0195 & ~pi0979;
assign w15652 = pi0194 & pi0979;
assign w15653 = ~w15651 & ~w15652;
assign w15654 = w14873 & w15653;
assign w15655 = w6339 & ~w14867;
assign w15656 = w6334 & w14867;
assign w15657 = ~w14841 & w38739;
assign w15658 = w14836 & w15657;
assign w15659 = w6324 & ~w14352;
assign w15660 = w6343 & w14352;
assign w15661 = ~w15659 & ~w15660;
assign w15662 = w14860 & w15661;
assign w15663 = ~w15658 & ~w15662;
assign w15664 = ~w15654 & w15663;
assign w15665 = ~w15650 & w15664;
assign w15666 = ~w14806 & ~w15665;
assign w15667 = (w6410 & w38740) | (w6410 & w38741) | (w38740 & w38741);
assign w15668 = (~pi0075 & w14807) | (~pi0075 & w38742) | (w14807 & w38742);
assign w15669 = ~w14882 & ~w15668;
assign w15670 = ~w15667 & w15669;
assign w15671 = ~w15666 & w15670;
assign w15672 = ~w15648 & ~w15671;
assign w15673 = (~w10099 & w10355) | (~w10099 & w38743) | (w10355 & w38743);
assign w15674 = ~w10210 & ~w10395;
assign w15675 = (w15674 & w15673) | (w15674 & w38744) | (w15673 & w38744);
assign w15676 = w10209 & w10593;
assign w15677 = ~w15674 & ~w15676;
assign w15678 = ~w15673 & w15677;
assign w15679 = ~w15675 & ~w15678;
assign w15680 = w14410 & w15679;
assign w15681 = (~w14638 & ~w14615) | (~w14638 & w38745) | (~w14615 & w38745);
assign w15682 = ~w14627 & ~w14763;
assign w15683 = pi3516 & ~w4323;
assign w15684 = w14704 & w38402;
assign w15685 = ~w15684 & w38746;
assign w15686 = ~w15682 & w15685;
assign w15687 = ~w14624 & ~w14680;
assign w15688 = ~w14631 & ~w14653;
assign w15689 = ~w15687 & ~w15688;
assign w15690 = w15686 & w15689;
assign w15691 = ~w14669 & ~w15484;
assign w15692 = ~w14658 & ~w15486;
assign w15693 = (w14662 & w14583) | (w14662 & w38747) | (w14583 & w38747);
assign w15694 = w14710 & w14772;
assign w15695 = ~w15693 & ~w15694;
assign w15696 = w14527 & ~w15695;
assign w15697 = w14586 & w38748;
assign w15698 = ~w15454 & ~w15697;
assign w15699 = ~w15696 & w15698;
assign w15700 = w15699 & w38749;
assign w15701 = w15690 & w15700;
assign w15702 = w15701 & w38750;
assign w15703 = w14606 & w15702;
assign w15704 = ~w15703 & w38538;
assign w15705 = (~w14731 & w4379) | (~w14731 & w38751) | (w4379 & w38751);
assign w15706 = (w14745 & w14738) | (w14745 & w38752) | (w14738 & w38752);
assign w15707 = ~w4339 & ~w14752;
assign w15708 = ~w4366 & ~w14749;
assign w15709 = ~w15707 & ~w15708;
assign w15710 = (w14735 & ~w15709) | (w14735 & w38753) | (~w15709 & w38753);
assign w15711 = ~w14734 & ~w15710;
assign w15712 = ~w15705 & ~w15711;
assign w15713 = ~w14658 & w14772;
assign w15714 = w14450 & ~w14622;
assign w15715 = w14454 & w38754;
assign w15716 = ~w14561 & ~w15715;
assign w15717 = w15714 & ~w15716;
assign w15718 = w14714 & ~w14763;
assign w15719 = ~w15518 & ~w15718;
assign w15720 = ~w14677 & w15510;
assign w15721 = ~w14648 & w15512;
assign w15722 = ~w15720 & ~w15721;
assign w15723 = w15719 & w15722;
assign w15724 = w15723 & w38755;
assign w15725 = ~w14666 & w14790;
assign w15726 = w14450 & ~w14651;
assign w15727 = w14564 & w15726;
assign w15728 = ~w14643 & ~w14689;
assign w15729 = pi3516 & ~w4331;
assign w15730 = (~w15729 & ~w15524) | (~w15729 & w38756) | (~w15524 & w38756);
assign w15731 = ~w14638 & w14761;
assign w15732 = w14640 & w14712;
assign w15733 = ~w15731 & w38757;
assign w15734 = w15733 & w38758;
assign w15735 = ~w15725 & w15734;
assign w15736 = w15724 & w15735;
assign w15737 = (w14758 & ~w15736) | (w14758 & w38705) | (~w15736 & w38705);
assign w15738 = w14798 & w40168;
assign w15739 = ~w7601 & w38759;
assign w15740 = (~w4323 & w14824) | (~w4323 & w38760) | (w14824 & w38760);
assign w15741 = ~w15739 & ~w15740;
assign w15742 = ~w4293 & ~w14816;
assign w15743 = (~w4331 & w14820) | (~w4331 & w38761) | (w14820 & w38761);
assign w15744 = ~w15742 & ~w15743;
assign w15745 = w15741 & w15744;
assign w15746 = w15100 & w15745;
assign w15747 = ~w15738 & w15746;
assign w15748 = ~w15737 & w38762;
assign w15749 = ~w15704 & w15748;
assign w15750 = ~w15680 & w15749;
assign w15751 = ~w14408 & w15750;
assign w15752 = w15750 & w38469;
assign w15753 = ~w4379 & w38763;
assign w15754 = ~w7601 & w38764;
assign w15755 = ~w14855 & w15754;
assign w15756 = pi0187 & pi0979;
assign w15757 = pi0188 & ~pi0979;
assign w15758 = ~w15756 & ~w15757;
assign w15759 = w14873 & w15758;
assign w15760 = w4347 & ~w14867;
assign w15761 = w4343 & w14867;
assign w15762 = ~w14841 & w38765;
assign w15763 = w14836 & w15762;
assign w15764 = w4353 & ~w14352;
assign w15765 = w4362 & w14352;
assign w15766 = ~w15764 & ~w15765;
assign w15767 = w14860 & w15766;
assign w15768 = ~w15763 & ~w15767;
assign w15769 = ~w15759 & w15768;
assign w15770 = ~w15755 & w15769;
assign w15771 = (~w14806 & w15753) | (~w14806 & w38766) | (w15753 & w38766);
assign w15772 = ~pi0076 & ~w14808;
assign w15773 = ~w14882 & ~w15772;
assign w15774 = ~w15771 & w15773;
assign w15775 = ~w15752 & ~w15774;
assign w15776 = ~w10603 & w38767;
assign w15777 = w14405 & w15776;
assign w15778 = ~w14407 & ~w15777;
assign w15779 = w14401 & w15778;
assign w15780 = w14495 & w38768;
assign w15781 = ~w14598 & ~w15780;
assign w15782 = w14610 & w38769;
assign w15783 = w15781 & ~w15782;
assign w15784 = ~w14630 & ~w15524;
assign w15785 = (~w15715 & w15784) | (~w15715 & w38770) | (w15784 & w38770);
assign w15786 = w15783 & w15785;
assign w15787 = ~w14499 & ~w15786;
assign w15788 = ~w14493 & w14500;
assign w15789 = ~w14700 & ~w15788;
assign w15790 = ~w14716 & w15789;
assign w15791 = ~w14611 & ~w14629;
assign w15792 = w14550 & ~w15791;
assign w15793 = ~w14603 & ~w15792;
assign w15794 = w15790 & w15793;
assign w15795 = w14590 & ~w15464;
assign w15796 = w15795 & w38771;
assign w15797 = w15794 & w15796;
assign w15798 = ~w15787 & w15797;
assign w15799 = w14518 & w14556;
assign w15800 = w14529 & w15459;
assign w15801 = w14495 & w14559;
assign w15802 = ~w14667 & ~w15801;
assign w15803 = ~w14568 & ~w15802;
assign w15804 = w14521 & w14531;
assign w15805 = ~w14519 & ~w14572;
assign w15806 = ~w15804 & w15805;
assign w15807 = w14656 & ~w15806;
assign w15808 = ~w15803 & ~w15807;
assign w15809 = ~w14499 & ~w15808;
assign w15810 = w14495 & w38772;
assign w15811 = ~w14542 & ~w15810;
assign w15812 = w14594 & w15811;
assign w15813 = ~w15457 & w15812;
assign w15814 = w14550 & w14613;
assign w15815 = ~w14494 & ~w15454;
assign w15816 = ~w15814 & w15815;
assign w15817 = w14537 & w15816;
assign w15818 = w15813 & w15817;
assign w15819 = w15818 & w38773;
assign w15820 = w15799 & w15819;
assign w15821 = w14583 & w38774;
assign w15822 = w14490 & ~w15056;
assign w15823 = w14534 & ~w15024;
assign w15824 = w14524 & ~w15041;
assign w15825 = ~w15823 & ~w15824;
assign w15826 = (w14710 & ~w15825) | (w14710 & w38775) | (~w15825 & w38775);
assign w15827 = w14583 & w38776;
assign w15828 = ~w15826 & w38777;
assign w15829 = w14504 & ~w15615;
assign w15830 = w14586 & ~w15051;
assign w15831 = ~w15829 & ~w15830;
assign w15832 = (w14526 & ~w15831) | (w14526 & w38778) | (~w15831 & w38778);
assign w15833 = pi3516 & ~w8195;
assign w15834 = (~w15833 & w14669) | (~w15833 & w38779) | (w14669 & w38779);
assign w15835 = ~w15832 & w15834;
assign w15836 = w15820 & w38780;
assign w15837 = ~w15836 & w38538;
assign w15838 = w14556 & w38365;
assign w15839 = (~w15037 & ~w14615) | (~w15037 & w38781) | (~w14615 & w38781);
assign w15840 = ~w14523 & ~w14536;
assign w15841 = ~w15032 & w15840;
assign w15842 = ~w14680 & ~w15024;
assign w15843 = ~w14627 & ~w15045;
assign w15844 = ~w15842 & ~w15843;
assign w15845 = ~w14631 & ~w15020;
assign w15846 = ~w14643 & ~w15029;
assign w15847 = ~w15845 & ~w15846;
assign w15848 = w15844 & w15847;
assign w15849 = w14522 & w15510;
assign w15850 = pi3516 & ~w8203;
assign w15851 = w14491 & w14511;
assign w15852 = ~w14588 & ~w15851;
assign w15853 = (~w15850 & w15852) | (~w15850 & w38782) | (w15852 & w38782);
assign w15854 = ~w15849 & w15853;
assign w15855 = w14594 & w15854;
assign w15856 = w14604 & w15855;
assign w15857 = w15848 & w15856;
assign w15858 = w15841 & w15857;
assign w15859 = w14575 & w38783;
assign w15860 = ~w14669 & ~w15056;
assign w15861 = ~w14789 & ~w15051;
assign w15862 = ~w14658 & ~w15041;
assign w15863 = ~w15861 & ~w15862;
assign w15864 = ~w15860 & w15863;
assign w15865 = w15859 & w15864;
assign w15866 = w15858 & w38784;
assign w15867 = (w14758 & ~w15866) | (w14758 & w38785) | (~w15866 & w38785);
assign w15868 = w14735 & w40169;
assign w15869 = ~w1143 & ~w14749;
assign w15870 = ~w14399 & w38787;
assign w15871 = w1143 & ~w14390;
assign w15872 = (w10747 & w1143) | (w10747 & w38309) | (w1143 & w38309);
assign w15873 = ~w15871 & w15872;
assign w15874 = (~pi0343 & w14399) | (~pi0343 & w38789) | (w14399 & w38789);
assign w15875 = ~w15869 & w15874;
assign w15876 = ~w8157 & ~w14752;
assign w15877 = ~w8172 & ~w14738;
assign w15878 = ~w15876 & ~w15877;
assign w15879 = w15875 & w15878;
assign w15880 = w15868 & ~w15879;
assign w15881 = ~w7699 & w38790;
assign w15882 = (~w15881 & w10746) | (~w15881 & w38791) | (w10746 & w38791);
assign w15883 = ~w8220 & ~w14816;
assign w15884 = ~w10746 & w14798;
assign w15885 = ~w8239 & w38792;
assign w15886 = ~w8265 & w38793;
assign w15887 = w14813 & ~w15886;
assign w15888 = ~w15885 & w15887;
assign w15889 = ~w15884 & w15888;
assign w15890 = (~w8195 & w14824) | (~w8195 & w38794) | (w14824 & w38794);
assign w15891 = (~w8203 & w14820) | (~w8203 & w38795) | (w14820 & w38795);
assign w15892 = ~w15890 & ~w15891;
assign w15893 = w15889 & w38796;
assign w15894 = w15893 & w38797;
assign w15895 = ~w15867 & w15894;
assign w15896 = ~w15837 & w15895;
assign w15897 = w14364 & w15896;
assign w15898 = ~w15779 & w15897;
assign w15899 = ~w8265 & w38798;
assign w15900 = ~w14855 & w15899;
assign w15901 = w8163 & ~w14352;
assign w15902 = w8149 & w14352;
assign w15903 = ~w15901 & ~w15902;
assign w15904 = w14860 & w15903;
assign w15905 = w8168 & ~w14867;
assign w15906 = w8153 & w14867;
assign w15907 = ~w14841 & w38799;
assign w15908 = w14836 & w15907;
assign w15909 = pi0089 & pi0979;
assign w15910 = pi0092 & ~pi0979;
assign w15911 = ~w15909 & ~w15910;
assign w15912 = w14873 & w15911;
assign w15913 = ~w15908 & ~w15912;
assign w15914 = ~w15904 & w15913;
assign w15915 = ~w15900 & w15914;
assign w15916 = ~w14806 & ~w15915;
assign w15917 = ~pi0077 & ~w14808;
assign w15918 = ~w14882 & ~w15917;
assign w15919 = (w15918 & w8239) | (w15918 & w38801) | (w8239 & w38801);
assign w15920 = ~w15916 & w15919;
assign w15921 = ~w15898 & ~w15920;
assign w15922 = ~w14887 & w38802;
assign w15923 = ~w14889 & ~w15557;
assign w15924 = (w15923 & ~w14325) | (w15923 & w38803) | (~w14325 & w38803);
assign w15925 = (~w14813 & w15924) | (~w14813 & w38804) | (w15924 & w38804);
assign w15926 = ~w15546 & ~w15925;
assign w15927 = ~w14887 & w38805;
assign w15928 = ~w14889 & ~w15657;
assign w15929 = (w15928 & ~w14962) | (w15928 & w38806) | (~w14962 & w38806);
assign w15930 = (~w14813 & w15929) | (~w14813 & w38807) | (w15929 & w38807);
assign w15931 = ~w15647 & ~w15930;
assign w15932 = w14841 & w40168;
assign w15933 = pi0080 & w14889;
assign w15934 = ~w14813 & ~w15933;
assign w15935 = w15934 & w40170;
assign w15936 = ~w15751 & ~w15935;
assign w15937 = (w15896 & ~w15778) | (w15896 & w38809) | (~w15778 & w38809);
assign w15938 = (~w15907 & w10746) | (~w15907 & w38810) | (w10746 & w38810);
assign w15939 = ~w14887 & w38811;
assign w15940 = ~w14813 & ~w15939;
assign w15941 = (w15940 & w15938) | (w15940 & w38812) | (w15938 & w38812);
assign w15942 = ~w15937 & ~w15941;
assign w15943 = ~pi0082 & ~w13946;
assign w15944 = (w13946 & w14941) | (w13946 & w38210) | (w14941 & w38210);
assign w15945 = ~w14984 & w15944;
assign w15946 = ~w15943 & ~w15945;
assign w15947 = pi0083 & ~w13946;
assign w15948 = w14959 & w38813;
assign w15949 = ~w15947 & ~w15948;
assign w15950 = pi0084 & ~w13946;
assign w15951 = (w13946 & ~w14901) | (w13946 & w38814) | (~w14901 & w38814);
assign w15952 = w14913 & w15951;
assign w15953 = ~w15950 & ~w15952;
assign w15954 = ~pi0868 & ~w13522;
assign w15955 = (w15954 & w13806) | (w15954 & w38815) | (w13806 & w38815);
assign w15956 = w15148 & w15954;
assign w15957 = ~w12505 & w15956;
assign w15958 = ~w15955 & ~w15957;
assign w15959 = w15151 & ~w15958;
assign w15960 = ~w13522 & ~w13537;
assign w15961 = w15148 & w15960;
assign w15962 = ~w12505 & w15961;
assign w15963 = (w15960 & w13806) | (w15960 & w38816) | (w13806 & w38816);
assign w15964 = pi0868 & ~w13532;
assign w15965 = ~w15963 & w15964;
assign w15966 = ~w15962 & w15965;
assign w15967 = (w13539 & w13806) | (w13539 & w38817) | (w13806 & w38817);
assign w15968 = pi0868 & w15967;
assign w15969 = ~w13192 & w13539;
assign w15970 = w13183 & w15969;
assign w15971 = w15969 & w38818;
assign w15972 = ~w12505 & w15971;
assign w15973 = ~w15968 & ~w15972;
assign w15974 = ~w15966 & w15973;
assign w15975 = ~w15959 & w15974;
assign w15976 = w10752 & ~w15975;
assign w15977 = (pi3245 & w7827) | (pi3245 & w38819) | (w7827 & w38819);
assign w15978 = (w5632 & w38822) | (w5632 & w38823) | (w38822 & w38823);
assign w15979 = pi0085 & w10759;
assign w15980 = w15173 & ~w15979;
assign w15981 = (w15980 & ~w15978) | (w15980 & w38824) | (~w15978 & w38824);
assign w15982 = ~w15976 & ~w15981;
assign w15983 = (~w11624 & w11508) | (~w11624 & w38825) | (w11508 & w38825);
assign w15984 = ~w11776 & w12088;
assign w15985 = ~w15983 & w15984;
assign w15986 = w15983 & ~w15984;
assign w15987 = ~w15985 & ~w15986;
assign w15988 = ~pi0868 & ~w15987;
assign w15989 = (w11777 & w11508) | (w11777 & w38826) | (w11508 & w38826);
assign w15990 = w12088 & ~w15989;
assign w15991 = ~w12034 & ~w12089;
assign w15992 = ~w15989 & w38827;
assign w15993 = (~w15991 & w15989) | (~w15991 & w38828) | (w15989 & w38828);
assign w15994 = ~w15992 & ~w15993;
assign w15995 = pi0868 & ~w15994;
assign w15996 = ~w15988 & ~w15995;
assign w15997 = pi0868 & w15987;
assign w15998 = (w11634 & ~w11507) | (w11634 & w38829) | (~w11507 & w38829);
assign w15999 = ~w11626 & ~w15998;
assign w16000 = ~w11636 & ~w15999;
assign w16001 = ~pi0868 & w16000;
assign w16002 = ~w15997 & ~w16001;
assign w16003 = ~w11401 & w11506;
assign w16004 = w11502 & w11634;
assign w16005 = ~w16003 & w16004;
assign w16006 = w16003 & ~w16004;
assign w16007 = ~w16005 & ~w16006;
assign w16008 = ~pi0868 & ~w16007;
assign w16009 = pi0868 & ~w16000;
assign w16010 = ~w16008 & ~w16009;
assign w16011 = ~w11298 & w11400;
assign w16012 = ~w11401 & ~w16011;
assign w16013 = ~pi0868 & w16012;
assign w16014 = (~w16013 & ~w16007) | (~w16013 & w38830) | (~w16007 & w38830);
assign w16015 = (~w11290 & w11294) | (~w11290 & w38831) | (w11294 & w38831);
assign w16016 = ~w11289 & w16015;
assign w16017 = w11289 & ~w16015;
assign w16018 = ~w16016 & ~w16017;
assign w16019 = ~pi0868 & w16018;
assign w16020 = (w11290 & w11288) | (w11290 & w38832) | (w11288 & w38832);
assign w16021 = ~w11297 & w38833;
assign w16022 = (~w11082 & w11297) | (~w11082 & w38834) | (w11297 & w38834);
assign w16023 = ~w16021 & ~w16022;
assign w16024 = pi0868 & ~w16023;
assign w16025 = ~w16019 & ~w16024;
assign w16026 = pi0868 & ~w16012;
assign w16027 = ~pi0868 & ~w16023;
assign w16028 = ~w11283 & w11287;
assign w16029 = ~w11288 & ~w16028;
assign w16030 = ~pi0868 & w16029;
assign w16031 = (~w16030 & w16018) | (~w16030 & w38835) | (w16018 & w38835);
assign w16032 = pi0868 & ~w16029;
assign w16033 = ~w11275 & w11279;
assign w16034 = ~w11181 & ~w11280;
assign w16035 = ~w16033 & w16034;
assign w16036 = w16033 & ~w16034;
assign w16037 = ~w16035 & ~w16036;
assign w16038 = ~pi0868 & ~w16037;
assign w16039 = ~w16032 & ~w16038;
assign w16040 = ~w11265 & w11274;
assign w16041 = ~w11275 & ~w16040;
assign w16042 = ~pi0868 & ~w16041;
assign w16043 = (~w16042 & w16037) | (~w16042 & w38836) | (w16037 & w38836);
assign w16044 = w11253 & w11264;
assign w16045 = ~w11265 & ~w16044;
assign w16046 = ~pi0868 & w16045;
assign w16047 = (~w16046 & ~w16041) | (~w16046 & w38837) | (~w16041 & w38837);
assign w16048 = pi0868 & w16045;
assign w16049 = ~w11215 & ~w11251;
assign w16050 = ~w11252 & ~w16049;
assign w16051 = ~pi0868 & w16050;
assign w16052 = ~w11240 & ~w11247;
assign w16053 = ~w11248 & ~w16052;
assign w16054 = ~pi0868 & ~w16053;
assign w16055 = (~w16054 & ~w16050) | (~w16054 & w38838) | (~w16050 & w38838);
assign w16056 = ~w11224 & w11235;
assign w16057 = ~w11236 & ~w16056;
assign w16058 = ~pi0868 & w16057;
assign w16059 = (~w16058 & w16053) | (~w16058 & w38839) | (w16053 & w38839);
assign w16060 = w10774 & ~w11216;
assign w16061 = ~w4685 & w16060;
assign w16062 = ~pi0868 & ~w16061;
assign w16063 = ~w11217 & w16062;
assign w16064 = (~w16063 & w16057) | (~w16063 & w38840) | (w16057 & w38840);
assign w16065 = ~pi0868 & pi1472;
assign w16066 = ~w16060 & ~w16065;
assign w16067 = ~w3631 & ~w16066;
assign w16068 = ~w11221 & ~w16067;
assign w16069 = ~pi1789 & ~pi1932;
assign w16070 = w16068 & w16069;
assign w16071 = w16070 & ~w16064;
assign w16072 = w16059 & w16071;
assign w16073 = w16072 & w16055;
assign w16074 = ~w16048 & w38841;
assign w16075 = w16047 & w16074;
assign w16076 = ~w16043 & w16075;
assign w16077 = ~w16039 & w16076;
assign w16078 = w16031 & w16077;
assign w16079 = (w16078 & w16026) | (w16078 & w38842) | (w16026 & w38842);
assign w16080 = ~w16025 & w16079;
assign w16081 = w16014 & w16080;
assign w16082 = ~w16010 & w16081;
assign w16083 = w16002 & w16082;
assign w16084 = ~w15996 & w16083;
assign w16085 = w10749 & w40171;
assign w16086 = pi0086 & w10759;
assign w16087 = w15173 & ~w16086;
assign w16088 = ~w16085 & w16087;
assign w16089 = (~w10752 & w16085) | (~w10752 & w38843) | (w16085 & w38843);
assign w16090 = ~pi0868 & ~w15994;
assign w16091 = w12064 & w38844;
assign w16092 = (~w12034 & ~w12064) | (~w12034 & w38845) | (~w12064 & w38845);
assign w16093 = (w16092 & w15989) | (w16092 & w38846) | (w15989 & w38846);
assign w16094 = ~w16091 & ~w16093;
assign w16095 = w12064 & w38847;
assign w16096 = ~w15990 & w16095;
assign w16097 = ~w16094 & ~w16096;
assign w16098 = ~w16090 & w16097;
assign w16099 = ~w16089 & ~w16098;
assign w16100 = w16084 & w16099;
assign w16101 = (~pi0868 & w15990) | (~pi0868 & w38848) | (w15990 & w38848);
assign w16102 = ~w16094 & w16101;
assign w16103 = ~w12502 & ~w13187;
assign w16104 = ~w12037 & w38849;
assign w16105 = (~w16103 & w12037) | (~w16103 & w38850) | (w12037 & w38850);
assign w16106 = ~w16104 & ~w16105;
assign w16107 = pi0868 & w16106;
assign w16108 = ~w16107 & w38851;
assign w16109 = ~w16088 & ~w16108;
assign w16110 = ~w16100 & w16109;
assign w16111 = w13923 & w15975;
assign w16112 = w13929 & ~w15978;
assign w16113 = ~pi0087 & w13933;
assign w16114 = w13927 & ~w16113;
assign w16115 = ~w16112 & w16114;
assign w16116 = ~w16111 & ~w16115;
assign w16117 = w13929 & w40171;
assign w16118 = pi0088 & w13933;
assign w16119 = w14336 & ~w16118;
assign w16120 = ~w16117 & w16119;
assign w16121 = (~w13923 & w16117) | (~w13923 & w38852) | (w16117 & w38852);
assign w16122 = ~w16098 & ~w16121;
assign w16123 = w16084 & w16122;
assign w16124 = ~w16107 & w38853;
assign w16125 = ~w16120 & ~w16124;
assign w16126 = ~w16123 & w16125;
assign w16127 = (~pi0089 & ~w15184) | (~pi0089 & w38854) | (~w15184 & w38854);
assign w16128 = (w15185 & ~w14901) | (w15185 & w38855) | (~w14901 & w38855);
assign w16129 = w14913 & w16128;
assign w16130 = ~w16127 & ~w16129;
assign w16131 = w15185 & ~w15975;
assign w16132 = (pi0090 & ~w15184) | (pi0090 & w38856) | (~w15184 & w38856);
assign w16133 = ~w16131 & ~w16132;
assign w16134 = (~pi0091 & ~w15184) | (~pi0091 & w38857) | (~w15184 & w38857);
assign w16135 = (w15185 & w16107) | (w15185 & w38858) | (w16107 & w38858);
assign w16136 = ~w16134 & ~w16135;
assign w16137 = ~w16098 & ~w16134;
assign w16138 = w16084 & w16137;
assign w16139 = ~w16136 & ~w16138;
assign w16140 = (~pi0092 & ~w15184) | (~pi0092 & w38859) | (~w15184 & w38859);
assign w16141 = (w15189 & ~w14901) | (w15189 & w38860) | (~w14901 & w38860);
assign w16142 = w14913 & w16141;
assign w16143 = ~w16140 & ~w16142;
assign w16144 = w15189 & ~w15975;
assign w16145 = (pi0093 & ~w15184) | (pi0093 & w38861) | (~w15184 & w38861);
assign w16146 = ~w16144 & ~w16145;
assign w16147 = (~pi0094 & ~w15184) | (~pi0094 & w38862) | (~w15184 & w38862);
assign w16148 = (w15189 & w16107) | (w15189 & w38863) | (w16107 & w38863);
assign w16149 = ~w16147 & ~w16148;
assign w16150 = ~w16098 & ~w16147;
assign w16151 = w16084 & w16150;
assign w16152 = ~w16149 & ~w16151;
assign w16153 = w10461 & w38865;
assign w16154 = (~w10594 & w10461) | (~w10594 & w38866) | (w10461 & w38866);
assign w16155 = ~w10546 & ~w16154;
assign w16156 = ~w16153 & ~w16155;
assign w16157 = (w10402 & w38867) | (w10402 & w38868) | (w38867 & w38868);
assign w16158 = w16156 & w40172;
assign w16159 = ~w16157 & ~w16158;
assign w16160 = w14410 & ~w16159;
assign w16161 = (w14640 & ~w14615) | (w14640 & w38869) | (~w14615 & w38869);
assign w16162 = w14522 & ~w15791;
assign w16163 = w14487 & w15463;
assign w16164 = ~w15814 & ~w16163;
assign w16165 = ~w16162 & w16164;
assign w16166 = w15455 & w16165;
assign w16167 = w14450 & ~w14648;
assign w16168 = ~w15580 & w16167;
assign w16169 = ~w14624 & w15589;
assign w16170 = ~w14638 & ~w14680;
assign w16171 = ~w16169 & ~w16170;
assign w16172 = ~w14627 & w14652;
assign w16173 = w14610 & w38870;
assign w16174 = w14487 & w16173;
assign w16175 = ~w16172 & ~w16174;
assign w16176 = w16171 & w16175;
assign w16177 = ~w14669 & ~w14763;
assign w16178 = w14704 & w38691;
assign w16179 = ~w14689 & w15469;
assign w16180 = ~w14666 & w15472;
assign w16181 = ~w16179 & ~w16180;
assign w16182 = ~w16178 & w16181;
assign w16183 = w14526 & w14583;
assign w16184 = w14469 & w14772;
assign w16185 = pi3516 & ~w6087;
assign w16186 = (~w16185 & ~w16183) | (~w16185 & w38871) | (~w16183 & w38871);
assign w16187 = ~w14700 & w16186;
assign w16188 = w16182 & w38872;
assign w16189 = w16176 & w16188;
assign w16190 = w16189 & w38873;
assign w16191 = ~w16161 & w16190;
assign w16192 = w16191 & w38874;
assign w16193 = ~w16192 & w38538;
assign w16194 = w15519 & w38875;
assign w16195 = w15505 & w16194;
assign w16196 = w15505 & w38876;
assign w16197 = ~w14658 & ~w14666;
assign w16198 = w14649 & w14714;
assign w16199 = ~w14763 & w15510;
assign w16200 = ~w14558 & ~w16199;
assign w16201 = ~w16198 & w16200;
assign w16202 = ~w16197 & w16201;
assign w16203 = ~w14624 & ~w14789;
assign w16204 = w14714 & w15726;
assign w16205 = ~w14536 & ~w16204;
assign w16206 = ~w14559 & ~w16205;
assign w16207 = ~w16203 & ~w16206;
assign w16208 = w16202 & w16207;
assign w16209 = ~w14614 & w38877;
assign w16210 = ~w14631 & ~w14689;
assign w16211 = ~w14643 & ~w15484;
assign w16212 = w14760 & w38878;
assign w16213 = pi3516 & ~w6091;
assign w16214 = (~w16213 & ~w15524) | (~w16213 & w38879) | (~w15524 & w38879);
assign w16215 = ~w16212 & w16214;
assign w16216 = ~w16211 & w16215;
assign w16217 = w16216 & w38880;
assign w16218 = w16208 & w16217;
assign w16219 = (w14758 & ~w16218) | (w14758 & w38881) | (~w16218 & w38881);
assign w16220 = (w14745 & w14749) | (w14745 & w38882) | (w14749 & w38882);
assign w16221 = ~w6060 & ~w14752;
assign w16222 = ~w6056 & ~w14738;
assign w16223 = ~w16221 & ~w16222;
assign w16224 = w16220 & w16223;
assign w16225 = w15868 & ~w16224;
assign w16226 = pi3245 & ~w7732;
assign w16227 = w14798 & w40191;
assign w16228 = ~w6111 & ~w14816;
assign w16229 = (~w6087 & w14824) | (~w6087 & w38887) | (w14824 & w38887);
assign w16230 = ~w16228 & ~w16229;
assign w16231 = (w16230 & w6176) | (w16230 & w38888) | (w6176 & w38888);
assign w16232 = ~w6091 & ~w14821;
assign w16233 = w7732 & w14803;
assign w16234 = ~w16232 & ~w16233;
assign w16235 = w15882 & w16234;
assign w16236 = w16231 & w16235;
assign w16237 = w16236 & w38889;
assign w16238 = ~w16219 & w16237;
assign w16239 = ~w16193 & w16238;
assign w16240 = ~w16160 & w16239;
assign w16241 = (w14882 & ~w16240) | (w14882 & w38890) | (~w16240 & w38890);
assign w16242 = ~w6176 & w38891;
assign w16243 = w7732 & ~w14856;
assign w16244 = ~w14855 & w16243;
assign w16245 = w6079 & ~w14352;
assign w16246 = w6075 & w14352;
assign w16247 = ~w16245 & ~w16246;
assign w16248 = w14860 & w16247;
assign w16249 = w6064 & ~w14867;
assign w16250 = w6070 & w14867;
assign w16251 = ~w14841 & w38892;
assign w16252 = w14836 & w16251;
assign w16253 = pi0147 & pi0979;
assign w16254 = pi0148 & ~pi0979;
assign w16255 = ~w16253 & ~w16254;
assign w16256 = w14873 & w16255;
assign w16257 = ~w16252 & ~w16256;
assign w16258 = ~w16248 & w16257;
assign w16259 = ~w16244 & w16258;
assign w16260 = (~w14806 & w16242) | (~w14806 & w38893) | (w16242 & w38893);
assign w16261 = ~pi0095 & ~w14808;
assign w16262 = ~w16260 & ~w16261;
assign w16263 = ~w16241 & w16262;
assign w16264 = w10126 & w38894;
assign w16265 = (~w10594 & ~w10126) | (~w10594 & w38895) | (~w10126 & w38895);
assign w16266 = ~w10399 & w16265;
assign w16267 = ~w16264 & ~w16266;
assign w16268 = (~w10099 & w10379) | (~w10099 & w38896) | (w10379 & w38896);
assign w16269 = (w10360 & w38897) | (w10360 & w38898) | (w38897 & w38898);
assign w16270 = ~w16267 & w16269;
assign w16271 = w16267 & ~w16269;
assign w16272 = ~w16270 & ~w16271;
assign w16273 = w14410 & w16272;
assign w16274 = w14538 & w38899;
assign w16275 = ~w14616 & ~w15051;
assign w16276 = w14770 & ~w15580;
assign w16277 = w14704 & w38900;
assign w16278 = pi3516 & ~w3108;
assign w16279 = (~w16278 & ~w15469) | (~w16278 & w38901) | (~w15469 & w38901);
assign w16280 = ~w16277 & w16279;
assign w16281 = ~w14716 & w16280;
assign w16282 = ~w14627 & w15027;
assign w16283 = ~w14680 & ~w15041;
assign w16284 = ~w16282 & ~w16283;
assign w16285 = w16281 & w16284;
assign w16286 = ~w14669 & ~w15020;
assign w16287 = w14527 & ~w15082;
assign w16288 = ~w14494 & ~w16173;
assign w16289 = ~w16287 & w16288;
assign w16290 = ~w16286 & w16289;
assign w16291 = w16285 & w16290;
assign w16292 = w16291 & w38902;
assign w16293 = w16274 & w16292;
assign w16294 = (~pi0709 & ~w16293) | (~pi0709 & w38725) | (~w16293 & w38725);
assign w16295 = w14422 & w16294;
assign w16296 = ~w14789 & w38903;
assign w16297 = ~w14658 & ~w15024;
assign w16298 = ~w14643 & ~w15045;
assign w16299 = ~w14631 & ~w15056;
assign w16300 = pi3516 & ~w3112;
assign w16301 = (~w16300 & ~w15524) | (~w16300 & w38904) | (~w15524 & w38904);
assign w16302 = w14761 & ~w15051;
assign w16303 = w14713 & ~w15615;
assign w16304 = ~w16302 & ~w16303;
assign w16305 = w16304 & w38905;
assign w16306 = w16305 & w38906;
assign w16307 = ~w16296 & w16306;
assign w16308 = (w14758 & ~w16307) | (w14758 & w38881) | (~w16307 & w38881);
assign w16309 = ~w3060 & ~w14738;
assign w16310 = ~w3075 & ~w14752;
assign w16311 = ~w16309 & ~w16310;
assign w16312 = w16220 & w16311;
assign w16313 = w15868 & ~w16312;
assign w16314 = w14798 & w40174;
assign w16315 = ~w3083 & ~w14816;
assign w16316 = (~w3112 & w14820) | (~w3112 & w38908) | (w14820 & w38908);
assign w16317 = ~w16315 & ~w16316;
assign w16318 = (w16317 & w3194) | (w16317 & w38909) | (w3194 & w38909);
assign w16319 = ~w3108 & ~w14825;
assign w16320 = ~w7699 & w38910;
assign w16321 = ~w16319 & ~w16320;
assign w16322 = w15100 & w16321;
assign w16323 = w16322 & w38911;
assign w16324 = ~w16313 & w16323;
assign w16325 = ~w16308 & w16324;
assign w16326 = ~w16295 & w16325;
assign w16327 = ~w16273 & w16326;
assign w16328 = ~w14408 & w16327;
assign w16329 = w16327 & w38469;
assign w16330 = ~w3194 & w38912;
assign w16331 = ~w7699 & w38913;
assign w16332 = ~w14855 & w16331;
assign w16333 = w3052 & ~w14352;
assign w16334 = w3066 & w14352;
assign w16335 = ~w16333 & ~w16334;
assign w16336 = w14860 & w16335;
assign w16337 = w3071 & ~w14867;
assign w16338 = w3056 & w14867;
assign w16339 = ~w14841 & w38914;
assign w16340 = w14836 & w16339;
assign w16341 = pi0140 & pi0979;
assign w16342 = pi0142 & ~pi0979;
assign w16343 = ~w16341 & ~w16342;
assign w16344 = w14873 & w16343;
assign w16345 = ~w16340 & ~w16344;
assign w16346 = ~w16336 & w16345;
assign w16347 = ~w16332 & w16346;
assign w16348 = (~w14806 & w16330) | (~w14806 & w38915) | (w16330 & w38915);
assign w16349 = ~pi0096 & ~w14808;
assign w16350 = ~w14882 & ~w16349;
assign w16351 = ~w16348 & w16350;
assign w16352 = ~w16329 & ~w16351;
assign w16353 = ~w10357 & w40175;
assign w16354 = (~w10594 & w10229) | (~w10594 & w38916) | (w10229 & w38916);
assign w16355 = ~w10356 & w16354;
assign w16356 = w10229 & w38917;
assign w16357 = ~w16355 & ~w16356;
assign w16358 = (w16357 & w16353) | (w16357 & w38918) | (w16353 & w38918);
assign w16359 = ~w16353 & w38919;
assign w16360 = ~w16358 & ~w16359;
assign w16361 = w14410 & w16360;
assign w16362 = (~w15041 & ~w14615) | (~w15041 & w38920) | (~w14615 & w38920);
assign w16363 = ~w14658 & ~w15051;
assign w16364 = ~w14669 & ~w15045;
assign w16365 = w14704 & w38536;
assign w16366 = pi3516 & ~w5204;
assign w16367 = ~w16365 & ~w16366;
assign w16368 = ~w14603 & w16367;
assign w16369 = w16368 & w38921;
assign w16370 = ~w14627 & ~w15020;
assign w16371 = ~w15024 & w15589;
assign w16372 = ~w16370 & ~w16371;
assign w16373 = ~w14631 & ~w15029;
assign w16374 = ~w14680 & ~w15037;
assign w16375 = ~w16373 & ~w16374;
assign w16376 = w16372 & w16375;
assign w16377 = w16376 & w38922;
assign w16378 = w16377 & w38923;
assign w16379 = w15017 & w16378;
assign w16380 = ~w16379 & w38538;
assign w16381 = ~w5319 & w38924;
assign w16382 = ~w14801 & ~w16381;
assign w16383 = (~pi0342 & ~w14733) | (~pi0342 & w38925) | (~w14733 & w38925);
assign w16384 = ~w16382 & w16383;
assign w16385 = w14798 & w40176;
assign w16386 = ~w5179 & ~w14816;
assign w16387 = ~w7569 & w38926;
assign w16388 = w14813 & ~w16387;
assign w16389 = ~w16386 & w16388;
assign w16390 = (~w5200 & w14820) | (~w5200 & w38927) | (w14820 & w38927);
assign w16391 = (~w5204 & w14824) | (~w5204 & w38928) | (w14824 & w38928);
assign w16392 = ~w16390 & ~w16391;
assign w16393 = w16389 & w16392;
assign w16394 = ~w16385 & w16393;
assign w16395 = ~w16384 & w16394;
assign w16396 = (w14745 & w14738) | (w14745 & w38929) | (w14738 & w38929);
assign w16397 = ~w5123 & ~w14752;
assign w16398 = ~w5119 & ~w14749;
assign w16399 = ~w16397 & ~w16398;
assign w16400 = w16396 & w16399;
assign w16401 = w14735 & w40177;
assign w16402 = ~w16400 & w16401;
assign w16403 = w14461 & w14507;
assign w16404 = w14495 & w38931;
assign w16405 = ~w14516 & ~w16404;
assign w16406 = w14712 & ~w15051;
assign w16407 = pi3516 & ~w5200;
assign w16408 = (~w16407 & ~w14541) | (~w16407 & w38932) | (~w14541 & w38932);
assign w16409 = ~w16406 & w16408;
assign w16410 = ~w15037 & w15524;
assign w16411 = w14760 & w38933;
assign w16412 = ~w16410 & ~w16411;
assign w16413 = w16409 & w16412;
assign w16414 = w16405 & w16413;
assign w16415 = w14564 & w16167;
assign w16416 = ~w14643 & ~w15056;
assign w16417 = ~w16415 & ~w16416;
assign w16418 = w16414 & w16417;
assign w16419 = w14714 & ~w15020;
assign w16420 = ~w15045 & w15510;
assign w16421 = ~w14636 & w15512;
assign w16422 = ~w16420 & ~w16421;
assign w16423 = ~w16419 & w16422;
assign w16424 = w14792 & w16423;
assign w16425 = ~w14789 & w38934;
assign w16426 = w14786 & ~w16425;
assign w16427 = w16418 & w38935;
assign w16428 = (~w16402 & w16427) | (~w16402 & w38936) | (w16427 & w38936);
assign w16429 = w16395 & w16428;
assign w16430 = ~w16380 & w16429;
assign w16431 = ~w16361 & w16430;
assign w16432 = ~w14408 & w16431;
assign w16433 = w16431 & w38469;
assign w16434 = ~w7569 & w38937;
assign w16435 = ~w14855 & w16434;
assign w16436 = w5138 & ~w14352;
assign w16437 = w5142 & w14352;
assign w16438 = ~w16436 & ~w16437;
assign w16439 = w14860 & w16438;
assign w16440 = w5115 & ~w14867;
assign w16441 = w5133 & w14867;
assign w16442 = ~w14841 & w38938;
assign w16443 = w14836 & w16442;
assign w16444 = pi0219 & pi0979;
assign w16445 = pi0221 & ~pi0979;
assign w16446 = ~w16444 & ~w16445;
assign w16447 = w14873 & w16446;
assign w16448 = ~w16443 & ~w16447;
assign w16449 = ~w16439 & w16448;
assign w16450 = ~w16435 & w16449;
assign w16451 = ~w14806 & ~w16450;
assign w16452 = (~pi0097 & w14807) | (~pi0097 & w38940) | (w14807 & w38940);
assign w16453 = ~w14882 & ~w16452;
assign w16454 = (w16453 & w5319) | (w16453 & w38941) | (w5319 & w38941);
assign w16455 = ~w16451 & w16454;
assign w16456 = ~w16433 & ~w16455;
assign w16457 = (~w10099 & w10461) | (~w10099 & w38943) | (w10461 & w38943);
assign w16458 = w10545 & ~w10593;
assign w16459 = (~w10594 & w10443) | (~w10594 & w38945) | (w10443 & w38945);
assign w16460 = ~w10545 & ~w16459;
assign w16461 = ~w16458 & ~w16460;
assign w16462 = (w10402 & w38946) | (w10402 & w38947) | (w38946 & w38947);
assign w16463 = w16461 & w40178;
assign w16464 = ~w16462 & ~w16463;
assign w16465 = w14410 & ~w16464;
assign w16466 = w14583 & w38948;
assign w16467 = ~w15024 & w15089;
assign w16468 = ~w16466 & ~w16467;
assign w16469 = ~w14474 & ~w14559;
assign w16470 = ~w16468 & ~w16469;
assign w16471 = w14586 & ~w15020;
assign w16472 = w14583 & w38949;
assign w16473 = w14711 & ~w15045;
assign w16474 = ~w10221 & w38950;
assign w16475 = w14600 & w16474;
assign w16476 = ~w16473 & ~w16475;
assign w16477 = ~w16472 & w16476;
assign w16478 = ~w16471 & w16477;
assign w16479 = (w14526 & ~w16478) | (w14526 & w38951) | (~w16478 & w38951);
assign w16480 = ~w14627 & ~w15051;
assign w16481 = ~w16163 & ~w16480;
assign w16482 = ~w14680 & ~w15029;
assign w16483 = w14610 & w15054;
assign w16484 = ~w14500 & ~w16483;
assign w16485 = w14484 & ~w16484;
assign w16486 = ~w16482 & ~w16485;
assign w16487 = w16481 & w16486;
assign w16488 = ~w14669 & ~w15041;
assign w16489 = pi3516 & ~w4083;
assign w16490 = w14454 & w38952;
assign w16491 = ~w16489 & ~w16490;
assign w16492 = ~w15792 & w16491;
assign w16493 = ~w16488 & w16492;
assign w16494 = w16487 & w16493;
assign w16495 = ~w16479 & w16494;
assign w16496 = (~pi0709 & ~w15466) | (~pi0709 & w38953) | (~w15466 & w38953);
assign w16497 = w14422 & w16496;
assign w16498 = ~w14615 & ~w15056;
assign w16499 = ~w14643 & ~w15037;
assign w16500 = ~w14631 & ~w15024;
assign w16501 = pi3516 & ~w4075;
assign w16502 = (~w16501 & ~w15524) | (~w16501 & w38954) | (~w15524 & w38954);
assign w16503 = ~w14536 & w16502;
assign w16504 = ~w16500 & w16503;
assign w16505 = ~w16499 & w16504;
assign w16506 = ~w14658 & ~w15045;
assign w16507 = ~w14789 & ~w15020;
assign w16508 = ~w15041 & w15510;
assign w16509 = w14454 & w38955;
assign w16510 = ~w16508 & ~w16509;
assign w16511 = w14611 & w15055;
assign w16512 = w14714 & ~w15051;
assign w16513 = ~w16511 & ~w16512;
assign w16514 = w16510 & w16513;
assign w16515 = w16514 & w38956;
assign w16516 = w16505 & w16515;
assign w16517 = ~w16498 & w16516;
assign w16518 = (w14758 & ~w16517) | (w14758 & w38881) | (~w16517 & w38881);
assign w16519 = ~w4023 & ~w14752;
assign w16520 = ~w4042 & ~w14738;
assign w16521 = ~w16519 & ~w16520;
assign w16522 = w16220 & w16521;
assign w16523 = w15868 & ~w16522;
assign w16524 = pi3245 & ~w7764;
assign w16525 = w14798 & w40189;
assign w16526 = (~w4075 & w14820) | (~w4075 & w38960) | (w14820 & w38960);
assign w16527 = (~w4083 & w14824) | (~w4083 & w38961) | (w14824 & w38961);
assign w16528 = (~w16527 & w4140) | (~w16527 & w38963) | (w4140 & w38963);
assign w16529 = ~w16526 & w16528;
assign w16530 = ~w4064 & ~w14816;
assign w16531 = w7764 & w14803;
assign w16532 = ~w16530 & ~w16531;
assign w16533 = (w10746 & w38964) | (w10746 & w38965) | (w38964 & w38965);
assign w16534 = w16529 & w16533;
assign w16535 = w16534 & w38966;
assign w16536 = ~w16518 & w16535;
assign w16537 = ~w16497 & w16536;
assign w16538 = ~w16465 & w16537;
assign w16539 = (w14882 & ~w16538) | (w14882 & w38890) | (~w16538 & w38890);
assign w16540 = w7764 & ~w14856;
assign w16541 = ~w14855 & w16540;
assign w16542 = w4046 & ~w14352;
assign w16543 = w4037 & w14352;
assign w16544 = ~w16542 & ~w16543;
assign w16545 = w14860 & w16544;
assign w16546 = w4031 & ~w14867;
assign w16547 = w4027 & w14867;
assign w16548 = ~w14841 & w38967;
assign w16549 = w14836 & w16548;
assign w16550 = pi0139 & pi0979;
assign w16551 = pi0141 & ~pi0979;
assign w16552 = ~w16550 & ~w16551;
assign w16553 = w14873 & w16552;
assign w16554 = ~w16549 & ~w16553;
assign w16555 = ~w16545 & w16554;
assign w16556 = ~w16541 & w16555;
assign w16557 = ~w14806 & ~w16556;
assign w16558 = (~pi0098 & w14807) | (~pi0098 & w38968) | (w14807 & w38968);
assign w16559 = (~w16558 & w4140) | (~w16558 & w38970) | (w4140 & w38970);
assign w16560 = ~w16557 & w16559;
assign w16561 = ~w16539 & w16560;
assign w16562 = ~w10099 & ~w10660;
assign w16563 = w10095 & w10105;
assign w16564 = (~w10099 & w10094) | (~w10099 & w38971) | (w10094 & w38971);
assign w16565 = (~w10594 & w9986) | (~w10594 & w38972) | (w9986 & w38972);
assign w16566 = ~w10097 & w16565;
assign w16567 = w9986 & w38973;
assign w16568 = ~w16566 & ~w16567;
assign w16569 = w16564 & ~w16568;
assign w16570 = ~w16564 & w16568;
assign w16571 = ~w16569 & ~w16570;
assign w16572 = w16562 & w38974;
assign w16573 = (~w16571 & ~w16562) | (~w16571 & w38975) | (~w16562 & w38975);
assign w16574 = ~w16572 & ~w16573;
assign w16575 = w14410 & w16574;
assign w16576 = w14640 & ~w14669;
assign w16577 = w14586 & ~w14653;
assign w16578 = w14534 & ~w15484;
assign w16579 = w14504 & ~w14638;
assign w16580 = ~w14776 & ~w16579;
assign w16581 = (w14583 & ~w16580) | (w14583 & w38976) | (~w16580 & w38976);
assign w16582 = w14534 & ~w14689;
assign w16583 = w14490 & w14772;
assign w16584 = w14504 & ~w14624;
assign w16585 = ~w16583 & ~w16584;
assign w16586 = ~w16582 & w16585;
assign w16587 = w14524 & ~w14763;
assign w16588 = w16585 & w38977;
assign w16589 = w14710 & ~w16588;
assign w16590 = ~w16589 & w38978;
assign w16591 = pi3516 & ~w7950;
assign w16592 = (~w16591 & w16590) | (~w16591 & w38979) | (w16590 & w38979);
assign w16593 = ~w16576 & w16592;
assign w16594 = w15820 & w38980;
assign w16595 = ~w16594 & w38538;
assign w16596 = ~w14716 & w14785;
assign w16597 = w15838 & w16596;
assign w16598 = w14576 & w16597;
assign w16599 = (w14673 & ~w14615) | (w14673 & w38981) | (~w14615 & w38981);
assign w16600 = ~w14653 & ~w14789;
assign w16601 = ~w14614 & w15483;
assign w16602 = ~w14658 & ~w14763;
assign w16603 = ~w16601 & ~w16602;
assign w16604 = ~w16600 & w16603;
assign w16605 = ~w14536 & w38982;
assign w16606 = ~w14587 & w16605;
assign w16607 = ~w14638 & ~w14643;
assign w16608 = ~w14680 & ~w14689;
assign w16609 = ~w14624 & ~w14631;
assign w16610 = ~w16608 & ~w16609;
assign w16611 = ~w16607 & w16610;
assign w16612 = ~w14669 & w14772;
assign w16613 = ~w14627 & ~w14666;
assign w16614 = pi3516 & ~w7958;
assign w16615 = (~w16614 & ~w15510) | (~w16614 & w38983) | (~w15510 & w38983);
assign w16616 = ~w16613 & w16615;
assign w16617 = ~w16612 & w16616;
assign w16618 = w16611 & w16617;
assign w16619 = w16618 & w38984;
assign w16620 = ~w16599 & w16619;
assign w16621 = (w14758 & ~w16620) | (w14758 & w38985) | (~w16620 & w38985);
assign w16622 = ~w7927 & ~w14738;
assign w16623 = ~w7942 & ~w14752;
assign w16624 = ~w16622 & ~w16623;
assign w16625 = w16220 & w16624;
assign w16626 = w15868 & ~w16625;
assign w16627 = (~w7950 & w14824) | (~w7950 & w38986) | (w14824 & w38986);
assign w16628 = pi3245 & ~w7994;
assign w16629 = ~w16628 & w40180;
assign w16630 = w14798 & w16629;
assign w16631 = ~w8080 & w38988;
assign w16632 = (w14813 & ~w7994) | (w14813 & w38989) | (~w7994 & w38989);
assign w16633 = ~w16631 & w16632;
assign w16634 = ~w16630 & w16633;
assign w16635 = ~w7982 & ~w14816;
assign w16636 = (~w7958 & w14820) | (~w7958 & w38990) | (w14820 & w38990);
assign w16637 = ~w16635 & ~w16636;
assign w16638 = w16634 & w38991;
assign w16639 = ~w16626 & w16638;
assign w16640 = ~w16621 & w16639;
assign w16641 = ~w16595 & w16640;
assign w16642 = ~w16575 & w16641;
assign w16643 = (w10746 & w38992) | (w10746 & w38993) | (w38992 & w38993);
assign w16644 = ~w14408 & w16643;
assign w16645 = w16642 & w16644;
assign w16646 = ~w8080 & w38994;
assign w16647 = w7994 & ~w14856;
assign w16648 = ~w14855 & w16647;
assign w16649 = w7919 & ~w14352;
assign w16650 = w7938 & w14352;
assign w16651 = ~w16649 & ~w16650;
assign w16652 = w14860 & w16651;
assign w16653 = w7923 & ~w14867;
assign w16654 = w7933 & w14867;
assign w16655 = ~w14841 & w38995;
assign w16656 = w14836 & w16655;
assign w16657 = pi0123 & pi0979;
assign w16658 = pi0124 & ~pi0979;
assign w16659 = ~w16657 & ~w16658;
assign w16660 = w14873 & w16659;
assign w16661 = ~w16656 & ~w16660;
assign w16662 = ~w16652 & w16661;
assign w16663 = ~w16648 & w16662;
assign w16664 = ~w16646 & w16663;
assign w16665 = (~pi0099 & w14807) | (~pi0099 & w38996) | (w14807 & w38996);
assign w16666 = ~w14882 & ~w16665;
assign w16667 = (w16666 & w16664) | (w16666 & w38997) | (w16664 & w38997);
assign w16668 = ~w16645 & ~w16667;
assign w16669 = ~w7891 & w38998;
assign w16670 = ~w14855 & w16669;
assign w16671 = w1513 & ~w14352;
assign w16672 = w1528 & w14352;
assign w16673 = ~w16671 & ~w16672;
assign w16674 = w14860 & w16673;
assign w16675 = w1532 & ~w14867;
assign w16676 = w1523 & w14867;
assign w16677 = ~w14841 & w38999;
assign w16678 = w14836 & w16677;
assign w16679 = pi0121 & pi0979;
assign w16680 = pi0125 & ~pi0979;
assign w16681 = ~w16679 & ~w16680;
assign w16682 = w14873 & w16681;
assign w16683 = ~w16678 & ~w16682;
assign w16684 = ~w16674 & w16683;
assign w16685 = ~w14852 & w16684;
assign w16686 = (~w14806 & ~w16685) | (~w14806 & w39000) | (~w16685 & w39000);
assign w16687 = ~pi0100 & ~w14808;
assign w16688 = (w1618 & w39001) | (w1618 & w39002) | (w39001 & w39002);
assign w16689 = (~w16688 & w16686) | (~w16688 & w39003) | (w16686 & w39003);
assign w16690 = ~w14882 & ~w16689;
assign w16691 = ~w14408 & w15882;
assign w16692 = w14610 & w39004;
assign w16693 = ~w14506 & ~w16692;
assign w16694 = w16405 & w16693;
assign w16695 = w14555 & w16694;
assign w16696 = w15817 & w39005;
assign w16697 = w15800 & w16696;
assign w16698 = w14583 & w39006;
assign w16699 = ~w15037 & w15089;
assign w16700 = w14583 & w39007;
assign w16701 = ~w16699 & ~w16700;
assign w16702 = ~w16698 & w16701;
assign w16703 = w14524 & ~w15615;
assign w16704 = w14583 & w39008;
assign w16705 = ~w15056 & w15085;
assign w16706 = ~w16704 & ~w16705;
assign w16707 = ~w16703 & w16706;
assign w16708 = (w14526 & ~w16707) | (w14526 & w39009) | (~w16707 & w39009);
assign w16709 = ~w14669 & ~w15051;
assign w16710 = pi3516 & ~w1540;
assign w16711 = (~w16710 & w14680) | (~w16710 & w39010) | (w14680 & w39010);
assign w16712 = ~w16709 & w16711;
assign w16713 = ~w16708 & w16712;
assign w16714 = w15798 & w16713;
assign w16715 = (~pi0709 & ~w16714) | (~pi0709 & w39011) | (~w16714 & w39011);
assign w16716 = w14422 & w16715;
assign w16717 = (~w15045 & ~w14615) | (~w15045 & w39012) | (~w14615 & w39012);
assign w16718 = ~w14658 & ~w15020;
assign w16719 = ~w14789 & ~w15029;
assign w16720 = ~w14643 & ~w15041;
assign w16721 = pi3516 & ~w1548;
assign w16722 = (~w16721 & ~w15510) | (~w16721 & w39013) | (~w15510 & w39013);
assign w16723 = ~w16720 & w16722;
assign w16724 = w16723 & w39014;
assign w16725 = ~w14631 & ~w15037;
assign w16726 = ~w14627 & ~w15024;
assign w16727 = ~w14680 & ~w15056;
assign w16728 = ~w16726 & ~w16727;
assign w16729 = ~w16725 & w16728;
assign w16730 = w16606 & w16729;
assign w16731 = w16730 & w39015;
assign w16732 = w16598 & w16731;
assign w16733 = ~w1509 & ~w14752;
assign w16734 = ~w1517 & ~w14738;
assign w16735 = ~w16733 & ~w16734;
assign w16736 = w16220 & w16735;
assign w16737 = w15868 & ~w16736;
assign w16738 = (pi3245 & w7891) | (pi3245 & w39016) | (w7891 & w39016);
assign w16739 = ~w16738 & w40181;
assign w16740 = w14798 & w16739;
assign w16741 = ~w7891 & w39019;
assign w16742 = (~w1540 & w14824) | (~w1540 & w39020) | (w14824 & w39020);
assign w16743 = ~w16741 & ~w16742;
assign w16744 = ~w1449 & ~w14816;
assign w16745 = (~w1548 & w14820) | (~w1548 & w39023) | (w14820 & w39023);
assign w16746 = (w1618 & w39024) | (w1618 & w39025) | (w39024 & w39025);
assign w16747 = w16746 & w39026;
assign w16748 = ~w16740 & w16747;
assign w16749 = ~w16737 & w16748;
assign w16750 = (w16749 & w16732) | (w16749 & w39027) | (w16732 & w39027);
assign w16751 = ~w16716 & w16750;
assign w16752 = ~w14410 & w16751;
assign w16753 = w10030 & w39028;
assign w16754 = (~w10594 & ~w10030) | (~w10594 & w39029) | (~w10030 & w39029);
assign w16755 = ~w10103 & w16754;
assign w16756 = ~w16753 & ~w16755;
assign w16757 = (w10403 & w39030) | (w10403 & w39031) | (w39030 & w39031);
assign w16758 = (~w10099 & w10079) | (~w10099 & w39032) | (w10079 & w39032);
assign w16759 = (~w16756 & w16757) | (~w16756 & w39033) | (w16757 & w39033);
assign w16760 = w16756 & w16758;
assign w16761 = ~w16757 & w16760;
assign w16762 = ~w16716 & w39034;
assign w16763 = ~w16759 & w16762;
assign w16764 = ~w16752 & ~w16763;
assign w16765 = ~w16764 & w39035;
assign w16766 = ~w16690 & ~w16765;
assign w16767 = (~w10594 & ~w10079) | (~w10594 & w39036) | (~w10079 & w39036);
assign w16768 = ~w10104 & w16767;
assign w16769 = w16562 & ~w16768;
assign w16770 = w10079 & w39037;
assign w16771 = ~w16768 & ~w16770;
assign w16772 = ~w16562 & ~w16771;
assign w16773 = ~w16769 & ~w16772;
assign w16774 = w14410 & ~w16773;
assign w16775 = w15838 & w39038;
assign w16776 = (w14662 & ~w14615) | (w14662 & w39039) | (~w14615 & w39039);
assign w16777 = ~w14631 & ~w15484;
assign w16778 = ~w14653 & w15510;
assign w16779 = pi3516 & ~w1191;
assign w16780 = (~w16779 & ~w15524) | (~w16779 & w39040) | (~w15524 & w39040);
assign w16781 = ~w16778 & w16780;
assign w16782 = ~w16777 & w16781;
assign w16783 = w14563 & w16782;
assign w16784 = ~w14614 & w14665;
assign w16785 = ~w14624 & ~w14658;
assign w16786 = ~w16784 & ~w16785;
assign w16787 = w16783 & w16786;
assign w16788 = ~w14789 & w39041;
assign w16789 = ~w14643 & ~w14763;
assign w16790 = w14550 & w15715;
assign w16791 = ~w16789 & ~w16790;
assign w16792 = ~w14680 & w14772;
assign w16793 = ~w14627 & ~w14689;
assign w16794 = ~w16792 & ~w16793;
assign w16795 = w16791 & w16794;
assign w16796 = w16795 & w39042;
assign w16797 = w16787 & w16796;
assign w16798 = w16797 & w39043;
assign w16799 = w14758 & ~w16798;
assign w16800 = w14586 & w14634;
assign w16801 = w14583 & w39044;
assign w16802 = ~w14677 & w15089;
assign w16803 = ~w16801 & ~w16802;
assign w16804 = w14583 & w39045;
assign w16805 = w14583 & w39046;
assign w16806 = ~w16804 & ~w16805;
assign w16807 = w16803 & w16806;
assign w16808 = ~w16800 & w16807;
assign w16809 = w14469 & ~w15695;
assign w16810 = ~w14543 & w39047;
assign w16811 = (~pi3518 & ~w14548) | (~pi3518 & w39048) | (~w14548 & w39048);
assign w16812 = ~w16810 & w16811;
assign w16813 = w14654 & w15714;
assign w16814 = (pi3518 & ~w14530) | (pi3518 & w39049) | (~w14530 & w39049);
assign w16815 = ~w16813 & w16814;
assign w16816 = w14521 & ~w16815;
assign w16817 = ~w16812 & w16816;
assign w16818 = ~w16809 & ~w16817;
assign w16819 = w16808 & w16818;
assign w16820 = w14526 & ~w16819;
assign w16821 = ~w14653 & ~w14669;
assign w16822 = w14640 & ~w14680;
assign w16823 = w14620 & w15472;
assign w16824 = pi3516 & ~w1187;
assign w16825 = ~w14589 & ~w16824;
assign w16826 = ~w16823 & w16825;
assign w16827 = ~w16822 & w16826;
assign w16828 = ~w16821 & w16827;
assign w16829 = w15794 & w16828;
assign w16830 = ~w16820 & w16829;
assign w16831 = w15781 & w39050;
assign w16832 = w14550 & ~w16831;
assign w16833 = w15859 & ~w16832;
assign w16834 = w16830 & w16833;
assign w16835 = (~pi0709 & ~w16834) | (~pi0709 & w39011) | (~w16834 & w39011);
assign w16836 = ~w1161 & ~w14752;
assign w16837 = ~w1147 & ~w14738;
assign w16838 = ~w16836 & ~w16837;
assign w16839 = w16220 & w16838;
assign w16840 = w15868 & ~w16839;
assign w16841 = pi3245 & w7860;
assign w16842 = (~w16841 & w1307) | (~w16841 & w39052) | (w1307 & w39052);
assign w16843 = w14798 & ~w16842;
assign w16844 = (~w1187 & w14824) | (~w1187 & w39053) | (w14824 & w39053);
assign w16845 = (~w1191 & w14820) | (~w1191 & w39055) | (w14820 & w39055);
assign w16846 = (~w16845 & w1307) | (~w16845 & w39056) | (w1307 & w39056);
assign w16847 = ~w16844 & w16846;
assign w16848 = ~w1136 & ~w14816;
assign w16849 = (w14813 & ~w7860) | (w14813 & w38989) | (~w7860 & w38989);
assign w16850 = ~w16848 & w16849;
assign w16851 = (w10746 & w39057) | (w10746 & w39058) | (w39057 & w39058);
assign w16852 = w16847 & w39059;
assign w16853 = ~w16840 & w16852;
assign w16854 = (w16853 & ~w16835) | (w16853 & w39060) | (~w16835 & w39060);
assign w16855 = ~w16799 & w16854;
assign w16856 = ~w16774 & w16855;
assign w16857 = ~w14408 & w16856;
assign w16858 = w16856 & w38469;
assign w16859 = ~w1307 & w39061;
assign w16860 = w7860 & ~w14856;
assign w16861 = ~w14855 & w16860;
assign w16862 = w1151 & ~w14352;
assign w16863 = w1157 & w14352;
assign w16864 = ~w16862 & ~w16863;
assign w16865 = w14860 & w16864;
assign w16866 = w1166 & ~w14867;
assign w16867 = w1170 & w14867;
assign w16868 = ~w14841 & w39062;
assign w16869 = w14836 & w16868;
assign w16870 = pi0122 & pi0979;
assign w16871 = pi0126 & ~pi0979;
assign w16872 = ~w16870 & ~w16871;
assign w16873 = w14873 & w16872;
assign w16874 = ~w16869 & ~w16873;
assign w16875 = ~w16865 & w16874;
assign w16876 = ~w16861 & w16875;
assign w16877 = (~w14806 & w16859) | (~w14806 & w39063) | (w16859 & w39063);
assign w16878 = ~pi0101 & ~w14808;
assign w16879 = ~w14882 & ~w16878;
assign w16880 = ~w16877 & w16879;
assign w16881 = ~w16858 & ~w16880;
assign w16882 = ~w7827 & w39064;
assign w16883 = ~w14855 & w16882;
assign w16884 = w5601 & ~w14352;
assign w16885 = w5582 & w14352;
assign w16886 = ~w16884 & ~w16885;
assign w16887 = w14860 & w16886;
assign w16888 = w5596 & ~w14867;
assign w16889 = w5586 & w14867;
assign w16890 = ~w14841 & w39067;
assign w16891 = w14836 & w16890;
assign w16892 = pi0090 & pi0979;
assign w16893 = pi0093 & ~pi0979;
assign w16894 = ~w16892 & ~w16893;
assign w16895 = w14873 & w16894;
assign w16896 = ~w16891 & ~w16895;
assign w16897 = ~w16887 & w16896;
assign w16898 = w16897 & w40182;
assign w16899 = ~pi0102 & ~w14808;
assign w16900 = (w16898 & w39069) | (w16898 & w39070) | (w39069 & w39070);
assign w16901 = ~w14882 & w16900;
assign w16902 = (w15022 & ~w14615) | (w15022 & w39071) | (~w14615 & w39071);
assign w16903 = ~w14789 & ~w15041;
assign w16904 = ~w15029 & w15510;
assign w16905 = pi3516 & ~w5617;
assign w16906 = (~w16905 & ~w15524) | (~w16905 & w39072) | (~w15524 & w39072);
assign w16907 = ~w14587 & w16906;
assign w16908 = ~w16904 & w16907;
assign w16909 = ~w16903 & w16908;
assign w16910 = ~w14614 & w15023;
assign w16911 = ~w14658 & ~w15037;
assign w16912 = ~w16910 & ~w16911;
assign w16913 = w16909 & w16912;
assign w16914 = ~w14558 & w16605;
assign w16915 = ~w14643 & ~w15020;
assign w16916 = ~w14627 & ~w15056;
assign w16917 = ~w14631 & ~w15045;
assign w16918 = ~w16916 & ~w16917;
assign w16919 = ~w16915 & w16918;
assign w16920 = w16914 & w16919;
assign w16921 = w16913 & w16920;
assign w16922 = w16921 & w39073;
assign w16923 = w14758 & ~w16922;
assign w16924 = ~w14680 & ~w15051;
assign w16925 = pi3516 & ~w5613;
assign w16926 = (~w16925 & ~w15472) | (~w16925 & w39074) | (~w15472 & w39074);
assign w16927 = w14504 & ~w15020;
assign w16928 = w15825 & w39075;
assign w16929 = w16183 & ~w16928;
assign w16930 = ~w15045 & w15469;
assign w16931 = ~w16929 & w39076;
assign w16932 = w16931 & w39077;
assign w16933 = w14555 & w16932;
assign w16934 = w14544 & w15801;
assign w16935 = w15781 & ~w16934;
assign w16936 = w14550 & ~w16935;
assign w16937 = w15794 & ~w16936;
assign w16938 = w16933 & w16937;
assign w16939 = (w14559 & ~w14541) | (w14559 & w39078) | (~w14541 & w39078);
assign w16940 = (~w16939 & w14545) | (~w16939 & w39079) | (w14545 & w39079);
assign w16941 = ~w14669 & ~w15029;
assign w16942 = w15816 & w39080;
assign w16943 = w14596 & w16942;
assign w16944 = w16938 & w16943;
assign w16945 = w15460 & w16274;
assign w16946 = (~pi0709 & ~w16944) | (~pi0709 & w39081) | (~w16944 & w39081);
assign w16947 = ~w5590 & ~w14752;
assign w16948 = ~w5605 & ~w14738;
assign w16949 = ~w16947 & ~w16948;
assign w16950 = w16220 & w16949;
assign w16951 = w15868 & ~w16950;
assign w16952 = (w5632 & w39082) | (w5632 & w39083) | (w39082 & w39083);
assign w16953 = (~w5617 & w14820) | (~w5617 & w39084) | (w14820 & w39084);
assign w16954 = ~w7827 & w39085;
assign w16955 = ~w16954 & w40183;
assign w16956 = ~w5566 & ~w14816;
assign w16957 = (~w5613 & w14824) | (~w5613 & w39088) | (w14824 & w39088);
assign w16958 = ~w16956 & ~w16957;
assign w16959 = w16955 & w39089;
assign w16960 = ~w16952 & w16959;
assign w16961 = ~w16951 & w16960;
assign w16962 = (w16961 & ~w16946) | (w16961 & w39090) | (~w16946 & w39090);
assign w16963 = ~w16923 & w16962;
assign w16964 = ~w14410 & w16963;
assign w16965 = w10493 & w39091;
assign w16966 = (~w10594 & ~w10493) | (~w10594 & w39092) | (~w10493 & w39092);
assign w16967 = ~w10541 & w16966;
assign w16968 = ~w16965 & ~w16967;
assign w16969 = w10548 & w40184;
assign w16970 = (~w10099 & w10524) | (~w10099 & w39096) | (w10524 & w39096);
assign w16971 = (w16969 & w39098) | (w16969 & w39099) | (w39098 & w39099);
assign w16972 = w16968 & w16970;
assign w16973 = (w16972 & ~w16969) | (w16972 & w39100) | (~w16969 & w39100);
assign w16974 = w16963 & w17669;
assign w16975 = ~w16964 & ~w16974;
assign w16976 = ~w16975 & w39101;
assign w16977 = ~w16901 & ~w16976;
assign w16978 = w10524 & w39104;
assign w16979 = (~w10594 & ~w10524) | (~w10594 & w39105) | (~w10524 & w39105);
assign w16980 = ~w10542 & w16979;
assign w16981 = ~w16978 & ~w16980;
assign w16982 = w16981 & w40185;
assign w16983 = (w10402 & w39106) | (w10402 & w39107) | (w39106 & w39107);
assign w16984 = ~w16982 & ~w16983;
assign w16985 = w14410 & w16984;
assign w16986 = ~w14653 & ~w14680;
assign w16987 = w14709 & ~w15791;
assign w16988 = ~w15464 & ~w16987;
assign w16989 = ~w16986 & w16988;
assign w16990 = pi3516 & ~w4941;
assign w16991 = (~w16990 & ~w15469) | (~w16990 & w39108) | (~w15469 & w39108);
assign w16992 = w16183 & ~w16586;
assign w16993 = w15472 & ~w15484;
assign w16994 = ~w16992 & w39109;
assign w16995 = w14610 & w39110;
assign w16996 = (~w16995 & ~w14690) | (~w16995 & w39111) | (~w14690 & w39111);
assign w16997 = w16994 & w16996;
assign w16998 = ~w15479 & ~w15780;
assign w16999 = w15621 & ~w16998;
assign w17000 = ~w14638 & ~w14669;
assign w17001 = ~w16999 & ~w17000;
assign w17002 = w16997 & w39112;
assign w17003 = w17002 & w39113;
assign w17004 = w14539 & w17003;
assign w17005 = (~pi0709 & ~w17004) | (~pi0709 & w39114) | (~w17004 & w39114);
assign w17006 = w14422 & w17005;
assign w17007 = ~w14614 & ~w14689;
assign w17008 = ~w14638 & w15510;
assign w17009 = w14612 & w14685;
assign w17010 = w14640 & w14714;
assign w17011 = ~w17009 & ~w17010;
assign w17012 = ~w17008 & w17011;
assign w17013 = ~w17007 & w17012;
assign w17014 = ~w14658 & ~w14677;
assign w17015 = ~w14763 & ~w14789;
assign w17016 = ~w17014 & ~w17015;
assign w17017 = w17013 & w17016;
assign w17018 = ~w14631 & ~w14666;
assign w17019 = pi3516 & ~w4933;
assign w17020 = (~w17019 & ~w15524) | (~w17019 & w39115) | (~w15524 & w39115);
assign w17021 = ~w14494 & w17020;
assign w17022 = ~w17018 & w17021;
assign w17023 = ~w14627 & w14772;
assign w17024 = ~w14624 & ~w14643;
assign w17025 = ~w17023 & ~w17024;
assign w17026 = w17022 & w17025;
assign w17027 = w16914 & w17026;
assign w17028 = w17017 & w17027;
assign w17029 = (w14758 & ~w17028) | (w14758 & w39116) | (~w17028 & w39116);
assign w17030 = ~w4977 & ~w14752;
assign w17031 = ~w4973 & ~w14738;
assign w17032 = ~w17030 & ~w17031;
assign w17033 = w16220 & w17032;
assign w17034 = w15868 & ~w17033;
assign w17035 = (~w4933 & w14820) | (~w4933 & w39117) | (w14820 & w39117);
assign w17036 = ~w7795 & w39118;
assign w17037 = (~w17036 & w5052) | (~w17036 & w39120) | (w5052 & w39120);
assign w17038 = ~w4962 & ~w14816;
assign w17039 = (~w4941 & w14824) | (~w4941 & w39121) | (w14824 & w39121);
assign w17040 = ~w17038 & ~w17039;
assign w17041 = w17037 & w39122;
assign w17042 = w14798 & w15171;
assign w17043 = w15882 & ~w17042;
assign w17044 = w17043 & w39123;
assign w17045 = ~w17029 & w17044;
assign w17046 = ~w17006 & w17045;
assign w17047 = ~w16985 & w17046;
assign w17048 = (w14882 & ~w17047) | (w14882 & w38890) | (~w17047 & w38890);
assign w17049 = ~w5052 & w39124;
assign w17050 = ~w7795 & w39125;
assign w17051 = ~w14855 & w17050;
assign w17052 = pi0070 & pi0979;
assign w17053 = pi0071 & ~pi0979;
assign w17054 = ~w17052 & ~w17053;
assign w17055 = w14873 & w17054;
assign w17056 = w4981 & ~w14867;
assign w17057 = w4996 & w14867;
assign w17058 = ~w14841 & w39126;
assign w17059 = w14836 & w17058;
assign w17060 = w4987 & ~w14352;
assign w17061 = w4992 & w14352;
assign w17062 = ~w17060 & ~w17061;
assign w17063 = w14860 & w17062;
assign w17064 = ~w17059 & ~w17063;
assign w17065 = ~w17055 & w17064;
assign w17066 = ~w17051 & w17065;
assign w17067 = (~w14806 & w17049) | (~w14806 & w39127) | (w17049 & w39127);
assign w17068 = ~pi0103 & ~w14808;
assign w17069 = ~w17067 & ~w17068;
assign w17070 = ~w17048 & w17069;
assign w17071 = ~w10099 & ~w10351;
assign w17072 = ~w10594 & ~w17071;
assign w17073 = (w17072 & ~w10330) | (w17072 & w39128) | (~w10330 & w39128);
assign w17074 = (pi1974 & w9956) | (pi1974 & w39129) | (w9956 & w39129);
assign w17075 = w10344 & w17074;
assign w17076 = (~w10353 & w17075) | (~w10353 & w39130) | (w17075 & w39130);
assign w17077 = w10344 & ~w10605;
assign w17078 = ~w10330 & w39131;
assign w17079 = (~w10351 & w17077) | (~w10351 & w39132) | (w17077 & w39132);
assign w17080 = ~w17076 & ~w17079;
assign w17081 = w14410 & ~w17080;
assign w17082 = ~w14614 & w39133;
assign w17083 = w15841 & w39134;
assign w17084 = w14640 & ~w14789;
assign w17085 = ~w14669 & ~w14689;
assign w17086 = ~w14720 & ~w17085;
assign w17087 = ~w17084 & w17086;
assign w17088 = ~w14631 & ~w14763;
assign w17089 = ~w14627 & ~w14677;
assign w17090 = ~w17088 & ~w17089;
assign w17091 = ~w14643 & w14652;
assign w17092 = (w14450 & ~w14527) | (w14450 & w14543) | (~w14527 & w14543);
assign w17093 = ~pi3518 & w14703;
assign w17094 = (~w14559 & w17093) | (~w14559 & w39135) | (w17093 & w39135);
assign w17095 = ~w17092 & w17094;
assign w17096 = ~w17091 & ~w17095;
assign w17097 = w17090 & w17096;
assign w17098 = ~w14638 & w14654;
assign w17099 = w14504 & ~w14648;
assign w17100 = w14469 & w39136;
assign w17101 = ~w17099 & ~w17100;
assign w17102 = w14483 & w14487;
assign w17103 = ~w17101 & w17102;
assign w17104 = (w14495 & w17103) | (w14495 & w39137) | (w17103 & w39137);
assign w17105 = pi3516 & ~w3576;
assign w17106 = (~w17105 & w15852) | (~w17105 & w39138) | (w15852 & w39138);
assign w17107 = ~w17104 & w17106;
assign w17108 = ~w14494 & w17107;
assign w17109 = ~w14666 & ~w14680;
assign w17110 = w14507 & ~w17101;
assign w17111 = w14548 & w15073;
assign w17112 = ~w17110 & ~w17111;
assign w17113 = (w14487 & w17110) | (w14487 & w39139) | (w17110 & w39139);
assign w17114 = w14548 & w14637;
assign w17115 = w14530 & w14772;
assign w17116 = ~w17114 & ~w17115;
assign w17117 = (w14610 & w17113) | (w14610 & w39140) | (w17113 & w39140);
assign w17118 = ~w17109 & ~w17117;
assign w17119 = w17108 & w17118;
assign w17120 = w17097 & w17119;
assign w17121 = w17120 & w39141;
assign w17122 = w14605 & w17121;
assign w17123 = ~w17122 & w38538;
assign w17124 = w14798 & w40171;
assign w17125 = ~w3588 & ~w14816;
assign w17126 = (~w3576 & w14824) | (~w3576 & w39143) | (w14824 & w39143);
assign w17127 = (~w17126 & w3710) | (~w17126 & w39144) | (w3710 & w39144);
assign w17128 = ~w17125 & w17127;
assign w17129 = (~w3580 & w14820) | (~w3580 & w39145) | (w14820 & w39145);
assign w17130 = w7473 & ~w14805;
assign w17131 = ~w17129 & ~w17130;
assign w17132 = (w10746 & w39146) | (w10746 & w39147) | (w39146 & w39147);
assign w17133 = w17128 & w39148;
assign w17134 = (w14745 & w14749) | (w14745 & w39149) | (w14749 & w39149);
assign w17135 = ~w3613 & ~w14752;
assign w17136 = ~w3631 & ~w14738;
assign w17137 = ~w17135 & ~w17136;
assign w17138 = w17134 & w17137;
assign w17139 = w14735 & w40186;
assign w17140 = ~w17138 & w17139;
assign w17141 = w14772 & ~w14789;
assign w17142 = w14792 & ~w16940;
assign w17143 = ~w17141 & w17142;
assign w17144 = w15801 & w39151;
assign w17145 = w14564 & w14698;
assign w17146 = w14583 & w39152;
assign w17147 = w14583 & w39153;
assign w17148 = w14548 & w39154;
assign w17149 = ~w17147 & ~w17148;
assign w17150 = (w14557 & ~w17149) | (w14557 & w39155) | (~w17149 & w39155);
assign w17151 = ~w17150 & w39156;
assign w17152 = ~w14677 & w14714;
assign w17153 = w15801 & ~w17112;
assign w17154 = ~w17152 & ~w17153;
assign w17155 = ~w14608 & w15512;
assign w17156 = w14530 & w14640;
assign w17157 = ~w17103 & w39157;
assign w17158 = w14454 & ~w17157;
assign w17159 = ~w17155 & ~w17158;
assign w17160 = w17154 & w17159;
assign w17161 = ~w14689 & w15510;
assign w17162 = pi3516 & ~w3580;
assign w17163 = (~w17162 & ~w15524) | (~w17162 & w39158) | (~w15524 & w39158);
assign w17164 = ~w17161 & w17163;
assign w17165 = w15075 & w17164;
assign w17166 = w17160 & w39159;
assign w17167 = (w14758 & ~w17166) | (w14758 & w39160) | (~w17166 & w39160);
assign w17168 = ~w17140 & ~w17167;
assign w17169 = w17133 & w17168;
assign w17170 = ~w17123 & w17169;
assign w17171 = ~w17081 & w17170;
assign w17172 = ~w14408 & w17171;
assign w17173 = w17171 & w38469;
assign w17174 = w7473 & ~w14856;
assign w17175 = ~w14855 & w17174;
assign w17176 = w3640 & ~w14352;
assign w17177 = w3617 & w14352;
assign w17178 = ~w17176 & ~w17177;
assign w17179 = w14860 & w17178;
assign w17180 = w3636 & ~w14867;
assign w17181 = w3621 & w14867;
assign w17182 = ~w14841 & w39161;
assign w17183 = w14836 & w17182;
assign w17184 = pi0091 & pi0979;
assign w17185 = pi0094 & ~pi0979;
assign w17186 = ~w17184 & ~w17185;
assign w17187 = w14873 & w17186;
assign w17188 = ~w17183 & ~w17187;
assign w17189 = ~w17179 & w17188;
assign w17190 = ~w17175 & w17189;
assign w17191 = ~w14806 & ~w17190;
assign w17192 = (~pi0104 & w14807) | (~pi0104 & w39163) | (w14807 & w39163);
assign w17193 = ~w14882 & ~w17192;
assign w17194 = (w17193 & w3710) | (w17193 & w39164) | (w3710 & w39164);
assign w17195 = ~w17191 & w17194;
assign w17196 = ~w17173 & ~w17195;
assign w17197 = (w14813 & ~w16538) | (w14813 & w39165) | (~w16538 & w39165);
assign w17198 = ~w14889 & ~w16548;
assign w17199 = ~pi0105 & w14889;
assign w17200 = ~w14813 & ~w17199;
assign w17201 = (w40189 & w39167) | (w40189 & w39168) | (w39167 & w39168);
assign w17202 = ~w17197 & ~w17201;
assign w17203 = w14841 & w40176;
assign w17204 = pi0106 & w14889;
assign w17205 = ~w14813 & ~w17204;
assign w17206 = w17205 & w40187;
assign w17207 = ~w16432 & ~w17206;
assign w17208 = (w14813 & ~w16240) | (w14813 & w39165) | (~w16240 & w39165);
assign w17209 = ~w14889 & ~w16251;
assign w17210 = ~pi0107 & w14889;
assign w17211 = ~w14813 & ~w17210;
assign w17212 = (w40191 & w39171) | (w40191 & w39172) | (w39171 & w39172);
assign w17213 = ~w17208 & ~w17212;
assign w17214 = ~w14887 & w39173;
assign w17215 = w14841 & w40174;
assign w17216 = ~w14889 & ~w16339;
assign w17217 = (~w17214 & w17215) | (~w17214 & w39174) | (w17215 & w39174);
assign w17218 = ~w14813 & ~w17217;
assign w17219 = ~w16328 & ~w17218;
assign w17220 = ~w14887 & w39175;
assign w17221 = ~w14889 & ~w16655;
assign w17222 = (w17221 & ~w16629) | (w17221 & w39176) | (~w16629 & w39176);
assign w17223 = (~w14813 & w17222) | (~w14813 & w39177) | (w17222 & w39177);
assign w17224 = w16642 & w16691;
assign w17225 = ~w17223 & ~w17224;
assign w17226 = ~w14887 & w39178;
assign w17227 = ~w14889 & ~w16677;
assign w17228 = (w17227 & ~w16739) | (w17227 & w39179) | (~w16739 & w39179);
assign w17229 = (~w14813 & w17228) | (~w14813 & w39180) | (w17228 & w39180);
assign w17230 = ~w16764 & w39181;
assign w17231 = ~w17229 & ~w17230;
assign w17232 = w14841 & ~w16842;
assign w17233 = pi0111 & w14889;
assign w17234 = ~w14813 & ~w17233;
assign w17235 = w17234 & w40188;
assign w17236 = ~w16857 & ~w17235;
assign w17237 = ~w14887 & w39183;
assign w17238 = (w5632 & w39184) | (w5632 & w39185) | (w39184 & w39185);
assign w17239 = ~w14889 & ~w16890;
assign w17240 = (~w17237 & w17238) | (~w17237 & w39186) | (w17238 & w39186);
assign w17241 = ~w14813 & ~w17240;
assign w17242 = ~w16975 & w39181;
assign w17243 = ~w17241 & ~w17242;
assign w17244 = (w14813 & ~w17047) | (w14813 & w39165) | (~w17047 & w39165);
assign w17245 = ~w14889 & ~w17058;
assign w17246 = ~pi0113 & w14889;
assign w17247 = ~w14813 & ~w17246;
assign w17248 = (w15171 & w39188) | (w15171 & w39189) | (w39188 & w39189);
assign w17249 = ~w17244 & ~w17248;
assign w17250 = ~w14887 & w39190;
assign w17251 = w14841 & w40171;
assign w17252 = ~w14889 & ~w17182;
assign w17253 = (~w17250 & w17251) | (~w17250 & w39191) | (w17251 & w39191);
assign w17254 = ~w14813 & ~w17253;
assign w17255 = ~w17172 & ~w17254;
assign w17256 = w13539 & w13806;
assign w17257 = w13539 & ~w13757;
assign w17258 = (w17257 & w13778) | (w17257 & w39192) | (w13778 & w39192);
assign w17259 = w13467 & ~w13768;
assign w17260 = w13764 & w17259;
assign w17261 = w13490 & w17259;
assign w17262 = (~w17261 & w17256) | (~w17261 & w39193) | (w17256 & w39193);
assign w17263 = w15969 & w40059;
assign w17264 = ~w12505 & w17263;
assign w17265 = ~w17262 & ~w17264;
assign w17266 = (pi0868 & ~w13730) | (pi0868 & w39194) | (~w13730 & w39194);
assign w17267 = ~w17264 & w39195;
assign w17268 = ~w13730 & w13768;
assign w17269 = ~w13467 & w14902;
assign w17270 = ~w17268 & ~w17269;
assign w17271 = ~w13765 & w17270;
assign w17272 = (w17271 & w14094) | (w17271 & w39196) | (w14094 & w39196);
assign w17273 = ~w13846 & w17272;
assign w17274 = w13467 & w14902;
assign w17275 = pi0868 & ~w17274;
assign w17276 = (w17275 & w14907) | (w17275 & w39197) | (w14907 & w39197);
assign w17277 = ~w17267 & ~w17276;
assign w17278 = ~w12505 & w15970;
assign w17279 = w13764 & ~w15967;
assign w17280 = ~w17278 & w17279;
assign w17281 = ~w17259 & w39198;
assign w17282 = (w10752 & w17280) | (w10752 & w39199) | (w17280 & w39199);
assign w17283 = w17277 & w17282;
assign w17284 = pi0115 & w10759;
assign w17285 = w15173 & ~w17284;
assign w17286 = (w17285 & ~w16629) | (w17285 & w39200) | (~w16629 & w39200);
assign w17287 = ~w17283 & ~w17286;
assign w17288 = pi0868 & w13764;
assign w17289 = ~w17258 & w17288;
assign w17290 = (pi0868 & w17259) | (pi0868 & w39201) | (w17259 & w39201);
assign w17291 = (~w17290 & w17256) | (~w17290 & w40060) | (w17256 & w40060);
assign w17292 = w15969 & w39202;
assign w17293 = ~w12505 & w17292;
assign w17294 = ~w17291 & ~w17293;
assign w17295 = ~w17265 & w17294;
assign w17296 = ~w13760 & ~w17258;
assign w17297 = ~w13490 & ~w13763;
assign w17298 = ~pi0868 & ~w17297;
assign w17299 = ~w17256 & w39203;
assign w17300 = ~w17278 & w17299;
assign w17301 = ~pi0868 & w17297;
assign w17302 = (~w17301 & w17256) | (~w17301 & w39204) | (w17256 & w39204);
assign w17303 = w15969 & w39205;
assign w17304 = ~w12505 & w17303;
assign w17305 = ~w17302 & ~w17304;
assign w17306 = ~w17300 & w17305;
assign w17307 = (w10752 & w17295) | (w10752 & w39206) | (w17295 & w39206);
assign w17308 = pi0116 & w10759;
assign w17309 = w15173 & ~w17308;
assign w17310 = (w17309 & ~w16739) | (w17309 & w39207) | (~w16739 & w39207);
assign w17311 = ~w17307 & ~w17310;
assign w17312 = ~w13532 & ~w15963;
assign w17313 = ~w15962 & w17312;
assign w17314 = ~pi0868 & ~w15967;
assign w17315 = ~w17278 & w17314;
assign w17316 = ~w17313 & w17315;
assign w17317 = pi0868 & w17297;
assign w17318 = ~w17256 & w39208;
assign w17319 = ~w17278 & w17318;
assign w17320 = pi0868 & ~w17297;
assign w17321 = (~w17320 & w17256) | (~w17320 & w39209) | (w17256 & w39209);
assign w17322 = w15969 & w40061;
assign w17323 = ~w12505 & w17322;
assign w17324 = ~w17321 & ~w17323;
assign w17325 = ~w17319 & w17324;
assign w17326 = ~w17325 & w39210;
assign w17327 = w10749 & ~w16842;
assign w17328 = pi0117 & w10759;
assign w17329 = w15173 & ~w17328;
assign w17330 = ~w17327 & w17329;
assign w17331 = ~w17326 & ~w17330;
assign w17332 = (w13923 & w17295) | (w13923 & w39211) | (w17295 & w39211);
assign w17333 = pi0118 & w13933;
assign w17334 = w14336 & ~w17333;
assign w17335 = (w17334 & ~w16739) | (w17334 & w39212) | (~w16739 & w39212);
assign w17336 = ~w17332 & ~w17335;
assign w17337 = (w13923 & w17280) | (w13923 & w39213) | (w17280 & w39213);
assign w17338 = w17277 & w17337;
assign w17339 = pi0119 & w13933;
assign w17340 = w14336 & ~w17339;
assign w17341 = (w17340 & ~w16629) | (w17340 & w39214) | (~w16629 & w39214);
assign w17342 = ~w17338 & ~w17341;
assign w17343 = ~w17325 & w39215;
assign w17344 = w13929 & ~w16842;
assign w17345 = pi0120 & w13933;
assign w17346 = w14336 & ~w17345;
assign w17347 = ~w17344 & w17346;
assign w17348 = ~w17343 & ~w17347;
assign w17349 = (w15185 & w17295) | (w15185 & w39216) | (w17295 & w39216);
assign w17350 = (pi0121 & ~w15184) | (pi0121 & w39217) | (~w15184 & w39217);
assign w17351 = ~w17349 & ~w17350;
assign w17352 = (pi0122 & ~w15184) | (pi0122 & w39218) | (~w15184 & w39218);
assign w17353 = ~w17325 & w39219;
assign w17354 = ~w17352 & ~w17353;
assign w17355 = (pi0123 & ~w15184) | (pi0123 & w39220) | (~w15184 & w39220);
assign w17356 = (w15185 & w17280) | (w15185 & w39221) | (w17280 & w39221);
assign w17357 = w17277 & w17356;
assign w17358 = ~w17355 & ~w17357;
assign w17359 = (pi0124 & ~w15184) | (pi0124 & w39222) | (~w15184 & w39222);
assign w17360 = (w15189 & w17280) | (w15189 & w39223) | (w17280 & w39223);
assign w17361 = w17277 & w17360;
assign w17362 = ~w17359 & ~w17361;
assign w17363 = (w15189 & w17295) | (w15189 & w39224) | (w17295 & w39224);
assign w17364 = pi0125 & ~w15189;
assign w17365 = ~w17363 & ~w17364;
assign w17366 = (pi0126 & ~w15184) | (pi0126 & w39225) | (~w15184 & w39225);
assign w17367 = ~w17325 & w39226;
assign w17368 = ~w17366 & ~w17367;
assign w17369 = ~w15353 & ~w15377;
assign w17370 = w15377 & ~w15410;
assign w17371 = w15325 & ~w17370;
assign w17372 = ~w17369 & w17371;
assign w17373 = w15407 & w15280;
assign w17374 = (w17373 & ~w15303) | (w17373 & w39227) | (~w15303 & w39227);
assign w17375 = w15303 & w39228;
assign w17376 = ~w17374 & ~w17375;
assign w17377 = w15326 & ~w17376;
assign w17378 = ~w15363 & ~w15433;
assign w17379 = w15300 & ~w15368;
assign w17380 = w17378 & ~w17379;
assign w17381 = ~w17377 & w17380;
assign w17382 = ~w17372 & w17381;
assign w17383 = ~w15303 & w15364;
assign w17384 = w15364 & w39229;
assign w17385 = ~w15297 & w15362;
assign w17386 = w15280 & w17385;
assign w17387 = ~w17384 & ~w17386;
assign w17388 = (w15380 & w17382) | (w15380 & w39230) | (w17382 & w39230);
assign w17389 = ~w15342 & w15379;
assign w17390 = (pi2555 & ~w15383) | (pi2555 & w39231) | (~w15383 & w39231);
assign w17391 = ~w17389 & w17390;
assign w17392 = ~w17388 & w17391;
assign w17393 = ~w15388 & w40133;
assign w17394 = (w6668 & w39234) | (w6668 & w39235) | (w39234 & w39235);
assign w17395 = ~w17393 & w17394;
assign w17396 = ~w17392 & ~w17395;
assign w17397 = ~w3710 & w39236;
assign w17398 = (w6668 & w39239) | (w6668 & w39240) | (w39239 & w39240);
assign w17399 = ~w17397 & w17398;
assign w17400 = w15378 & w39241;
assign w17401 = (pi2555 & ~w15383) | (pi2555 & w39242) | (~w15383 & w39242);
assign w17402 = (~w17399 & w17400) | (~w17399 & w39243) | (w17400 & w39243);
assign w17403 = pi0128 & ~w15208;
assign w17404 = ~w15228 & ~w17403;
assign w17405 = w15228 & w17403;
assign w17406 = ~w17404 & ~w17405;
assign w17407 = (w17406 & ~w15303) | (w17406 & w39244) | (~w15303 & w39244);
assign w17408 = w15303 & w39245;
assign w17409 = w15326 & w39246;
assign w17410 = w15325 & w17376;
assign w17411 = (w15280 & ~w15300) | (w15280 & w15353) | (~w15300 & w15353);
assign w17412 = ~w17410 & w17411;
assign w17413 = (w17378 & ~w17412) | (w17378 & w39247) | (~w17412 & w39247);
assign w17414 = w15362 & w15368;
assign w17415 = w15364 & w39248;
assign w17416 = ~w17414 & ~w17415;
assign w17417 = w15380 & ~w17399;
assign w17418 = (w17417 & w17413) | (w17417 & w39249) | (w17413 & w39249);
assign w17419 = ~w17402 & ~w17418;
assign w17420 = pi0599 & w9958;
assign w17421 = ~w17420 & w40209;
assign w17422 = (w341 & w39252) | (w341 & w39253) | (w39252 & w39253);
assign w17423 = (~pi2758 & w10058) | (~pi2758 & w39254) | (w10058 & w39254);
assign w17424 = (~w17423 & w15776) | (~w17423 & w39255) | (w15776 & w39255);
assign w17425 = ~pi3426 & ~w9958;
assign w17426 = (~w17174 & w3710) | (~w17174 & w39257) | (w3710 & w39257);
assign w17427 = ~w9954 & w17425;
assign w17428 = (~w17427 & ~w17426) | (~w17427 & w39258) | (~w17426 & w39258);
assign w17429 = (w15776 & w39259) | (w15776 & w39260) | (w39259 & w39260);
assign w17430 = w9954 & w17425;
assign w17431 = (~w17430 & ~w17426) | (~w17430 & w39261) | (~w17426 & w39261);
assign w17432 = ~w17424 & ~w17431;
assign w17433 = ~w17432 & w39262;
assign w17434 = ~w17422 & ~w17433;
assign w17435 = w12503 & w39263;
assign w17436 = (w17435 & w12037) | (w17435 & w39264) | (w12037 & w39264);
assign w17437 = w13192 & ~w13799;
assign w17438 = ~w13797 & ~w13802;
assign w17439 = w12760 & w17438;
assign w17440 = w17438 & w17837;
assign w17441 = ~w17436 & w17440;
assign w17442 = ~w12973 & ~w13774;
assign w17443 = (w12981 & ~w17442) | (w12981 & w39266) | (~w17442 & w39266);
assign w17444 = pi0868 & ~w17442;
assign w17445 = (w13775 & w17442) | (w13775 & w39267) | (w17442 & w39267);
assign w17446 = ~w17443 & ~w17445;
assign w17447 = ~w12749 & ~w17446;
assign w17448 = ~w12749 & ~w13775;
assign w17449 = ~w17442 & w17448;
assign w17450 = pi0868 & w17449;
assign w17451 = ~w17447 & ~w17450;
assign w17452 = ~w17441 & ~w17451;
assign w17453 = ~w12981 & ~w13775;
assign w17454 = ~w17444 & w17453;
assign w17455 = ~w17436 & w39268;
assign w17456 = pi0868 & ~w17446;
assign w17457 = ~w17444 & w39269;
assign w17458 = ~w17456 & ~w17457;
assign w17459 = ~w17455 & w17458;
assign w17460 = ~w17452 & w17459;
assign w17461 = w10752 & ~w17460;
assign w17462 = pi0130 & w10759;
assign w17463 = w15173 & ~w17462;
assign w17464 = (w17463 & ~w14325) | (w17463 & w39270) | (~w14325 & w39270);
assign w17465 = ~w17461 & ~w17464;
assign w17466 = w13923 & ~w17460;
assign w17467 = pi0131 & w13933;
assign w17468 = w14336 & ~w17467;
assign w17469 = (w17468 & ~w14325) | (w17468 & w39271) | (~w14325 & w39271);
assign w17470 = ~w17466 & ~w17469;
assign w17471 = w15185 & ~w17460;
assign w17472 = (pi0132 & ~w15184) | (pi0132 & w39272) | (~w15184 & w39272);
assign w17473 = ~w17471 & ~w17472;
assign w17474 = w15189 & ~w17460;
assign w17475 = (pi0133 & ~w15184) | (pi0133 & w39273) | (~w15184 & w39273);
assign w17476 = ~w17474 & ~w17475;
assign w17477 = ~w10652 & ~w10719;
assign w17478 = w10689 & w39274;
assign w17479 = pi0936 & pi1909;
assign w17480 = pi3586 & w17479;
assign w17481 = w10741 & ~w17480;
assign w17482 = ~w17478 & w17481;
assign w17483 = ~w17477 & w17482;
assign w17484 = w10749 & w40189;
assign w17485 = pi0135 & w10759;
assign w17486 = w15173 & ~w17485;
assign w17487 = ~w17484 & w17486;
assign w17488 = (~w10752 & w17484) | (~w10752 & w39275) | (w17484 & w39275);
assign w17489 = ~w12982 & ~w13774;
assign w17490 = (~w13075 & w12982) | (~w13075 & w17492) | (w12982 & w17492);
assign w17491 = ~w13779 & ~w17490;
assign w17492 = ~w13075 & w13774;
assign w17493 = ~w13779 & w17448;
assign w17494 = ~w17492 & w17493;
assign w17495 = ~w17491 & ~w17494;
assign w17496 = w17440 & ~w17491;
assign w17497 = ~w17436 & w17496;
assign w17498 = ~w13179 & ~w13780;
assign w17499 = ~pi0868 & ~w17498;
assign w17500 = ~w17497 & w39276;
assign w17501 = ~pi0868 & w17498;
assign w17502 = (w17501 & w17497) | (w17501 & w39277) | (w17497 & w39277);
assign w17503 = ~w17500 & ~w17502;
assign w17504 = (pi0868 & w13806) | (pi0868 & w40087) | (w13806 & w40087);
assign w17505 = pi0868 & w15148;
assign w17506 = ~w12505 & w17505;
assign w17507 = ~w17504 & ~w17506;
assign w17508 = w15162 & ~w17507;
assign w17509 = ~w17487 & ~w17508;
assign w17510 = w17503 & w17509;
assign w17511 = ~w17488 & ~w17510;
assign w17512 = w12981 & ~w17442;
assign w17513 = ~w17449 & ~w17512;
assign w17514 = ~w17512 & w40190;
assign w17515 = (~w17513 & w17436) | (~w17513 & w40079) | (w17436 & w40079);
assign w17516 = w12982 & ~w13774;
assign w17517 = (~pi0868 & ~w12982) | (~pi0868 & w39278) | (~w12982 & w39278);
assign w17518 = ~w17517 & w40190;
assign w17519 = (~pi0868 & ~w17516) | (~pi0868 & w39279) | (~w17516 & w39279);
assign w17520 = (w17519 & w17436) | (w17519 & w40080) | (w17436 & w40080);
assign w17521 = ~w17515 & w17520;
assign w17522 = w17439 & ~w17489;
assign w17523 = ~w13774 & w17448;
assign w17524 = ~w17489 & ~w17523;
assign w17525 = (~w17524 & w17437) | (~w17524 & w39280) | (w17437 & w39280);
assign w17526 = w17435 & ~w17524;
assign w17527 = ~w12093 & w17526;
assign w17528 = ~w13075 & ~w13779;
assign w17529 = pi0868 & ~w17528;
assign w17530 = ~w17527 & w39281;
assign w17531 = pi0868 & w17528;
assign w17532 = (w17531 & w17527) | (w17531 & w39282) | (w17527 & w39282);
assign w17533 = ~w17530 & ~w17532;
assign w17534 = w17533 & w40081;
assign w17535 = w10749 & w40174;
assign w17536 = pi0136 & w10759;
assign w17537 = w15173 & ~w17536;
assign w17538 = ~w17535 & w17537;
assign w17539 = ~w17534 & ~w17538;
assign w17540 = w13929 & w40189;
assign w17541 = pi0137 & w13933;
assign w17542 = w14336 & ~w17541;
assign w17543 = ~w17540 & w17542;
assign w17544 = (~w13923 & w17540) | (~w13923 & w39283) | (w17540 & w39283);
assign w17545 = ~w17508 & ~w17543;
assign w17546 = w17503 & w17545;
assign w17547 = ~w17544 & ~w17546;
assign w17548 = w17533 & w40082;
assign w17549 = w13929 & w40174;
assign w17550 = pi0138 & w13933;
assign w17551 = w14336 & ~w17550;
assign w17552 = ~w17549 & w17551;
assign w17553 = ~w17548 & ~w17552;
assign w17554 = (~pi0139 & ~w15184) | (~pi0139 & w39284) | (~w15184 & w39284);
assign w17555 = w15185 & ~w17508;
assign w17556 = w17503 & w17555;
assign w17557 = ~w17554 & ~w17556;
assign w17558 = (pi0140 & ~w15184) | (pi0140 & w39285) | (~w15184 & w39285);
assign w17559 = w17533 & w40083;
assign w17560 = ~w17558 & ~w17559;
assign w17561 = (~pi0141 & ~w15184) | (~pi0141 & w39286) | (~w15184 & w39286);
assign w17562 = w15189 & ~w17508;
assign w17563 = w17503 & w17562;
assign w17564 = ~w17561 & ~w17563;
assign w17565 = (pi0142 & ~w15184) | (pi0142 & w39287) | (~w15184 & w39287);
assign w17566 = w17533 & w40084;
assign w17567 = ~w17565 & ~w17566;
assign w17568 = (~w17423 & ~w15776) | (~w17423 & w39255) | (~w15776 & w39255);
assign w17569 = ~pi1041 & pi1042;
assign w17570 = ~pi1479 & w17569;
assign w17571 = ~pi1042 & pi1533;
assign w17572 = pi1042 & pi1551;
assign w17573 = pi1041 & ~w17572;
assign w17574 = ~w17571 & w17573;
assign w17575 = (~pi1093 & w17574) | (~pi1093 & w39288) | (w17574 & w39288);
assign w17576 = ~pi1041 & pi1497;
assign w17577 = pi1041 & pi1568;
assign w17578 = w10566 & ~w17577;
assign w17579 = ~w17576 & w17578;
assign w17580 = pi1041 & pi1613;
assign w17581 = ~pi1041 & pi1612;
assign w17582 = w10559 & ~w17581;
assign w17583 = ~w17580 & w17582;
assign w17584 = ~w17579 & ~w17583;
assign w17585 = ~w17575 & w17584;
assign w17586 = w10558 & w39289;
assign w17587 = (~w17586 & ~w6413) | (~w17586 & w39290) | (~w6413 & w39290);
assign w17588 = (w9954 & w17587) | (w9954 & w39291) | (w17587 & w39291);
assign w17589 = (w15776 & w39292) | (w15776 & w39293) | (w39292 & w39293);
assign w17590 = (~w9954 & w17587) | (~w9954 & w39294) | (w17587 & w39294);
assign w17591 = w17568 & w17590;
assign w17592 = w17425 & w17481;
assign w17593 = (w17592 & ~w341) | (w17592 & w39296) | (~w341 & w39296);
assign w17594 = ~w17591 & w39297;
assign w17595 = w6668 & ~w9958;
assign w17596 = w10689 & ~w17595;
assign w17597 = ~w17596 & w17587;
assign w17598 = (w17481 & ~w10689) | (w17481 & w39298) | (~w10689 & w39298);
assign w17599 = ~w17597 & w17598;
assign w17600 = ~w17594 & ~w17599;
assign w17601 = ~w17420 & w40144;
assign w17602 = (w341 & w39301) | (w341 & w39302) | (w39301 & w39302);
assign w17603 = ~w17432 & w39303;
assign w17604 = ~w17602 & ~w17603;
assign w17605 = w10749 & w40191;
assign w17606 = pi0145 & w10759;
assign w17607 = w15173 & ~w17606;
assign w17608 = ~w17605 & w17607;
assign w17609 = (~w10752 & w17605) | (~w10752 & w39304) | (w17605 & w39304);
assign w17610 = pi0868 & ~w17498;
assign w17611 = ~w17497 & w39305;
assign w17612 = pi0868 & w17498;
assign w17613 = (w17612 & w17497) | (w17612 & w39306) | (w17497 & w39306);
assign w17614 = ~w17611 & ~w17613;
assign w17615 = ~pi0868 & w17528;
assign w17616 = ~w17527 & w39307;
assign w17617 = ~pi0868 & ~w17528;
assign w17618 = (w17617 & w17527) | (w17617 & w39308) | (w17527 & w39308);
assign w17619 = ~w17616 & ~w17618;
assign w17620 = ~w17608 & w17619;
assign w17621 = w17614 & w17620;
assign w17622 = ~w17609 & ~w17621;
assign w17623 = w13929 & w40191;
assign w17624 = pi0146 & w13933;
assign w17625 = w14336 & ~w17624;
assign w17626 = ~w17623 & w17625;
assign w17627 = (~w13923 & w17623) | (~w13923 & w39309) | (w17623 & w39309);
assign w17628 = w17619 & ~w17626;
assign w17629 = w17614 & w17628;
assign w17630 = ~w17627 & ~w17629;
assign w17631 = (~pi0147 & ~w15184) | (~pi0147 & w39310) | (~w15184 & w39310);
assign w17632 = w15185 & w17619;
assign w17633 = w17614 & w17632;
assign w17634 = ~w17631 & ~w17633;
assign w17635 = (~pi0148 & ~w15184) | (~pi0148 & w39311) | (~w15184 & w39311);
assign w17636 = w15189 & w17619;
assign w17637 = w17614 & w17636;
assign w17638 = ~w17635 & ~w17637;
assign w17639 = w10689 & w39312;
assign w17640 = w17481 & ~w17639;
assign w17641 = ~pi1493 & w10564;
assign w17642 = ~pi1420 & w10559;
assign w17643 = ~pi1511 & w10566;
assign w17644 = ~w17642 & ~w17643;
assign w17645 = (~pi1041 & ~w17644) | (~pi1041 & w39314) | (~w17644 & w39314);
assign w17646 = (pi1041 & ~w10564) | (pi1041 & w39315) | (~w10564 & w39315);
assign w17647 = pi1547 & w10561;
assign w17648 = pi1580 & w10566;
assign w17649 = pi1414 & w10559;
assign w17650 = ~w17648 & ~w17649;
assign w17651 = w17650 & w39316;
assign w17652 = ~w17645 & ~w17651;
assign w17653 = w10558 & w39317;
assign w17654 = ~w10719 & ~w17653;
assign w17655 = (w17654 & w3710) | (w17654 & w39318) | (w3710 & w39318);
assign w17656 = w17640 & ~w17655;
assign w17657 = w10615 & w17080;
assign w17658 = ~w15014 & w17657;
assign w17659 = w17640 & w17658;
assign w17660 = ~w16360 & w17659;
assign w17661 = w17660 & w39319;
assign w17662 = w17661 & w39320;
assign w17663 = w17662 & w39321;
assign w17664 = w15776 & w16464;
assign w17665 = w17663 & w17664;
assign w17666 = w16773 & ~w16984;
assign w17667 = w17665 & w17666;
assign w17668 = ~w16759 & ~w16761;
assign w17669 = ~w16971 & ~w16973;
assign w17670 = ~w16574 & w17669;
assign w17671 = w17668 & w17670;
assign w17672 = w17667 & w17671;
assign w17673 = ~w17656 & ~w17672;
assign w17674 = ~pi0715 & pi2020;
assign w17675 = ~w10613 & w39322;
assign w17676 = w10750 & w17675;
assign w17677 = (pi0150 & ~w17675) | (pi0150 & w39323) | (~w17675 & w39323);
assign w17678 = ~pi0715 & ~w15778;
assign w17679 = (w17676 & ~w10746) | (w17676 & w39324) | (~w10746 & w39324);
assign w17680 = (w17679 & w15778) | (w17679 & w39325) | (w15778 & w39325);
assign w17681 = ~w17677 & ~w17680;
assign w17682 = w13922 & w17675;
assign w17683 = (pi0151 & ~w17675) | (pi0151 & w39326) | (~w17675 & w39326);
assign w17684 = (w17682 & ~w10746) | (w17682 & w39327) | (~w10746 & w39327);
assign w17685 = ~w17678 & w17684;
assign w17686 = ~w17683 & ~w17685;
assign w17687 = w10641 & ~w10719;
assign w17688 = (w17687 & w10625) | (w17687 & w39328) | (w10625 & w39328);
assign w17689 = (w17481 & ~w10719) | (w17481 & w39329) | (~w10719 & w39329);
assign w17690 = ~w17688 & w17689;
assign w17691 = (~pi0153 & ~w17675) | (~pi0153 & w39330) | (~w17675 & w39330);
assign w17692 = ~w14405 & w39331;
assign w17693 = w17676 & ~w17692;
assign w17694 = pi0715 & w40189;
assign w17695 = ~pi0715 & w14405;
assign w17696 = (~w17694 & ~w14405) | (~w17694 & w39333) | (~w14405 & w39333);
assign w17697 = w17693 & w17696;
assign w17698 = ~w17691 & ~w17697;
assign w17699 = (~pi0154 & ~w17675) | (~pi0154 & w39334) | (~w17675 & w39334);
assign w17700 = pi0715 & w40191;
assign w17701 = (~w17700 & ~w14405) | (~w17700 & w39336) | (~w14405 & w39336);
assign w17702 = w17693 & w17701;
assign w17703 = ~w17699 & ~w17702;
assign w17704 = (~pi0155 & ~w17675) | (~pi0155 & w39337) | (~w17675 & w39337);
assign w17705 = pi0715 & w40174;
assign w17706 = (~w17705 & ~w14405) | (~w17705 & w39339) | (~w14405 & w39339);
assign w17707 = w17693 & w17706;
assign w17708 = ~w17704 & ~w17707;
assign w17709 = (pi0156 & ~w17675) | (pi0156 & w39340) | (~w17675 & w39340);
assign w17710 = ~w14405 & w39341;
assign w17711 = w17676 & ~w17710;
assign w17712 = pi0715 & ~w14325;
assign w17713 = w14405 & w39342;
assign w17714 = ~w17712 & ~w17713;
assign w17715 = w17711 & w17714;
assign w17716 = ~w17709 & ~w17715;
assign w17717 = (~pi0157 & ~w17675) | (~pi0157 & w39343) | (~w17675 & w39343);
assign w17718 = pi0715 & w14962;
assign w17719 = (~w17718 & ~w14405) | (~w17718 & w39345) | (~w14405 & w39345);
assign w17720 = w17693 & w17719;
assign w17721 = ~w17717 & ~w17720;
assign w17722 = (~pi0158 & ~w17675) | (~pi0158 & w39346) | (~w17675 & w39346);
assign w17723 = pi0715 & w40168;
assign w17724 = (~w17723 & ~w14405) | (~w17723 & w39348) | (~w14405 & w39348);
assign w17725 = w17693 & w17724;
assign w17726 = ~w17722 & ~w17725;
assign w17727 = (pi0159 & ~w17675) | (pi0159 & w39349) | (~w17675 & w39349);
assign w17728 = (w5319 & w39350) | (w5319 & w39351) | (w39350 & w39351);
assign w17729 = (~w17728 & ~w14405) | (~w17728 & w39353) | (~w14405 & w39353);
assign w17730 = w17711 & w17729;
assign w17731 = ~w17727 & ~w17730;
assign w17732 = (pi0160 & ~w17675) | (pi0160 & w39354) | (~w17675 & w39354);
assign w17733 = pi0715 & ~w13916;
assign w17734 = (~w17733 & ~w14405) | (~w17733 & w39356) | (~w14405 & w39356);
assign w17735 = w17711 & w17734;
assign w17736 = ~w17732 & ~w17735;
assign w17737 = (pi0161 & ~w17675) | (pi0161 & w39357) | (~w17675 & w39357);
assign w17738 = (w4748 & w39358) | (w4748 & w39359) | (w39358 & w39359);
assign w17739 = (~w17738 & ~w14405) | (~w17738 & w39361) | (~w14405 & w39361);
assign w17740 = w17711 & w17739;
assign w17741 = ~w17737 & ~w17740;
assign w17742 = (~pi0162 & ~w17675) | (~pi0162 & w39362) | (~w17675 & w39362);
assign w17743 = pi0715 & w16629;
assign w17744 = (~w17743 & ~w17695) | (~w17743 & w39363) | (~w17695 & w39363);
assign w17745 = w17693 & w17744;
assign w17746 = ~w17742 & ~w17745;
assign w17747 = (~pi0163 & ~w17675) | (~pi0163 & w39364) | (~w17675 & w39364);
assign w17748 = pi0715 & w16739;
assign w17749 = (~w17748 & ~w17695) | (~w17748 & w39365) | (~w17695 & w39365);
assign w17750 = w17693 & w17749;
assign w17751 = ~w17747 & ~w17750;
assign w17752 = (~pi0164 & ~w17675) | (~pi0164 & w39366) | (~w17675 & w39366);
assign w17753 = pi0715 & ~w16842;
assign w17754 = (~w17753 & ~w17695) | (~w17753 & w39367) | (~w17695 & w39367);
assign w17755 = w17693 & w17754;
assign w17756 = ~w17752 & ~w17755;
assign w17757 = (~pi0165 & ~w17675) | (~pi0165 & w39368) | (~w17675 & w39368);
assign w17758 = (w5632 & w39369) | (w5632 & w39370) | (w39369 & w39370);
assign w17759 = w14405 & w39371;
assign w17760 = ~w17758 & ~w17759;
assign w17761 = w17693 & w17760;
assign w17762 = ~w17757 & ~w17761;
assign w17763 = (~pi0166 & ~w17675) | (~pi0166 & w39372) | (~w17675 & w39372);
assign w17764 = pi0715 & w40192;
assign w17765 = (~w17764 & ~w14405) | (~w17764 & w39374) | (~w14405 & w39374);
assign w17766 = w17693 & w17765;
assign w17767 = ~w17763 & ~w17766;
assign w17768 = (~pi0167 & ~w17675) | (~pi0167 & w39375) | (~w17675 & w39375);
assign w17769 = w17682 & ~w17692;
assign w17770 = w17696 & w17769;
assign w17771 = ~w17768 & ~w17770;
assign w17772 = (~pi0168 & ~w17675) | (~pi0168 & w39376) | (~w17675 & w39376);
assign w17773 = w17701 & w17769;
assign w17774 = ~w17772 & ~w17773;
assign w17775 = (~pi0169 & ~w17675) | (~pi0169 & w39377) | (~w17675 & w39377);
assign w17776 = w17706 & w17769;
assign w17777 = ~w17775 & ~w17776;
assign w17778 = (pi0170 & ~w17675) | (pi0170 & w39378) | (~w17675 & w39378);
assign w17779 = w17682 & ~w17710;
assign w17780 = w17714 & w17779;
assign w17781 = ~w17778 & ~w17780;
assign w17782 = (~pi0171 & ~w17675) | (~pi0171 & w39379) | (~w17675 & w39379);
assign w17783 = w17719 & w17769;
assign w17784 = ~w17782 & ~w17783;
assign w17785 = (~pi0172 & ~w17675) | (~pi0172 & w39380) | (~w17675 & w39380);
assign w17786 = w17724 & w17769;
assign w17787 = ~w17785 & ~w17786;
assign w17788 = (pi0173 & ~w17675) | (pi0173 & w39381) | (~w17675 & w39381);
assign w17789 = w17729 & w17779;
assign w17790 = ~w17788 & ~w17789;
assign w17791 = (pi0174 & ~w17675) | (pi0174 & w39382) | (~w17675 & w39382);
assign w17792 = (w3710 & w39383) | (w3710 & w39384) | (w39383 & w39384);
assign w17793 = (~w17792 & ~w14405) | (~w17792 & w39386) | (~w14405 & w39386);
assign w17794 = w17711 & w17793;
assign w17795 = ~w17791 & ~w17794;
assign w17796 = (pi0175 & ~w17675) | (pi0175 & w39387) | (~w17675 & w39387);
assign w17797 = w17734 & w17779;
assign w17798 = ~w17796 & ~w17797;
assign w17799 = (pi0176 & ~w17675) | (pi0176 & w39388) | (~w17675 & w39388);
assign w17800 = w17739 & w17779;
assign w17801 = ~w17799 & ~w17800;
assign w17802 = (~pi0177 & ~w17675) | (~pi0177 & w39389) | (~w17675 & w39389);
assign w17803 = w17744 & w17769;
assign w17804 = ~w17802 & ~w17803;
assign w17805 = (~pi0178 & ~w17675) | (~pi0178 & w39390) | (~w17675 & w39390);
assign w17806 = w17749 & w17769;
assign w17807 = ~w17805 & ~w17806;
assign w17808 = (~pi0179 & ~w17675) | (~pi0179 & w39391) | (~w17675 & w39391);
assign w17809 = w17754 & w17769;
assign w17810 = ~w17808 & ~w17809;
assign w17811 = (~pi0180 & ~w17675) | (~pi0180 & w39392) | (~w17675 & w39392);
assign w17812 = w17760 & w17769;
assign w17813 = ~w17811 & ~w17812;
assign w17814 = (~pi0181 & ~w17675) | (~pi0181 & w39393) | (~w17675 & w39393);
assign w17815 = w17765 & w17769;
assign w17816 = ~w17814 & ~w17815;
assign w17817 = (pi0182 & ~w17675) | (pi0182 & w39394) | (~w17675 & w39394);
assign w17818 = w17779 & w17793;
assign w17819 = ~w17817 & ~w17818;
assign w17820 = ~pi0709 & pi2140;
assign w17821 = ~w10613 & w39395;
assign w17822 = w10750 & w17821;
assign w17823 = pi0709 & ~w16842;
assign w17824 = (w17822 & w16835) | (w17822 & w39396) | (w16835 & w39396);
assign w17825 = (pi0183 & ~w17821) | (pi0183 & w39397) | (~w17821 & w39397);
assign w17826 = ~w17824 & ~w17825;
assign w17827 = w13922 & w17821;
assign w17828 = (w17827 & w16835) | (w17827 & w39398) | (w16835 & w39398);
assign w17829 = pi0184 & ~w17827;
assign w17830 = ~w17828 & ~w17829;
assign w17831 = w10749 & w40168;
assign w17832 = pi0185 & w10759;
assign w17833 = w15173 & ~w17832;
assign w17834 = ~w17831 & w17833;
assign w17835 = (~w10752 & w17831) | (~w10752 & w39399) | (w17831 & w39399);
assign w17836 = pi0868 & ~w17438;
assign w17837 = (w12760 & ~w13192) | (w12760 & w39400) | (~w13192 & w39400);
assign w17838 = (~w17836 & w17436) | (~w17836 & w39401) | (w17436 & w39401);
assign w17839 = (~w13799 & w12505) | (~w13799 & w39403) | (w12505 & w39403);
assign w17840 = ~w17838 & w17839;
assign w17841 = w12760 & ~w13799;
assign w17842 = ~pi0868 & ~w17841;
assign w17843 = w12760 & ~w17438;
assign w17844 = (pi0868 & ~w13803) | (pi0868 & w39405) | (~w13803 & w39405);
assign w17845 = ~w17843 & w17844;
assign w17846 = ~w17845 & w40193;
assign w17847 = ~w17834 & w17846;
assign w17848 = ~w17840 & w17847;
assign w17849 = ~w17835 & ~w17848;
assign w17850 = w13929 & w40168;
assign w17851 = pi0186 & w13933;
assign w17852 = w14336 & ~w17851;
assign w17853 = ~w17850 & w17852;
assign w17854 = (~w13923 & w17850) | (~w13923 & w39406) | (w17850 & w39406);
assign w17855 = w17846 & ~w17853;
assign w17856 = ~w17840 & w17855;
assign w17857 = ~w17854 & ~w17856;
assign w17858 = (~pi0187 & ~w15184) | (~pi0187 & w39407) | (~w15184 & w39407);
assign w17859 = w15185 & w17846;
assign w17860 = ~w17840 & w17859;
assign w17861 = ~w17858 & ~w17860;
assign w17862 = (~pi0188 & ~w15184) | (~pi0188 & w39408) | (~w15184 & w39408);
assign w17863 = w15189 & w17846;
assign w17864 = ~w17840 & w17863;
assign w17865 = ~w17862 & ~w17864;
assign w17866 = ~pi0248 & pi1017;
assign w17867 = ~pi0278 & pi0329;
assign w17868 = pi1017 & ~w17867;
assign w17869 = ~w17866 & ~w17868;
assign w17870 = ~pi0278 & pi1017;
assign w17871 = pi0278 & ~pi1017;
assign w17872 = ~w17870 & ~w17871;
assign w17873 = ~pi0248 & ~pi0329;
assign w17874 = ~pi0329 & pi0350;
assign w17875 = pi0331 & ~pi1017;
assign w17876 = ~pi0331 & pi1017;
assign w17877 = ~w17875 & ~w17876;
assign w17878 = (~w17874 & w17877) | (~w17874 & w39409) | (w17877 & w39409);
assign w17879 = (~w17873 & w17878) | (~w17873 & w39410) | (w17878 & w39410);
assign w17880 = w17872 & w17879;
assign w17881 = pi0370 & ~pi1017;
assign w17882 = ~pi0370 & pi1017;
assign w17883 = pi0329 & ~w17882;
assign w17884 = w17883 & w39411;
assign w17885 = ~pi0329 & ~pi0479;
assign w17886 = pi0248 & ~pi0329;
assign w17887 = ~w17885 & ~w17886;
assign w17888 = ~w17872 & ~w17887;
assign w17889 = ~w17884 & ~w17888;
assign w17890 = (~w17869 & w17880) | (~w17869 & w39412) | (w17880 & w39412);
assign w17891 = pi0278 & ~w17882;
assign w17892 = ~w17875 & w17891;
assign w17893 = ~pi0278 & ~w17881;
assign w17894 = (~pi0329 & ~w17893) | (~pi0329 & w39413) | (~w17893 & w39413);
assign w17895 = ~w17892 & w17894;
assign w17896 = pi0329 & pi0350;
assign w17897 = w17872 & w17896;
assign w17898 = ~w17895 & w39414;
assign w17899 = pi0329 & pi0479;
assign w17900 = ~w17899 & w39415;
assign w17901 = (~pi1017 & w17898) | (~pi1017 & w39416) | (w17898 & w39416);
assign w17902 = ~w17890 & ~w17901;
assign w17903 = w17870 & ~w17899;
assign w17904 = ~pi0248 & ~w17903;
assign w17905 = (w17878 & w39417) | (w17878 & w39418) | (w39417 & w39418);
assign w17906 = (~w17885 & ~w17883) | (~w17885 & w39419) | (~w17883 & w39419);
assign w17907 = ~w17906 & w39420;
assign w17908 = ~w17905 & ~w17907;
assign w17909 = w17904 & w17908;
assign w17910 = ~w17902 & ~w17909;
assign w17911 = (~pi1017 & w17902) | (~pi1017 & w39421) | (w17902 & w39421);
assign w17912 = ~pi0329 & ~w17877;
assign w17913 = (pi0248 & w17912) | (pi0248 & w39422) | (w17912 & w39422);
assign w17914 = w17872 & w17899;
assign w17915 = w17872 & w39423;
assign w17916 = ~pi0329 & ~pi0370;
assign w17917 = ~w17896 & ~w17916;
assign w17918 = w17870 & ~w17917;
assign w17919 = pi0329 & ~pi0350;
assign w17920 = w17871 & ~w17916;
assign w17921 = ~w17919 & w17920;
assign w17922 = ~w17918 & ~w17921;
assign w17923 = ~w17915 & w17922;
assign w17924 = w17923 & w39424;
assign w17925 = (w17869 & w17880) | (w17869 & w39425) | (w17880 & w39425);
assign w17926 = ~w17924 & ~w17925;
assign w17927 = w17911 & w17926;
assign w17928 = ~w17911 & ~w17926;
assign w17929 = ~w17927 & ~w17928;
assign w17930 = ~pi0248 & ~pi0278;
assign w17931 = (~w17890 & ~w17911) | (~w17890 & w39426) | (~w17911 & w39426);
assign w17932 = ~w17867 & ~w17871;
assign w17933 = pi0248 & ~w17932;
assign w17934 = (~w17933 & ~w17908) | (~w17933 & w39427) | (~w17908 & w39427);
assign w17935 = pi0248 & ~w17914;
assign w17936 = w17922 & w17935;
assign w17937 = pi0350 & pi0370;
assign w17938 = pi1017 & ~w17937;
assign w17939 = ~pi0278 & w17886;
assign w17940 = ~w17938 & w17939;
assign w17941 = pi0278 & pi1017;
assign w17942 = (w17941 & w17906) | (w17941 & w39428) | (w17906 & w39428);
assign w17943 = ~w17940 & ~w17942;
assign w17944 = (w17943 & w17934) | (w17943 & w39429) | (w17934 & w39429);
assign w17945 = w17872 & w17887;
assign w17946 = w17906 & ~w17945;
assign w17947 = w17933 & ~w17946;
assign w17948 = ~w17869 & w17936;
assign w17949 = ~w17947 & ~w17948;
assign w17950 = (~pi1017 & w17899) | (~pi1017 & w39430) | (w17899 & w39430);
assign w17951 = pi0278 & pi0329;
assign w17952 = ~w17950 & w17951;
assign w17953 = pi0248 & pi0278;
assign w17954 = ~pi0329 & w17871;
assign w17955 = w17953 & ~w17954;
assign w17956 = ~w17952 & w17955;
assign w17957 = ~w17948 & w39431;
assign w17958 = ~pi0247 & ~w17866;
assign w17959 = ~w17957 & w17958;
assign w17960 = (~pi0247 & w17959) | (~pi0247 & w39432) | (w17959 & w39432);
assign w17961 = pi1017 & w17895;
assign w17962 = ~w17868 & w17908;
assign w17963 = (pi0248 & w17962) | (pi0248 & w39433) | (w17962 & w39433);
assign w17964 = w17904 & ~w17908;
assign w17965 = ~w17898 & w17941;
assign w17966 = ~w17964 & ~w17965;
assign w17967 = ~w17963 & w17966;
assign w17968 = ~w17960 & ~w17967;
assign w17969 = (~pi0247 & ~w17968) | (~pi0247 & w39434) | (~w17968 & w39434);
assign w17970 = w17929 & ~w17969;
assign w17971 = (~pi0247 & w17969) | (~pi0247 & w39435) | (w17969 & w39435);
assign w17972 = w17872 & w17873;
assign w17973 = ~w17884 & w17945;
assign w17974 = ~pi0248 & w17878;
assign w17975 = (~w17872 & ~w17878) | (~w17872 & w39422) | (~w17878 & w39422);
assign w17976 = ~w17973 & ~w17975;
assign w17977 = ~pi1017 & w17976;
assign w17978 = ~w17895 & w39436;
assign w17979 = pi1017 & w17978;
assign w17980 = ~w17977 & ~w17979;
assign w17981 = (w17869 & ~w17923) | (w17869 & w39437) | (~w17923 & w39437);
assign w17982 = ~w17869 & ~w17976;
assign w17983 = ~w17981 & ~w17982;
assign w17984 = w17980 & ~w17983;
assign w17985 = (~w17941 & w17912) | (~w17941 & w39438) | (w17912 & w39438);
assign w17986 = pi0278 & ~w17876;
assign w17987 = ~pi0350 & ~pi1017;
assign w17988 = ~pi0329 & ~w17987;
assign w17989 = ~w17986 & w17988;
assign w17990 = ~w17989 & w40194;
assign w17991 = (w17868 & w17974) | (w17868 & w39441) | (w17974 & w39441);
assign w17992 = ~pi1017 & w17978;
assign w17993 = ~w17991 & ~w17992;
assign w17994 = ~w17992 & w39442;
assign w17995 = w17984 & w39443;
assign w17996 = (~w17972 & ~w17995) | (~w17972 & w39444) | (~w17995 & w39444);
assign w17997 = ~w17971 & w17996;
assign w17998 = (~pi1017 & ~w17971) | (~pi1017 & w39445) | (~w17971 & w39445);
assign w17999 = ~w17997 & w17998;
assign w18000 = ~pi0247 & pi1017;
assign w18001 = pi0955 & ~w18000;
assign w18002 = ~pi0189 & ~pi0955;
assign w18003 = ~pi0582 & pi3530;
assign w18004 = ~pi2599 & ~w18003;
assign w18005 = ~w18002 & w18004;
assign w18006 = (w18005 & w17999) | (w18005 & w39446) | (w17999 & w39446);
assign w18007 = ~pi0831 & w6668;
assign w18008 = pi2599 & ~w18003;
assign w18009 = w6668 & w39447;
assign w18010 = ~w1307 & w39448;
assign w18011 = ~pi0610 & w18003;
assign w18012 = (w18008 & ~w6668) | (w18008 & w39449) | (~w6668 & w39449);
assign w18013 = (w6668 & w39452) | (w6668 & w39453) | (w39452 & w39453);
assign w18014 = ~w18010 & w18013;
assign w18015 = ~w18006 & w18014;
assign w18016 = pi0868 & ~w17453;
assign w18017 = pi0868 & w12749;
assign w18018 = (~w18017 & w17436) | (~w18017 & w39454) | (w17436 & w39454);
assign w18019 = ~w18016 & ~w18018;
assign w18020 = ~pi0868 & ~w17438;
assign w18021 = ~w18016 & ~w18020;
assign w18022 = ~w18017 & ~w18021;
assign w18023 = (w18022 & w17436) | (w18022 & w39455) | (w17436 & w39455);
assign w18024 = w12983 & w18016;
assign w18025 = ~w18023 & ~w18024;
assign w18026 = ~w18019 & w18025;
assign w18027 = w10752 & ~w18026;
assign w18028 = pi0190 & w10759;
assign w18029 = w15173 & ~w18028;
assign w18030 = (w18029 & ~w14962) | (w18029 & w39456) | (~w14962 & w39456);
assign w18031 = ~w18027 & ~w18030;
assign w18032 = w13923 & ~w18026;
assign w18033 = pi0191 & w13933;
assign w18034 = w14336 & ~w18033;
assign w18035 = (w18034 & ~w14962) | (w18034 & w39457) | (~w14962 & w39457);
assign w18036 = ~w18032 & ~w18035;
assign w18037 = pi0868 & ~w16097;
assign w18038 = (w10752 & w18037) | (w10752 & w39458) | (w18037 & w39458);
assign w18039 = ~pi0695 & w40209;
assign w18040 = (w341 & w39461) | (w341 & w39462) | (w39461 & w39462);
assign w18041 = ~w10753 & ~w18040;
assign w18042 = (w18041 & ~w10746) | (w18041 & w39463) | (~w10746 & w39463);
assign w18043 = w15173 & ~w18042;
assign w18044 = ~w18038 & ~w18043;
assign w18045 = (w13923 & w18037) | (w13923 & w39464) | (w18037 & w39464);
assign w18046 = ~pi0695 & w40144;
assign w18047 = (~pi0193 & ~w40144) | (~pi0193 & w39465) | (~w40144 & w39465);
assign w18048 = ~w13925 & ~w18047;
assign w18049 = (w18048 & ~w10746) | (w18048 & w39466) | (~w10746 & w39466);
assign w18050 = w14336 & ~w18049;
assign w18051 = ~w18045 & ~w18050;
assign w18052 = w15185 & ~w18026;
assign w18053 = (pi0194 & ~w15184) | (pi0194 & w39467) | (~w15184 & w39467);
assign w18054 = ~w18052 & ~w18053;
assign w18055 = w15189 & ~w18026;
assign w18056 = (pi0195 & ~w15184) | (pi0195 & w39468) | (~w15184 & w39468);
assign w18057 = ~w18055 & ~w18056;
assign w18058 = ~w10667 & w39469;
assign w18059 = w10689 & w39470;
assign w18060 = w17481 & ~w18059;
assign w18061 = ~w18058 & w18060;
assign w18062 = pi0709 & w40189;
assign w18063 = (w17822 & w16496) | (w17822 & w39471) | (w16496 & w39471);
assign w18064 = (pi0197 & ~w17821) | (pi0197 & w39472) | (~w17821 & w39472);
assign w18065 = ~w18063 & ~w18064;
assign w18066 = (w17827 & w16496) | (w17827 & w39473) | (w16496 & w39473);
assign w18067 = pi0198 & ~w17827;
assign w18068 = ~w18066 & ~w18067;
assign w18069 = ~pi0586 & w14424;
assign w18070 = pi0586 & ~w14424;
assign w18071 = ~w18069 & ~w18070;
assign w18072 = ~pi2021 & w14449;
assign w18073 = pi0152 & w10005;
assign w18074 = w18072 & ~w18073;
assign w18075 = (w18074 & ~w18071) | (w18074 & w39474) | (~w18071 & w39474);
assign w18076 = ~w14424 & w14651;
assign w18077 = w14424 & ~w14651;
assign w18078 = ~w18076 & ~w18077;
assign w18079 = ~w14424 & w14648;
assign w18080 = w14424 & ~w14648;
assign w18081 = ~w18079 & ~w18080;
assign w18082 = w14684 & w14702;
assign w18083 = w14687 & ~w18082;
assign w18084 = (w14664 & w18083) | (w14664 & w39475) | (w18083 & w39475);
assign w18085 = (~w14675 & w18084) | (~w14675 & w39476) | (w18084 & w39476);
assign w18086 = w14424 & w14608;
assign w18087 = w14633 & w18086;
assign w18088 = w18087 & w40195;
assign w18089 = ~w14684 & ~w14702;
assign w18090 = ~w14687 & ~w18089;
assign w18091 = (~w14664 & w18090) | (~w14664 & w39478) | (w18090 & w39478);
assign w18092 = (w14675 & w18091) | (w14675 & w39479) | (w18091 & w39479);
assign w18093 = ~w14424 & ~w14608;
assign w18094 = ~w14633 & w18093;
assign w18095 = w18094 & w40196;
assign w18096 = w14636 & ~w14648;
assign w18097 = ~w14636 & w14648;
assign w18098 = ~w18096 & ~w18097;
assign w18099 = ~w14424 & w14633;
assign w18100 = w14424 & ~w14633;
assign w18101 = ~w18099 & ~w18100;
assign w18102 = w14633 & ~w14697;
assign w18103 = ~w14633 & w14697;
assign w18104 = ~w18102 & ~w18103;
assign w18105 = w18101 & ~w18104;
assign w18106 = w18098 & ~w18105;
assign w18107 = ~w18095 & w18106;
assign w18108 = (w18081 & ~w18107) | (w18081 & w39481) | (~w18107 & w39481);
assign w18109 = (w18075 & w18108) | (w18075 & w39482) | (w18108 & w39482);
assign w18110 = w18075 & w18078;
assign w18111 = w18081 & w18098;
assign w18112 = w18101 & w18104;
assign w18113 = ~w14622 & w18093;
assign w18114 = w14622 & w18086;
assign w18115 = ~w18113 & ~w18114;
assign w18116 = w14619 & ~w14675;
assign w18117 = w14424 & ~w18116;
assign w18118 = ~w14619 & w14675;
assign w18119 = ~w14424 & ~w18118;
assign w18120 = ~w18117 & ~w18119;
assign w18121 = ~w14424 & ~w14687;
assign w18122 = w14661 & w18121;
assign w18123 = ~w14684 & w14702;
assign w18124 = w18122 & ~w18123;
assign w18125 = ~w14424 & ~w14664;
assign w18126 = w14672 & w18125;
assign w18127 = w14424 & w14664;
assign w18128 = ~w14672 & w18127;
assign w18129 = ~w18126 & ~w18128;
assign w18130 = w14424 & w14687;
assign w18131 = ~w14661 & w18130;
assign w18132 = w14684 & ~w14702;
assign w18133 = w18131 & ~w18132;
assign w18134 = ~w18129 & ~w18133;
assign w18135 = (w18120 & ~w18134) | (w18120 & w39483) | (~w18134 & w39483);
assign w18136 = (w18112 & w18135) | (w18112 & w39484) | (w18135 & w39484);
assign w18137 = (w18110 & w18136) | (w18110 & w39485) | (w18136 & w39485);
assign w18138 = (w3563 & w18137) | (w3563 & w39486) | (w18137 & w39486);
assign w18139 = ~w18109 & w18138;
assign w18140 = (w18136 & w39487) | (w18136 & w39488) | (w39487 & w39488);
assign w18141 = w18111 & w18112;
assign w18142 = ~w18115 & w18120;
assign w18143 = ~w18122 & ~w18131;
assign w18144 = ~w18129 & ~w18143;
assign w18145 = w18142 & ~w18144;
assign w18146 = (w18110 & w18145) | (w18110 & w39489) | (w18145 & w39489);
assign w18147 = w5754 & w18146;
assign w18148 = ~w18140 & ~w18147;
assign w18149 = w18141 & w18142;
assign w18150 = w18110 & ~w18149;
assign w18151 = (~w5217 & w18149) | (~w5217 & w39490) | (w18149 & w39490);
assign w18152 = ~w5754 & ~w18146;
assign w18153 = ~w18151 & ~w18152;
assign w18154 = (w18153 & w18139) | (w18153 & w39491) | (w18139 & w39491);
assign w18155 = ~w18073 & w18078;
assign w18156 = (~w9999 & ~w18078) | (~w9999 & w39492) | (~w18078 & w39492);
assign w18157 = w9999 & w18078;
assign w18158 = ~w18071 & w18157;
assign w18159 = (w18072 & w18158) | (w18072 & w39493) | (w18158 & w39493);
assign w18160 = ~w1178 & w18159;
assign w18161 = ~w18149 & w39494;
assign w18162 = ~w18160 & ~w18161;
assign w18163 = ~w18158 & w39495;
assign w18164 = ~w9999 & w18072;
assign w18165 = w18072 & w39496;
assign w18166 = ~w10613 & w39497;
assign w18167 = ~w18163 & w18166;
assign w18168 = pi0867 & ~pi3426;
assign w18169 = ~w18168 & w40197;
assign w18170 = w10750 & ~w18169;
assign w18171 = ~pi0867 & w18159;
assign w18172 = ~w18171 & w40198;
assign w18173 = w18170 & ~w18172;
assign w18174 = (~pi0199 & w18169) | (~pi0199 & w39502) | (w18169 & w39502);
assign w18175 = ~w18173 & ~w18174;
assign w18176 = (pi0200 & w18169) | (pi0200 & w39503) | (w18169 & w39503);
assign w18177 = (~pi0867 & w18149) | (~pi0867 & w39505) | (w18149 & w39505);
assign w18178 = ~w18177 & w40199;
assign w18179 = w18170 & w18178;
assign w18180 = ~w18176 & ~w18179;
assign w18181 = (pi0201 & w18169) | (pi0201 & w39506) | (w18169 & w39506);
assign w18182 = (w5893 & w39507) | (w5893 & w39508) | (w39507 & w39508);
assign w18183 = ~pi0867 & ~w18146;
assign w18184 = ~w18182 & ~w18183;
assign w18185 = ~w18169 & w39509;
assign w18186 = ~w18181 & ~w18185;
assign w18187 = (pi0202 & w18169) | (pi0202 & w39510) | (w18169 & w39510);
assign w18188 = (pi0867 & w4748) | (pi0867 & w39511) | (w4748 & w39511);
assign w18189 = ~pi0867 & ~w18137;
assign w18190 = ~w18188 & ~w18189;
assign w18191 = ~w18169 & w39512;
assign w18192 = ~w18187 & ~w18191;
assign w18193 = (w18154 & w39513) | (w18154 & w39514) | (w39513 & w39514);
assign w18194 = ~w18172 & w18193;
assign w18195 = ~pi0203 & ~w18193;
assign w18196 = ~w18194 & ~w18195;
assign w18197 = pi0204 & ~w18193;
assign w18198 = w18178 & w18193;
assign w18199 = ~w18197 & ~w18198;
assign w18200 = (pi0867 & w3710) | (pi0867 & w39515) | (w3710 & w39515);
assign w18201 = (w18108 & w39516) | (w18108 & w39517) | (w39516 & w39517);
assign w18202 = ~w18200 & ~w18201;
assign w18203 = ~w18169 & w39518;
assign w18204 = (~pi0205 & w18169) | (~pi0205 & w39519) | (w18169 & w39519);
assign w18205 = ~w18203 & ~w18204;
assign w18206 = pi0206 & ~w18193;
assign w18207 = w18190 & w18193;
assign w18208 = ~w18206 & ~w18207;
assign w18209 = pi0207 & ~w18193;
assign w18210 = w18184 & w18193;
assign w18211 = ~w18209 & ~w18210;
assign w18212 = w18193 & ~w18202;
assign w18213 = ~pi0208 & ~w18193;
assign w18214 = ~w18212 & ~w18213;
assign w18215 = ~pi0868 & w16106;
assign w18216 = w13185 & ~w13187;
assign w18217 = (~w12502 & w12037) | (~w12502 & w39520) | (w12037 & w39520);
assign w18218 = w18216 & ~w18217;
assign w18219 = ~w12502 & ~w13185;
assign w18220 = ~w16104 & w18219;
assign w18221 = ~w18218 & ~w18220;
assign w18222 = pi0868 & w18221;
assign w18223 = ~w18222 & w39521;
assign w18224 = w10749 & w40159;
assign w18225 = pi0209 & w10759;
assign w18226 = w15173 & ~w18225;
assign w18227 = ~w18224 & w18226;
assign w18228 = ~w18223 & ~w18227;
assign w18229 = ~w18222 & w39522;
assign w18230 = w13929 & w40159;
assign w18231 = pi0210 & w13933;
assign w18232 = w14336 & ~w18231;
assign w18233 = ~w18230 & w18232;
assign w18234 = ~w18229 & ~w18233;
assign w18235 = w10752 & ~w15996;
assign w18236 = (w341 & w39523) | (w341 & w39524) | (w39523 & w39524);
assign w18237 = ~w10753 & ~w18236;
assign w18238 = (w18237 & w16629) | (w18237 & w39525) | (w16629 & w39525);
assign w18239 = w15173 & ~w18238;
assign w18240 = ~w18235 & ~w18239;
assign w18241 = w13923 & ~w15996;
assign w18242 = (~pi0212 & ~w40144) | (~pi0212 & w39526) | (~w40144 & w39526);
assign w18243 = ~w13925 & ~w18242;
assign w18244 = (w18243 & w16629) | (w18243 & w39527) | (w16629 & w39527);
assign w18245 = w14336 & ~w18244;
assign w18246 = ~w18241 & ~w18245;
assign w18247 = (w15185 & w18222) | (w15185 & w39528) | (w18222 & w39528);
assign w18248 = (~pi0213 & ~w15184) | (~pi0213 & w39529) | (~w15184 & w39529);
assign w18249 = ~w18247 & ~w18248;
assign w18250 = (w15189 & w18222) | (w15189 & w39530) | (w18222 & w39530);
assign w18251 = ~pi0214 & ~w15189;
assign w18252 = ~w18250 & ~w18251;
assign w18253 = pi0868 & ~w17841;
assign w18254 = ~w12505 & w39531;
assign w18255 = (~w12495 & ~w13185) | (~w12495 & w39532) | (~w13185 & w39532);
assign w18256 = (w12503 & w12037) | (w12503 & w39533) | (w12037 & w39533);
assign w18257 = ~w12479 & ~w13186;
assign w18258 = ~pi0868 & w18257;
assign w18259 = (w18258 & w18256) | (w18258 & w39534) | (w18256 & w39534);
assign w18260 = pi0868 & w17841;
assign w18261 = (w18260 & w12505) | (w18260 & w39535) | (w12505 & w39535);
assign w18262 = ~w18259 & ~w18261;
assign w18263 = ~w18254 & w18262;
assign w18264 = ~pi0868 & ~w18257;
assign w18265 = (w10752 & w18256) | (w10752 & w39537) | (w18256 & w39537);
assign w18266 = w18262 & w39538;
assign w18267 = w10749 & w40176;
assign w18268 = pi0215 & w10759;
assign w18269 = w15173 & ~w18268;
assign w18270 = ~w18267 & w18269;
assign w18271 = ~w18266 & ~w18270;
assign w18272 = ~pi0868 & w18221;
assign w18273 = pi0868 & ~w18257;
assign w18274 = ~w18256 & w39539;
assign w18275 = pi0868 & w18257;
assign w18276 = (w18275 & w18256) | (w18275 & w39540) | (w18256 & w39540);
assign w18277 = ~w18274 & ~w18276;
assign w18278 = ~w18272 & w39541;
assign w18279 = pi0216 & w10759;
assign w18280 = w15173 & ~w18279;
assign w18281 = (w18280 & ~w13916) | (w18280 & w39542) | (~w13916 & w39542);
assign w18282 = ~w18278 & ~w18281;
assign w18283 = ~w18272 & w39543;
assign w18284 = pi0217 & w13933;
assign w18285 = w14336 & ~w18284;
assign w18286 = (w18285 & ~w13916) | (w18285 & w39544) | (~w13916 & w39544);
assign w18287 = ~w18283 & ~w18286;
assign w18288 = (w13923 & w18256) | (w13923 & w39545) | (w18256 & w39545);
assign w18289 = w18262 & w39546;
assign w18290 = w13929 & w40176;
assign w18291 = pi0218 & w13933;
assign w18292 = w14336 & ~w18291;
assign w18293 = ~w18290 & w18292;
assign w18294 = ~w18289 & ~w18293;
assign w18295 = (pi0219 & ~w15184) | (pi0219 & w39547) | (~w15184 & w39547);
assign w18296 = (w15185 & w18256) | (w15185 & w39548) | (w18256 & w39548);
assign w18297 = w18262 & w39549;
assign w18298 = ~w18295 & ~w18297;
assign w18299 = (pi0220 & ~w15184) | (pi0220 & w39550) | (~w15184 & w39550);
assign w18300 = ~w18272 & w39551;
assign w18301 = ~w18299 & ~w18300;
assign w18302 = (pi0221 & ~w15184) | (pi0221 & w39552) | (~w15184 & w39552);
assign w18303 = (w15189 & w18256) | (w15189 & w39553) | (w18256 & w39553);
assign w18304 = w18263 & w18303;
assign w18305 = ~w18302 & ~w18304;
assign w18306 = (pi0222 & ~w15184) | (pi0222 & w39554) | (~w15184 & w39554);
assign w18307 = ~w18272 & w39555;
assign w18308 = ~w18306 & ~w18307;
assign w18309 = pi1426 & ~w7;
assign w18310 = (~pi1426 & ~w9) | (~pi1426 & w39556) | (~w9 & w39556);
assign w18311 = ~w18309 & ~w18310;
assign w18312 = ~pi3438 & ~pi3472;
assign w18313 = ~pi3681 & w18312;
assign w18314 = w18312 & w39557;
assign w18315 = pi3641 & pi3681;
assign w18316 = pi1605 & pi1606;
assign w18317 = pi1681 & pi1704;
assign w18318 = w18316 & w18317;
assign w18319 = pi3641 & w18318;
assign w18320 = (~w18315 & ~w18318) | (~w18315 & w39558) | (~w18318 & w39558);
assign w18321 = pi0619 & pi0620;
assign w18322 = pi0691 & pi1370;
assign w18323 = w18321 & w18322;
assign w18324 = ~w18320 & w18323;
assign w18325 = ~w18320 & w39559;
assign w18326 = ~w18315 & ~w18325;
assign w18327 = (~pi0849 & w18325) | (~pi0849 & w39560) | (w18325 & w39560);
assign w18328 = (w18325 & w39561) | (w18325 & w39562) | (w39561 & w39562);
assign w18329 = (w18325 & w39563) | (w18325 & w39564) | (w39563 & w39564);
assign w18330 = ~pi0822 & w18329;
assign w18331 = (~w18315 & ~w18329) | (~w18315 & w39565) | (~w18329 & w39565);
assign w18332 = (w18329 & w39566) | (w18329 & w39567) | (w39566 & w39567);
assign w18333 = (w18329 & w39568) | (w18329 & w39569) | (w39568 & w39569);
assign w18334 = (w18329 & w39570) | (w18329 & w39571) | (w39570 & w39571);
assign w18335 = ~pi0496 & w18334;
assign w18336 = (~w18315 & ~w18334) | (~w18315 & w39572) | (~w18334 & w39572);
assign w18337 = (w18334 & w39573) | (w18334 & w39574) | (w39573 & w39574);
assign w18338 = (w18334 & w39575) | (w18334 & w39576) | (w39575 & w39576);
assign w18339 = (w18334 & w39577) | (w18334 & w39578) | (w39577 & w39578);
assign w18340 = (w18334 & w39579) | (w18334 & w39580) | (w39579 & w39580);
assign w18341 = (~pi0303 & w18340) | (~pi0303 & w39581) | (w18340 & w39581);
assign w18342 = (w18340 & w39585) | (w18340 & w39586) | (w39585 & w39586);
assign w18343 = ~pi0336 & ~pi0367;
assign w18344 = ~pi0398 & ~pi0458;
assign w18345 = w18343 & w18344;
assign w18346 = ~pi0223 & ~pi0246;
assign w18347 = ~pi0277 & ~pi0303;
assign w18348 = w18346 & w18347;
assign w18349 = w18345 & w18348;
assign w18350 = ~pi0728 & ~pi0822;
assign w18351 = ~pi0849 & ~pi0863;
assign w18352 = w18350 & w18351;
assign w18353 = ~pi0496 & ~pi0577;
assign w18354 = ~pi0653 & ~pi0699;
assign w18355 = w18353 & w18354;
assign w18356 = w18352 & w18355;
assign w18357 = w18349 & w18356;
assign w18358 = pi0827 & ~pi3681;
assign w18359 = w18357 & w18358;
assign w18360 = (w18340 & w39589) | (w18340 & w39590) | (w39589 & w39590);
assign w18361 = ~w18342 & w18360;
assign w18362 = (~w18313 & ~w18357) | (~w18313 & w39592) | (~w18357 & w39592);
assign w18363 = ~w18361 & w18362;
assign w18364 = ~w18314 & ~w18363;
assign w18365 = ~w17985 & w39593;
assign w18366 = pi0955 & ~pi2599;
assign w18367 = ~w18003 & w18366;
assign w18368 = w17971 & w18367;
assign w18369 = w17971 & w39594;
assign w18370 = ~w17985 & w39595;
assign w18371 = ~w17971 & w18370;
assign w18372 = (w5632 & w39596) | (w5632 & w39597) | (w39596 & w39597);
assign w18373 = ~pi0622 & w18003;
assign w18374 = ~w18003 & w39598;
assign w18375 = (w6668 & w39599) | (w6668 & w39600) | (w39599 & w39600);
assign w18376 = (w6668 & w39603) | (w6668 & w39604) | (w39603 & w39604);
assign w18377 = ~w18372 & w39605;
assign w18378 = ~w18369 & w18377;
assign w18379 = w17911 & w39606;
assign w18380 = ~w17976 & w18379;
assign w18381 = w18379 & w39607;
assign w18382 = (w17990 & ~w18379) | (w17990 & w39608) | (~w18379 & w39608);
assign w18383 = w17971 & w18382;
assign w18384 = (w18367 & w17971) | (w18367 & w39609) | (w17971 & w39609);
assign w18385 = ~w18383 & w18384;
assign w18386 = ~w5052 & w39610;
assign w18387 = ~pi0621 & w18003;
assign w18388 = (w6668 & w39613) | (w6668 & w39614) | (w39613 & w39614);
assign w18389 = ~w18386 & w18388;
assign w18390 = ~w18385 & w18389;
assign w18391 = pi0709 & w40192;
assign w18392 = (w17822 & w17005) | (w17822 & w39615) | (w17005 & w39615);
assign w18393 = (pi0226 & ~w17821) | (pi0226 & w39616) | (~w17821 & w39616);
assign w18394 = ~w18392 & ~w18393;
assign w18395 = (w17827 & w17005) | (w17827 & w39617) | (w17005 & w39617);
assign w18396 = pi0227 & ~w17827;
assign w18397 = ~w18395 & ~w18396;
assign w18398 = ~w15997 & w39618;
assign w18399 = (w341 & w39619) | (w341 & w39620) | (w39619 & w39620);
assign w18400 = ~w10753 & ~w18399;
assign w18401 = (w18400 & w16739) | (w18400 & w39621) | (w16739 & w39621);
assign w18402 = w15173 & ~w18401;
assign w18403 = ~w18398 & ~w18402;
assign w18404 = ~w15997 & w39622;
assign w18405 = (~pi0229 & ~w40144) | (~pi0229 & w39623) | (~w40144 & w39623);
assign w18406 = ~w13925 & ~w18405;
assign w18407 = (w18406 & w16739) | (w18406 & w39624) | (w16739 & w39624);
assign w18408 = w14336 & ~w18407;
assign w18409 = ~w18404 & ~w18408;
assign w18410 = pi1953 & w9958;
assign w18411 = ~w10613 & w39625;
assign w18412 = w10750 & w18411;
assign w18413 = (pi0230 & ~w18411) | (pi0230 & w39626) | (~w18411 & w39626);
assign w18414 = w15776 & ~w17425;
assign w18415 = ~w16574 & w17425;
assign w18416 = ~w18414 & ~w18415;
assign w18417 = w18412 & ~w18416;
assign w18418 = ~w18413 & ~w18417;
assign w18419 = w13922 & w18411;
assign w18420 = (pi0231 & ~w18411) | (pi0231 & w39627) | (~w18411 & w39627);
assign w18421 = ~w18416 & w18419;
assign w18422 = ~w18420 & ~w18421;
assign w18423 = pi0232 & ~w18375;
assign w18424 = ~w17980 & ~w18379;
assign w18425 = ~w18380 & ~w18424;
assign w18426 = ~w17971 & w18425;
assign w18427 = (w18366 & ~w17971) | (w18366 & w39628) | (~w17971 & w39628);
assign w18428 = ~w18426 & w18427;
assign w18429 = (~w18003 & w6176) | (~w18003 & w39630) | (w6176 & w39630);
assign w18430 = ~w18428 & w18429;
assign w18431 = pi0631 & w18003;
assign w18432 = (w6668 & w39631) | (w6668 & w39632) | (w39631 & w39632);
assign w18433 = ~w18430 & w18432;
assign w18434 = ~w18423 & ~w18433;
assign w18435 = (w5632 & w39633) | (w5632 & w39634) | (w39633 & w39634);
assign w18436 = (w16944 & w39635) | (w16944 & w39636) | (w39635 & w39636);
assign w18437 = w17822 & ~w18436;
assign w18438 = (pi0233 & ~w17821) | (pi0233 & w39637) | (~w17821 & w39637);
assign w18439 = ~w18437 & ~w18438;
assign w18440 = w17827 & ~w18436;
assign w18441 = (pi0234 & ~w17821) | (pi0234 & w39638) | (~w17821 & w39638);
assign w18442 = ~w18440 & ~w18441;
assign w18443 = ~pi0710 & pi2140;
assign w18444 = ~w10613 & w39639;
assign w18445 = w10750 & w18444;
assign w18446 = (w6176 & w39640) | (w6176 & w39641) | (w39640 & w39641);
assign w18447 = w16218 & w39642;
assign w18448 = (w18445 & w18447) | (w18445 & w39643) | (w18447 & w39643);
assign w18449 = (~pi0235 & ~w18444) | (~pi0235 & w39644) | (~w18444 & w39644);
assign w18450 = ~w18448 & ~w18449;
assign w18451 = w13922 & w18444;
assign w18452 = (w18451 & w18447) | (w18451 & w39645) | (w18447 & w39645);
assign w18453 = ~pi0236 & ~w18451;
assign w18454 = ~w18452 & ~w18453;
assign w18455 = ~pi0237 & ~w18375;
assign w18456 = (~w17993 & ~w18379) | (~w17993 & w39646) | (~w18379 & w39646);
assign w18457 = ~w18381 & ~w18456;
assign w18458 = ~w17971 & ~w18457;
assign w18459 = (w18366 & ~w17971) | (w18366 & w39647) | (~w17971 & w39647);
assign w18460 = ~w18458 & w18459;
assign w18461 = ~w18003 & w40200;
assign w18462 = ~w18460 & w18461;
assign w18463 = ~pi0608 & w18003;
assign w18464 = (w6668 & w39649) | (w6668 & w39650) | (w39649 & w39650);
assign w18465 = ~w18462 & w18464;
assign w18466 = ~w18455 & ~w18465;
assign w18467 = pi0709 & w40191;
assign w18468 = (~w18467 & w16192) | (~w18467 & w39651) | (w16192 & w39651);
assign w18469 = w17822 & ~w18468;
assign w18470 = (pi0238 & ~w17821) | (pi0238 & w39652) | (~w17821 & w39652);
assign w18471 = ~w18469 & ~w18470;
assign w18472 = w17827 & ~w18468;
assign w18473 = (pi0239 & ~w17821) | (pi0239 & w39653) | (~w17821 & w39653);
assign w18474 = ~w18472 & ~w18473;
assign w18475 = (w10752 & w16009) | (w10752 & w39654) | (w16009 & w39654);
assign w18476 = (w1307 & w39655) | (w1307 & w39656) | (w39655 & w39656);
assign w18477 = (w341 & w39657) | (w341 & w39658) | (w39657 & w39658);
assign w18478 = ~w10753 & ~w18477;
assign w18479 = (w15173 & w18476) | (w15173 & w39659) | (w18476 & w39659);
assign w18480 = ~w18475 & ~w18479;
assign w18481 = (w13923 & w16009) | (w13923 & w39660) | (w16009 & w39660);
assign w18482 = (w1307 & w39661) | (w1307 & w39662) | (w39661 & w39662);
assign w18483 = (~pi0241 & ~w40144) | (~pi0241 & w39663) | (~w40144 & w39663);
assign w18484 = ~w13925 & ~w18483;
assign w18485 = (w14336 & w18482) | (w14336 & w39664) | (w18482 & w39664);
assign w18486 = ~w18481 & ~w18485;
assign w18487 = (pi0242 & ~w18411) | (pi0242 & w39665) | (~w18411 & w39665);
assign w18488 = ~w16574 & ~w17425;
assign w18489 = w17425 & w17668;
assign w18490 = ~w18488 & ~w18489;
assign w18491 = w18412 & ~w18490;
assign w18492 = ~w18487 & ~w18491;
assign w18493 = (pi0243 & ~w18411) | (pi0243 & w39666) | (~w18411 & w39666);
assign w18494 = ~w17425 & ~w17668;
assign w18495 = ~w16773 & w17425;
assign w18496 = ~w18494 & ~w18495;
assign w18497 = w18412 & w18496;
assign w18498 = ~w18493 & ~w18497;
assign w18499 = (pi0244 & ~w18411) | (pi0244 & w39667) | (~w18411 & w39667);
assign w18500 = w18419 & ~w18490;
assign w18501 = ~w18499 & ~w18500;
assign w18502 = (pi0245 & ~w18411) | (pi0245 & w39668) | (~w18411 & w39668);
assign w18503 = w18419 & w18496;
assign w18504 = ~w18502 & ~w18503;
assign w18505 = w18312 & w39669;
assign w18506 = pi0246 & w40201;
assign w18507 = ~w18359 & w40202;
assign w18508 = ~w18506 & w18507;
assign w18509 = (~w18313 & ~w18357) | (~w18313 & w39671) | (~w18357 & w39671);
assign w18510 = ~w18508 & w18509;
assign w18511 = ~w18505 & ~w18510;
assign w18512 = ~pi0247 & w18012;
assign w18513 = (w17983 & ~w17911) | (w17983 & w39672) | (~w17911 & w39672);
assign w18514 = ~w18379 & ~w18513;
assign w18515 = ~w17971 & ~w18514;
assign w18516 = (pi0955 & ~w17971) | (pi0955 & w39673) | (~w17971 & w39673);
assign w18517 = ~w18515 & w18516;
assign w18518 = ~pi0247 & ~pi0955;
assign w18519 = w18004 & ~w18518;
assign w18520 = ~w18517 & w18519;
assign w18521 = ~pi0630 & w18003;
assign w18522 = (w6668 & w39675) | (w6668 & w39676) | (w39675 & w39676);
assign w18523 = (w18522 & w3194) | (w18522 & w39677) | (w3194 & w39677);
assign w18524 = ~w18520 & w18523;
assign w18525 = ~w18512 & ~w18524;
assign w18526 = ~w17929 & w17969;
assign w18527 = ~w17970 & ~w18526;
assign w18528 = w18367 & ~w18527;
assign w18529 = pi0629 & w18003;
assign w18530 = ~w18529 & w40203;
assign w18531 = (~w18012 & w18528) | (~w18012 & w39680) | (w18528 & w39680);
assign w18532 = ~pi0248 & ~w18375;
assign w18533 = ~w18531 & ~w18532;
assign w18534 = (w4140 & w39681) | (w4140 & w39682) | (w39681 & w39682);
assign w18535 = w16517 & w39642;
assign w18536 = (w18445 & w18535) | (w18445 & w39683) | (w18535 & w39683);
assign w18537 = (~pi0249 & ~w18444) | (~pi0249 & w39684) | (~w18444 & w39684);
assign w18538 = ~w18536 & ~w18537;
assign w18539 = (w3194 & w39685) | (w3194 & w39686) | (w39685 & w39686);
assign w18540 = w16307 & w39642;
assign w18541 = (w18445 & w18540) | (w18445 & w39687) | (w18540 & w39687);
assign w18542 = (~pi0250 & ~w18444) | (~pi0250 & w39688) | (~w18444 & w39688);
assign w18543 = ~w18541 & ~w18542;
assign w18544 = (pi0251 & ~w18444) | (pi0251 & w39689) | (~w18444 & w39689);
assign w18545 = pi0710 & ~w10746;
assign w18546 = (~pi0710 & ~w15866) | (~pi0710 & w39690) | (~w15866 & w39690);
assign w18547 = (w18445 & w18546) | (w18445 & w39691) | (w18546 & w39691);
assign w18548 = ~w18544 & ~w18547;
assign w18549 = (w18451 & w18535) | (w18451 & w39692) | (w18535 & w39692);
assign w18550 = ~pi0252 & ~w18451;
assign w18551 = ~w18549 & ~w18550;
assign w18552 = (w18451 & w18540) | (w18451 & w39693) | (w18540 & w39693);
assign w18553 = ~pi0253 & ~w18451;
assign w18554 = ~w18552 & ~w18553;
assign w18555 = (pi0254 & ~w18444) | (pi0254 & w39694) | (~w18444 & w39694);
assign w18556 = (w18451 & w18546) | (w18451 & w39695) | (w18546 & w39695);
assign w18557 = ~w18555 & ~w18556;
assign w18558 = w10752 & w16014;
assign w18559 = w18039 & ~w15978;
assign w18560 = (w341 & w39696) | (w341 & w39697) | (w39696 & w39697);
assign w18561 = ~w10753 & ~w18560;
assign w18562 = (w15173 & w18559) | (w15173 & w39698) | (w18559 & w39698);
assign w18563 = ~w18558 & ~w18562;
assign w18564 = (w10752 & w16026) | (w10752 & w39699) | (w16026 & w39699);
assign w18565 = (w5052 & w39700) | (w5052 & w39701) | (w39700 & w39701);
assign w18566 = (w341 & w39702) | (w341 & w39703) | (w39702 & w39703);
assign w18567 = ~w10753 & ~w18566;
assign w18568 = (w15173 & w18565) | (w15173 & w39704) | (w18565 & w39704);
assign w18569 = ~w18564 & ~w18568;
assign w18570 = w13923 & w16014;
assign w18571 = w18046 & ~w15978;
assign w18572 = (~pi0257 & ~w40144) | (~pi0257 & w39705) | (~w40144 & w39705);
assign w18573 = ~w13925 & ~w18572;
assign w18574 = (w14336 & w18571) | (w14336 & w39706) | (w18571 & w39706);
assign w18575 = ~w18570 & ~w18574;
assign w18576 = (w13923 & w16026) | (w13923 & w39707) | (w16026 & w39707);
assign w18577 = (~pi0258 & ~w40144) | (~pi0258 & w39708) | (~w40144 & w39708);
assign w18578 = ~w13925 & ~w18577;
assign w18579 = (w18578 & w15171) | (w18578 & w39709) | (w15171 & w39709);
assign w18580 = w14336 & ~w18579;
assign w18581 = ~w18576 & ~w18580;
assign w18582 = pi0709 & w14962;
assign w18583 = (w17822 & w15600) | (w17822 & w39710) | (w15600 & w39710);
assign w18584 = (pi0259 & ~w17821) | (pi0259 & w39711) | (~w17821 & w39711);
assign w18585 = ~w18583 & ~w18584;
assign w18586 = pi0709 & w14325;
assign w18587 = (w17822 & w15494) | (w17822 & w39712) | (w15494 & w39712);
assign w18588 = (pi0260 & ~w17821) | (pi0260 & w39713) | (~w17821 & w39713);
assign w18589 = ~w18587 & ~w18588;
assign w18590 = pi0709 & w16739;
assign w18591 = (w17822 & w16715) | (w17822 & w39714) | (w16715 & w39714);
assign w18592 = (pi0261 & ~w17821) | (pi0261 & w39715) | (~w17821 & w39715);
assign w18593 = ~w18591 & ~w18592;
assign w18594 = pi0709 & w40171;
assign w18595 = (~w18594 & w17122) | (~w18594 & w39716) | (w17122 & w39716);
assign w18596 = w17822 & ~w18595;
assign w18597 = (pi0262 & ~w17821) | (pi0262 & w39717) | (~w17821 & w39717);
assign w18598 = ~w18596 & ~w18597;
assign w18599 = (w17827 & w15600) | (w17827 & w39718) | (w15600 & w39718);
assign w18600 = pi0263 & ~w17827;
assign w18601 = ~w18599 & ~w18600;
assign w18602 = (w17827 & w15494) | (w17827 & w39719) | (w15494 & w39719);
assign w18603 = pi0264 & ~w17827;
assign w18604 = ~w18602 & ~w18603;
assign w18605 = (w17827 & w16715) | (w17827 & w39720) | (w16715 & w39720);
assign w18606 = pi0265 & ~w17827;
assign w18607 = ~w18605 & ~w18606;
assign w18608 = w17827 & ~w18595;
assign w18609 = (pi0266 & ~w17821) | (pi0266 & w39721) | (~w17821 & w39721);
assign w18610 = ~w18608 & ~w18609;
assign w18611 = (w10752 & w16024) | (w10752 & w39722) | (w16024 & w39722);
assign w18612 = (w4140 & w39723) | (w4140 & w39724) | (w39723 & w39724);
assign w18613 = (w341 & w39725) | (w341 & w39726) | (w39725 & w39726);
assign w18614 = ~w10753 & ~w18613;
assign w18615 = (w15173 & w18612) | (w15173 & w39727) | (w18612 & w39727);
assign w18616 = ~w18611 & ~w18615;
assign w18617 = (w13923 & w16024) | (w13923 & w39728) | (w16024 & w39728);
assign w18618 = (w4140 & w39729) | (w4140 & w39730) | (w39729 & w39730);
assign w18619 = (~pi0268 & ~w40144) | (~pi0268 & w39731) | (~w40144 & w39731);
assign w18620 = ~w13925 & ~w18619;
assign w18621 = (w14336 & w18618) | (w14336 & w39732) | (w18618 & w39732);
assign w18622 = ~w18617 & ~w18621;
assign w18623 = pi0709 & w40168;
assign w18624 = (~w18623 & w15703) | (~w18623 & w39733) | (w15703 & w39733);
assign w18625 = w17822 & ~w18624;
assign w18626 = (pi0269 & ~w17821) | (pi0269 & w39734) | (~w17821 & w39734);
assign w18627 = ~w18625 & ~w18626;
assign w18628 = w17827 & ~w18624;
assign w18629 = (pi0270 & ~w17821) | (pi0270 & w39735) | (~w17821 & w39735);
assign w18630 = ~w18628 & ~w18629;
assign w18631 = pi0710 & ~w16842;
assign w18632 = (~w18631 & w16798) | (~w18631 & w39736) | (w16798 & w39736);
assign w18633 = w18445 & ~w18632;
assign w18634 = (pi0271 & ~w18444) | (pi0271 & w39737) | (~w18444 & w39737);
assign w18635 = ~w18633 & ~w18634;
assign w18636 = w18451 & ~w18632;
assign w18637 = (pi0272 & ~w18444) | (pi0272 & w39738) | (~w18444 & w39738);
assign w18638 = ~w18636 & ~w18637;
assign w18639 = (pi0273 & ~w18411) | (pi0273 & w39739) | (~w18411 & w39739);
assign w18640 = w16773 & ~w17425;
assign w18641 = w17425 & w17669;
assign w18642 = (w18412 & w18640) | (w18412 & w39740) | (w18640 & w39740);
assign w18643 = ~w18639 & ~w18642;
assign w18644 = (pi0274 & ~w18411) | (pi0274 & w39741) | (~w18411 & w39741);
assign w18645 = ~w16984 & w17425;
assign w18646 = ~w17425 & w17669;
assign w18647 = (w18412 & w18646) | (w18412 & w39742) | (w18646 & w39742);
assign w18648 = ~w18644 & ~w18647;
assign w18649 = (pi0275 & ~w18411) | (pi0275 & w39743) | (~w18411 & w39743);
assign w18650 = (w18419 & w18640) | (w18419 & w39744) | (w18640 & w39744);
assign w18651 = ~w18649 & ~w18650;
assign w18652 = (pi0276 & ~w18411) | (pi0276 & w39745) | (~w18411 & w39745);
assign w18653 = (w18419 & w18646) | (w18419 & w39746) | (w18646 & w39746);
assign w18654 = ~w18652 & ~w18653;
assign w18655 = w18312 & w39747;
assign w18656 = pi0277 & ~w18341;
assign w18657 = ~w18359 & w40201;
assign w18658 = ~w18656 & w18657;
assign w18659 = (~w18313 & ~w18357) | (~w18313 & w39749) | (~w18357 & w39749);
assign w18660 = ~w18658 & w18659;
assign w18661 = ~w18655 & ~w18660;
assign w18662 = (~pi0247 & w17960) | (~pi0247 & w39750) | (w17960 & w39750);
assign w18663 = w17931 & w18662;
assign w18664 = (w18367 & w18662) | (w18367 & w39751) | (w18662 & w39751);
assign w18665 = ~w18663 & w18664;
assign w18666 = w18009 & ~w6413;
assign w18667 = pi0611 & w18003;
assign w18668 = (w6668 & w39754) | (w6668 & w39755) | (w39754 & w39755);
assign w18669 = ~w18666 & w18668;
assign w18670 = ~w18665 & w18669;
assign w18671 = pi0709 & w40174;
assign w18672 = (w17822 & w16294) | (w17822 & w39756) | (w16294 & w39756);
assign w18673 = (pi0279 & ~w17821) | (pi0279 & w39757) | (~w17821 & w39757);
assign w18674 = ~w18672 & ~w18673;
assign w18675 = (w17827 & w16294) | (w17827 & w39758) | (w16294 & w39758);
assign w18676 = pi0280 & ~w17827;
assign w18677 = ~w18675 & ~w18676;
assign w18678 = pi0710 & ~w15978;
assign w18679 = (~w18678 & ~w16922) | (~w18678 & w39759) | (~w16922 & w39759);
assign w18680 = w18445 & ~w18679;
assign w18681 = (~pi0281 & ~w18444) | (~pi0281 & w39760) | (~w18444 & w39760);
assign w18682 = ~w18680 & ~w18681;
assign w18683 = (w5052 & w39761) | (w5052 & w39762) | (w39761 & w39762);
assign w18684 = w17028 & w39763;
assign w18685 = (w18445 & w18684) | (w18445 & w39764) | (w18684 & w39764);
assign w18686 = (~pi0282 & ~w18444) | (~pi0282 & w39765) | (~w18444 & w39765);
assign w18687 = ~w18685 & ~w18686;
assign w18688 = (w16922 & w39766) | (w16922 & w39767) | (w39766 & w39767);
assign w18689 = (~pi0283 & ~w18444) | (~pi0283 & w39768) | (~w18444 & w39768);
assign w18690 = ~w18688 & ~w18689;
assign w18691 = (w18451 & w18684) | (w18451 & w39769) | (w18684 & w39769);
assign w18692 = ~pi0284 & ~w18451;
assign w18693 = ~w18691 & ~w18692;
assign w18694 = pi0709 & ~w10746;
assign w18695 = (~w18694 & w15836) | (~w18694 & w39770) | (w15836 & w39770);
assign w18696 = w17822 & ~w18695;
assign w18697 = (pi0285 & ~w17821) | (pi0285 & w39771) | (~w17821 & w39771);
assign w18698 = ~w18696 & ~w18697;
assign w18699 = w17827 & ~w18695;
assign w18700 = (pi0286 & ~w17821) | (pi0286 & w39772) | (~w17821 & w39772);
assign w18701 = ~w18699 & ~w18700;
assign w18702 = pi0710 & ~w14325;
assign w18703 = w15531 & w39773;
assign w18704 = (w18445 & w18703) | (w18445 & w39774) | (w18703 & w39774);
assign w18705 = (~pi0287 & ~w18444) | (~pi0287 & w39775) | (~w18444 & w39775);
assign w18706 = ~w18704 & ~w18705;
assign w18707 = pi0710 & ~w14962;
assign w18708 = w15632 & w39776;
assign w18709 = (w18445 & w18708) | (w18445 & w39777) | (w18708 & w39777);
assign w18710 = (~pi0288 & ~w18444) | (~pi0288 & w39778) | (~w18444 & w39778);
assign w18711 = ~w18709 & ~w18710;
assign w18712 = (w4748 & w39779) | (w4748 & w39780) | (w39779 & w39780);
assign w18713 = w15097 & w39781;
assign w18714 = (w18445 & w18713) | (w18445 & w39782) | (w18713 & w39782);
assign w18715 = (~pi0289 & ~w18444) | (~pi0289 & w39783) | (~w18444 & w39783);
assign w18716 = ~w18714 & ~w18715;
assign w18717 = (w18451 & w18703) | (w18451 & w39784) | (w18703 & w39784);
assign w18718 = ~pi0290 & ~w18451;
assign w18719 = ~w18717 & ~w18718;
assign w18720 = (w18451 & w18708) | (w18451 & w39785) | (w18708 & w39785);
assign w18721 = ~pi0291 & ~w18451;
assign w18722 = ~w18720 & ~w18721;
assign w18723 = (w18451 & w18713) | (w18451 & w39786) | (w18713 & w39786);
assign w18724 = ~pi0292 & ~w18451;
assign w18725 = ~w18723 & ~w18724;
assign w18726 = w10752 & w16031;
assign w18727 = (w6176 & w39787) | (w6176 & w39788) | (w39787 & w39788);
assign w18728 = (w341 & w39789) | (w341 & w39790) | (w39789 & w39790);
assign w18729 = ~w10753 & ~w18728;
assign w18730 = (w15173 & w18727) | (w15173 & w39791) | (w18727 & w39791);
assign w18731 = ~w18726 & ~w18730;
assign w18732 = w13923 & w16031;
assign w18733 = (w6176 & w39792) | (w6176 & w39793) | (w39792 & w39793);
assign w18734 = (~pi0294 & ~w40144) | (~pi0294 & w39794) | (~w40144 & w39794);
assign w18735 = ~w13925 & ~w18734;
assign w18736 = (w14336 & w18733) | (w14336 & w39795) | (w18733 & w39795);
assign w18737 = ~w18732 & ~w18736;
assign w18738 = (pi0295 & ~w18411) | (pi0295 & w39796) | (~w18411 & w39796);
assign w18739 = ~w16984 & ~w17425;
assign w18740 = w16464 & w17425;
assign w18741 = ~w18739 & ~w18740;
assign w18742 = w18412 & ~w18741;
assign w18743 = ~w18738 & ~w18742;
assign w18744 = (pi0296 & ~w18411) | (pi0296 & w39797) | (~w18411 & w39797);
assign w18745 = w18419 & ~w18741;
assign w18746 = ~w18744 & ~w18745;
assign w18747 = pi0709 & w16629;
assign w18748 = (~w18747 & w16594) | (~w18747 & w39798) | (w16594 & w39798);
assign w18749 = w17822 & ~w18748;
assign w18750 = (pi0297 & ~w17821) | (pi0297 & w39799) | (~w17821 & w39799);
assign w18751 = ~w18749 & ~w18750;
assign w18752 = w17827 & ~w18748;
assign w18753 = (pi0298 & ~w17821) | (pi0298 & w39800) | (~w17821 & w39800);
assign w18754 = ~w18752 & ~w18753;
assign w18755 = pi0710 & ~w13916;
assign w18756 = (~w18755 & ~w14796) | (~w18755 & w39801) | (~w14796 & w39801);
assign w18757 = w18445 & ~w18756;
assign w18758 = (~pi0299 & ~w18444) | (~pi0299 & w39802) | (~w18444 & w39802);
assign w18759 = ~w18757 & ~w18758;
assign w18760 = (w14796 & w39803) | (w14796 & w39804) | (w39803 & w39804);
assign w18761 = (~pi0300 & ~w18444) | (~pi0300 & w39805) | (~w18444 & w39805);
assign w18762 = ~w18760 & ~w18761;
assign w18763 = (pi0301 & ~w18411) | (pi0301 & w39806) | (~w18411 & w39806);
assign w18764 = w16159 & w17425;
assign w18765 = w16464 & ~w17425;
assign w18766 = ~w18764 & ~w18765;
assign w18767 = w18412 & ~w18766;
assign w18768 = ~w18763 & ~w18767;
assign w18769 = (pi0302 & ~w18411) | (pi0302 & w39807) | (~w18411 & w39807);
assign w18770 = w18419 & ~w18766;
assign w18771 = ~w18769 & ~w18770;
assign w18772 = w18312 & w39808;
assign w18773 = ~w18340 & w39809;
assign w18774 = ~w18341 & ~w18359;
assign w18775 = ~w18773 & w18774;
assign w18776 = (~w18313 & ~w18357) | (~w18313 & w39811) | (~w18357 & w39811);
assign w18777 = ~w18775 & w18776;
assign w18778 = ~w18772 & ~w18777;
assign w18779 = pi0709 & w40176;
assign w18780 = (~w18779 & w16379) | (~w18779 & w39812) | (w16379 & w39812);
assign w18781 = w17822 & ~w18780;
assign w18782 = (pi0304 & ~w17821) | (pi0304 & w39813) | (~w17821 & w39813);
assign w18783 = ~w18781 & ~w18782;
assign w18784 = pi0709 & w40159;
assign w18785 = (~w18784 & w15063) | (~w18784 & w39814) | (w15063 & w39814);
assign w18786 = w17822 & ~w18785;
assign w18787 = (pi0305 & ~w17821) | (pi0305 & w39815) | (~w17821 & w39815);
assign w18788 = ~w18786 & ~w18787;
assign w18789 = w17827 & ~w18780;
assign w18790 = (pi0306 & ~w17821) | (pi0306 & w39816) | (~w17821 & w39816);
assign w18791 = ~w18789 & ~w18790;
assign w18792 = w17827 & ~w18785;
assign w18793 = (pi0307 & ~w17821) | (pi0307 & w39817) | (~w17821 & w39817);
assign w18794 = ~w18792 & ~w18793;
assign w18795 = pi0710 & ~w16739;
assign w18796 = (~w18795 & ~w16732) | (~w18795 & w39818) | (~w16732 & w39818);
assign w18797 = w18445 & ~w18796;
assign w18798 = (~pi0308 & ~w18444) | (~pi0308 & w39819) | (~w18444 & w39819);
assign w18799 = ~w18797 & ~w18798;
assign w18800 = (w3710 & w39820) | (w3710 & w39821) | (w39820 & w39821);
assign w18801 = w17166 & w39822;
assign w18802 = (w18445 & w18801) | (w18445 & w39823) | (w18801 & w39823);
assign w18803 = (~pi0309 & ~w18444) | (~pi0309 & w39824) | (~w18444 & w39824);
assign w18804 = ~w18802 & ~w18803;
assign w18805 = (w16732 & w39825) | (w16732 & w39826) | (w39825 & w39826);
assign w18806 = (~pi0310 & ~w18444) | (~pi0310 & w39827) | (~w18444 & w39827);
assign w18807 = ~w18805 & ~w18806;
assign w18808 = (w18451 & w18801) | (w18451 & w39828) | (w18801 & w39828);
assign w18809 = ~pi0311 & ~w18451;
assign w18810 = ~w18808 & ~w18809;
assign w18811 = (w10752 & w16032) | (w10752 & w39829) | (w16032 & w39829);
assign w18812 = (w3194 & w39830) | (w3194 & w39831) | (w39830 & w39831);
assign w18813 = (w341 & w39832) | (w341 & w39833) | (w39832 & w39833);
assign w18814 = ~w10753 & ~w18813;
assign w18815 = (w15173 & w18812) | (w15173 & w39834) | (w18812 & w39834);
assign w18816 = ~w18811 & ~w18815;
assign w18817 = (w13923 & w16032) | (w13923 & w39835) | (w16032 & w39835);
assign w18818 = (w3194 & w39836) | (w3194 & w39837) | (w39836 & w39837);
assign w18819 = (~pi0313 & ~w40144) | (~pi0313 & w39838) | (~w40144 & w39838);
assign w18820 = ~w13925 & ~w18819;
assign w18821 = (w14336 & w18818) | (w14336 & w39839) | (w18818 & w39839);
assign w18822 = ~w18817 & ~w18821;
assign w18823 = (w15277 & ~w15303) | (w15277 & w39840) | (~w15303 & w39840);
assign w18824 = w15394 & ~w18823;
assign w18825 = (w6410 & w39841) | (w6410 & w39842) | (w39841 & w39842);
assign w18826 = (w6668 & w39845) | (w6668 & w39846) | (w39845 & w39846);
assign w18827 = ~w18825 & w18826;
assign w18828 = (~w18827 & ~w18823) | (~w18827 & w39847) | (~w18823 & w39847);
assign w18829 = ~w18824 & w18828;
assign w18830 = pi0709 & w13916;
assign w18831 = (w17822 & w14729) | (w17822 & w39848) | (w14729 & w39848);
assign w18832 = (pi0315 & ~w17821) | (pi0315 & w39849) | (~w17821 & w39849);
assign w18833 = ~w18831 & ~w18832;
assign w18834 = (w17827 & w14729) | (w17827 & w39850) | (w14729 & w39850);
assign w18835 = pi0316 & ~w17827;
assign w18836 = ~w18834 & ~w18835;
assign w18837 = (w4379 & w39851) | (w4379 & w39852) | (w39851 & w39852);
assign w18838 = w15736 & w39773;
assign w18839 = (w18445 & w18838) | (w18445 & w39853) | (w18838 & w39853);
assign w18840 = (~pi0317 & ~w18444) | (~pi0317 & w39854) | (~w18444 & w39854);
assign w18841 = ~w18839 & ~w18840;
assign w18842 = pi0710 & ~w16629;
assign w18843 = w16620 & w39855;
assign w18844 = (w18445 & w18843) | (w18445 & w39856) | (w18843 & w39856);
assign w18845 = (~pi0318 & ~w18444) | (~pi0318 & w39857) | (~w18444 & w39857);
assign w18846 = ~w18844 & ~w18845;
assign w18847 = (w18451 & w18838) | (w18451 & w39858) | (w18838 & w39858);
assign w18848 = ~pi0319 & ~w18451;
assign w18849 = ~w18847 & ~w18848;
assign w18850 = (w18451 & w18843) | (w18451 & w39859) | (w18843 & w39859);
assign w18851 = ~pi0320 & ~w18451;
assign w18852 = ~w18850 & ~w18851;
assign w18853 = (pi0321 & ~w18411) | (pi0321 & w39860) | (~w18411 & w39860);
assign w18854 = ~w16272 & w17425;
assign w18855 = w16159 & ~w17425;
assign w18856 = ~w18854 & ~w18855;
assign w18857 = w18412 & ~w18856;
assign w18858 = ~w18853 & ~w18857;
assign w18859 = (pi0322 & ~w18411) | (pi0322 & w39861) | (~w18411 & w39861);
assign w18860 = w18419 & ~w18856;
assign w18861 = ~w18859 & ~w18860;
assign w18862 = (w5319 & w39862) | (w5319 & w39863) | (w39862 & w39863);
assign w18863 = (~w18862 & ~w16427) | (~w18862 & w39864) | (~w16427 & w39864);
assign w18864 = w18445 & ~w18863;
assign w18865 = (~pi0323 & ~w18444) | (~pi0323 & w39865) | (~w18444 & w39865);
assign w18866 = ~w18864 & ~w18865;
assign w18867 = (w16427 & w39866) | (w16427 & w39867) | (w39866 & w39867);
assign w18868 = (~pi0324 & ~w18444) | (~pi0324 & w39868) | (~w18444 & w39868);
assign w18869 = ~w18867 & ~w18868;
assign w18870 = (w17425 & w15451) | (w17425 & w39869) | (w15451 & w39869);
assign w18871 = w16272 & ~w17425;
assign w18872 = ~w18870 & ~w18871;
assign w18873 = w18412 & ~w18872;
assign w18874 = (~pi0325 & ~w18411) | (~pi0325 & w39870) | (~w18411 & w39870);
assign w18875 = ~w18873 & ~w18874;
assign w18876 = w18419 & ~w18872;
assign w18877 = (~pi0326 & ~w18411) | (~pi0326 & w39871) | (~w18411 & w39871);
assign w18878 = ~w18876 & ~w18877;
assign w18879 = w10752 & ~w16043;
assign w18880 = (w341 & w39872) | (w341 & w39873) | (w39872 & w39873);
assign w18881 = ~w10753 & ~w18880;
assign w18882 = (w18881 & w14325) | (w18881 & w39874) | (w14325 & w39874);
assign w18883 = w15173 & ~w18882;
assign w18884 = ~w18879 & ~w18883;
assign w18885 = w13923 & ~w16043;
assign w18886 = (~pi0328 & ~w40144) | (~pi0328 & w39875) | (~w40144 & w39875);
assign w18887 = ~w13925 & ~w18886;
assign w18888 = (w18887 & w14325) | (w18887 & w39876) | (w14325 & w39876);
assign w18889 = w14336 & ~w18888;
assign w18890 = ~w18885 & ~w18889;
assign w18891 = pi0329 & w18012;
assign w18892 = (w18008 & w4379) | (w18008 & w39877) | (w4379 & w39877);
assign w18893 = w17960 & w17967;
assign w18894 = (pi0955 & w17960) | (pi0955 & w39878) | (w17960 & w39878);
assign w18895 = ~w18893 & w18894;
assign w18896 = pi0329 & ~pi0955;
assign w18897 = w18004 & ~w18896;
assign w18898 = pi0628 & w18003;
assign w18899 = (w6668 & w39879) | (w6668 & w39880) | (w39879 & w39880);
assign w18900 = (w18899 & w18895) | (w18899 & w39881) | (w18895 & w39881);
assign w18901 = ~w18892 & w18900;
assign w18902 = ~w18891 & ~w18901;
assign w18903 = (pi2555 & w17383) | (pi2555 & w39882) | (w17383 & w39882);
assign w18904 = w4380 & ~w15388;
assign w18905 = (w6668 & w39885) | (w6668 & w39886) | (w39885 & w39886);
assign w18906 = ~w18904 & w18905;
assign w18907 = ~w18903 & ~w18906;
assign w18908 = ~pi0627 & w18003;
assign w18909 = w17944 & w17959;
assign w18910 = (w18367 & w17959) | (w18367 & w39888) | (w17959 & w39888);
assign w18911 = ~w18909 & w18910;
assign w18912 = ~w18908 & ~w18911;
assign w18913 = (w18912 & w5319) | (w18912 & w39889) | (w5319 & w39889);
assign w18914 = ~w18012 & ~w18913;
assign w18915 = pi0331 & ~w18375;
assign w18916 = ~w18914 & ~w18915;
assign w18917 = w5209 & w5763;
assign w18918 = ~w6295 & w18072;
assign w18919 = w18917 & w18918;
assign w18920 = ~pi3516 & ~w1182;
assign w18921 = ~w3392 & ~w3567;
assign w18922 = ~w4327 & w4670;
assign w18923 = w18921 & w18922;
assign w18924 = w18920 & w18923;
assign w18925 = w14449 & w39890;
assign w18926 = pi0712 & ~w18925;
assign w18927 = (w18926 & ~w18924) | (w18926 & w39891) | (~w18924 & w39891);
assign w18928 = w10614 & w39892;
assign w18929 = pi0332 & ~w18928;
assign w18930 = pi0712 & ~w18109;
assign w18931 = ~pi0712 & w40171;
assign w18932 = ~w18930 & ~w18931;
assign w18933 = w18928 & ~w18932;
assign w18934 = ~w18929 & ~w18933;
assign w18935 = w10614 & w39893;
assign w18936 = pi0333 & ~w18935;
assign w18937 = ~w18932 & w18935;
assign w18938 = ~w18936 & ~w18937;
assign w18939 = w10752 & w16047;
assign w18940 = (w341 & w39894) | (w341 & w39895) | (w39894 & w39895);
assign w18941 = ~w10753 & ~w18940;
assign w18942 = (w18941 & w14962) | (w18941 & w39896) | (w14962 & w39896);
assign w18943 = w15173 & ~w18942;
assign w18944 = ~w18939 & ~w18943;
assign w18945 = w13923 & w16047;
assign w18946 = (~pi0335 & ~w40144) | (~pi0335 & w39897) | (~w40144 & w39897);
assign w18947 = ~w13925 & ~w18946;
assign w18948 = (w18947 & w14962) | (w18947 & w39898) | (w14962 & w39898);
assign w18949 = w14336 & ~w18948;
assign w18950 = ~w18945 & ~w18949;
assign w18951 = w18312 & w39899;
assign w18952 = pi0336 & ~w18339;
assign w18953 = ~w18340 & ~w18359;
assign w18954 = ~w18952 & w18953;
assign w18955 = (~w18313 & ~w18357) | (~w18313 & w39901) | (~w18357 & w39901);
assign w18956 = ~w18954 & w18955;
assign w18957 = ~w18951 & ~w18956;
assign w18958 = (pi0337 & ~w18411) | (pi0337 & w39902) | (~w18411 & w39902);
assign w18959 = ~w15451 & w39903;
assign w18960 = w15577 & w17425;
assign w18961 = (w18412 & w18959) | (w18412 & w39904) | (w18959 & w39904);
assign w18962 = ~w18958 & ~w18961;
assign w18963 = (pi0338 & ~w18411) | (pi0338 & w39905) | (~w18411 & w39905);
assign w18964 = ~w15679 & w17425;
assign w18965 = w15577 & ~w17425;
assign w18966 = ~w18964 & ~w18965;
assign w18967 = w18412 & ~w18966;
assign w18968 = ~w18963 & ~w18967;
assign w18969 = (pi0339 & ~w18411) | (pi0339 & w39906) | (~w18411 & w39906);
assign w18970 = (w18419 & w18959) | (w18419 & w39907) | (w18959 & w39907);
assign w18971 = ~w18969 & ~w18970;
assign w18972 = (pi0340 & ~w18411) | (pi0340 & w39908) | (~w18411 & w39908);
assign w18973 = w18419 & ~w18966;
assign w18974 = ~w18972 & ~w18973;
assign w18975 = w14387 & w39909;
assign w18976 = ~pi0713 & w18975;
assign w18977 = w15870 & w18976;
assign w18978 = ~pi0713 & ~pi0714;
assign w18979 = pi3245 & w14396;
assign w18980 = (~w18978 & w18979) | (~w18978 & w39910) | (w18979 & w39910);
assign w18981 = w15870 & w18980;
assign w18982 = w14392 & ~w18979;
assign w18983 = w15870 & ~w18982;
assign w18984 = ~pi3245 & w14395;
assign w18985 = ~pi3245 & ~w14376;
assign w18986 = (~w18985 & ~w14392) | (~w18985 & w39911) | (~w14392 & w39911);
assign w18987 = w15870 & w18986;
assign w18988 = ~w16048 & w39912;
assign w18989 = (w4379 & w39913) | (w4379 & w39914) | (w39913 & w39914);
assign w18990 = (w341 & w39915) | (w341 & w39916) | (w39915 & w39916);
assign w18991 = ~w10753 & ~w18990;
assign w18992 = (w15173 & w18989) | (w15173 & w39917) | (w18989 & w39917);
assign w18993 = ~w18988 & ~w18992;
assign w18994 = ~w16048 & w39918;
assign w18995 = (~pi0345 & ~w40144) | (~pi0345 & w39919) | (~w40144 & w39919);
assign w18996 = ~w13925 & ~w18995;
assign w18997 = (w18996 & w40168) | (w18996 & w39920) | (w40168 & w39920);
assign w18998 = w14336 & ~w18997;
assign w18999 = ~w18994 & ~w18998;
assign w19000 = w15679 & ~w17425;
assign w19001 = w16360 & w17425;
assign w19002 = (w18412 & w19000) | (w18412 & w39921) | (w19000 & w39921);
assign w19003 = (~pi0346 & ~w18411) | (~pi0346 & w39922) | (~w18411 & w39922);
assign w19004 = ~w19002 & ~w19003;
assign w19005 = (pi0347 & ~w18411) | (pi0347 & w39923) | (~w18411 & w39923);
assign w19006 = ~w16360 & ~w17425;
assign w19007 = (w14417 & w39924) | (w14417 & w39925) | (w39924 & w39925);
assign w19008 = ~w19006 & ~w19007;
assign w19009 = w18412 & ~w19008;
assign w19010 = ~w19005 & ~w19009;
assign w19011 = (w18419 & w19000) | (w18419 & w39926) | (w19000 & w39926);
assign w19012 = ~pi0348 & ~w18419;
assign w19013 = ~w19011 & ~w19012;
assign w19014 = (pi0349 & ~w18411) | (pi0349 & w39927) | (~w18411 & w39927);
assign w19015 = w18419 & ~w19008;
assign w19016 = ~w19014 & ~w19015;
assign w19017 = ~pi0626 & w18003;
assign w19018 = pi0247 & ~pi1017;
assign w19019 = ~w17953 & w19018;
assign w19020 = ~pi0247 & pi0248;
assign w19021 = ~w17950 & w19020;
assign w19022 = ~pi0329 & w17941;
assign w19023 = (~w19022 & w19021) | (~w19022 & w39930) | (w19021 & w39930);
assign w19024 = ~w17949 & w19023;
assign w19025 = ~w17948 & w39931;
assign w19026 = w18367 & ~w19025;
assign w19027 = ~w19024 & w19026;
assign w19028 = ~w19017 & ~w19027;
assign w19029 = (w5893 & w39932) | (w5893 & w39933) | (w39932 & w39933);
assign w19030 = ~w18012 & ~w19029;
assign w19031 = pi0350 & ~w18375;
assign w19032 = ~w19030 & ~w19031;
assign w19033 = pi0975 & ~pi1422;
assign w19034 = pi1770 & pi1855;
assign w19035 = pi1937 & w19034;
assign w19036 = w19033 & ~w19035;
assign w19037 = pi3428 & ~w19033;
assign w19038 = ~w19036 & ~w19037;
assign w19039 = ~w19036 & w39934;
assign w19040 = ~pi3147 & pi3578;
assign w19041 = pi3580 & w19040;
assign w19042 = (~w19033 & w19039) | (~w19033 & w39935) | (w19039 & w39935);
assign w19043 = pi0351 & ~w19042;
assign w19044 = w2251 & ~w7764;
assign w19045 = pi3567 & pi3574;
assign w19046 = pi3566 & w19045;
assign w19047 = pi3553 & pi3560;
assign w19048 = w19046 & w39937;
assign w19049 = pi3565 & pi3577;
assign w19050 = ~pi3564 & w19049;
assign w19051 = w19048 & w19050;
assign w19052 = pi3564 & pi3577;
assign w19053 = ~pi3565 & w19052;
assign w19054 = w19048 & w19053;
assign w19055 = ~w19051 & ~w19054;
assign w19056 = pi3563 & pi3564;
assign w19057 = pi3553 & w19056;
assign w19058 = w19049 & w19057;
assign w19059 = w19057 & w39938;
assign w19060 = ~pi3566 & w19045;
assign w19061 = w19059 & w19060;
assign w19062 = w19046 & w39939;
assign w19063 = ~pi3563 & w19052;
assign w19064 = w19062 & w19063;
assign w19065 = ~w19061 & ~w19064;
assign w19066 = w19055 & w19065;
assign w19067 = ~pi3567 & pi3574;
assign w19068 = w19059 & w39940;
assign w19069 = pi3567 & ~pi3574;
assign w19070 = w19059 & w39941;
assign w19071 = ~pi3577 & w19056;
assign w19072 = w19062 & w19071;
assign w19073 = w19045 & w39942;
assign w19074 = w19058 & w19073;
assign w19075 = ~w19072 & ~w19074;
assign w19076 = w19075 & w39943;
assign w19077 = w19066 & w19076;
assign w19078 = pi4024 & w19077;
assign w19079 = w19048 & w39944;
assign w19080 = w19048 & w39945;
assign w19081 = ~w19079 & ~w19080;
assign w19082 = w19059 & w39946;
assign w19083 = w19062 & w39947;
assign w19084 = ~w19082 & ~w19083;
assign w19085 = w19081 & w19084;
assign w19086 = w19059 & w39948;
assign w19087 = w19059 & w39949;
assign w19088 = w19062 & w39950;
assign w19089 = w19058 & w39951;
assign w19090 = ~w19088 & ~w19089;
assign w19091 = w19090 & w39952;
assign w19092 = w19085 & w19091;
assign w19093 = ~w19078 & w19092;
assign w19094 = ~w2249 & w2250;
assign w19095 = ~w19078 & w39953;
assign w19096 = ~pi2515 & pi3445;
assign w19097 = (w19039 & w39954) | (w19039 & w39955) | (w39954 & w39955);
assign w19098 = ~w19095 & w19097;
assign w19099 = ~w19044 & w19098;
assign w19100 = w19099 & w40204;
assign w19101 = ~w19043 & ~w19100;
assign w19102 = pi0352 & ~w19042;
assign w19103 = w2251 & ~w7732;
assign w19104 = pi4023 & w19077;
assign w19105 = w19062 & w39957;
assign w19106 = w19048 & w39958;
assign w19107 = ~w19105 & ~w19106;
assign w19108 = w19062 & w39959;
assign w19109 = w19048 & w39960;
assign w19110 = ~w19108 & ~w19109;
assign w19111 = w19107 & w19110;
assign w19112 = w19059 & w39961;
assign w19113 = w19059 & w39962;
assign w19114 = w19059 & w39963;
assign w19115 = w19058 & w39964;
assign w19116 = ~w19114 & ~w19115;
assign w19117 = w19116 & w39965;
assign w19118 = w19111 & w19117;
assign w19119 = ~w19104 & w19118;
assign w19120 = ~w19104 & w39966;
assign w19121 = ~pi2515 & pi3474;
assign w19122 = (w19039 & w39967) | (w19039 & w39968) | (w39967 & w39968);
assign w19123 = ~w19120 & w19122;
assign w19124 = ~w19103 & w19123;
assign w19125 = w19124 & w40205;
assign w19126 = ~w19102 & ~w19125;
assign w19127 = pi0353 & ~w19042;
assign w19128 = (w2251 & w7699) | (w2251 & w39970) | (w7699 & w39970);
assign w19129 = pi4022 & w19077;
assign w19130 = w19059 & w39971;
assign w19131 = w19048 & w39972;
assign w19132 = ~w19130 & ~w19131;
assign w19133 = w19062 & w39973;
assign w19134 = w19048 & w39974;
assign w19135 = ~w19133 & ~w19134;
assign w19136 = w19132 & w19135;
assign w19137 = w19059 & w39975;
assign w19138 = w19059 & w39976;
assign w19139 = w19062 & w39977;
assign w19140 = w19058 & w39978;
assign w19141 = ~w19139 & ~w19140;
assign w19142 = w19141 & w39979;
assign w19143 = w19136 & w19142;
assign w19144 = ~w19129 & w19143;
assign w19145 = ~w19129 & w39980;
assign w19146 = ~pi2515 & pi3477;
assign w19147 = (w19039 & w39981) | (w19039 & w39982) | (w39981 & w39982);
assign w19148 = ~w19145 & w19147;
assign w19149 = ~w19128 & w19148;
assign w19150 = w19149 & w40206;
assign w19151 = ~w19127 & ~w19150;
assign w19152 = ~pi0354 & ~w19042;
assign w19153 = (w3412 & w39983) | (w3412 & w39984) | (w39983 & w39984);
assign w19154 = (w2257 & w7667) | (w2257 & w39985) | (w7667 & w39985);
assign w19155 = pi4021 & w19077;
assign w19156 = w19048 & w39986;
assign w19157 = w19062 & w39987;
assign w19158 = ~w19156 & ~w19157;
assign w19159 = w19059 & w39988;
assign w19160 = w19062 & w39989;
assign w19161 = ~w19159 & ~w19160;
assign w19162 = w19158 & w19161;
assign w19163 = w19059 & w39990;
assign w19164 = w19059 & w39991;
assign w19165 = w19048 & w39992;
assign w19166 = w19058 & w39993;
assign w19167 = ~w19165 & ~w19166;
assign w19168 = w19167 & w39994;
assign w19169 = w19162 & w19168;
assign w19170 = ~w19155 & w19169;
assign w19171 = ~w19155 & w39995;
assign w19172 = pi2515 & ~w19171;
assign w19173 = ~w19154 & w19172;
assign w19174 = ~pi2515 & ~pi3476;
assign w19175 = (w19039 & w39996) | (w19039 & w39997) | (w39996 & w39997);
assign w19176 = (w19175 & w19153) | (w19175 & w39998) | (w19153 & w39998);
assign w19177 = ~w19152 & ~w19176;
assign w19178 = pi0355 & ~w19042;
assign w19179 = w6609 & ~w6413;
assign w19180 = (w2251 & w7634) | (w2251 & w39999) | (w7634 & w39999);
assign w19181 = pi4020 & w19077;
assign w19182 = w19048 & w40000;
assign w19183 = w19048 & w40001;
assign w19184 = ~w19182 & ~w19183;
assign w19185 = w19059 & w40002;
assign w19186 = w19062 & w40003;
assign w19187 = ~w19185 & ~w19186;
assign w19188 = w19184 & w19187;
assign w19189 = w19059 & w40004;
assign w19190 = w19059 & w40005;
assign w19191 = w19062 & w40006;
assign w19192 = w19058 & w40007;
assign w19193 = ~w19191 & ~w19192;
assign w19194 = w19193 & w40008;
assign w19195 = w19188 & w19194;
assign w19196 = ~w19181 & w19195;
assign w19197 = ~w19181 & w40009;
assign w19198 = ~pi2515 & pi3475;
assign w19199 = (w19039 & w40010) | (w19039 & w40011) | (w40010 & w40011);
assign w19200 = ~w19197 & w19199;
assign w19201 = ~w19180 & w19200;
assign w19202 = ~w19179 & w19201;
assign w19203 = ~w19178 & ~w19202;
assign w19204 = pi0356 & ~w19042;
assign w19205 = (w2251 & w7601) | (w2251 & w40013) | (w7601 & w40013);
assign w19206 = pi4019 & w19077;
assign w19207 = w19062 & w40014;
assign w19208 = w19059 & w40015;
assign w19209 = ~w19207 & ~w19208;
assign w19210 = w19062 & w40016;
assign w19211 = w19048 & w40017;
assign w19212 = ~w19210 & ~w19211;
assign w19213 = w19209 & w19212;
assign w19214 = w19059 & w40018;
assign w19215 = w19059 & w40019;
assign w19216 = w19048 & w40020;
assign w19217 = w19058 & w40021;
assign w19218 = ~w19216 & ~w19217;
assign w19219 = w19218 & w40022;
assign w19220 = w19213 & w19219;
assign w19221 = ~w19206 & w19220;
assign w19222 = ~w19206 & w40023;
assign w19223 = ~pi2515 & pi3470;
assign w19224 = (w19039 & w40024) | (w19039 & w40025) | (w40024 & w40025);
assign w19225 = ~w19222 & w19224;
assign w19226 = ~w19205 & w19225;
assign w19227 = w19226 & w40207;
assign w19228 = ~w19204 & ~w19227;
assign w19229 = pi0357 & ~w19042;
assign w19230 = (w2251 & w7569) | (w2251 & w40027) | (w7569 & w40027);
assign w19231 = pi4018 & w19077;
assign w19232 = w19048 & w40028;
assign w19233 = w19062 & w40029;
assign w19234 = ~w19232 & ~w19233;
assign w19235 = w19062 & w40030;
assign w19236 = w19059 & w40031;
assign w19237 = ~w19235 & ~w19236;
assign w19238 = w19234 & w19237;
assign w19239 = w19059 & w40032;
assign w19240 = w19059 & w40033;
assign w19241 = w19048 & w40034;
assign w19242 = w19058 & w40035;
assign w19243 = ~w19241 & ~w19242;
assign w19244 = w19243 & w40036;
assign w19245 = w19238 & w19244;
assign w19246 = ~w19231 & w19245;
assign w19247 = ~w19231 & w40037;
assign w19248 = ~pi2515 & pi3446;
assign w19249 = (w19039 & w40038) | (w19039 & w40039) | (w40038 & w40039);
assign w19250 = ~w19247 & w19249;
assign w19251 = ~w19230 & w19250;
assign w19252 = w19251 & w40208;
assign w19253 = ~w19229 & ~w19252;
assign w19254 = ~pi0358 & ~w19042;
assign w19255 = (w5893 & w40040) | (w5893 & w40041) | (w40040 & w40041);
assign w19256 = w2257 & ~w7537;
assign w19257 = pi4017 & w19077;
assign w19258 = w19048 & w40042;
assign w19259 = w19062 & w40043;
assign w19260 = ~w19258 & ~w19259;
assign w19261 = w19059 & w40044;
assign w19262 = w19062 & w40045;
assign w19263 = ~w19261 & ~w19262;
assign w19264 = w19260 & w19263;
assign w19265 = w19059 & w40046;
assign w19266 = w19059 & w40047;
assign w19267 = w19048 & w40048;
assign w19268 = pi4113 & w19074;
assign w19269 = ~w19267 & ~w19268;
assign w19270 = ~w19266 & w19269;
assign w19271 = ~w19265 & w19270;
assign w19272 = w19264 & w19271;
assign w19273 = ~w19257 & w19272;
assign w19274 = w7230 & w19273;
assign w19275 = pi2515 & ~w19274;
assign w19276 = ~w19256 & w19275;
assign w19277 = ~w19255 & w19276;
assign w19278 = ~pi2515 & ~pi3462;
assign w19279 = w19042 & ~w19278;
assign w19280 = ~w19277 & w19279;
assign w19281 = ~w19254 & ~w19280;
assign w19282 = ~pi0359 & ~w19042;
assign w19283 = pi1422 & ~w4749;
assign w19284 = w2257 & ~w7505;
assign w19285 = pi4016 & w19077;
assign w19286 = pi4040 & w19054;
assign w19287 = pi4208 & w19072;
assign w19288 = ~w19286 & ~w19287;
assign w19289 = pi4088 & w19064;
assign w19290 = pi4064 & w19051;
assign w19291 = ~w19289 & ~w19290;
assign w19292 = w19288 & w19291;
assign w19293 = pi4184 & w19070;
assign w19294 = pi4160 & w19068;
assign w19295 = pi4136 & w19061;
assign w19296 = pi4112 & w19074;
assign w19297 = ~w19295 & ~w19296;
assign w19298 = ~w19294 & w19297;
assign w19299 = ~w19293 & w19298;
assign w19300 = w19292 & w19299;
assign w19301 = ~w19285 & w19300;
assign w19302 = w7230 & w19301;
assign w19303 = pi2515 & ~w19302;
assign w19304 = ~w19284 & w19303;
assign w19305 = ~w19283 & w19304;
assign w19306 = ~pi2515 & ~pi3468;
assign w19307 = w19042 & ~w19306;
assign w19308 = ~w19305 & w19307;
assign w19309 = ~w19282 & ~w19308;
assign w19310 = pi0360 & ~w19042;
assign w19311 = w6609 & ~w8240;
assign w19312 = w2251 & ~w8266;
assign w19313 = pi4030 & w19077;
assign w19314 = pi4078 & w19051;
assign w19315 = pi4150 & w19061;
assign w19316 = ~w19314 & ~w19315;
assign w19317 = pi4102 & w19064;
assign w19318 = pi4222 & w19072;
assign w19319 = ~w19317 & ~w19318;
assign w19320 = w19316 & w19319;
assign w19321 = pi4198 & w19070;
assign w19322 = pi4174 & w19068;
assign w19323 = pi4054 & w19054;
assign w19324 = pi4126 & w19074;
assign w19325 = ~w19323 & ~w19324;
assign w19326 = ~w19322 & w19325;
assign w19327 = ~w19321 & w19326;
assign w19328 = w19320 & w19327;
assign w19329 = ~w19313 & w19328;
assign w19330 = w19094 & w19329;
assign w19331 = ~pi2515 & pi3467;
assign w19332 = w19042 & ~w19331;
assign w19333 = ~w19330 & w19332;
assign w19334 = ~w19312 & w19333;
assign w19335 = ~w19311 & w19334;
assign w19336 = ~w19310 & ~w19335;
assign w19337 = ~pi0361 & ~w19042;
assign w19338 = w6609 & w8081;
assign w19339 = w2251 & w7994;
assign w19340 = pi4029 & w19077;
assign w19341 = pi4077 & w19051;
assign w19342 = pi4053 & w19054;
assign w19343 = ~w19341 & ~w19342;
assign w19344 = pi4149 & w19061;
assign w19345 = pi4101 & w19064;
assign w19346 = ~w19344 & ~w19345;
assign w19347 = w19343 & w19346;
assign w19348 = pi4173 & w19068;
assign w19349 = pi4197 & w19070;
assign w19350 = pi4221 & w19072;
assign w19351 = pi4125 & w19074;
assign w19352 = ~w19350 & ~w19351;
assign w19353 = ~w19349 & w19352;
assign w19354 = ~w19348 & w19353;
assign w19355 = w19347 & w19354;
assign w19356 = ~w19340 & w19355;
assign w19357 = w19094 & ~w19356;
assign w19358 = ~pi2515 & ~pi3465;
assign w19359 = w19042 & ~w19358;
assign w19360 = ~w19357 & w19359;
assign w19361 = ~w19339 & w19360;
assign w19362 = ~w19338 & w19361;
assign w19363 = ~w19337 & ~w19362;
assign w19364 = pi0362 & ~w19042;
assign w19365 = ~w1639 & w6609;
assign w19366 = w2251 & ~w7892;
assign w19367 = pi4028 & w19077;
assign w19368 = pi4076 & w19051;
assign w19369 = pi4052 & w19054;
assign w19370 = ~w19368 & ~w19369;
assign w19371 = pi4100 & w19064;
assign w19372 = pi4220 & w19072;
assign w19373 = ~w19371 & ~w19372;
assign w19374 = w19370 & w19373;
assign w19375 = pi4196 & w19070;
assign w19376 = pi4172 & w19068;
assign w19377 = pi4148 & w19061;
assign w19378 = pi4124 & w19074;
assign w19379 = ~w19377 & ~w19378;
assign w19380 = ~w19376 & w19379;
assign w19381 = ~w19375 & w19380;
assign w19382 = w19374 & w19381;
assign w19383 = ~w19367 & w19382;
assign w19384 = w19094 & w19383;
assign w19385 = ~pi2515 & pi3466;
assign w19386 = w19042 & ~w19385;
assign w19387 = ~w19384 & w19386;
assign w19388 = ~w19366 & w19387;
assign w19389 = ~w19365 & w19388;
assign w19390 = ~w19364 & ~w19389;
assign w19391 = ~pi2515 & ~pi3447;
assign w19392 = pi1422 & ~w1308;
assign w19393 = w2257 & ~w7860;
assign w19394 = pi4027 & w19077;
assign w19395 = pi4147 & w19061;
assign w19396 = pi4051 & w19054;
assign w19397 = ~w19395 & ~w19396;
assign w19398 = pi4099 & w19064;
assign w19399 = pi4075 & w19051;
assign w19400 = ~w19398 & ~w19399;
assign w19401 = w19397 & w19400;
assign w19402 = pi4171 & w19068;
assign w19403 = pi4195 & w19070;
assign w19404 = pi4219 & w19072;
assign w19405 = pi4123 & w19074;
assign w19406 = ~w19404 & ~w19405;
assign w19407 = ~w19403 & w19406;
assign w19408 = ~w19402 & w19407;
assign w19409 = w19401 & w19408;
assign w19410 = ~w19394 & w19409;
assign w19411 = w7230 & w19410;
assign w19412 = pi2515 & ~w19411;
assign w19413 = ~w19393 & w19412;
assign w19414 = ~w19392 & w19413;
assign w19415 = ~w19391 & ~w19414;
assign w19416 = w19042 & ~w19415;
assign w19417 = pi0363 & ~w19042;
assign w19418 = ~w19416 & ~w19417;
assign w19419 = pi0364 & ~w19042;
assign w19420 = ~w5635 & w6609;
assign w19421 = w2251 & ~w7828;
assign w19422 = pi4026 & w19077;
assign w19423 = pi4146 & w19061;
assign w19424 = pi4098 & w19064;
assign w19425 = ~w19423 & ~w19424;
assign w19426 = pi4218 & w19072;
assign w19427 = pi4050 & w19054;
assign w19428 = ~w19426 & ~w19427;
assign w19429 = w19425 & w19428;
assign w19430 = pi4194 & w19070;
assign w19431 = pi4170 & w19068;
assign w19432 = pi4074 & w19051;
assign w19433 = pi4122 & w19074;
assign w19434 = ~w19432 & ~w19433;
assign w19435 = ~w19431 & w19434;
assign w19436 = ~w19430 & w19435;
assign w19437 = w19429 & w19436;
assign w19438 = ~w19422 & w19437;
assign w19439 = w19094 & w19438;
assign w19440 = ~pi2515 & pi3463;
assign w19441 = w19042 & ~w19440;
assign w19442 = ~w19439 & w19441;
assign w19443 = ~w19421 & w19442;
assign w19444 = ~w19420 & w19443;
assign w19445 = ~w19419 & ~w19444;
assign w19446 = pi0365 & ~w19042;
assign w19447 = ~w5053 & w6609;
assign w19448 = w2251 & ~w7796;
assign w19449 = pi4025 & w19077;
assign w19450 = pi4145 & w19061;
assign w19451 = pi4073 & w19051;
assign w19452 = ~w19450 & ~w19451;
assign w19453 = pi4049 & w19054;
assign w19454 = pi4097 & w19064;
assign w19455 = ~w19453 & ~w19454;
assign w19456 = w19452 & w19455;
assign w19457 = pi4169 & w19068;
assign w19458 = pi4193 & w19070;
assign w19459 = pi4217 & w19072;
assign w19460 = pi4121 & w19074;
assign w19461 = ~w19459 & ~w19460;
assign w19462 = ~w19458 & w19461;
assign w19463 = ~w19457 & w19462;
assign w19464 = w19456 & w19463;
assign w19465 = ~w19449 & w19464;
assign w19466 = w19094 & w19465;
assign w19467 = ~pi2515 & pi3448;
assign w19468 = w19042 & ~w19467;
assign w19469 = ~w19466 & w19468;
assign w19470 = ~w19448 & w19469;
assign w19471 = ~w19447 & w19470;
assign w19472 = ~w19446 & ~w19471;
assign w19473 = pi0366 & ~w19042;
assign w19474 = ~w3711 & w6609;
assign w19475 = w2251 & ~w7473;
assign w19476 = pi4015 & w19077;
assign w19477 = pi4039 & w19054;
assign w19478 = pi4063 & w19051;
assign w19479 = ~w19477 & ~w19478;
assign w19480 = pi4087 & w19064;
assign w19481 = pi4207 & w19072;
assign w19482 = ~w19480 & ~w19481;
assign w19483 = w19479 & w19482;
assign w19484 = pi4159 & w19068;
assign w19485 = pi4183 & w19070;
assign w19486 = pi4135 & w19061;
assign w19487 = pi4111 & w19074;
assign w19488 = ~w19486 & ~w19487;
assign w19489 = ~w19485 & w19488;
assign w19490 = ~w19484 & w19489;
assign w19491 = w19483 & w19490;
assign w19492 = ~w19476 & w19491;
assign w19493 = w19094 & w19492;
assign w19494 = ~pi2515 & pi3464;
assign w19495 = w19042 & ~w19494;
assign w19496 = ~w19493 & w19495;
assign w19497 = ~w19475 & w19496;
assign w19498 = ~w19474 & w19497;
assign w19499 = ~w19473 & ~w19498;
assign w19500 = ~pi2395 & w18313;
assign w19501 = pi0367 & ~w18338;
assign w19502 = ~w18339 & ~w18359;
assign w19503 = ~w19501 & w19502;
assign w19504 = ~pi1725 & w18359;
assign w19505 = ~w18313 & ~w19504;
assign w19506 = ~w19503 & w19505;
assign w19507 = ~w19500 & ~w19506;
assign w19508 = pi2555 & ~w15303;
assign w19509 = w40134 & ~w15388;
assign w19510 = pi0368 & w15388;
assign w19511 = ~pi2555 & ~w19510;
assign w19512 = ~w19509 & w19511;
assign w19513 = ~w19508 & ~w19512;
assign w19514 = pi3266 & ~pi3271;
assign w19515 = ~pi3246 & ~pi3255;
assign w19516 = w19514 & w19515;
assign w19517 = ~pi2567 & pi3142;
assign w19518 = w19516 & w19517;
assign w19519 = ~pi1008 & ~pi3426;
assign w19520 = ~pi3305 & ~w19519;
assign w19521 = ~w370 & ~w19520;
assign w19522 = ~w19518 & ~w19521;
assign w19523 = pi3305 & ~w19522;
assign w19524 = ~pi3682 & ~w19383;
assign w19525 = ~pi3261 & pi3682;
assign w19526 = ~w19524 & ~w19525;
assign w19527 = w19523 & ~w19526;
assign w19528 = pi0785 & w19518;
assign w19529 = pi0369 & w19522;
assign w19530 = ~w19528 & ~w19529;
assign w19531 = ~w19527 & w19530;
assign w19532 = ~w4749 & w18009;
assign w19533 = ~pi0370 & ~w18375;
assign w19534 = pi0479 & w17870;
assign w19535 = ~w17954 & ~w19534;
assign w19536 = ~pi0247 & ~w19535;
assign w19537 = pi0247 & ~pi0278;
assign w19538 = ~pi0479 & w19537;
assign w19539 = ~w17952 & ~w19538;
assign w19540 = ~w19536 & w19539;
assign w19541 = pi0248 & ~w19540;
assign w19542 = w18367 & ~w19019;
assign w19543 = ~w19541 & w19542;
assign w19544 = pi0694 & w18003;
assign w19545 = ~w19543 & ~w19544;
assign w19546 = ~w19533 & w19545;
assign w19547 = ~w19532 & w19546;
assign w19548 = ~pi3682 & ~w19410;
assign w19549 = ~pi3283 & pi3682;
assign w19550 = ~w19548 & ~w19549;
assign w19551 = w19523 & ~w19550;
assign w19552 = pi0825 & w19518;
assign w19553 = pi0371 & w19522;
assign w19554 = ~w19552 & ~w19553;
assign w19555 = ~w19551 & w19554;
assign w19556 = ~pi3682 & ~w19438;
assign w19557 = ~pi3273 & pi3682;
assign w19558 = ~w19556 & ~w19557;
assign w19559 = w19523 & ~w19558;
assign w19560 = pi0855 & w19518;
assign w19561 = pi0372 & w19522;
assign w19562 = ~w19560 & ~w19561;
assign w19563 = ~w19559 & w19562;
assign w19564 = ~pi3682 & ~w19465;
assign w19565 = ~pi3263 & pi3682;
assign w19566 = ~w19564 & ~w19565;
assign w19567 = w19523 & ~w19566;
assign w19568 = pi0856 & w19518;
assign w19569 = pi0373 & w19522;
assign w19570 = ~w19568 & ~w19569;
assign w19571 = ~w19567 & w19570;
assign w19572 = ~pi3682 & ~w19093;
assign w19573 = ~pi3282 & pi3682;
assign w19574 = ~w19572 & ~w19573;
assign w19575 = w19523 & ~w19574;
assign w19576 = pi0857 & w19518;
assign w19577 = pi0374 & w19522;
assign w19578 = ~w19576 & ~w19577;
assign w19579 = ~w19575 & w19578;
assign w19580 = ~pi3682 & ~w19119;
assign w19581 = ~pi3264 & pi3682;
assign w19582 = ~w19580 & ~w19581;
assign w19583 = w19523 & ~w19582;
assign w19584 = pi0858 & w19518;
assign w19585 = pi0375 & w19522;
assign w19586 = ~w19584 & ~w19585;
assign w19587 = ~w19583 & w19586;
assign w19588 = w19519 & ~w19522;
assign w19589 = w8240 & w19588;
assign w19590 = ~pi3682 & ~w19144;
assign w19591 = ~pi3274 & pi3682;
assign w19592 = ~w19590 & ~w19591;
assign w19593 = w19523 & ~w19592;
assign w19594 = pi0824 & w19518;
assign w19595 = pi0376 & w19522;
assign w19596 = ~w19594 & ~w19595;
assign w19597 = ~w19593 & w19596;
assign w19598 = ~w19589 & w19597;
assign w19599 = w8081 & w19588;
assign w19600 = ~pi3682 & ~w19170;
assign w19601 = ~pi3280 & pi3682;
assign w19602 = ~w19600 & ~w19601;
assign w19603 = w19523 & ~w19602;
assign w19604 = pi0823 & w19518;
assign w19605 = pi0377 & w19522;
assign w19606 = ~w19604 & ~w19605;
assign w19607 = ~w19603 & w19606;
assign w19608 = ~w19599 & w19607;
assign w19609 = w1639 & w19588;
assign w19610 = ~pi3682 & ~w19196;
assign w19611 = ~pi3279 & pi3682;
assign w19612 = ~w19610 & ~w19611;
assign w19613 = w19523 & ~w19612;
assign w19614 = pi0859 & w19518;
assign w19615 = pi0378 & w19522;
assign w19616 = ~w19614 & ~w19615;
assign w19617 = ~w19613 & w19616;
assign w19618 = ~w19609 & w19617;
assign w19619 = ~pi3682 & ~w19329;
assign w19620 = ~pi3253 & pi3682;
assign w19621 = ~w19619 & ~w19620;
assign w19622 = w19523 & ~w19621;
assign w19623 = pi0853 & w19518;
assign w19624 = pi0379 & w19522;
assign w19625 = ~w19623 & ~w19624;
assign w19626 = ~w19622 & w19625;
assign w19627 = ~pi3682 & ~w19356;
assign w19628 = ~pi3272 & pi3682;
assign w19629 = ~w19627 & ~w19628;
assign w19630 = w19523 & ~w19629;
assign w19631 = pi0854 & w19518;
assign w19632 = pi0380 & w19522;
assign w19633 = ~w19631 & ~w19632;
assign w19634 = ~w19630 & w19633;
assign w19635 = w1308 & w19588;
assign w19636 = ~pi3682 & ~w19221;
assign w19637 = ~pi3275 & pi3682;
assign w19638 = ~w19636 & ~w19637;
assign w19639 = w19523 & ~w19638;
assign w19640 = pi0730 & w19518;
assign w19641 = pi0381 & w19522;
assign w19642 = ~w19640 & ~w19641;
assign w19643 = ~w19639 & w19642;
assign w19644 = ~w19635 & w19643;
assign w19645 = w4141 & w19588;
assign w19646 = ~pi3682 & ~w19301;
assign w19647 = ~pi3258 & pi3682;
assign w19648 = ~w19646 & ~w19647;
assign w19649 = w19523 & ~w19648;
assign w19650 = pi0851 & w19518;
assign w19651 = pi0382 & w19522;
assign w19652 = ~w19650 & ~w19651;
assign w19653 = ~w19649 & w19652;
assign w19654 = ~w19645 & w19653;
assign w19655 = w6177 & w19588;
assign w19656 = ~pi3682 & ~w19492;
assign w19657 = ~pi3259 & pi3682;
assign w19658 = ~w19656 & ~w19657;
assign w19659 = w19523 & ~w19658;
assign w19660 = pi0860 & w19518;
assign w19661 = pi0383 & w19522;
assign w19662 = ~w19660 & ~w19661;
assign w19663 = ~w19659 & w19662;
assign w19664 = ~w19655 & w19663;
assign w19665 = w3195 & w19588;
assign w19666 = pi4014 & w19077;
assign w19667 = pi4134 & w19061;
assign w19668 = pi4086 & w19064;
assign w19669 = ~w19667 & ~w19668;
assign w19670 = pi4206 & w19072;
assign w19671 = pi4038 & w19054;
assign w19672 = ~w19670 & ~w19671;
assign w19673 = w19669 & w19672;
assign w19674 = pi4182 & w19070;
assign w19675 = pi4158 & w19068;
assign w19676 = pi4062 & w19051;
assign w19677 = pi4110 & w19074;
assign w19678 = ~w19676 & ~w19677;
assign w19679 = ~w19675 & w19678;
assign w19680 = ~w19674 & w19679;
assign w19681 = w19673 & w19680;
assign w19682 = ~w19666 & w19681;
assign w19683 = ~pi3682 & ~w19682;
assign w19684 = ~pi3286 & pi3682;
assign w19685 = ~w19683 & ~w19684;
assign w19686 = w19523 & ~w19685;
assign w19687 = pi0852 & w19518;
assign w19688 = pi0384 & w19522;
assign w19689 = ~w19687 & ~w19688;
assign w19690 = ~w19686 & w19689;
assign w19691 = ~w19665 & w19690;
assign w19692 = w40134 & w19588;
assign w19693 = pi4013 & w19077;
assign w19694 = pi4061 & w19051;
assign w19695 = pi4133 & w19061;
assign w19696 = ~w19694 & ~w19695;
assign w19697 = pi4085 & w19064;
assign w19698 = pi4205 & w19072;
assign w19699 = ~w19697 & ~w19698;
assign w19700 = w19696 & w19699;
assign w19701 = pi4181 & w19070;
assign w19702 = pi4157 & w19068;
assign w19703 = pi4037 & w19054;
assign w19704 = pi4109 & w19074;
assign w19705 = ~w19703 & ~w19704;
assign w19706 = ~w19702 & w19705;
assign w19707 = ~w19701 & w19706;
assign w19708 = w19700 & w19707;
assign w19709 = ~w19693 & w19708;
assign w19710 = ~pi3682 & ~w19709;
assign w19711 = ~pi3287 & pi3682;
assign w19712 = ~w19710 & ~w19711;
assign w19713 = w19523 & ~w19712;
assign w19714 = pi0821 & w19518;
assign w19715 = pi0385 & w19522;
assign w19716 = ~w19714 & ~w19715;
assign w19717 = ~w19713 & w19716;
assign w19718 = ~w19692 & w19717;
assign w19719 = w6413 & w19588;
assign w19720 = pi4012 & w19077;
assign w19721 = pi4036 & w19054;
assign w19722 = pi4084 & w19064;
assign w19723 = ~w19721 & ~w19722;
assign w19724 = pi4132 & w19061;
assign w19725 = pi4060 & w19051;
assign w19726 = ~w19724 & ~w19725;
assign w19727 = w19723 & w19726;
assign w19728 = pi4156 & w19068;
assign w19729 = pi4180 & w19070;
assign w19730 = pi4204 & w19072;
assign w19731 = pi4108 & w19074;
assign w19732 = ~w19730 & ~w19731;
assign w19733 = ~w19729 & w19732;
assign w19734 = ~w19728 & w19733;
assign w19735 = w19727 & w19734;
assign w19736 = ~w19720 & w19735;
assign w19737 = ~pi3682 & ~w19736;
assign w19738 = ~pi3289 & pi3682;
assign w19739 = ~w19737 & ~w19738;
assign w19740 = w19523 & ~w19739;
assign w19741 = ~pi0937 & w19518;
assign w19742 = pi0386 & w19522;
assign w19743 = ~w19741 & ~w19742;
assign w19744 = ~w19740 & w19743;
assign w19745 = ~w19719 & w19744;
assign w19746 = w4380 & w19588;
assign w19747 = pi4011 & w19077;
assign w19748 = pi4035 & w19054;
assign w19749 = pi4059 & w19051;
assign w19750 = ~w19748 & ~w19749;
assign w19751 = pi4083 & w19064;
assign w19752 = pi4203 & w19072;
assign w19753 = ~w19751 & ~w19752;
assign w19754 = w19750 & w19753;
assign w19755 = pi4179 & w19070;
assign w19756 = pi4155 & w19068;
assign w19757 = pi4131 & w19061;
assign w19758 = pi4107 & w19074;
assign w19759 = ~w19757 & ~w19758;
assign w19760 = ~w19756 & w19759;
assign w19761 = ~w19755 & w19760;
assign w19762 = w19754 & w19761;
assign w19763 = ~w19747 & w19762;
assign w19764 = ~pi3682 & ~w19763;
assign w19765 = ~pi3288 & pi3682;
assign w19766 = ~w19764 & ~w19765;
assign w19767 = w19523 & ~w19766;
assign w19768 = ~pi1045 & w19518;
assign w19769 = pi0387 & w19522;
assign w19770 = ~w19768 & ~w19769;
assign w19771 = ~w19767 & w19770;
assign w19772 = ~w19746 & w19771;
assign w19773 = w5320 & w19588;
assign w19774 = pi4010 & w19077;
assign w19775 = pi4202 & w19072;
assign w19776 = pi4130 & w19061;
assign w19777 = ~w19775 & ~w19776;
assign w19778 = pi4082 & w19064;
assign w19779 = pi4058 & w19051;
assign w19780 = ~w19778 & ~w19779;
assign w19781 = w19777 & w19780;
assign w19782 = pi4154 & w19068;
assign w19783 = pi4178 & w19070;
assign w19784 = pi4034 & w19054;
assign w19785 = pi4106 & w19074;
assign w19786 = ~w19784 & ~w19785;
assign w19787 = ~w19783 & w19786;
assign w19788 = ~w19782 & w19787;
assign w19789 = w19781 & w19788;
assign w19790 = ~w19774 & w19789;
assign w19791 = ~pi3682 & ~w19790;
assign w19792 = ~pi3260 & pi3682;
assign w19793 = ~w19791 & ~w19792;
assign w19794 = w19523 & ~w19793;
assign w19795 = ~pi1082 & w19518;
assign w19796 = pi0388 & w19522;
assign w19797 = ~w19795 & ~w19796;
assign w19798 = ~w19794 & w19797;
assign w19799 = ~w19773 & w19798;
assign w19800 = w5914 & w19588;
assign w19801 = pi4009 & w19077;
assign w19802 = pi4033 & w19054;
assign w19803 = pi4201 & w19072;
assign w19804 = ~w19802 & ~w19803;
assign w19805 = pi4081 & w19064;
assign w19806 = pi4057 & w19051;
assign w19807 = ~w19805 & ~w19806;
assign w19808 = w19804 & w19807;
assign w19809 = pi4177 & w19070;
assign w19810 = pi4153 & w19068;
assign w19811 = pi4129 & w19061;
assign w19812 = pi4105 & w19074;
assign w19813 = ~w19811 & ~w19812;
assign w19814 = ~w19810 & w19813;
assign w19815 = ~w19809 & w19814;
assign w19816 = w19808 & w19815;
assign w19817 = ~w19801 & w19816;
assign w19818 = ~pi3682 & ~w19817;
assign w19819 = ~pi3284 & pi3682;
assign w19820 = ~w19818 & ~w19819;
assign w19821 = w19523 & ~w19820;
assign w19822 = ~pi1080 & w19518;
assign w19823 = pi0389 & w19522;
assign w19824 = ~w19822 & ~w19823;
assign w19825 = ~w19821 & w19824;
assign w19826 = ~w19800 & w19825;
assign w19827 = w4749 & w19588;
assign w19828 = pi4008 & w19077;
assign w19829 = pi4032 & w19054;
assign w19830 = pi4080 & w19064;
assign w19831 = ~w19829 & ~w19830;
assign w19832 = pi4200 & w19072;
assign w19833 = pi4128 & w19061;
assign w19834 = ~w19832 & ~w19833;
assign w19835 = w19831 & w19834;
assign w19836 = pi4176 & w19070;
assign w19837 = pi4152 & w19068;
assign w19838 = pi4056 & w19051;
assign w19839 = pi4104 & w19074;
assign w19840 = ~w19838 & ~w19839;
assign w19841 = ~w19837 & w19840;
assign w19842 = ~w19836 & w19841;
assign w19843 = w19835 & w19842;
assign w19844 = ~w19828 & w19843;
assign w19845 = ~pi3682 & ~w19844;
assign w19846 = ~pi3262 & pi3682;
assign w19847 = ~w19845 & ~w19846;
assign w19848 = w19523 & ~w19847;
assign w19849 = ~pi1052 & w19518;
assign w19850 = pi0390 & w19522;
assign w19851 = ~w19849 & ~w19850;
assign w19852 = ~w19848 & w19851;
assign w19853 = ~w19827 & w19852;
assign w19854 = w5635 & w19588;
assign w19855 = ~pi3682 & ~w19246;
assign w19856 = ~pi3276 & pi3682;
assign w19857 = ~w19855 & ~w19856;
assign w19858 = w19523 & ~w19857;
assign w19859 = pi0731 & w19518;
assign w19860 = pi0391 & w19522;
assign w19861 = ~w19859 & ~w19860;
assign w19862 = ~w19858 & w19861;
assign w19863 = ~w19854 & w19862;
assign w19864 = w5053 & w19588;
assign w19865 = ~pi3682 & ~w19273;
assign w19866 = ~pi3265 & pi3682;
assign w19867 = ~w19865 & ~w19866;
assign w19868 = w19523 & ~w19867;
assign w19869 = pi0938 & w19518;
assign w19870 = pi0392 & w19522;
assign w19871 = ~w19869 & ~w19870;
assign w19872 = ~w19868 & w19871;
assign w19873 = ~w19864 & w19872;
assign w19874 = w3711 & w19588;
assign w19875 = pi4007 & w19077;
assign w19876 = pi4055 & w19051;
assign w19877 = pi4127 & w19061;
assign w19878 = ~w19876 & ~w19877;
assign w19879 = pi4079 & w19064;
assign w19880 = pi4199 & w19072;
assign w19881 = ~w19879 & ~w19880;
assign w19882 = w19878 & w19881;
assign w19883 = pi4151 & w19068;
assign w19884 = pi4175 & w19070;
assign w19885 = pi4031 & w19054;
assign w19886 = pi4103 & w19074;
assign w19887 = ~w19885 & ~w19886;
assign w19888 = ~w19884 & w19887;
assign w19889 = ~w19883 & w19888;
assign w19890 = w19882 & w19889;
assign w19891 = ~w19875 & w19890;
assign w19892 = ~pi3682 & ~w19891;
assign w19893 = ~pi3277 & pi3682;
assign w19894 = ~w19892 & ~w19893;
assign w19895 = w19523 & ~w19894;
assign w19896 = ~pi0911 & w19518;
assign w19897 = pi0393 & w19522;
assign w19898 = ~w19896 & ~w19897;
assign w19899 = ~w19895 & w19898;
assign w19900 = ~w19874 & w19899;
assign w19901 = pi0394 & ~w18928;
assign w19902 = pi0712 & ~w18137;
assign w19903 = ~pi0712 & ~w40159;
assign w19904 = ~w19902 & ~w19903;
assign w19905 = w18928 & w19904;
assign w19906 = ~w19901 & ~w19905;
assign w19907 = pi0395 & ~w18935;
assign w19908 = w18935 & w19904;
assign w19909 = ~w19907 & ~w19908;
assign w19910 = w10752 & w16055;
assign w19911 = ~w40176 & w18039;
assign w19912 = ~pi0396 & ~w18039;
assign w19913 = ~w10753 & ~w19912;
assign w19914 = ~w19911 & w19913;
assign w19915 = w15173 & ~w19914;
assign w19916 = ~w19910 & ~w19915;
assign w19917 = w13923 & w16055;
assign w19918 = ~w40176 & w18046;
assign w19919 = ~pi0397 & ~w18046;
assign w19920 = ~w13925 & ~w19919;
assign w19921 = ~w19918 & w19920;
assign w19922 = w14336 & ~w19921;
assign w19923 = ~w19917 & ~w19922;
assign w19924 = ~pi2090 & w18313;
assign w19925 = pi0398 & ~w18337;
assign w19926 = ~w18338 & ~w18359;
assign w19927 = ~w19925 & w19926;
assign w19928 = ~pi1877 & w18359;
assign w19929 = ~w18313 & ~w19928;
assign w19930 = ~w19927 & w19929;
assign w19931 = ~w19924 & ~w19930;
assign w19932 = pi0399 & ~w18928;
assign w19933 = pi0712 & ~w18146;
assign w19934 = ~pi0712 & ~w13916;
assign w19935 = ~w19933 & ~w19934;
assign w19936 = w18928 & w19935;
assign w19937 = ~w19932 & ~w19936;
assign w19938 = pi0400 & ~w18935;
assign w19939 = w18935 & w19935;
assign w19940 = ~w19938 & ~w19939;
assign w19941 = pi0401 & ~w18412;
assign w19942 = ~w15014 & w17425;
assign w19943 = w14420 & ~w17425;
assign w19944 = ~w19942 & ~w19943;
assign w19945 = w18412 & ~w19944;
assign w19946 = ~w19941 & ~w19945;
assign w19947 = pi0402 & ~w18419;
assign w19948 = w18419 & ~w19944;
assign w19949 = ~w19947 & ~w19948;
assign w19950 = pi2813 & ~pi3552;
assign w19951 = ~pi0565 & pi3362;
assign w19952 = w909 & w19951;
assign w19953 = ~w19950 & ~w19952;
assign w19954 = w342 & w19953;
assign w19955 = ~w19526 & ~w19954;
assign w19956 = pi3246 & ~pi3255;
assign w19957 = w19514 & w19956;
assign w19958 = w19517 & w19957;
assign w19959 = ~pi0403 & ~w19958;
assign w19960 = ~pi0785 & w19958;
assign w19961 = ~w19959 & ~w19960;
assign w19962 = w19954 & w19961;
assign w19963 = ~w19955 & ~w19962;
assign w19964 = ~w342 & w2230;
assign w19965 = ~pi2549 & pi3042;
assign w19966 = pi2549 & ~pi3042;
assign w19967 = pi3028 & ~w19966;
assign w19968 = ~w19965 & w19967;
assign w19969 = pi2409 & pi3043;
assign w19970 = ~pi2409 & ~pi3043;
assign w19971 = pi2902 & ~pi3083;
assign w19972 = ~w19970 & w19971;
assign w19973 = ~w19969 & w19972;
assign w19974 = ~w19968 & w19973;
assign w19975 = ~pi2647 & pi3045;
assign w19976 = pi2647 & ~pi3045;
assign w19977 = pi3070 & ~w19976;
assign w19978 = ~w19975 & w19977;
assign w19979 = ~pi2540 & pi3047;
assign w19980 = pi2540 & ~pi3047;
assign w19981 = pi3032 & ~w19980;
assign w19982 = ~w19979 & w19981;
assign w19983 = ~w19978 & ~w19982;
assign w19984 = ~pi2788 & pi3061;
assign w19985 = pi2788 & ~pi3061;
assign w19986 = pi3031 & ~w19985;
assign w19987 = ~w19984 & w19986;
assign w19988 = ~pi2794 & pi3040;
assign w19989 = pi2794 & ~pi3040;
assign w19990 = pi3026 & ~w19989;
assign w19991 = ~w19988 & w19990;
assign w19992 = ~w19987 & ~w19991;
assign w19993 = w19983 & w19992;
assign w19994 = w19974 & w19993;
assign w19995 = pi2529 & ~pi3088;
assign w19996 = ~pi2529 & pi3088;
assign w19997 = pi3030 & ~w19996;
assign w19998 = ~w19995 & w19997;
assign w19999 = ~pi2797 & pi3092;
assign w20000 = pi2797 & ~pi3092;
assign w20001 = pi3090 & ~w20000;
assign w20002 = ~w19999 & w20001;
assign w20003 = ~w19998 & ~w20002;
assign w20004 = pi2796 & ~pi3103;
assign w20005 = ~pi2796 & pi3103;
assign w20006 = pi3081 & ~w20005;
assign w20007 = ~w20004 & w20006;
assign w20008 = pi2405 & ~pi2904;
assign w20009 = ~pi2405 & pi2904;
assign w20010 = pi3058 & ~w20009;
assign w20011 = ~w20008 & w20010;
assign w20012 = ~w20007 & ~w20011;
assign w20013 = w20003 & w20012;
assign w20014 = pi2553 & ~pi2970;
assign w20015 = ~pi2553 & pi2970;
assign w20016 = pi3062 & ~w20015;
assign w20017 = ~w20014 & w20016;
assign w20018 = pi2551 & ~pi3041;
assign w20019 = ~pi2551 & pi3041;
assign w20020 = pi3060 & ~w20019;
assign w20021 = ~w20018 & w20020;
assign w20022 = ~w20017 & ~w20021;
assign w20023 = pi2646 & ~pi2811;
assign w20024 = ~pi2646 & pi2811;
assign w20025 = pi2859 & ~w20024;
assign w20026 = ~w20023 & w20025;
assign w20027 = pi2404 & ~pi3044;
assign w20028 = ~pi2404 & pi3044;
assign w20029 = pi3057 & ~w20028;
assign w20030 = ~w20027 & w20029;
assign w20031 = ~w20026 & ~w20030;
assign w20032 = w20022 & w20031;
assign w20033 = pi2644 & ~pi2898;
assign w20034 = ~pi2644 & pi2898;
assign w20035 = pi3087 & ~w20034;
assign w20036 = ~w20033 & w20035;
assign w20037 = pi2473 & ~pi2806;
assign w20038 = ~pi2473 & pi2806;
assign w20039 = pi3029 & ~w20038;
assign w20040 = ~w20037 & w20039;
assign w20041 = ~w20036 & ~w20040;
assign w20042 = pi2645 & ~pi2791;
assign w20043 = ~pi2645 & pi2791;
assign w20044 = pi3027 & ~w20043;
assign w20045 = ~w20042 & w20044;
assign w20046 = pi2953 & ~pi3046;
assign w20047 = ~pi2953 & pi3046;
assign w20048 = pi3078 & ~w20047;
assign w20049 = ~w20046 & w20048;
assign w20050 = ~w20045 & ~w20049;
assign w20051 = w20041 & w20050;
assign w20052 = w20032 & w20051;
assign w20053 = w20013 & w20052;
assign w20054 = w19994 & w20053;
assign w20055 = ~pi2473 & pi3053;
assign w20056 = pi2473 & ~pi3053;
assign w20057 = pi3038 & ~w20056;
assign w20058 = ~w20055 & w20057;
assign w20059 = pi2409 & pi3052;
assign w20060 = ~pi2409 & ~pi3052;
assign w20061 = pi3051 & ~pi3082;
assign w20062 = ~w20060 & w20061;
assign w20063 = ~w20059 & w20062;
assign w20064 = ~w20058 & w20063;
assign w20065 = pi2551 & ~pi2957;
assign w20066 = ~pi2551 & pi2957;
assign w20067 = pi3036 & ~w20066;
assign w20068 = ~w20065 & w20067;
assign w20069 = pi2796 & ~pi3048;
assign w20070 = ~pi2796 & pi3048;
assign w20071 = pi2792 & ~w20070;
assign w20072 = ~w20069 & w20071;
assign w20073 = ~w20068 & ~w20072;
assign w20074 = pi2775 & ~pi2788;
assign w20075 = ~pi2775 & pi2788;
assign w20076 = pi2883 & ~w20075;
assign w20077 = ~w20074 & w20076;
assign w20078 = ~pi2953 & pi3069;
assign w20079 = pi2953 & ~pi3069;
assign w20080 = pi2823 & ~w20079;
assign w20081 = ~w20078 & w20080;
assign w20082 = ~w20077 & ~w20081;
assign w20083 = w20073 & w20082;
assign w20084 = w20064 & w20083;
assign w20085 = pi2553 & ~pi2971;
assign w20086 = ~pi2553 & pi2971;
assign w20087 = pi2903 & ~w20086;
assign w20088 = ~w20085 & w20087;
assign w20089 = pi2646 & ~pi2958;
assign w20090 = ~pi2646 & pi2958;
assign w20091 = pi2905 & ~w20090;
assign w20092 = ~w20089 & w20091;
assign w20093 = ~w20088 & ~w20092;
assign w20094 = pi2549 & ~pi2818;
assign w20095 = ~pi2549 & pi2818;
assign w20096 = pi3037 & ~w20095;
assign w20097 = ~w20094 & w20096;
assign w20098 = ~pi2540 & pi2882;
assign w20099 = pi2540 & ~pi2882;
assign w20100 = pi2973 & ~w20099;
assign w20101 = ~w20098 & w20100;
assign w20102 = ~w20097 & ~w20101;
assign w20103 = w20093 & w20102;
assign w20104 = ~pi2404 & pi2930;
assign w20105 = pi2404 & ~pi2930;
assign w20106 = pi3089 & ~w20105;
assign w20107 = ~w20104 & w20106;
assign w20108 = ~pi2405 & pi3054;
assign w20109 = pi2405 & ~pi3054;
assign w20110 = pi3039 & ~w20109;
assign w20111 = ~w20108 & w20110;
assign w20112 = ~w20107 & ~w20111;
assign w20113 = ~pi2797 & pi3050;
assign w20114 = pi2797 & ~pi3050;
assign w20115 = pi2881 & ~w20114;
assign w20116 = ~w20113 & w20115;
assign w20117 = pi2645 & ~pi3110;
assign w20118 = ~pi2645 & pi3110;
assign w20119 = pi3035 & ~w20118;
assign w20120 = ~w20117 & w20119;
assign w20121 = ~w20116 & ~w20120;
assign w20122 = w20112 & w20121;
assign w20123 = pi2529 & ~pi2915;
assign w20124 = ~pi2529 & pi2915;
assign w20125 = pi3071 & ~w20124;
assign w20126 = ~w20123 & w20125;
assign w20127 = ~pi2644 & pi3049;
assign w20128 = pi2644 & ~pi3049;
assign w20129 = pi3034 & ~w20128;
assign w20130 = ~w20127 & w20129;
assign w20131 = ~w20126 & ~w20130;
assign w20132 = ~pi2794 & pi2899;
assign w20133 = pi2794 & ~pi2899;
assign w20134 = pi3033 & ~w20133;
assign w20135 = ~w20132 & w20134;
assign w20136 = pi2647 & ~pi3080;
assign w20137 = ~pi2647 & pi3080;
assign w20138 = pi3064 & ~w20137;
assign w20139 = ~w20136 & w20138;
assign w20140 = ~w20135 & ~w20139;
assign w20141 = w20131 & w20140;
assign w20142 = w20122 & w20141;
assign w20143 = w20103 & w20142;
assign w20144 = w20084 & w20143;
assign w20145 = ~w20054 & ~w20144;
assign w20146 = ~pi2802 & ~pi3426;
assign w20147 = ~w20145 & w20146;
assign w20148 = pi1032 & ~pi2971;
assign w20149 = ~pi1032 & pi2971;
assign w20150 = pi2903 & ~w20149;
assign w20151 = ~w20148 & w20150;
assign w20152 = ~pi2978 & pi3052;
assign w20153 = pi2978 & ~pi3052;
assign w20154 = ~w20152 & ~w20153;
assign w20155 = ~pi2417 & ~pi3426;
assign w20156 = ~pi3051 & ~pi3082;
assign w20157 = w20155 & w20156;
assign w20158 = ~w20154 & w20157;
assign w20159 = ~w20151 & w20158;
assign w20160 = pi1013 & ~pi3110;
assign w20161 = ~pi1013 & pi3110;
assign w20162 = pi3035 & ~w20161;
assign w20163 = ~w20160 & w20162;
assign w20164 = pi1039 & ~pi2882;
assign w20165 = ~pi1039 & pi2882;
assign w20166 = pi2973 & ~w20165;
assign w20167 = ~w20164 & w20166;
assign w20168 = ~w20163 & ~w20167;
assign w20169 = ~pi2979 & pi3053;
assign w20170 = pi2979 & ~pi3053;
assign w20171 = pi3038 & ~w20170;
assign w20172 = ~w20169 & w20171;
assign w20173 = ~pi1036 & pi2915;
assign w20174 = pi1036 & ~pi2915;
assign w20175 = pi3071 & ~w20174;
assign w20176 = ~w20173 & w20175;
assign w20177 = ~w20172 & ~w20176;
assign w20178 = w20168 & w20177;
assign w20179 = w20159 & w20178;
assign w20180 = pi1031 & ~pi3050;
assign w20181 = ~pi1031 & pi3050;
assign w20182 = pi2881 & ~w20181;
assign w20183 = ~w20180 & w20182;
assign w20184 = ~pi1028 & pi2899;
assign w20185 = pi1028 & ~pi2899;
assign w20186 = pi3033 & ~w20185;
assign w20187 = ~w20184 & w20186;
assign w20188 = ~w20183 & ~w20187;
assign w20189 = ~pi1012 & pi2818;
assign w20190 = pi1012 & ~pi2818;
assign w20191 = pi3037 & ~w20190;
assign w20192 = ~w20189 & w20191;
assign w20193 = pi1029 & ~pi3048;
assign w20194 = ~pi1029 & pi3048;
assign w20195 = pi2792 & ~w20194;
assign w20196 = ~w20193 & w20195;
assign w20197 = ~w20192 & ~w20196;
assign w20198 = w20188 & w20197;
assign w20199 = ~pi2930 & pi2980;
assign w20200 = pi2930 & ~pi2980;
assign w20201 = pi3089 & ~w20200;
assign w20202 = ~w20199 & w20201;
assign w20203 = ~pi1030 & pi3049;
assign w20204 = pi1030 & ~pi3049;
assign w20205 = pi3034 & ~w20204;
assign w20206 = ~w20203 & w20205;
assign w20207 = ~w20202 & ~w20206;
assign w20208 = pi1035 & ~pi3080;
assign w20209 = ~pi1035 & pi3080;
assign w20210 = pi3064 & ~w20209;
assign w20211 = ~w20208 & w20210;
assign w20212 = pi1033 & ~pi2957;
assign w20213 = ~pi1033 & pi2957;
assign w20214 = pi3036 & ~w20213;
assign w20215 = ~w20212 & w20214;
assign w20216 = ~w20211 & ~w20215;
assign w20217 = w20207 & w20216;
assign w20218 = pi2981 & ~pi3054;
assign w20219 = ~pi2981 & pi3054;
assign w20220 = pi3039 & ~w20219;
assign w20221 = ~w20218 & w20220;
assign w20222 = ~pi1038 & pi2775;
assign w20223 = pi1038 & ~pi2775;
assign w20224 = pi2883 & ~w20223;
assign w20225 = ~w20222 & w20224;
assign w20226 = ~w20221 & ~w20225;
assign w20227 = ~pi1034 & pi2958;
assign w20228 = pi1034 & ~pi2958;
assign w20229 = pi2905 & ~w20228;
assign w20230 = ~w20227 & w20229;
assign w20231 = ~pi1037 & pi3069;
assign w20232 = pi1037 & ~pi3069;
assign w20233 = pi2823 & ~w20232;
assign w20234 = ~w20231 & w20233;
assign w20235 = ~w20230 & ~w20234;
assign w20236 = w20226 & w20235;
assign w20237 = w20217 & w20236;
assign w20238 = w20198 & w20237;
assign w20239 = w20179 & w20238;
assign w20240 = ~pi2806 & pi2979;
assign w20241 = pi2806 & ~pi2979;
assign w20242 = pi3029 & ~w20241;
assign w20243 = ~w20240 & w20242;
assign w20244 = ~pi2978 & pi3043;
assign w20245 = pi2978 & ~pi3043;
assign w20246 = ~w20244 & ~w20245;
assign w20247 = ~pi2902 & ~pi3083;
assign w20248 = w20155 & w20247;
assign w20249 = ~w20246 & w20248;
assign w20250 = ~w20243 & w20249;
assign w20251 = ~pi2904 & pi2981;
assign w20252 = pi2904 & ~pi2981;
assign w20253 = pi3058 & ~w20252;
assign w20254 = ~w20251 & w20253;
assign w20255 = pi1038 & ~pi3061;
assign w20256 = ~pi1038 & pi3061;
assign w20257 = pi3031 & ~w20256;
assign w20258 = ~w20255 & w20257;
assign w20259 = ~w20254 & ~w20258;
assign w20260 = ~pi1029 & pi3103;
assign w20261 = pi1029 & ~pi3103;
assign w20262 = pi3081 & ~w20261;
assign w20263 = ~w20260 & w20262;
assign w20264 = pi1033 & ~pi3041;
assign w20265 = ~pi1033 & pi3041;
assign w20266 = pi3060 & ~w20265;
assign w20267 = ~w20264 & w20266;
assign w20268 = ~w20263 & ~w20267;
assign w20269 = w20259 & w20268;
assign w20270 = w20250 & w20269;
assign w20271 = pi1034 & ~pi2811;
assign w20272 = ~pi1034 & pi2811;
assign w20273 = pi2859 & ~w20272;
assign w20274 = ~w20271 & w20273;
assign w20275 = pi1013 & ~pi2791;
assign w20276 = ~pi1013 & pi2791;
assign w20277 = pi3027 & ~w20276;
assign w20278 = ~w20275 & w20277;
assign w20279 = ~w20274 & ~w20278;
assign w20280 = pi2980 & ~pi3044;
assign w20281 = ~pi2980 & pi3044;
assign w20282 = pi3057 & ~w20281;
assign w20283 = ~w20280 & w20282;
assign w20284 = pi1028 & ~pi3040;
assign w20285 = ~pi1028 & pi3040;
assign w20286 = pi3026 & ~w20285;
assign w20287 = ~w20284 & w20286;
assign w20288 = ~w20283 & ~w20287;
assign w20289 = w20279 & w20288;
assign w20290 = pi1032 & ~pi2970;
assign w20291 = ~pi1032 & pi2970;
assign w20292 = pi3062 & ~w20291;
assign w20293 = ~w20290 & w20292;
assign w20294 = pi1031 & ~pi3092;
assign w20295 = ~pi1031 & pi3092;
assign w20296 = pi3090 & ~w20295;
assign w20297 = ~w20294 & w20296;
assign w20298 = ~w20293 & ~w20297;
assign w20299 = ~pi1036 & pi3088;
assign w20300 = pi1036 & ~pi3088;
assign w20301 = pi3030 & ~w20300;
assign w20302 = ~w20299 & w20301;
assign w20303 = pi1039 & ~pi3047;
assign w20304 = ~pi1039 & pi3047;
assign w20305 = pi3032 & ~w20304;
assign w20306 = ~w20303 & w20305;
assign w20307 = ~w20302 & ~w20306;
assign w20308 = w20298 & w20307;
assign w20309 = ~pi1030 & pi2898;
assign w20310 = pi1030 & ~pi2898;
assign w20311 = pi3087 & ~w20310;
assign w20312 = ~w20309 & w20311;
assign w20313 = pi1012 & ~pi3042;
assign w20314 = ~pi1012 & pi3042;
assign w20315 = pi3028 & ~w20314;
assign w20316 = ~w20313 & w20315;
assign w20317 = ~w20312 & ~w20316;
assign w20318 = pi1035 & ~pi3045;
assign w20319 = ~pi1035 & pi3045;
assign w20320 = pi3070 & ~w20319;
assign w20321 = ~w20318 & w20320;
assign w20322 = pi1037 & ~pi3046;
assign w20323 = ~pi1037 & pi3046;
assign w20324 = pi3078 & ~w20323;
assign w20325 = ~w20322 & w20324;
assign w20326 = ~w20321 & ~w20325;
assign w20327 = w20317 & w20326;
assign w20328 = w20308 & w20327;
assign w20329 = w20289 & w20328;
assign w20330 = w20270 & w20329;
assign w20331 = ~w20239 & ~w20330;
assign w20332 = ~w20147 & w20331;
assign w20333 = ~pi2761 & ~w20332;
assign w20334 = pi2482 & ~pi3012;
assign w20335 = ~pi2482 & pi3012;
assign w20336 = pi3073 & ~w20335;
assign w20337 = ~w20334 & w20336;
assign w20338 = pi2472 & pi3013;
assign w20339 = ~pi2472 & ~pi3013;
assign w20340 = ~pi2643 & ~pi2996;
assign w20341 = ~w20339 & w20340;
assign w20342 = ~w20338 & w20341;
assign w20343 = ~w20337 & w20342;
assign w20344 = pi2479 & ~pi3056;
assign w20345 = ~pi2479 & pi3056;
assign w20346 = pi2900 & ~w20345;
assign w20347 = ~w20344 & w20346;
assign w20348 = pi2400 & ~pi3014;
assign w20349 = ~pi2400 & pi3014;
assign w20350 = pi2997 & ~w20349;
assign w20351 = ~w20348 & w20350;
assign w20352 = ~w20347 & ~w20351;
assign w20353 = ~pi2483 & pi2977;
assign w20354 = pi2483 & ~pi2977;
assign w20355 = pi2907 & ~w20354;
assign w20356 = ~w20353 & w20355;
assign w20357 = pi2484 & ~pi3015;
assign w20358 = ~pi2484 & pi3015;
assign w20359 = pi2998 & ~w20358;
assign w20360 = ~w20357 & w20359;
assign w20361 = ~w20356 & ~w20360;
assign w20362 = w20352 & w20361;
assign w20363 = w20343 & w20362;
assign w20364 = ~pi2478 & pi3011;
assign w20365 = pi2478 & ~pi3011;
assign w20366 = pi2995 & ~w20365;
assign w20367 = ~w20364 & w20366;
assign w20368 = ~pi2517 & pi2786;
assign w20369 = pi2517 & ~pi2786;
assign w20370 = pi3000 & ~w20369;
assign w20371 = ~w20368 & w20370;
assign w20372 = ~w20367 & ~w20371;
assign w20373 = pi2516 & ~pi3016;
assign w20374 = ~pi2516 & pi3016;
assign w20375 = pi3001 & ~w20374;
assign w20376 = ~w20373 & w20375;
assign w20377 = pi2481 & ~pi2991;
assign w20378 = ~pi2481 & pi2991;
assign w20379 = pi3067 & ~w20378;
assign w20380 = ~w20377 & w20379;
assign w20381 = ~w20376 & ~w20380;
assign w20382 = w20372 & w20381;
assign w20383 = pi2475 & ~pi3009;
assign w20384 = ~pi2475 & pi3009;
assign w20385 = pi2954 & ~w20384;
assign w20386 = ~w20383 & w20385;
assign w20387 = pi2408 & ~pi2972;
assign w20388 = ~pi2408 & pi2972;
assign w20389 = pi2887 & ~w20388;
assign w20390 = ~w20387 & w20389;
assign w20391 = ~w20386 & ~w20390;
assign w20392 = pi2518 & ~pi2959;
assign w20393 = ~pi2518 & pi2959;
assign w20394 = pi2999 & ~w20393;
assign w20395 = ~w20392 & w20394;
assign w20396 = ~pi2480 & pi3108;
assign w20397 = pi2480 & ~pi3108;
assign w20398 = pi3072 & ~w20397;
assign w20399 = ~w20396 & w20398;
assign w20400 = ~w20395 & ~w20399;
assign w20401 = w20391 & w20400;
assign w20402 = pi2476 & ~pi3010;
assign w20403 = ~pi2476 & pi3010;
assign w20404 = pi2994 & ~w20403;
assign w20405 = ~w20402 & w20404;
assign w20406 = pi2485 & ~pi2886;
assign w20407 = ~pi2485 & pi2886;
assign w20408 = pi2901 & ~w20407;
assign w20409 = ~w20406 & w20408;
assign w20410 = ~w20405 & ~w20409;
assign w20411 = ~pi2514 & pi2984;
assign w20412 = pi2514 & ~pi2984;
assign w20413 = pi2908 & ~w20412;
assign w20414 = ~w20411 & w20413;
assign w20415 = pi2477 & ~pi3095;
assign w20416 = ~pi2477 & pi3095;
assign w20417 = pi2955 & ~w20416;
assign w20418 = ~w20415 & w20417;
assign w20419 = ~w20414 & ~w20418;
assign w20420 = w20410 & w20419;
assign w20421 = w20401 & w20420;
assign w20422 = w20382 & w20421;
assign w20423 = w20363 & w20422;
assign w20424 = pi2408 & ~pi2910;
assign w20425 = ~pi2408 & pi2910;
assign w20426 = pi2857 & ~w20425;
assign w20427 = ~w20424 & w20426;
assign w20428 = pi2472 & pi3022;
assign w20429 = ~pi2472 & ~pi3022;
assign w20430 = ~pi2643 & ~pi3005;
assign w20431 = ~w20429 & w20430;
assign w20432 = ~w20428 & w20431;
assign w20433 = ~w20427 & w20432;
assign w20434 = pi2477 & ~pi3066;
assign w20435 = ~pi2477 & pi3066;
assign w20436 = pi3003 & ~w20435;
assign w20437 = ~w20434 & w20436;
assign w20438 = ~pi2517 & pi3024;
assign w20439 = pi2517 & ~pi3024;
assign w20440 = pi3085 & ~w20439;
assign w20441 = ~w20438 & w20440;
assign w20442 = ~w20437 & ~w20441;
assign w20443 = ~pi2483 & pi3021;
assign w20444 = pi2483 & ~pi3021;
assign w20445 = pi2838 & ~w20444;
assign w20446 = ~w20443 & w20445;
assign w20447 = pi2484 & ~pi2906;
assign w20448 = ~pi2484 & pi2906;
assign w20449 = pi3007 & ~w20448;
assign w20450 = ~w20447 & w20449;
assign w20451 = ~w20446 & ~w20450;
assign w20452 = w20442 & w20451;
assign w20453 = w20433 & w20452;
assign w20454 = pi2476 & ~pi3017;
assign w20455 = ~pi2476 & pi3017;
assign w20456 = pi3002 & ~w20455;
assign w20457 = ~w20454 & w20456;
assign w20458 = pi2514 & ~pi2909;
assign w20459 = ~pi2514 & pi2909;
assign w20460 = pi2858 & ~w20459;
assign w20461 = ~w20458 & w20460;
assign w20462 = ~w20457 & ~w20461;
assign w20463 = pi2516 & ~pi3025;
assign w20464 = ~pi2516 & pi3025;
assign w20465 = pi3008 & ~w20464;
assign w20466 = ~w20463 & w20465;
assign w20467 = pi2480 & ~pi3019;
assign w20468 = ~pi2480 & pi3019;
assign w20469 = pi2821 & ~w20468;
assign w20470 = ~w20467 & w20469;
assign w20471 = ~w20466 & ~w20470;
assign w20472 = w20462 & w20471;
assign w20473 = ~pi2482 & pi3020;
assign w20474 = pi2482 & ~pi3020;
assign w20475 = pi2839 & ~w20474;
assign w20476 = ~w20473 & w20475;
assign w20477 = pi2400 & ~pi2837;
assign w20478 = ~pi2400 & pi2837;
assign w20479 = pi3006 & ~w20478;
assign w20480 = ~w20477 & w20479;
assign w20481 = ~w20476 & ~w20480;
assign w20482 = pi2478 & ~pi3018;
assign w20483 = ~pi2478 & pi3018;
assign w20484 = pi3004 & ~w20483;
assign w20485 = ~w20482 & w20484;
assign w20486 = pi2479 & ~pi2956;
assign w20487 = ~pi2479 & pi2956;
assign w20488 = pi2884 & ~w20487;
assign w20489 = ~w20486 & w20488;
assign w20490 = ~w20485 & ~w20489;
assign w20491 = w20481 & w20490;
assign w20492 = pi2518 & ~pi3023;
assign w20493 = ~pi2518 & pi3023;
assign w20494 = pi3077 & ~w20493;
assign w20495 = ~w20492 & w20494;
assign w20496 = ~pi2481 & pi2790;
assign w20497 = pi2481 & ~pi2790;
assign w20498 = pi2822 & ~w20497;
assign w20499 = ~w20496 & w20498;
assign w20500 = ~w20495 & ~w20499;
assign w20501 = pi2485 & ~pi2885;
assign w20502 = ~pi2485 & pi2885;
assign w20503 = pi3094 & ~w20502;
assign w20504 = ~w20501 & w20503;
assign w20505 = ~pi2475 & pi2815;
assign w20506 = pi2475 & ~pi2815;
assign w20507 = pi2880 & ~w20506;
assign w20508 = ~w20505 & w20507;
assign w20509 = ~w20504 & ~w20508;
assign w20510 = w20500 & w20509;
assign w20511 = w20491 & w20510;
assign w20512 = w20472 & w20511;
assign w20513 = w20453 & w20512;
assign w20514 = pi2800 & ~pi3362;
assign w20515 = ~pi3643 & ~pi3644;
assign w20516 = w20514 & w20515;
assign w20517 = pi0408 & ~pi2762;
assign w20518 = w2231 & w20517;
assign w20519 = w381 & w20518;
assign w20520 = ~w20516 & ~w20519;
assign w20521 = ~w20513 & w20520;
assign w20522 = ~w20423 & w20521;
assign w20523 = ~w20333 & w20522;
assign w20524 = w19964 & ~w20523;
assign w20525 = ~pi0404 & ~w20524;
assign w20526 = w323 & w932;
assign w20527 = w6681 & w20526;
assign w20528 = w0 & w20527;
assign w20529 = ~w20525 & w20528;
assign w20530 = ~w19582 & ~w19954;
assign w20531 = ~pi0405 & ~w19958;
assign w20532 = ~pi0858 & w19958;
assign w20533 = ~w20531 & ~w20532;
assign w20534 = w19954 & w20533;
assign w20535 = ~w20530 & ~w20534;
assign w20536 = ~w19638 & ~w19954;
assign w20537 = ~pi0406 & ~w19958;
assign w20538 = ~pi0730 & w19958;
assign w20539 = ~w20537 & ~w20538;
assign w20540 = w19954 & w20539;
assign w20541 = ~w20536 & ~w20540;
assign w20542 = ~w19847 & ~w19954;
assign w20543 = pi0407 & ~w19958;
assign w20544 = pi1052 & w19958;
assign w20545 = ~w20543 & ~w20544;
assign w20546 = w19954 & w20545;
assign w20547 = ~w20542 & ~w20546;
assign w20548 = ~w19766 & ~w19954;
assign w20549 = ~pi0408 & ~w19958;
assign w20550 = pi1045 & w19958;
assign w20551 = ~w20549 & ~w20550;
assign w20552 = w19954 & w20551;
assign w20553 = ~w20548 & ~w20552;
assign w20554 = ~w19648 & ~w19954;
assign w20555 = ~pi0409 & ~w19958;
assign w20556 = ~pi0851 & w19958;
assign w20557 = ~w20555 & ~w20556;
assign w20558 = w19954 & w20557;
assign w20559 = ~w20554 & ~w20558;
assign w20560 = ~w19658 & ~w19954;
assign w20561 = ~pi0410 & ~w19958;
assign w20562 = ~pi0860 & w19958;
assign w20563 = ~w20561 & ~w20562;
assign w20564 = w19954 & w20563;
assign w20565 = ~w20560 & ~w20564;
assign w20566 = ~w19685 & ~w19954;
assign w20567 = ~pi0411 & ~w19958;
assign w20568 = ~pi0852 & w19958;
assign w20569 = ~w20567 & ~w20568;
assign w20570 = w19954 & w20569;
assign w20571 = ~w20566 & ~w20570;
assign w20572 = ~w19712 & ~w19954;
assign w20573 = ~pi0412 & ~w19958;
assign w20574 = ~pi0821 & w19958;
assign w20575 = ~w20573 & ~w20574;
assign w20576 = w19954 & w20575;
assign w20577 = ~w20572 & ~w20576;
assign w20578 = ~w19739 & ~w19954;
assign w20579 = ~pi0413 & ~w19958;
assign w20580 = pi0937 & w19958;
assign w20581 = ~w20579 & ~w20580;
assign w20582 = w19954 & w20581;
assign w20583 = ~w20578 & ~w20582;
assign w20584 = ~w19793 & ~w19954;
assign w20585 = ~pi0414 & ~w19958;
assign w20586 = pi1082 & w19958;
assign w20587 = ~w20585 & ~w20586;
assign w20588 = w19954 & w20587;
assign w20589 = ~w20584 & ~w20588;
assign w20590 = ~w19820 & ~w19954;
assign w20591 = ~pi0415 & ~w19958;
assign w20592 = pi1080 & w19958;
assign w20593 = ~w20591 & ~w20592;
assign w20594 = w19954 & w20593;
assign w20595 = ~w20590 & ~w20594;
assign w20596 = ~w19621 & ~w19954;
assign w20597 = ~pi0416 & ~w19958;
assign w20598 = ~pi0853 & w19958;
assign w20599 = ~w20597 & ~w20598;
assign w20600 = w19954 & w20599;
assign w20601 = ~w20596 & ~w20600;
assign w20602 = ~w19629 & ~w19954;
assign w20603 = ~pi0417 & ~w19958;
assign w20604 = ~pi0854 & w19958;
assign w20605 = ~w20603 & ~w20604;
assign w20606 = w19954 & w20605;
assign w20607 = ~w20602 & ~w20606;
assign w20608 = ~w19550 & ~w19954;
assign w20609 = ~pi0418 & ~w19958;
assign w20610 = ~pi0825 & w19958;
assign w20611 = ~w20609 & ~w20610;
assign w20612 = w19954 & w20611;
assign w20613 = ~w20608 & ~w20612;
assign w20614 = ~w19558 & ~w19954;
assign w20615 = ~pi0419 & ~w19958;
assign w20616 = ~pi0855 & w19958;
assign w20617 = ~w20615 & ~w20616;
assign w20618 = w19954 & w20617;
assign w20619 = ~w20614 & ~w20618;
assign w20620 = ~w19566 & ~w19954;
assign w20621 = ~pi0420 & ~w19958;
assign w20622 = ~pi0856 & w19958;
assign w20623 = ~w20621 & ~w20622;
assign w20624 = w19954 & w20623;
assign w20625 = ~w20620 & ~w20624;
assign w20626 = ~w19574 & ~w19954;
assign w20627 = ~pi0421 & ~w19958;
assign w20628 = ~pi0857 & w19958;
assign w20629 = ~w20627 & ~w20628;
assign w20630 = w19954 & w20629;
assign w20631 = ~w20626 & ~w20630;
assign w20632 = ~w19592 & ~w19954;
assign w20633 = ~pi0422 & ~w19958;
assign w20634 = ~pi0824 & w19958;
assign w20635 = ~w20633 & ~w20634;
assign w20636 = w19954 & w20635;
assign w20637 = ~w20632 & ~w20636;
assign w20638 = ~w19602 & ~w19954;
assign w20639 = ~pi0423 & ~w19958;
assign w20640 = ~pi0823 & w19958;
assign w20641 = ~w20639 & ~w20640;
assign w20642 = w19954 & w20641;
assign w20643 = ~w20638 & ~w20642;
assign w20644 = ~w19612 & ~w19954;
assign w20645 = ~pi0424 & ~w19958;
assign w20646 = ~pi0859 & w19958;
assign w20647 = ~w20645 & ~w20646;
assign w20648 = w19954 & w20647;
assign w20649 = ~w20644 & ~w20648;
assign w20650 = ~w19857 & ~w19954;
assign w20651 = ~pi0425 & ~w19958;
assign w20652 = ~pi0731 & w19958;
assign w20653 = ~w20651 & ~w20652;
assign w20654 = w19954 & w20653;
assign w20655 = ~w20650 & ~w20654;
assign w20656 = ~w19867 & ~w19954;
assign w20657 = ~pi0426 & ~w19958;
assign w20658 = ~pi0938 & w19958;
assign w20659 = ~w20657 & ~w20658;
assign w20660 = w19954 & w20659;
assign w20661 = ~w20656 & ~w20660;
assign w20662 = ~w19894 & ~w19954;
assign w20663 = pi0427 & ~w19958;
assign w20664 = pi0911 & w19958;
assign w20665 = ~w20663 & ~w20664;
assign w20666 = w19954 & w20665;
assign w20667 = ~w20662 & ~w20666;
assign w20668 = w19033 & w19041;
assign w20669 = ~pi0975 & ~pi1422;
assign w20670 = ~pi1771 & ~pi3580;
assign w20671 = pi3581 & w20670;
assign w20672 = w20669 & ~w20671;
assign w20673 = w19039 & w20672;
assign w20674 = ~w20668 & ~w20673;
assign w20675 = ~pi0428 & w20674;
assign w20676 = w19094 & ~w19709;
assign w20677 = ~w19174 & ~w20674;
assign w20678 = ~w20676 & w20677;
assign w20679 = ~w20675 & ~w20678;
assign w20680 = ~pi0429 & w20674;
assign w20681 = w19094 & ~w19736;
assign w20682 = ~pi3475 & ~w2250;
assign w20683 = ~w20674 & ~w20682;
assign w20684 = ~w20681 & w20683;
assign w20685 = ~w20680 & ~w20684;
assign w20686 = ~pi0430 & w20674;
assign w20687 = w19094 & ~w19763;
assign w20688 = ~pi3470 & ~w2250;
assign w20689 = ~w20674 & ~w20688;
assign w20690 = ~w20687 & w20689;
assign w20691 = ~w20686 & ~w20690;
assign w20692 = ~pi0431 & w20674;
assign w20693 = w19094 & ~w19790;
assign w20694 = ~pi3446 & ~w2250;
assign w20695 = ~w20674 & ~w20694;
assign w20696 = ~w20693 & w20695;
assign w20697 = ~w20692 & ~w20696;
assign w20698 = ~pi0432 & w20674;
assign w20699 = w19094 & ~w19817;
assign w20700 = ~w19278 & ~w20674;
assign w20701 = ~w20699 & w20700;
assign w20702 = ~w20698 & ~w20701;
assign w20703 = ~pi0433 & w20674;
assign w20704 = w19094 & ~w19844;
assign w20705 = ~w19306 & ~w20674;
assign w20706 = ~w20704 & w20705;
assign w20707 = ~w20703 & ~w20706;
assign w20708 = ~pi0434 & w20674;
assign w20709 = w19094 & ~w19891;
assign w20710 = ~pi3464 & ~w2250;
assign w20711 = ~w20674 & ~w20710;
assign w20712 = ~w20709 & w20711;
assign w20713 = ~w20708 & ~w20712;
assign w20714 = ~pi0435 & w20674;
assign w20715 = w19094 & ~w19682;
assign w20716 = ~pi3477 & ~w2250;
assign w20717 = ~w20674 & ~w20716;
assign w20718 = ~w20715 & w20717;
assign w20719 = ~w20714 & ~w20718;
assign w20720 = pi0436 & ~w18412;
assign w20721 = ~w15014 & ~w17425;
assign w20722 = w17080 & w17425;
assign w20723 = ~w20721 & ~w20722;
assign w20724 = w18412 & ~w20723;
assign w20725 = ~w20720 & ~w20724;
assign w20726 = pi0437 & ~w18419;
assign w20727 = w18419 & ~w20723;
assign w20728 = ~w20726 & ~w20727;
assign w20729 = pi0438 & ~pi3419;
assign w20730 = w2896 & w4141;
assign w20731 = w898 & w7505;
assign w20732 = ~w891 & w897;
assign w20733 = ~w19301 & w20732;
assign w20734 = pi3419 & ~w20733;
assign w20735 = ~w20731 & w20734;
assign w20736 = ~w20730 & w20735;
assign w20737 = ~w20729 & ~w20736;
assign w20738 = pi0439 & ~pi3419;
assign w20739 = w2896 & w6177;
assign w20740 = w898 & w7473;
assign w20741 = ~w19492 & w20732;
assign w20742 = pi3419 & ~w20741;
assign w20743 = ~w20740 & w20742;
assign w20744 = ~w20739 & w20743;
assign w20745 = ~w20738 & ~w20744;
assign w20746 = pi0440 & ~pi3419;
assign w20747 = w2896 & w3195;
assign w20748 = ~w19682 & w20732;
assign w20749 = pi3419 & ~w20748;
assign w20750 = ~w20747 & w20749;
assign w20751 = ~w20746 & ~w20750;
assign w20752 = pi0441 & ~pi3419;
assign w20753 = w2896 & w40134;
assign w20754 = ~w19709 & w20732;
assign w20755 = pi3419 & ~w20754;
assign w20756 = ~w20753 & w20755;
assign w20757 = ~w20752 & ~w20756;
assign w20758 = pi0442 & ~pi3419;
assign w20759 = w2896 & w6413;
assign w20760 = ~w19736 & w20732;
assign w20761 = pi3419 & ~w20760;
assign w20762 = ~w20759 & w20761;
assign w20763 = ~w20758 & ~w20762;
assign w20764 = pi0443 & ~pi3419;
assign w20765 = w2896 & w4380;
assign w20766 = ~w19763 & w20732;
assign w20767 = pi3419 & ~w20766;
assign w20768 = ~w20765 & w20767;
assign w20769 = ~w20764 & ~w20768;
assign w20770 = pi0444 & ~pi3419;
assign w20771 = w2896 & w5320;
assign w20772 = ~w19790 & w20732;
assign w20773 = pi3419 & ~w20772;
assign w20774 = ~w20771 & w20773;
assign w20775 = ~w20770 & ~w20774;
assign w20776 = pi0445 & ~pi3419;
assign w20777 = w898 & w8266;
assign w20778 = ~w19329 & w20732;
assign w20779 = pi3419 & ~w20778;
assign w20780 = ~w20777 & w20779;
assign w20781 = ~w20776 & ~w20780;
assign w20782 = pi0446 & ~pi3419;
assign w20783 = w898 & w7994;
assign w20784 = ~w19356 & w20732;
assign w20785 = pi3419 & ~w20784;
assign w20786 = ~w20783 & w20785;
assign w20787 = ~w20782 & ~w20786;
assign w20788 = pi0447 & ~pi3419;
assign w20789 = w898 & w7892;
assign w20790 = ~w19383 & w20732;
assign w20791 = pi3419 & ~w20790;
assign w20792 = ~w20789 & w20791;
assign w20793 = ~w20788 & ~w20792;
assign w20794 = pi0448 & ~pi3419;
assign w20795 = w898 & w7860;
assign w20796 = ~w19410 & w20732;
assign w20797 = pi3419 & ~w20796;
assign w20798 = ~w20795 & w20797;
assign w20799 = ~w20794 & ~w20798;
assign w20800 = pi0449 & ~pi3419;
assign w20801 = w2896 & w4749;
assign w20802 = ~w19844 & w20732;
assign w20803 = pi3419 & ~w20802;
assign w20804 = ~w20801 & w20803;
assign w20805 = ~w20800 & ~w20804;
assign w20806 = pi0450 & ~pi3419;
assign w20807 = w898 & w7828;
assign w20808 = ~w19438 & w20732;
assign w20809 = pi3419 & ~w20808;
assign w20810 = ~w20807 & w20809;
assign w20811 = ~w20806 & ~w20810;
assign w20812 = pi0451 & ~pi3419;
assign w20813 = w898 & w7796;
assign w20814 = ~w19465 & w20732;
assign w20815 = pi3419 & ~w20814;
assign w20816 = ~w20813 & w20815;
assign w20817 = ~w20812 & ~w20816;
assign w20818 = pi0452 & ~pi3419;
assign w20819 = w898 & w7732;
assign w20820 = ~w19119 & w20732;
assign w20821 = pi3419 & ~w20820;
assign w20822 = ~w20819 & w20821;
assign w20823 = ~w20818 & ~w20822;
assign w20824 = pi0453 & ~pi3419;
assign w20825 = w2896 & w8240;
assign w20826 = w898 & w7700;
assign w20827 = ~w19144 & w20732;
assign w20828 = pi3419 & ~w20827;
assign w20829 = ~w20826 & w20828;
assign w20830 = ~w20825 & w20829;
assign w20831 = ~w20824 & ~w20830;
assign w20832 = pi0454 & ~pi3419;
assign w20833 = w2896 & w8081;
assign w20834 = w898 & w7668;
assign w20835 = ~w19170 & w20732;
assign w20836 = pi3419 & ~w20835;
assign w20837 = ~w20834 & w20836;
assign w20838 = ~w20833 & w20837;
assign w20839 = ~w20832 & ~w20838;
assign w20840 = pi0455 & ~pi3419;
assign w20841 = w1308 & w2896;
assign w20842 = w898 & w7602;
assign w20843 = ~w19221 & w20732;
assign w20844 = pi3419 & ~w20843;
assign w20845 = ~w20842 & w20844;
assign w20846 = ~w20841 & w20845;
assign w20847 = ~w20840 & ~w20846;
assign w20848 = pi0456 & ~pi3419;
assign w20849 = w2896 & w5635;
assign w20850 = w898 & w7570;
assign w20851 = ~w19246 & w20732;
assign w20852 = pi3419 & ~w20851;
assign w20853 = ~w20850 & w20852;
assign w20854 = ~w20849 & w20853;
assign w20855 = ~w20848 & ~w20854;
assign w20856 = pi0457 & ~pi3419;
assign w20857 = w2896 & w5053;
assign w20858 = w898 & w7537;
assign w20859 = ~w19273 & w20732;
assign w20860 = pi3419 & ~w20859;
assign w20861 = ~w20858 & w20860;
assign w20862 = ~w20857 & w20861;
assign w20863 = ~w20856 & ~w20862;
assign w20864 = ~pi2091 & w18313;
assign w20865 = pi0458 & w18336;
assign w20866 = ~w18337 & ~w18359;
assign w20867 = ~w20865 & w20866;
assign w20868 = ~pi1878 & w18359;
assign w20869 = ~w18313 & ~w20868;
assign w20870 = ~w20867 & w20869;
assign w20871 = ~w20864 & ~w20870;
assign w20872 = pi0459 & ~pi3419;
assign w20873 = w2896 & w5914;
assign w20874 = ~w19817 & w20732;
assign w20875 = pi3419 & ~w20874;
assign w20876 = ~w20873 & w20875;
assign w20877 = ~w20872 & ~w20876;
assign w20878 = pi0460 & ~pi3419;
assign w20879 = w2896 & w3711;
assign w20880 = ~w19891 & w20732;
assign w20881 = pi3419 & ~w20880;
assign w20882 = ~w20879 & w20881;
assign w20883 = ~w20878 & ~w20882;
assign w20884 = pi0461 & ~pi3419;
assign w20885 = w1639 & w2896;
assign w20886 = w898 & w7635;
assign w20887 = ~w19196 & w20732;
assign w20888 = pi3419 & ~w20887;
assign w20889 = ~w20886 & w20888;
assign w20890 = ~w20885 & w20889;
assign w20891 = ~w20884 & ~w20890;
assign w20892 = pi0462 & ~pi3419;
assign w20893 = w898 & w7764;
assign w20894 = ~w19093 & w20732;
assign w20895 = pi3419 & ~w20894;
assign w20896 = ~w20893 & w20895;
assign w20897 = ~w20892 & ~w20896;
assign w20898 = pi0463 & ~w18412;
assign w20899 = w17080 & ~w17425;
assign w20900 = w8211 & w17425;
assign w20901 = ~w20899 & ~w20900;
assign w20902 = w18412 & ~w20901;
assign w20903 = ~w20898 & ~w20902;
assign w20904 = pi0464 & ~w18419;
assign w20905 = w18419 & ~w20901;
assign w20906 = ~w20904 & ~w20905;
assign w20907 = pi0887 & pi1739;
assign w20908 = pi0888 & pi3667;
assign w20909 = ~pi0888 & ~pi3667;
assign w20910 = ~pi0887 & ~w20909;
assign w20911 = ~w20908 & w20910;
assign w20912 = ~w20907 & ~w20911;
assign w20913 = pi0790 & ~w314;
assign w20914 = ~pi0790 & pi3670;
assign w20915 = ~w20913 & ~w20914;
assign w20916 = ~pi0881 & w20915;
assign w20917 = pi0881 & ~w20915;
assign w20918 = ~w20916 & ~w20917;
assign w20919 = pi3249 & pi3647;
assign w20920 = w20918 & w20919;
assign w20921 = ~pi0889 & ~w20920;
assign w20922 = pi0889 & ~pi3550;
assign w20923 = ~pi0791 & ~w20922;
assign w20924 = ~w20921 & w20923;
assign w20925 = pi0889 & ~pi3493;
assign w20926 = ~pi0889 & pi2387;
assign w20927 = pi0791 & ~w20926;
assign w20928 = ~w20925 & w20927;
assign w20929 = ~pi0654 & ~w20928;
assign w20930 = ~w20924 & w20929;
assign w20931 = pi0526 & pi0531;
assign w20932 = pi0525 & pi0527;
assign w20933 = pi0554 & w20932;
assign w20934 = w20931 & w20933;
assign w20935 = ~w20930 & ~w20934;
assign w20936 = ~pi0696 & w20935;
assign w20937 = ~pi0882 & ~pi0883;
assign w20938 = ~pi0543 & ~w20937;
assign w20939 = w20936 & w20938;
assign w20940 = ~pi0474 & pi0543;
assign w20941 = w20935 & w20940;
assign w20942 = ~pi0465 & ~w20935;
assign w20943 = ~w20941 & ~w20942;
assign w20944 = ~w20939 & w20943;
assign w20945 = ~pi0478 & pi0543;
assign w20946 = w20935 & w20945;
assign w20947 = ~pi0466 & ~w20935;
assign w20948 = ~w20946 & ~w20947;
assign w20949 = ~w20939 & w20948;
assign w20950 = ~pi0466 & pi0543;
assign w20951 = w20935 & w20950;
assign w20952 = ~pi0467 & ~w20935;
assign w20953 = ~w20951 & ~w20952;
assign w20954 = ~w20939 & w20953;
assign w20955 = ~pi0467 & pi0543;
assign w20956 = w20935 & w20955;
assign w20957 = ~pi0468 & ~w20935;
assign w20958 = ~w20956 & ~w20957;
assign w20959 = ~w20939 & w20958;
assign w20960 = ~pi0468 & pi0543;
assign w20961 = w20935 & w20960;
assign w20962 = ~pi0469 & ~w20935;
assign w20963 = ~w20961 & ~w20962;
assign w20964 = ~w20939 & w20963;
assign w20965 = ~pi0469 & pi0543;
assign w20966 = w20935 & w20965;
assign w20967 = ~pi0470 & ~w20935;
assign w20968 = ~w20966 & ~w20967;
assign w20969 = ~w20939 & w20968;
assign w20970 = ~pi0470 & pi0543;
assign w20971 = w20935 & w20970;
assign w20972 = ~pi0471 & ~w20935;
assign w20973 = ~w20971 & ~w20972;
assign w20974 = ~w20939 & w20973;
assign w20975 = pi0543 & ~pi0697;
assign w20976 = w20935 & w20975;
assign w20977 = ~pi0472 & ~w20935;
assign w20978 = ~w20976 & ~w20977;
assign w20979 = ~w20939 & w20978;
assign w20980 = ~pi0472 & pi0543;
assign w20981 = w20935 & w20980;
assign w20982 = ~pi0473 & ~w20935;
assign w20983 = ~w20981 & ~w20982;
assign w20984 = ~w20939 & w20983;
assign w20985 = ~pi0473 & pi0543;
assign w20986 = w20935 & w20985;
assign w20987 = ~pi0474 & ~w20935;
assign w20988 = ~w20986 & ~w20987;
assign w20989 = ~w20939 & w20988;
assign w20990 = ~pi0465 & pi0543;
assign w20991 = w20935 & w20990;
assign w20992 = ~pi0475 & ~w20935;
assign w20993 = ~w20991 & ~w20992;
assign w20994 = ~w20939 & w20993;
assign w20995 = ~pi0475 & pi0543;
assign w20996 = w20935 & w20995;
assign w20997 = ~pi0476 & ~w20935;
assign w20998 = ~w20996 & ~w20997;
assign w20999 = ~w20939 & w20998;
assign w21000 = ~pi0476 & pi0543;
assign w21001 = w20935 & w21000;
assign w21002 = ~pi0477 & ~w20935;
assign w21003 = ~w21001 & ~w21002;
assign w21004 = ~w20939 & w21003;
assign w21005 = ~pi0477 & pi0543;
assign w21006 = w20935 & w21005;
assign w21007 = ~pi0478 & ~w20935;
assign w21008 = ~w21006 & ~w21007;
assign w21009 = ~w20939 & w21008;
assign w21010 = pi0479 & ~w18375;
assign w21011 = pi2599 & w3711;
assign w21012 = ~w17866 & w18366;
assign w21013 = ~w17955 & w21012;
assign w21014 = ~w18003 & ~w21013;
assign w21015 = ~w21011 & w21014;
assign w21016 = pi0693 & w18003;
assign w21017 = ~w18012 & ~w21016;
assign w21018 = ~w21015 & w21017;
assign w21019 = ~w21010 & ~w21018;
assign w21020 = pi0480 & ~w18928;
assign w21021 = pi0712 & ~w18150;
assign w21022 = ~pi0712 & ~w40176;
assign w21023 = ~w21021 & ~w21022;
assign w21024 = w18928 & w21023;
assign w21025 = ~w21020 & ~w21024;
assign w21026 = pi0481 & ~w18935;
assign w21027 = w18935 & w21023;
assign w21028 = ~w21026 & ~w21027;
assign w21029 = w13981 & w13989;
assign w21030 = w14002 & w21029;
assign w21031 = w6689 & w21030;
assign w21032 = ~pi3330 & pi3394;
assign w21033 = pi2763 & w2307;
assign w21034 = w21032 & w21033;
assign w21035 = pi0832 & pi0921;
assign w21036 = ~pi2487 & pi3392;
assign w21037 = w21035 & ~w21036;
assign w21038 = ~w21034 & w21037;
assign w21039 = ~w21031 & w21038;
assign w21040 = ~w370 & ~w21039;
assign w21041 = pi0482 & ~w21040;
assign w21042 = w6413 & ~w21035;
assign w21043 = ~w2195 & w21031;
assign w21044 = pi0482 & w21034;
assign w21045 = ~w21036 & ~w21044;
assign w21046 = ~w21043 & w21045;
assign w21047 = pi0615 & ~w21046;
assign w21048 = ~pi0585 & ~pi0632;
assign w21049 = ~pi0592 & w21048;
assign w21050 = ~pi0603 & w21049;
assign w21051 = ~pi0591 & w21050;
assign w21052 = ~pi0578 & w21051;
assign w21053 = pi0578 & ~w21051;
assign w21054 = ~w21052 & ~w21053;
assign w21055 = ~w21047 & w21054;
assign w21056 = pi0647 & pi1709;
assign w21057 = ~pi0647 & pi1865;
assign w21058 = ~pi0616 & ~w21057;
assign w21059 = ~w21056 & w21058;
assign w21060 = pi0616 & pi0647;
assign w21061 = ~pi1864 & w21060;
assign w21062 = pi0616 & ~pi0647;
assign w21063 = ~pi1811 & w21062;
assign w21064 = ~w21061 & ~w21063;
assign w21065 = ~w21059 & w21064;
assign w21066 = w21047 & w21065;
assign w21067 = w21035 & ~w21066;
assign w21068 = ~w21055 & w21067;
assign w21069 = ~w21042 & ~w21068;
assign w21070 = w5635 & ~w21035;
assign w21071 = pi0647 & pi1664;
assign w21072 = ~pi0647 & pi1809;
assign w21073 = ~pi0616 & ~w21072;
assign w21074 = ~w21071 & w21073;
assign w21075 = ~pi1819 & w21060;
assign w21076 = ~pi1656 & w21062;
assign w21077 = ~w21075 & ~w21076;
assign w21078 = ~w21074 & w21077;
assign w21079 = w21047 & w21078;
assign w21080 = ~pi0572 & w21052;
assign w21081 = ~pi0571 & w21080;
assign w21082 = ~pi0602 & w21081;
assign w21083 = ~pi0590 & w21082;
assign w21084 = ~pi0594 & w21083;
assign w21085 = ~pi0595 & w21084;
assign w21086 = pi0595 & ~w21084;
assign w21087 = ~w21085 & ~w21086;
assign w21088 = ~w21047 & w21087;
assign w21089 = w21035 & ~w21088;
assign w21090 = ~w21079 & w21089;
assign w21091 = ~w21070 & ~w21090;
assign w21092 = w5053 & ~w21035;
assign w21093 = pi0647 & pi1632;
assign w21094 = ~pi0647 & pi1710;
assign w21095 = ~pi0616 & ~w21094;
assign w21096 = ~w21093 & w21095;
assign w21097 = ~pi1820 & w21060;
assign w21098 = ~pi1634 & w21062;
assign w21099 = ~w21097 & ~w21098;
assign w21100 = ~w21096 & w21099;
assign w21101 = w21047 & w21100;
assign w21102 = pi0594 & ~w21083;
assign w21103 = ~w21084 & ~w21102;
assign w21104 = ~w21047 & w21103;
assign w21105 = w21035 & ~w21104;
assign w21106 = ~w21101 & w21105;
assign w21107 = ~w21092 & ~w21106;
assign w21108 = w21091 & w21107;
assign w21109 = w21069 & w21108;
assign w21110 = ~w3711 & ~w21035;
assign w21111 = pi0647 & ~pi1665;
assign w21112 = ~pi0647 & ~pi1810;
assign w21113 = ~pi0616 & ~w21112;
assign w21114 = ~w21111 & w21113;
assign w21115 = pi1657 & w21062;
assign w21116 = pi1821 & w21060;
assign w21117 = ~w21115 & ~w21116;
assign w21118 = ~w21114 & w21117;
assign w21119 = w21047 & w21118;
assign w21120 = ~pi0585 & ~w21047;
assign w21121 = w21035 & ~w21120;
assign w21122 = ~w21119 & w21121;
assign w21123 = w21040 & ~w21122;
assign w21124 = ~w21110 & w21123;
assign w21125 = ~w4749 & ~w21035;
assign w21126 = pi0647 & ~pi1630;
assign w21127 = ~pi0647 & ~pi1711;
assign w21128 = ~pi0616 & ~w21127;
assign w21129 = ~w21126 & w21128;
assign w21130 = pi1817 & w21060;
assign w21131 = pi1638 & w21062;
assign w21132 = ~w21130 & ~w21131;
assign w21133 = ~w21129 & w21132;
assign w21134 = w21047 & w21133;
assign w21135 = pi0585 & pi0632;
assign w21136 = ~w21048 & ~w21135;
assign w21137 = ~w21047 & ~w21136;
assign w21138 = w21035 & ~w21137;
assign w21139 = ~w21134 & w21138;
assign w21140 = ~w21125 & ~w21139;
assign w21141 = w21124 & ~w21140;
assign w21142 = w5914 & ~w21035;
assign w21143 = pi0647 & pi1662;
assign w21144 = ~pi0647 & pi1806;
assign w21145 = ~pi0616 & ~w21144;
assign w21146 = ~w21143 & w21145;
assign w21147 = ~pi1816 & w21060;
assign w21148 = ~pi1654 & w21062;
assign w21149 = ~w21147 & ~w21148;
assign w21150 = ~w21146 & w21149;
assign w21151 = w21047 & w21150;
assign w21152 = pi0592 & ~w21048;
assign w21153 = ~w21049 & ~w21152;
assign w21154 = ~w21047 & w21153;
assign w21155 = w21035 & ~w21154;
assign w21156 = ~w21151 & w21155;
assign w21157 = ~w21142 & ~w21156;
assign w21158 = w40134 & ~w21035;
assign w21159 = pi0647 & pi1659;
assign w21160 = ~pi0647 & pi1803;
assign w21161 = ~pi0616 & ~w21160;
assign w21162 = ~w21159 & w21161;
assign w21163 = ~pi1814 & w21060;
assign w21164 = ~pi1652 & w21062;
assign w21165 = ~w21163 & ~w21164;
assign w21166 = ~w21162 & w21165;
assign w21167 = w21047 & w21166;
assign w21168 = pi0572 & ~w21052;
assign w21169 = ~w21080 & ~w21168;
assign w21170 = ~w21047 & w21169;
assign w21171 = w21035 & ~w21170;
assign w21172 = ~w21167 & w21171;
assign w21173 = ~w21158 & ~w21172;
assign w21174 = w21157 & w21173;
assign w21175 = w21141 & w21174;
assign w21176 = w21109 & w21175;
assign w21177 = w6177 & ~w21035;
assign w21178 = pi0647 & pi1658;
assign w21179 = ~pi0647 & pi1801;
assign w21180 = ~pi0616 & ~w21179;
assign w21181 = ~w21178 & w21180;
assign w21182 = ~pi1813 & w21060;
assign w21183 = ~pi1651 & w21062;
assign w21184 = ~w21182 & ~w21183;
assign w21185 = ~w21181 & w21184;
assign w21186 = w21047 & w21185;
assign w21187 = pi0602 & ~w21081;
assign w21188 = ~w21082 & ~w21187;
assign w21189 = ~w21047 & w21188;
assign w21190 = w21035 & ~w21189;
assign w21191 = ~w21186 & w21190;
assign w21192 = ~w21177 & ~w21191;
assign w21193 = w4380 & ~w21035;
assign w21194 = pi0591 & ~w21050;
assign w21195 = ~w21051 & ~w21194;
assign w21196 = ~w21047 & w21195;
assign w21197 = pi0647 & pi1660;
assign w21198 = ~pi0647 & pi1804;
assign w21199 = ~pi0616 & ~w21198;
assign w21200 = ~w21197 & w21199;
assign w21201 = ~pi1815 & w21060;
assign w21202 = ~pi1653 & w21062;
assign w21203 = ~w21201 & ~w21202;
assign w21204 = ~w21200 & w21203;
assign w21205 = w21047 & w21204;
assign w21206 = w21035 & ~w21205;
assign w21207 = ~w21196 & w21206;
assign w21208 = ~w21193 & ~w21207;
assign w21209 = w3195 & ~w21035;
assign w21210 = pi0647 & pi1633;
assign w21211 = ~pi0647 & pi1802;
assign w21212 = ~pi0616 & ~w21211;
assign w21213 = ~w21210 & w21212;
assign w21214 = ~pi1708 & w21060;
assign w21215 = ~pi1639 & w21062;
assign w21216 = ~w21214 & ~w21215;
assign w21217 = ~w21213 & w21216;
assign w21218 = w21047 & w21217;
assign w21219 = pi0571 & ~w21080;
assign w21220 = ~w21081 & ~w21219;
assign w21221 = ~w21047 & w21220;
assign w21222 = w21035 & ~w21221;
assign w21223 = ~w21218 & w21222;
assign w21224 = ~w21209 & ~w21223;
assign w21225 = w21208 & w21224;
assign w21226 = w21192 & w21225;
assign w21227 = w1308 & ~w21035;
assign w21228 = pi0647 & pi1631;
assign w21229 = ~pi0647 & pi1808;
assign w21230 = ~pi0616 & ~w21229;
assign w21231 = ~w21228 & w21230;
assign w21232 = ~pi1859 & w21060;
assign w21233 = ~pi1636 & w21062;
assign w21234 = ~w21232 & ~w21233;
assign w21235 = ~w21231 & w21234;
assign w21236 = w21047 & w21235;
assign w21237 = pi0593 & ~w21085;
assign w21238 = ~pi0593 & w21085;
assign w21239 = ~w21237 & ~w21238;
assign w21240 = ~w21047 & w21239;
assign w21241 = w21035 & ~w21240;
assign w21242 = ~w21236 & w21241;
assign w21243 = ~w21227 & ~w21242;
assign w21244 = w5320 & ~w21035;
assign w21245 = pi0603 & ~w21049;
assign w21246 = ~w21050 & ~w21245;
assign w21247 = ~w21047 & w21246;
assign w21248 = pi0647 & pi1661;
assign w21249 = ~pi0647 & pi1805;
assign w21250 = ~pi0616 & ~w21249;
assign w21251 = ~w21248 & w21250;
assign w21252 = ~pi1707 & w21060;
assign w21253 = ~pi1637 & w21062;
assign w21254 = ~w21252 & ~w21253;
assign w21255 = ~w21251 & w21254;
assign w21256 = w21047 & w21255;
assign w21257 = w21035 & ~w21256;
assign w21258 = ~w21247 & w21257;
assign w21259 = ~w21244 & ~w21258;
assign w21260 = w21243 & w21259;
assign w21261 = ~w1639 & ~w21035;
assign w21262 = pi0573 & w21238;
assign w21263 = ~pi0573 & ~w21238;
assign w21264 = ~w21262 & ~w21263;
assign w21265 = ~w21047 & w21264;
assign w21266 = pi0647 & pi1663;
assign w21267 = ~pi0647 & pi1807;
assign w21268 = ~pi0616 & ~w21267;
assign w21269 = ~w21266 & w21268;
assign w21270 = ~pi1818 & w21060;
assign w21271 = ~pi1655 & w21062;
assign w21272 = ~w21270 & ~w21271;
assign w21273 = ~w21269 & w21272;
assign w21274 = w21047 & ~w21273;
assign w21275 = w21035 & ~w21274;
assign w21276 = ~w21265 & w21275;
assign w21277 = ~w21261 & ~w21276;
assign w21278 = w4141 & ~w21035;
assign w21279 = pi0590 & ~w21082;
assign w21280 = ~w21083 & ~w21279;
assign w21281 = ~w21047 & w21280;
assign w21282 = pi0647 & pi1635;
assign w21283 = ~pi0647 & pi1712;
assign w21284 = ~pi0616 & ~w21283;
assign w21285 = ~w21282 & w21284;
assign w21286 = ~pi1812 & w21060;
assign w21287 = ~pi1650 & w21062;
assign w21288 = ~w21286 & ~w21287;
assign w21289 = ~w21285 & w21288;
assign w21290 = w21047 & w21289;
assign w21291 = w21035 & ~w21290;
assign w21292 = ~w21281 & w21291;
assign w21293 = ~w21278 & ~w21292;
assign w21294 = ~w21277 & w21293;
assign w21295 = w21260 & w21294;
assign w21296 = w21226 & w21295;
assign w21297 = w21176 & w21296;
assign w21298 = ~w21041 & ~w21297;
assign w21299 = ~w18155 & w18164;
assign w21300 = pi0712 & ~w21299;
assign w21301 = ~pi0712 & w40174;
assign w21302 = ~w21300 & ~w21301;
assign w21303 = w18928 & ~w21302;
assign w21304 = pi0483 & ~w18928;
assign w21305 = ~w21303 & ~w21304;
assign w21306 = ~pi0712 & w14325;
assign w21307 = ~w21300 & ~w21306;
assign w21308 = w18928 & ~w21307;
assign w21309 = pi0484 & ~w18928;
assign w21310 = ~w21308 & ~w21309;
assign w21311 = ~pi0712 & w14962;
assign w21312 = ~w21300 & ~w21311;
assign w21313 = w18928 & ~w21312;
assign w21314 = pi0485 & ~w18928;
assign w21315 = ~w21313 & ~w21314;
assign w21316 = w18935 & ~w21302;
assign w21317 = pi0486 & ~w18935;
assign w21318 = ~w21316 & ~w21317;
assign w21319 = w18935 & ~w21307;
assign w21320 = pi0487 & ~w18935;
assign w21321 = ~w21319 & ~w21320;
assign w21322 = w18935 & ~w21312;
assign w21323 = pi0488 & ~w18935;
assign w21324 = ~w21322 & ~w21323;
assign w21325 = w10752 & w16059;
assign w21326 = ~w13916 & w18039;
assign w21327 = ~pi0489 & ~w18039;
assign w21328 = ~w10753 & ~w21327;
assign w21329 = ~w21326 & w21328;
assign w21330 = w15173 & ~w21329;
assign w21331 = ~w21325 & ~w21330;
assign w21332 = w13923 & w16059;
assign w21333 = ~w13916 & w18046;
assign w21334 = ~pi0490 & ~w18046;
assign w21335 = ~w13925 & ~w21334;
assign w21336 = ~w21333 & w21335;
assign w21337 = w14336 & ~w21336;
assign w21338 = ~w21332 & ~w21337;
assign w21339 = pi0604 & ~pi3377;
assign w21340 = pi0491 & ~w21339;
assign w21341 = ~pi0491 & ~pi3377;
assign w21342 = pi1771 & w21341;
assign w21343 = ~w21340 & ~w21342;
assign w21344 = pi0654 & pi2765;
assign w21345 = ~pi0729 & w21344;
assign w21346 = pi0498 & pi0504;
assign w21347 = pi0497 & w21346;
assign w21348 = pi0493 & w21347;
assign w21349 = pi0492 & w21348;
assign w21350 = pi0547 & pi0548;
assign w21351 = pi0549 & pi0550;
assign w21352 = pi0551 & w21351;
assign w21353 = w21350 & w21352;
assign w21354 = pi0552 & pi0553;
assign w21355 = pi0563 & w21354;
assign w21356 = w21353 & w21355;
assign w21357 = w21349 & w21356;
assign w21358 = w21345 & ~w21357;
assign w21359 = ~pi0654 & ~pi2765;
assign w21360 = pi0729 & ~w21344;
assign w21361 = ~w21359 & w21360;
assign w21362 = ~w20930 & w21361;
assign w21363 = ~w21358 & ~w21362;
assign w21364 = w21345 & w21349;
assign w21365 = ~w21356 & w21364;
assign w21366 = ~w21363 & ~w21365;
assign w21367 = ~pi0893 & ~w21366;
assign w21368 = ~pi0492 & ~w21348;
assign w21369 = ~w21349 & ~w21368;
assign w21370 = ~w21363 & w21369;
assign w21371 = pi1697 & ~w21370;
assign w21372 = ~w21367 & w21371;
assign w21373 = ~pi0493 & ~w21347;
assign w21374 = ~w21348 & ~w21373;
assign w21375 = w21366 & ~w21374;
assign w21376 = pi0884 & ~w21366;
assign w21377 = pi1697 & ~w21376;
assign w21378 = ~w21375 & w21377;
assign w21379 = pi0494 & ~w18928;
assign w21380 = pi0712 & ~w18159;
assign w21381 = ~pi0712 & w40168;
assign w21382 = ~w21380 & ~w21381;
assign w21383 = w18928 & ~w21382;
assign w21384 = ~w21379 & ~w21383;
assign w21385 = pi0495 & ~w18935;
assign w21386 = w18935 & ~w21382;
assign w21387 = ~w21385 & ~w21386;
assign w21388 = ~pi2398 & w18313;
assign w21389 = pi0496 & ~w18334;
assign w21390 = ~w18335 & ~w18359;
assign w21391 = ~w21389 & w21390;
assign w21392 = ~pi1706 & w18359;
assign w21393 = ~w18313 & ~w21392;
assign w21394 = ~w21391 & w21393;
assign w21395 = ~w21388 & ~w21394;
assign w21396 = ~pi0497 & ~w21346;
assign w21397 = ~w21347 & ~w21396;
assign w21398 = w21366 & ~w21397;
assign w21399 = pi0885 & ~w21366;
assign w21400 = pi1697 & ~w21399;
assign w21401 = ~w21398 & w21400;
assign w21402 = pi0498 & w21366;
assign w21403 = pi0741 & ~w21366;
assign w21404 = pi1697 & ~w21403;
assign w21405 = ~w21402 & w21404;
assign w21406 = pi0959 & pi1746;
assign w21407 = pi0960 & pi3666;
assign w21408 = ~pi0960 & ~pi3666;
assign w21409 = ~pi0959 & ~w21408;
assign w21410 = ~w21407 & w21409;
assign w21411 = ~w21406 & ~w21410;
assign w21412 = pi0941 & ~w305;
assign w21413 = ~pi0941 & pi3668;
assign w21414 = ~w21412 & ~w21413;
assign w21415 = ~pi0954 & w21414;
assign w21416 = pi0954 & ~w21414;
assign w21417 = ~w21415 & ~w21416;
assign w21418 = pi3251 & pi3635;
assign w21419 = w21417 & w21418;
assign w21420 = ~pi0961 & ~w21419;
assign w21421 = pi0961 & ~pi3549;
assign w21422 = ~pi0899 & ~w21421;
assign w21423 = ~w21420 & w21422;
assign w21424 = ~pi0961 & pi2399;
assign w21425 = pi0961 & ~pi3480;
assign w21426 = pi0899 & ~w21425;
assign w21427 = ~w21424 & w21426;
assign w21428 = ~pi0655 & ~w21427;
assign w21429 = ~w21423 & w21428;
assign w21430 = ~pi0655 & ~pi2521;
assign w21431 = pi0655 & pi2521;
assign w21432 = pi0700 & ~w21431;
assign w21433 = ~w21430 & w21432;
assign w21434 = ~w21429 & w21433;
assign w21435 = pi0557 & pi0558;
assign w21436 = pi0560 & w21435;
assign w21437 = pi0499 & pi0500;
assign w21438 = pi0555 & pi0556;
assign w21439 = w21437 & w21438;
assign w21440 = w21436 & w21439;
assign w21441 = pi0502 & pi0503;
assign w21442 = pi0501 & w21441;
assign w21443 = pi0559 & pi0561;
assign w21444 = pi0564 & w21443;
assign w21445 = w21442 & w21444;
assign w21446 = w21440 & w21445;
assign w21447 = ~pi0700 & w21431;
assign w21448 = ~w21446 & w21447;
assign w21449 = ~w21434 & ~w21448;
assign w21450 = w21437 & w21442;
assign w21451 = w21448 & w21450;
assign w21452 = ~w21449 & ~w21451;
assign w21453 = ~pi0799 & ~w21452;
assign w21454 = pi0500 & w21442;
assign w21455 = ~pi0499 & ~w21454;
assign w21456 = ~w21450 & ~w21455;
assign w21457 = ~w21449 & w21456;
assign w21458 = pi1696 & ~w21457;
assign w21459 = ~w21453 & w21458;
assign w21460 = ~pi0500 & ~w21442;
assign w21461 = ~w21454 & ~w21460;
assign w21462 = w21452 & ~w21461;
assign w21463 = pi0957 & ~w21452;
assign w21464 = pi1696 & ~w21463;
assign w21465 = ~w21462 & w21464;
assign w21466 = ~pi0501 & ~w21441;
assign w21467 = ~w21442 & ~w21466;
assign w21468 = w21452 & ~w21467;
assign w21469 = pi1009 & ~w21452;
assign w21470 = pi1696 & ~w21469;
assign w21471 = ~w21468 & w21470;
assign w21472 = ~pi0502 & ~pi0503;
assign w21473 = ~w21441 & ~w21472;
assign w21474 = w21452 & ~w21473;
assign w21475 = pi0793 & ~w21452;
assign w21476 = pi1696 & ~w21475;
assign w21477 = ~w21474 & w21476;
assign w21478 = pi0503 & w21452;
assign w21479 = pi0795 & ~w21452;
assign w21480 = pi1696 & ~w21479;
assign w21481 = ~w21478 & w21480;
assign w21482 = ~pi0498 & ~pi0504;
assign w21483 = ~w21346 & ~w21482;
assign w21484 = w21366 & ~w21483;
assign w21485 = pi0739 & ~w21366;
assign w21486 = pi1697 & ~w21485;
assign w21487 = ~w21484 & w21486;
assign w21488 = ~w363 & w926;
assign w21489 = ~w343 & ~w2239;
assign w21490 = pi0421 & w379;
assign w21491 = ~pi0405 & w21490;
assign w21492 = w6971 & w21491;
assign w21493 = pi0408 & w21492;
assign w21494 = w2377 & ~w21493;
assign w21495 = ~w343 & ~w21494;
assign w21496 = ~w21489 & ~w21495;
assign w21497 = w21488 & w21496;
assign w21498 = ~pi0505 & w21497;
assign w21499 = pi1734 & w822;
assign w21500 = pi1438 & w830;
assign w21501 = w926 & ~w21500;
assign w21502 = pi1729 & w828;
assign w21503 = pi1443 & w825;
assign w21504 = ~w21502 & ~w21503;
assign w21505 = w21501 & w21504;
assign w21506 = ~w21499 & w21505;
assign w21507 = pi0427 & ~w375;
assign w21508 = ~pi0408 & w375;
assign w21509 = ~w21507 & ~w21508;
assign w21510 = ~w354 & w21509;
assign w21511 = w21506 & ~w21510;
assign w21512 = pi3244 & ~w926;
assign w21513 = ~w21511 & ~w21512;
assign w21514 = pi1733 & w822;
assign w21515 = pi1437 & w830;
assign w21516 = w926 & ~w21515;
assign w21517 = pi1728 & w828;
assign w21518 = pi1442 & w825;
assign w21519 = ~w21517 & ~w21518;
assign w21520 = w21516 & w21519;
assign w21521 = ~w21514 & w21520;
assign w21522 = ~pi0413 & w375;
assign w21523 = pi0407 & ~w375;
assign w21524 = ~w21522 & ~w21523;
assign w21525 = ~w354 & w21524;
assign w21526 = w21521 & ~w21525;
assign w21527 = pi3292 & ~w926;
assign w21528 = ~w21526 & ~w21527;
assign w21529 = w21513 & ~w21528;
assign w21530 = ~pi1011 & w6668;
assign w21531 = w21529 & ~w21530;
assign w21532 = ~w21513 & w21528;
assign w21533 = ~pi0983 & w6668;
assign w21534 = w21532 & ~w21533;
assign w21535 = ~w21531 & ~w21534;
assign w21536 = ~pi1050 & w6668;
assign w21537 = w21513 & w21528;
assign w21538 = ~w21536 & w21537;
assign w21539 = ~pi0984 & w6668;
assign w21540 = ~w21513 & ~w21528;
assign w21541 = ~w21539 & w21540;
assign w21542 = ~w21538 & ~w21541;
assign w21543 = w21535 & w21542;
assign w21544 = w40134 & w21543;
assign w21545 = pi2232 & w21531;
assign w21546 = pi2218 & w21534;
assign w21547 = ~w21545 & ~w21546;
assign w21548 = pi2204 & w21538;
assign w21549 = pi2246 & w21541;
assign w21550 = ~w21548 & ~w21549;
assign w21551 = w21547 & w21550;
assign w21552 = ~w21497 & w21551;
assign w21553 = ~w21544 & w21552;
assign w21554 = ~w21498 & ~w21553;
assign w21555 = ~pi0506 & w21497;
assign w21556 = w6413 & w21543;
assign w21557 = pi2247 & w21541;
assign w21558 = pi2219 & w21534;
assign w21559 = ~w21557 & ~w21558;
assign w21560 = pi2233 & ~w21530;
assign w21561 = w21529 & w21560;
assign w21562 = pi2205 & w21538;
assign w21563 = ~w21561 & ~w21562;
assign w21564 = w21559 & w21563;
assign w21565 = ~w21497 & w21564;
assign w21566 = ~w21556 & w21565;
assign w21567 = ~w21555 & ~w21566;
assign w21568 = ~pi0507 & w21497;
assign w21569 = w4380 & w21543;
assign w21570 = pi2248 & w21541;
assign w21571 = pi2220 & w21534;
assign w21572 = ~w21570 & ~w21571;
assign w21573 = pi2234 & ~w21530;
assign w21574 = w21529 & w21573;
assign w21575 = pi2206 & w21538;
assign w21576 = ~w21574 & ~w21575;
assign w21577 = w21572 & w21576;
assign w21578 = ~w21497 & w21577;
assign w21579 = ~w21569 & w21578;
assign w21580 = ~w21568 & ~w21579;
assign w21581 = ~pi0508 & w21497;
assign w21582 = w5320 & w21543;
assign w21583 = pi2221 & w21534;
assign w21584 = pi2235 & w21531;
assign w21585 = ~w21583 & ~w21584;
assign w21586 = pi2207 & w21538;
assign w21587 = pi2249 & w21541;
assign w21588 = ~w21586 & ~w21587;
assign w21589 = w21585 & w21588;
assign w21590 = ~w21497 & w21589;
assign w21591 = ~w21582 & w21590;
assign w21592 = ~w21581 & ~w21591;
assign w21593 = ~pi0509 & w21497;
assign w21594 = w5914 & w21543;
assign w21595 = pi2222 & w21534;
assign w21596 = pi2208 & w21538;
assign w21597 = ~w21595 & ~w21596;
assign w21598 = pi2236 & ~w21530;
assign w21599 = w21529 & w21598;
assign w21600 = pi2250 & w21541;
assign w21601 = ~w21599 & ~w21600;
assign w21602 = w21597 & w21601;
assign w21603 = ~w21497 & w21602;
assign w21604 = ~w21594 & w21603;
assign w21605 = ~w21593 & ~w21604;
assign w21606 = ~pi0510 & w21497;
assign w21607 = w4749 & w21543;
assign w21608 = pi2237 & w21531;
assign w21609 = pi2223 & w21534;
assign w21610 = ~w21608 & ~w21609;
assign w21611 = pi2251 & w21541;
assign w21612 = pi2209 & w21538;
assign w21613 = ~w21611 & ~w21612;
assign w21614 = w21610 & w21613;
assign w21615 = ~w21497 & w21614;
assign w21616 = ~w21607 & w21615;
assign w21617 = ~w21606 & ~w21616;
assign w21618 = ~pi0408 & w21492;
assign w21619 = w2358 & ~w21618;
assign w21620 = ~w343 & ~w21619;
assign w21621 = w21488 & ~w21620;
assign w21622 = ~pi0511 & w21621;
assign w21623 = ~pi0427 & ~w354;
assign w21624 = w21506 & ~w21623;
assign w21625 = pi3394 & ~w926;
assign w21626 = ~w21624 & ~w21625;
assign w21627 = ~pi0407 & ~w354;
assign w21628 = w21521 & ~w21627;
assign w21629 = pi3330 & ~w926;
assign w21630 = ~w21628 & ~w21629;
assign w21631 = ~w21626 & ~w21630;
assign w21632 = ~pi0945 & w6668;
assign w21633 = w21631 & ~w21632;
assign w21634 = ~pi0986 & w6668;
assign w21635 = w21626 & w21630;
assign w21636 = ~w21634 & w21635;
assign w21637 = ~w21633 & ~w21636;
assign w21638 = ~pi0985 & w6668;
assign w21639 = ~w21626 & w21630;
assign w21640 = ~w21638 & w21639;
assign w21641 = w21626 & ~w21630;
assign w21642 = ~pi0760 & w6668;
assign w21643 = w21641 & ~w21642;
assign w21644 = ~w21640 & ~w21643;
assign w21645 = w21637 & w21644;
assign w21646 = w4141 & w21645;
assign w21647 = pi2314 & w21633;
assign w21648 = pi2279 & w21636;
assign w21649 = ~w21647 & ~w21648;
assign w21650 = pi2303 & ~w21642;
assign w21651 = w21641 & w21650;
assign w21652 = pi2292 & w21640;
assign w21653 = ~w21651 & ~w21652;
assign w21654 = w21649 & w21653;
assign w21655 = ~w21621 & w21654;
assign w21656 = ~w21646 & w21655;
assign w21657 = ~w21622 & ~w21656;
assign w21658 = ~pi0512 & w21621;
assign w21659 = w6177 & w21645;
assign w21660 = pi2315 & w21633;
assign w21661 = pi2089 & w21643;
assign w21662 = ~w21660 & ~w21661;
assign w21663 = pi2280 & w21636;
assign w21664 = pi2067 & w21640;
assign w21665 = ~w21663 & ~w21664;
assign w21666 = w21662 & w21665;
assign w21667 = ~w21621 & w21666;
assign w21668 = ~w21659 & w21667;
assign w21669 = ~w21658 & ~w21668;
assign w21670 = ~pi0513 & w21621;
assign w21671 = w40134 & w21645;
assign w21672 = pi2294 & w21640;
assign w21673 = pi2305 & w21643;
assign w21674 = ~w21672 & ~w21673;
assign w21675 = pi2317 & w21633;
assign w21676 = pi2282 & w21636;
assign w21677 = ~w21675 & ~w21676;
assign w21678 = w21674 & w21677;
assign w21679 = ~w21621 & w21678;
assign w21680 = ~w21671 & w21679;
assign w21681 = ~w21670 & ~w21680;
assign w21682 = ~pi0514 & w21621;
assign w21683 = w6413 & w21645;
assign w21684 = pi2084 & w21643;
assign w21685 = pi2318 & w21633;
assign w21686 = ~w21684 & ~w21685;
assign w21687 = pi2283 & w21636;
assign w21688 = pi2295 & w21640;
assign w21689 = ~w21687 & ~w21688;
assign w21690 = w21686 & w21689;
assign w21691 = ~w21621 & w21690;
assign w21692 = ~w21683 & w21691;
assign w21693 = ~w21682 & ~w21692;
assign w21694 = ~pi0515 & w21621;
assign w21695 = w4380 & w21645;
assign w21696 = pi2296 & w21640;
assign w21697 = pi2087 & w21643;
assign w21698 = ~w21696 & ~w21697;
assign w21699 = pi2319 & w21633;
assign w21700 = pi2284 & w21636;
assign w21701 = ~w21699 & ~w21700;
assign w21702 = w21698 & w21701;
assign w21703 = ~w21621 & w21702;
assign w21704 = ~w21695 & w21703;
assign w21705 = ~w21694 & ~w21704;
assign w21706 = ~pi0516 & w21621;
assign w21707 = w5914 & w21645;
assign w21708 = pi2307 & w21643;
assign w21709 = pi2286 & w21636;
assign w21710 = ~w21708 & ~w21709;
assign w21711 = pi2321 & ~w21632;
assign w21712 = w21631 & w21711;
assign w21713 = pi2298 & w21640;
assign w21714 = ~w21712 & ~w21713;
assign w21715 = w21710 & w21714;
assign w21716 = ~w21621 & w21715;
assign w21717 = ~w21707 & w21716;
assign w21718 = ~w21706 & ~w21717;
assign w21719 = ~pi0517 & w21621;
assign w21720 = w4749 & w21645;
assign w21721 = pi2322 & w21633;
assign w21722 = pi2068 & w21636;
assign w21723 = ~w21721 & ~w21722;
assign w21724 = pi2308 & ~w21642;
assign w21725 = w21641 & w21724;
assign w21726 = pi2299 & w21640;
assign w21727 = ~w21725 & ~w21726;
assign w21728 = w21723 & w21727;
assign w21729 = ~w21621 & w21728;
assign w21730 = ~w21720 & w21729;
assign w21731 = ~w21719 & ~w21730;
assign w21732 = ~pi0518 & w21621;
assign w21733 = w1639 & w21645;
assign w21734 = pi2323 & w21633;
assign w21735 = pi2287 & w21636;
assign w21736 = ~w21734 & ~w21735;
assign w21737 = pi2309 & ~w21642;
assign w21738 = w21641 & w21737;
assign w21739 = pi2300 & w21640;
assign w21740 = ~w21738 & ~w21739;
assign w21741 = w21736 & w21740;
assign w21742 = ~w21621 & w21741;
assign w21743 = ~w21733 & w21742;
assign w21744 = ~w21732 & ~w21743;
assign w21745 = ~pi0519 & w21621;
assign w21746 = w5635 & w21645;
assign w21747 = pi2325 & w21633;
assign w21748 = pi2311 & w21643;
assign w21749 = ~w21747 & ~w21748;
assign w21750 = pi2289 & w21636;
assign w21751 = pi2088 & w21640;
assign w21752 = ~w21750 & ~w21751;
assign w21753 = w21749 & w21752;
assign w21754 = ~w21621 & w21753;
assign w21755 = ~w21746 & w21754;
assign w21756 = ~w21745 & ~w21755;
assign w21757 = ~pi0520 & w21621;
assign w21758 = w5053 & w21645;
assign w21759 = pi2326 & w21633;
assign w21760 = pi2312 & w21643;
assign w21761 = ~w21759 & ~w21760;
assign w21762 = pi2290 & w21636;
assign w21763 = pi2301 & w21640;
assign w21764 = ~w21762 & ~w21763;
assign w21765 = w21761 & w21764;
assign w21766 = ~w21621 & w21765;
assign w21767 = ~w21758 & w21766;
assign w21768 = ~w21757 & ~w21767;
assign w21769 = ~pi0521 & w21621;
assign w21770 = w3711 & w21645;
assign w21771 = pi2313 & w21643;
assign w21772 = pi2291 & w21636;
assign w21773 = ~w21771 & ~w21772;
assign w21774 = pi2327 & ~w21632;
assign w21775 = w21631 & w21774;
assign w21776 = pi2302 & w21640;
assign w21777 = ~w21775 & ~w21776;
assign w21778 = w21773 & w21777;
assign w21779 = ~w21621 & w21778;
assign w21780 = ~w21770 & w21779;
assign w21781 = ~w21769 & ~w21780;
assign w21782 = pi1597 & ~w6682;
assign w21783 = ~pi1444 & pi3141;
assign w21784 = ~pi3300 & w21783;
assign w21785 = ~pi0875 & pi1444;
assign w21786 = pi0522 & pi3372;
assign w21787 = ~w21785 & w21786;
assign w21788 = ~w21784 & w21787;
assign w21789 = pi3237 & ~w21788;
assign w21790 = ~w21782 & w21789;
assign w21791 = pi0523 & w343;
assign w21792 = ~w343 & ~w2238;
assign w21793 = pi0418 & w2901;
assign w21794 = ~pi0420 & w21793;
assign w21795 = w376 & w21491;
assign w21796 = ~pi0410 & w21795;
assign w21797 = ~w21794 & ~w21796;
assign w21798 = pi0420 & w21491;
assign w21799 = ~pi0409 & w21798;
assign w21800 = pi0419 & ~w21799;
assign w21801 = ~w21797 & w21800;
assign w21802 = pi0405 & pi0422;
assign w21803 = w2374 & w21802;
assign w21804 = pi0419 & w2355;
assign w21805 = ~w21793 & ~w21804;
assign w21806 = ~w21803 & w21805;
assign w21807 = pi0422 & w2235;
assign w21808 = w2241 & w2242;
assign w21809 = ~w21807 & ~w21808;
assign w21810 = w376 & w21490;
assign w21811 = pi0418 & w14357;
assign w21812 = ~w21810 & ~w21811;
assign w21813 = w21809 & w21812;
assign w21814 = w21806 & w21813;
assign w21815 = pi0410 & w21795;
assign w21816 = ~w2231 & w2901;
assign w21817 = ~w21815 & ~w21816;
assign w21818 = ~w21814 & w21817;
assign w21819 = ~w21801 & w21818;
assign w21820 = w2231 & w21491;
assign w21821 = ~pi0422 & w21820;
assign w21822 = w21812 & ~w21821;
assign w21823 = ~w2901 & w21822;
assign w21824 = pi0414 & ~w21823;
assign w21825 = pi0411 & w21823;
assign w21826 = ~w21824 & ~w21825;
assign w21827 = w21819 & ~w21826;
assign w21828 = pi0427 & ~w21823;
assign w21829 = ~pi0408 & w21823;
assign w21830 = ~w21828 & ~w21829;
assign w21831 = w21827 & w21830;
assign w21832 = ~w10712 & ~w21823;
assign w21833 = ~pi0412 & pi0413;
assign w21834 = w21823 & ~w21833;
assign w21835 = ~w21832 & ~w21834;
assign w21836 = w21831 & w21835;
assign w21837 = ~pi0413 & w21823;
assign w21838 = pi0412 & w21837;
assign w21839 = pi0407 & ~w21823;
assign w21840 = pi0415 & w21839;
assign w21841 = ~w21838 & ~w21840;
assign w21842 = w21827 & ~w21841;
assign w21843 = w21819 & w21826;
assign w21844 = ~w21837 & ~w21839;
assign w21845 = w21843 & w21844;
assign w21846 = ~w21842 & ~w21845;
assign w21847 = ~w21836 & w21846;
assign w21848 = w21792 & ~w21847;
assign w21849 = ~w21791 & ~w21848;
assign w21850 = pi0524 & w343;
assign w21851 = ~w343 & w2238;
assign w21852 = ~w21847 & w21851;
assign w21853 = ~w21850 & ~w21852;
assign w21854 = pi0525 & w20931;
assign w21855 = ~pi0525 & ~w20931;
assign w21856 = ~w21854 & ~w21855;
assign w21857 = ~w20933 & ~w21856;
assign w21858 = w21366 & w21857;
assign w21859 = ~pi0526 & pi0531;
assign w21860 = pi0531 & ~w20933;
assign w21861 = pi0526 & ~w21860;
assign w21862 = ~w21859 & ~w21861;
assign w21863 = w21366 & w21862;
assign w21864 = ~pi0527 & ~w21854;
assign w21865 = pi0527 & w21854;
assign w21866 = ~pi0554 & w21865;
assign w21867 = ~w21864 & ~w21866;
assign w21868 = w21366 & ~w21867;
assign w21869 = ~pi0528 & pi0529;
assign w21870 = pi0530 & pi0542;
assign w21871 = pi0532 & w21870;
assign w21872 = pi0529 & ~w21871;
assign w21873 = pi0528 & ~w21872;
assign w21874 = ~w21869 & ~w21873;
assign w21875 = w21452 & w21874;
assign w21876 = ~w21869 & ~w21872;
assign w21877 = w21452 & ~w21876;
assign w21878 = pi0528 & pi0529;
assign w21879 = pi0532 & w21878;
assign w21880 = ~w21870 & w21879;
assign w21881 = pi0530 & w21880;
assign w21882 = ~pi0530 & ~w21879;
assign w21883 = ~w21881 & ~w21882;
assign w21884 = w21452 & ~w21883;
assign w21885 = ~w21859 & ~w21860;
assign w21886 = w21366 & ~w21885;
assign w21887 = ~pi0532 & ~w21878;
assign w21888 = ~w21880 & ~w21887;
assign w21889 = w21452 & ~w21888;
assign w21890 = ~pi0533 & w21497;
assign w21891 = w4141 & w21543;
assign w21892 = pi2229 & w21531;
assign w21893 = pi2201 & w21538;
assign w21894 = ~w21892 & ~w21893;
assign w21895 = pi2215 & ~w21533;
assign w21896 = w21532 & w21895;
assign w21897 = pi2243 & w21541;
assign w21898 = ~w21896 & ~w21897;
assign w21899 = w21894 & w21898;
assign w21900 = ~w21497 & w21899;
assign w21901 = ~w21891 & w21900;
assign w21902 = ~w21890 & ~w21901;
assign w21903 = ~pi0534 & w21497;
assign w21904 = w1308 & w21543;
assign w21905 = pi2239 & w21531;
assign w21906 = pi2225 & w21534;
assign w21907 = ~w21905 & ~w21906;
assign w21908 = pi2211 & w21538;
assign w21909 = pi2253 & w21541;
assign w21910 = ~w21908 & ~w21909;
assign w21911 = w21907 & w21910;
assign w21912 = ~w21497 & w21911;
assign w21913 = ~w21904 & w21912;
assign w21914 = ~w21903 & ~w21913;
assign w21915 = ~pi0535 & w21497;
assign w21916 = w5635 & w21543;
assign w21917 = pi2254 & w21541;
assign w21918 = pi2226 & w21534;
assign w21919 = ~w21917 & ~w21918;
assign w21920 = pi2240 & ~w21530;
assign w21921 = w21529 & w21920;
assign w21922 = pi2212 & w21538;
assign w21923 = ~w21921 & ~w21922;
assign w21924 = w21919 & w21923;
assign w21925 = ~w21497 & w21924;
assign w21926 = ~w21916 & w21925;
assign w21927 = ~w21915 & ~w21926;
assign w21928 = ~pi0536 & w21497;
assign w21929 = w5053 & w21543;
assign w21930 = pi2255 & w21541;
assign w21931 = pi2241 & w21531;
assign w21932 = ~w21930 & ~w21931;
assign w21933 = pi2227 & w21534;
assign w21934 = pi2213 & w21538;
assign w21935 = ~w21933 & ~w21934;
assign w21936 = w21932 & w21935;
assign w21937 = ~w21497 & w21936;
assign w21938 = ~w21929 & w21937;
assign w21939 = ~w21928 & ~w21938;
assign w21940 = pi0537 & w343;
assign w21941 = pi0407 & pi0415;
assign w21942 = w21832 & ~w21941;
assign w21943 = ~pi0412 & ~pi0413;
assign w21944 = pi0412 & pi0413;
assign w21945 = ~w21943 & ~w21944;
assign w21946 = w21823 & ~w21945;
assign w21947 = ~w21942 & ~w21946;
assign w21948 = w21827 & ~w21947;
assign w21949 = pi0420 & w21793;
assign w21950 = ~w21815 & ~w21949;
assign w21951 = w21800 & ~w21950;
assign w21952 = ~pi0407 & pi0427;
assign w21953 = w397 & w21952;
assign w21954 = w21951 & w21953;
assign w21955 = ~w21948 & ~w21954;
assign w21956 = w21792 & ~w21955;
assign w21957 = ~w21940 & ~w21956;
assign w21958 = pi0538 & w343;
assign w21959 = w21851 & ~w21955;
assign w21960 = ~w21958 & ~w21959;
assign w21961 = pi0539 & w343;
assign w21962 = w397 & w10685;
assign w21963 = ~w2343 & ~w21800;
assign w21964 = ~w21962 & ~w21963;
assign w21965 = ~w343 & ~w21950;
assign w21966 = ~w21964 & w21965;
assign w21967 = ~w21961 & ~w21966;
assign w21968 = ~w343 & w6682;
assign w21969 = w2230 & w21968;
assign w21970 = w2343 & w10685;
assign w21971 = w21951 & w21970;
assign w21972 = w21969 & w21971;
assign w21973 = w2241 & w14357;
assign w21974 = ~w21795 & ~w21973;
assign w21975 = ~w6602 & w21974;
assign w21976 = pi0426 & w21795;
assign w21977 = pi0411 & w21976;
assign w21978 = pi0420 & ~w21795;
assign w21979 = pi0414 & w21978;
assign w21980 = ~w21977 & ~w21979;
assign w21981 = ~w21975 & ~w21980;
assign w21982 = ~pi0415 & ~w21795;
assign w21983 = ~pi0412 & w21795;
assign w21984 = ~w21982 & ~w21983;
assign w21985 = ~pi0413 & w21795;
assign w21986 = pi0407 & ~w21795;
assign w21987 = ~w21985 & ~w21986;
assign w21988 = w21984 & w21987;
assign w21989 = w21981 & w21988;
assign w21990 = ~pi0425 & w21798;
assign w21991 = pi0419 & ~w21990;
assign w21992 = pi0427 & ~w21795;
assign w21993 = ~pi0408 & w21795;
assign w21994 = ~w21992 & ~w21993;
assign w21995 = w21991 & ~w21994;
assign w21996 = w21989 & ~w21995;
assign w21997 = ~pi0414 & w21978;
assign w21998 = ~pi0411 & w21976;
assign w21999 = ~w21997 & ~w21998;
assign w22000 = ~w21975 & ~w21999;
assign w22001 = w21987 & ~w21994;
assign w22002 = ~w21984 & w21991;
assign w22003 = ~w22001 & w22002;
assign w22004 = w22000 & w22003;
assign w22005 = pi0419 & w2233;
assign w22006 = pi0405 & w21490;
assign w22007 = ~pi0411 & ~pi0413;
assign w22008 = pi0419 & ~pi0424;
assign w22009 = w22007 & w22008;
assign w22010 = ~pi0420 & ~w22009;
assign w22011 = w22006 & w22010;
assign w22012 = ~w22005 & ~w22011;
assign w22013 = ~w22004 & w22012;
assign w22014 = ~w21996 & w22013;
assign w22015 = w21969 & ~w22014;
assign w22016 = pi0540 & w6684;
assign w22017 = ~w22015 & ~w22016;
assign w22018 = ~w21972 & w22017;
assign w22019 = pi0541 & w6684;
assign w22020 = w6682 & w14887;
assign w22021 = w10751 & ~w14393;
assign w22022 = w14360 & w14369;
assign w22023 = pi0406 & ~pi0425;
assign w22024 = ~w22022 & w22023;
assign w22025 = w15184 & w22024;
assign w22026 = ~w22021 & ~w22025;
assign w22027 = w22020 & ~w22026;
assign w22028 = ~w22019 & ~w22027;
assign w22029 = ~pi0542 & ~w21881;
assign w22030 = w21452 & ~w22029;
assign w22031 = pi2018 & ~w6682;
assign w22032 = pi0877 & pi1447;
assign w22033 = ~pi1447 & pi2820;
assign w22034 = ~w22032 & ~w22033;
assign w22035 = pi0544 & ~pi3373;
assign w22036 = ~w22034 & w22035;
assign w22037 = pi3068 & ~w22036;
assign w22038 = ~w22031 & w22037;
assign w22039 = w13 & ~w111;
assign w22040 = w109 & w22039;
assign w22041 = ~w903 & ~w2891;
assign w22042 = ~w7233 & w22041;
assign w22043 = w22040 & ~w22042;
assign w22044 = pi0787 & ~w22043;
assign w22045 = ~pi0687 & ~pi0723;
assign w22046 = ~pi0724 & ~pi0725;
assign w22047 = ~pi0726 & ~pi0732;
assign w22048 = w22046 & w22047;
assign w22049 = w22045 & w22048;
assign w22050 = ~pi0772 & ~pi0782;
assign w22051 = ~pi0786 & w22050;
assign w22052 = ~pi0733 & ~pi0769;
assign w22053 = ~pi0770 & ~pi0771;
assign w22054 = w22052 & w22053;
assign w22055 = w22051 & w22054;
assign w22056 = w22049 & w22055;
assign w22057 = ~w22044 & w22056;
assign w22058 = pi0787 & w22057;
assign w22059 = w347 & w22058;
assign w22060 = pi3490 & pi3544;
assign w22061 = pi0545 & pi3186;
assign w22062 = ~w22060 & w22061;
assign w22063 = ~w22059 & w22062;
assign w22064 = pi1598 & ~w6682;
assign w22065 = pi2975 & ~w22064;
assign w22066 = ~w22063 & w22065;
assign w22067 = pi1049 & ~w6682;
assign w22068 = pi2976 & ~w22067;
assign w22069 = ~pi1738 & ~pi3302;
assign w22070 = ~pi0879 & pi1738;
assign w22071 = pi3189 & ~w22070;
assign w22072 = ~w22069 & w22071;
assign w22073 = pi1931 & ~w22072;
assign w22074 = pi0546 & ~w22073;
assign w22075 = w22068 & ~w22074;
assign w22076 = pi0553 & w21365;
assign w22077 = pi0552 & w22076;
assign w22078 = pi0551 & w22077;
assign w22079 = pi0563 & w22078;
assign w22080 = pi0550 & w22079;
assign w22081 = pi0549 & w22080;
assign w22082 = pi0548 & w22081;
assign w22083 = ~w21363 & ~w22082;
assign w22084 = ~pi0547 & w22083;
assign w22085 = pi0948 & w21363;
assign w22086 = ~w22084 & ~w22085;
assign w22087 = ~pi0548 & ~w22081;
assign w22088 = w22083 & ~w22087;
assign w22089 = ~pi0949 & w21363;
assign w22090 = ~w22088 & ~w22089;
assign w22091 = ~pi0950 & w21363;
assign w22092 = ~pi0549 & ~w22080;
assign w22093 = ~w22081 & ~w22092;
assign w22094 = ~w21363 & w22093;
assign w22095 = ~w22091 & ~w22094;
assign w22096 = ~pi0951 & w21363;
assign w22097 = ~pi0550 & ~w22079;
assign w22098 = ~w22080 & ~w22097;
assign w22099 = ~w21363 & w22098;
assign w22100 = ~w22096 & ~w22099;
assign w22101 = ~pi0892 & w21363;
assign w22102 = ~pi0551 & ~w22077;
assign w22103 = ~w22078 & ~w22102;
assign w22104 = ~w21363 & w22103;
assign w22105 = ~w22101 & ~w22104;
assign w22106 = ~pi0952 & w21363;
assign w22107 = ~pi0552 & ~w22076;
assign w22108 = ~w22077 & ~w22107;
assign w22109 = ~w21363 & w22108;
assign w22110 = ~w22106 & ~w22109;
assign w22111 = ~pi0953 & w21363;
assign w22112 = ~pi0553 & ~w21364;
assign w22113 = ~w22076 & ~w22112;
assign w22114 = ~w21363 & w22113;
assign w22115 = ~w22111 & ~w22114;
assign w22116 = ~pi0554 & ~w21865;
assign w22117 = w21366 & ~w22116;
assign w22118 = pi0561 & w21451;
assign w22119 = pi0564 & w22118;
assign w22120 = pi0560 & w22119;
assign w22121 = pi0559 & w22120;
assign w22122 = pi0558 & w22121;
assign w22123 = pi0557 & w22122;
assign w22124 = pi0556 & w22123;
assign w22125 = ~w21449 & ~w22124;
assign w22126 = ~pi0555 & w22125;
assign w22127 = pi0963 & w21449;
assign w22128 = ~w22126 & ~w22127;
assign w22129 = ~pi0556 & ~w22123;
assign w22130 = w22125 & ~w22129;
assign w22131 = ~pi0964 & w21449;
assign w22132 = ~w22130 & ~w22131;
assign w22133 = ~pi0965 & w21449;
assign w22134 = ~pi0557 & ~w22122;
assign w22135 = ~w22123 & ~w22134;
assign w22136 = ~w21449 & w22135;
assign w22137 = ~w22133 & ~w22136;
assign w22138 = ~pi0900 & w21449;
assign w22139 = ~pi0558 & ~w22121;
assign w22140 = ~w22122 & ~w22139;
assign w22141 = ~w21449 & w22140;
assign w22142 = ~w22138 & ~w22141;
assign w22143 = ~pi0797 & w21449;
assign w22144 = ~pi0559 & ~w22120;
assign w22145 = ~w22121 & ~w22144;
assign w22146 = ~w21449 & w22145;
assign w22147 = ~w22143 & ~w22146;
assign w22148 = ~pi0798 & w21449;
assign w22149 = ~pi0560 & ~w22119;
assign w22150 = ~w22120 & ~w22149;
assign w22151 = ~w21449 & w22150;
assign w22152 = ~w22148 & ~w22151;
assign w22153 = ~pi0561 & w21452;
assign w22154 = pi0967 & w21449;
assign w22155 = ~w22118 & ~w22154;
assign w22156 = ~w22153 & w22155;
assign w22157 = ~pi0891 & w21363;
assign w22158 = ~pi0563 & ~w22078;
assign w22159 = ~w22079 & ~w22158;
assign w22160 = ~w21363 & w22159;
assign w22161 = ~w22157 & ~w22160;
assign w22162 = ~pi0966 & w21449;
assign w22163 = ~pi0564 & ~w22118;
assign w22164 = ~w22119 & ~w22163;
assign w22165 = ~w21449 & w22164;
assign w22166 = ~w22162 & ~w22165;
assign w22167 = ~pi3479 & ~pi3682;
assign w22168 = ~pi3479 & pi3682;
assign w22169 = ~w343 & w2230;
assign w22170 = ~w2356 & w21806;
assign w22171 = w6606 & w22170;
assign w22172 = pi2978 & ~w22171;
assign w22173 = ~w21821 & ~w22172;
assign w22174 = ~w874 & ~w2377;
assign w22175 = w422 & w22174;
assign w22176 = ~w2383 & ~w22175;
assign w22177 = w2349 & ~w2358;
assign w22178 = ~w2382 & w22177;
assign w22179 = ~w422 & ~w2377;
assign w22180 = ~w2379 & ~w22179;
assign w22181 = ~w22178 & w22180;
assign w22182 = w22176 & ~w22181;
assign w22183 = ~w3465 & w22182;
assign w22184 = ~w22176 & ~w22181;
assign w22185 = ~w3814 & w22184;
assign w22186 = w422 & w2378;
assign w22187 = ~w22177 & ~w22186;
assign w22188 = w22176 & ~w22187;
assign w22189 = ~w1639 & w22188;
assign w22190 = ~w22176 & ~w22187;
assign w22191 = ~w3711 & w22190;
assign w22192 = ~w22178 & ~w22191;
assign w22193 = ~w22189 & w22192;
assign w22194 = ~w22185 & ~w22193;
assign w22195 = ~w22183 & w22194;
assign w22196 = ~w22176 & w22181;
assign w22197 = w3761 & w22196;
assign w22198 = ~w3721 & w22181;
assign w22199 = w22176 & ~w22198;
assign w22200 = ~w22197 & ~w22199;
assign w22201 = ~w1377 & w22179;
assign w22202 = ~w3746 & w22187;
assign w22203 = ~w22201 & w22202;
assign w22204 = ~w22200 & w22203;
assign w22205 = ~w22176 & w22187;
assign w22206 = ~w3761 & w22181;
assign w22207 = w22205 & ~w22206;
assign w22208 = w1369 & w22207;
assign w22209 = ~w22204 & ~w22208;
assign w22210 = ~w22195 & w22209;
assign w22211 = ~w22173 & ~w22210;
assign w22212 = ~w874 & w1369;
assign w22213 = w874 & ~w1639;
assign w22214 = ~w22212 & ~w22213;
assign w22215 = w422 & w22214;
assign w22216 = w1377 & ~w22215;
assign w22217 = ~pi3680 & w883;
assign w22218 = pi2409 & ~w2239;
assign w22219 = ~w22217 & w22218;
assign w22220 = ~w819 & ~w874;
assign w22221 = w874 & w1308;
assign w22222 = ~w22220 & ~w22221;
assign w22223 = w422 & w22218;
assign w22224 = ~w22222 & w22223;
assign w22225 = ~w22219 & ~w22224;
assign w22226 = ~w22216 & ~w22225;
assign w22227 = ~w22211 & ~w22226;
assign w22228 = w22169 & ~w22227;
assign w22229 = ~pi0565 & w343;
assign w22230 = ~pi3682 & ~w343;
assign w22231 = ~w22229 & ~w22230;
assign w22232 = ~w22228 & ~w22231;
assign w22233 = ~pi0566 & w21497;
assign w22234 = w6177 & w21543;
assign w22235 = pi2244 & w21541;
assign w22236 = pi2230 & w21531;
assign w22237 = ~w22235 & ~w22236;
assign w22238 = pi2216 & w21534;
assign w22239 = pi2202 & w21538;
assign w22240 = ~w22238 & ~w22239;
assign w22241 = w22237 & w22240;
assign w22242 = ~w21497 & w22241;
assign w22243 = ~w22234 & w22242;
assign w22244 = ~w22233 & ~w22243;
assign w22245 = ~pi0567 & w21497;
assign w22246 = w3195 & w21543;
assign w22247 = pi2217 & w21534;
assign w22248 = pi2245 & w21541;
assign w22249 = ~w22247 & ~w22248;
assign w22250 = pi2231 & ~w21530;
assign w22251 = w21529 & w22250;
assign w22252 = pi2203 & w21538;
assign w22253 = ~w22251 & ~w22252;
assign w22254 = w22249 & w22253;
assign w22255 = ~w21497 & w22254;
assign w22256 = ~w22246 & w22255;
assign w22257 = ~w22245 & ~w22256;
assign w22258 = ~pi0568 & w21497;
assign w22259 = w1639 & w21543;
assign w22260 = pi2238 & w21531;
assign w22261 = pi2224 & w21534;
assign w22262 = ~w22260 & ~w22261;
assign w22263 = pi2252 & w21541;
assign w22264 = pi2210 & w21538;
assign w22265 = ~w22263 & ~w22264;
assign w22266 = w22262 & w22265;
assign w22267 = ~w21497 & w22266;
assign w22268 = ~w22259 & w22267;
assign w22269 = ~w22258 & ~w22268;
assign w22270 = ~pi0569 & w21497;
assign w22271 = w3711 & w21543;
assign w22272 = pi2256 & w21541;
assign w22273 = pi2228 & w21534;
assign w22274 = ~w22272 & ~w22273;
assign w22275 = pi2242 & ~w21530;
assign w22276 = w21529 & w22275;
assign w22277 = pi2214 & w21538;
assign w22278 = ~w22276 & ~w22277;
assign w22279 = w22274 & w22278;
assign w22280 = ~w21497 & w22279;
assign w22281 = ~w22271 & w22280;
assign w22282 = ~w22270 & ~w22281;
assign w22283 = pi1048 & ~w6682;
assign w22284 = pi3239 & ~w22283;
assign w22285 = ~pi1735 & ~pi3144;
assign w22286 = ~pi3303 & w22285;
assign w22287 = pi0878 & pi1735;
assign w22288 = pi3226 & ~w22287;
assign w22289 = ~w22286 & w22288;
assign w22290 = pi1931 & ~w22289;
assign w22291 = pi0570 & ~w22290;
assign w22292 = w22284 & ~w22291;
assign w22293 = w21040 & ~w21224;
assign w22294 = pi0571 & ~w21040;
assign w22295 = ~w22293 & ~w22294;
assign w22296 = w21040 & ~w21173;
assign w22297 = pi0572 & ~w21040;
assign w22298 = ~w22296 & ~w22297;
assign w22299 = pi0573 & ~w21040;
assign w22300 = w21040 & w21277;
assign w22301 = ~w22299 & ~w22300;
assign w22302 = pi0574 & w343;
assign w22303 = w21827 & ~w21830;
assign w22304 = w21835 & w22303;
assign w22305 = w21843 & ~w21844;
assign w22306 = w2332 & w10653;
assign w22307 = w21951 & w22306;
assign w22308 = ~w22305 & ~w22307;
assign w22309 = ~w22304 & w22308;
assign w22310 = w21792 & ~w22309;
assign w22311 = ~w22302 & ~w22310;
assign w22312 = ~pi0426 & ~w21991;
assign w22313 = ~w21974 & ~w22312;
assign w22314 = w2244 & w6605;
assign w22315 = w21822 & w22314;
assign w22316 = ~w21816 & ~w22315;
assign w22317 = ~w22313 & w22316;
assign w22318 = ~w2236 & ~w14370;
assign w22319 = ~w378 & ~w22318;
assign w22320 = ~w21821 & ~w22319;
assign w22321 = pi0427 & ~w22320;
assign w22322 = ~pi0408 & w22320;
assign w22323 = ~w22321 & ~w22322;
assign w22324 = w22317 & ~w22323;
assign w22325 = pi0414 & ~w22320;
assign w22326 = pi0411 & w22320;
assign w22327 = ~w22325 & ~w22326;
assign w22328 = w21968 & w22327;
assign w22329 = w22324 & w22328;
assign w22330 = pi0407 & w21982;
assign w22331 = ~w22320 & w22330;
assign w22332 = w21943 & w22320;
assign w22333 = ~w22331 & ~w22332;
assign w22334 = w22329 & ~w22333;
assign w22335 = ~pi0575 & w6684;
assign w22336 = w375 & w21968;
assign w22337 = w2231 & w22336;
assign w22338 = ~w22335 & ~w22337;
assign w22339 = ~w22334 & w22338;
assign w22340 = pi0576 & w343;
assign w22341 = w21851 & ~w22309;
assign w22342 = ~w22340 & ~w22341;
assign w22343 = ~pi2092 & w18313;
assign w22344 = pi0577 & ~w18333;
assign w22345 = ~w18334 & ~w18359;
assign w22346 = ~w22344 & w22345;
assign w22347 = ~pi1716 & w18359;
assign w22348 = ~w18313 & ~w22347;
assign w22349 = ~w22346 & w22348;
assign w22350 = ~w22343 & ~w22349;
assign w22351 = w21040 & ~w21069;
assign w22352 = pi0578 & ~w21040;
assign w22353 = ~w22351 & ~w22352;
assign w22354 = w10712 & ~w22320;
assign w22355 = w21833 & w22320;
assign w22356 = ~w22354 & ~w22355;
assign w22357 = w22329 & ~w22356;
assign w22358 = ~pi0579 & w6684;
assign w22359 = w6971 & w22336;
assign w22360 = ~w22358 & ~w22359;
assign w22361 = ~w22357 & w22360;
assign w22362 = ~pi0407 & pi0415;
assign w22363 = ~w22320 & w22362;
assign w22364 = w21944 & w22320;
assign w22365 = ~w22363 & ~w22364;
assign w22366 = w22329 & ~w22365;
assign w22367 = ~pi0580 & w6684;
assign w22368 = ~pi0418 & w22336;
assign w22369 = ~w22367 & ~w22368;
assign w22370 = ~w22366 & w22369;
assign w22371 = w10752 & ~w16064;
assign w22372 = ~w40159 & w18039;
assign w22373 = ~pi0583 & ~w18039;
assign w22374 = ~w10753 & ~w22373;
assign w22375 = ~w22372 & w22374;
assign w22376 = w15173 & ~w22375;
assign w22377 = ~w22371 & ~w22376;
assign w22378 = w13923 & ~w16064;
assign w22379 = ~w40159 & w18046;
assign w22380 = ~pi0584 & ~w18046;
assign w22381 = ~w13925 & ~w22380;
assign w22382 = ~w22379 & w22381;
assign w22383 = w14336 & ~w22382;
assign w22384 = ~w22378 & ~w22383;
assign w22385 = pi0585 & ~w21040;
assign w22386 = ~w21124 & ~w22385;
assign w22387 = ~pi0835 & w3195;
assign w22388 = w13945 & w18925;
assign w22389 = w10689 & ~w22388;
assign w22390 = ~w14424 & w18073;
assign w22391 = w14424 & ~w18073;
assign w22392 = w18925 & ~w22391;
assign w22393 = ~w22390 & w22392;
assign w22394 = w10614 & w22393;
assign w22395 = ~pi1402 & w10564;
assign w22396 = ~pi1513 & w10559;
assign w22397 = ~pi1495 & w10566;
assign w22398 = ~w22396 & ~w22397;
assign w22399 = ~w22395 & w22398;
assign w22400 = ~pi1041 & ~w22399;
assign w22401 = pi1410 & w10564;
assign w22402 = pi1041 & ~w22401;
assign w22403 = pi1614 & w10559;
assign w22404 = pi1532 & w10561;
assign w22405 = pi1566 & w10566;
assign w22406 = ~w22404 & ~w22405;
assign w22407 = ~w22403 & w22406;
assign w22408 = w22402 & w22407;
assign w22409 = ~w22400 & ~w22408;
assign w22410 = w10627 & ~w22409;
assign w22411 = ~w22394 & ~w22410;
assign w22412 = ~w22389 & w22411;
assign w22413 = ~w22387 & w22412;
assign w22414 = ~pi0586 & w22389;
assign w22415 = w17481 & ~w22414;
assign w22416 = ~w22413 & w22415;
assign w22417 = ~pi0587 & w21621;
assign w22418 = w3195 & w21645;
assign w22419 = pi2316 & w21633;
assign w22420 = pi2304 & w21643;
assign w22421 = ~w22419 & ~w22420;
assign w22422 = pi2293 & w21640;
assign w22423 = pi2281 & w21636;
assign w22424 = ~w22422 & ~w22423;
assign w22425 = w22421 & w22424;
assign w22426 = ~w21621 & w22425;
assign w22427 = ~w22418 & w22426;
assign w22428 = ~w22417 & ~w22427;
assign w22429 = ~pi0588 & w21621;
assign w22430 = w5320 & w21645;
assign w22431 = pi2306 & w21643;
assign w22432 = pi2320 & w21633;
assign w22433 = ~w22431 & ~w22432;
assign w22434 = pi2297 & w21640;
assign w22435 = pi2285 & w21636;
assign w22436 = ~w22434 & ~w22435;
assign w22437 = w22433 & w22436;
assign w22438 = ~w21621 & w22437;
assign w22439 = ~w22430 & w22438;
assign w22440 = ~w22429 & ~w22439;
assign w22441 = ~pi0589 & w21621;
assign w22442 = w1308 & w21645;
assign w22443 = pi2122 & w21640;
assign w22444 = pi2324 & ~w21632;
assign w22445 = w21631 & w22444;
assign w22446 = ~w22443 & ~w22445;
assign w22447 = pi2310 & ~w21642;
assign w22448 = w21641 & w22447;
assign w22449 = pi2288 & w21636;
assign w22450 = ~w22448 & ~w22449;
assign w22451 = w22446 & w22450;
assign w22452 = ~w21621 & w22451;
assign w22453 = ~w22442 & w22452;
assign w22454 = ~w22441 & ~w22453;
assign w22455 = w21040 & ~w21293;
assign w22456 = pi0590 & ~w21040;
assign w22457 = ~w22455 & ~w22456;
assign w22458 = w21040 & ~w21208;
assign w22459 = pi0591 & ~w21040;
assign w22460 = ~w22458 & ~w22459;
assign w22461 = w21040 & ~w21157;
assign w22462 = pi0592 & ~w21040;
assign w22463 = ~w22461 & ~w22462;
assign w22464 = w21040 & ~w21243;
assign w22465 = pi0593 & ~w21040;
assign w22466 = ~w22464 & ~w22465;
assign w22467 = w21040 & ~w21107;
assign w22468 = pi0594 & ~w21040;
assign w22469 = ~w22467 & ~w22468;
assign w22470 = w21040 & ~w21091;
assign w22471 = pi0595 & ~w21040;
assign w22472 = ~w22470 & ~w22471;
assign w22473 = w22317 & w22323;
assign w22474 = w22328 & w22473;
assign w22475 = ~w22365 & w22474;
assign w22476 = ~pi0596 & w6684;
assign w22477 = pi0418 & w22336;
assign w22478 = ~w22476 & ~w22477;
assign w22479 = ~w22475 & w22478;
assign w22480 = ~w22356 & w22474;
assign w22481 = ~pi0597 & w6684;
assign w22482 = w376 & w22336;
assign w22483 = ~w22481 & ~w22482;
assign w22484 = ~w22480 & w22483;
assign w22485 = ~pi0598 & w6684;
assign w22486 = w21941 & ~w22320;
assign w22487 = pi0412 & ~pi0413;
assign w22488 = w22320 & w22487;
assign w22489 = ~w22486 & ~w22488;
assign w22490 = w22474 & ~w22489;
assign w22491 = ~w22485 & ~w22490;
assign w22492 = ~pi0599 & w6684;
assign w22493 = w22329 & ~w22489;
assign w22494 = ~w22492 & ~w22493;
assign w22495 = pi3575 & pi3647;
assign w22496 = pi0895 & w22495;
assign w22497 = ~pi0931 & pi3647;
assign w22498 = ~pi1067 & w22497;
assign w22499 = ~pi1069 & ~pi1088;
assign w22500 = w22498 & w22499;
assign w22501 = ~pi1068 & w22500;
assign w22502 = ~pi1083 & w22501;
assign w22503 = ~pi0932 & w22502;
assign w22504 = ~pi0940 & w22503;
assign w22505 = ~pi0847 & w22504;
assign w22506 = ~pi1085 & w22505;
assign w22507 = ~pi0689 & w22506;
assign w22508 = ~pi0651 & w22507;
assign w22509 = ~pi0727 & w22508;
assign w22510 = ~pi1087 & w22509;
assign w22511 = ~pi0617 & w22510;
assign w22512 = ~pi0600 & w22511;
assign w22513 = pi0600 & ~w22511;
assign w22514 = ~pi0738 & ~pi0790;
assign w22515 = pi0737 & pi1088;
assign w22516 = pi0651 & pi0872;
assign w22517 = ~w22515 & ~w22516;
assign w22518 = pi0743 & pi0932;
assign w22519 = ~pi0743 & ~pi0932;
assign w22520 = ~w22518 & ~w22519;
assign w22521 = w22517 & w22520;
assign w22522 = ~pi0689 & ~pi0871;
assign w22523 = ~pi0744 & ~pi1083;
assign w22524 = ~w22522 & ~w22523;
assign w22525 = ~pi0742 & ~pi0940;
assign w22526 = pi0870 & pi1087;
assign w22527 = ~w22525 & ~w22526;
assign w22528 = w22524 & w22527;
assign w22529 = w22521 & w22528;
assign w22530 = pi0689 & pi0871;
assign w22531 = ~pi0747 & ~pi1067;
assign w22532 = ~w22530 & ~w22531;
assign w22533 = ~pi0651 & ~pi0872;
assign w22534 = pi0747 & pi1067;
assign w22535 = ~w22533 & ~w22534;
assign w22536 = w22532 & w22535;
assign w22537 = pi0847 & pi0894;
assign w22538 = ~pi0746 & ~pi1069;
assign w22539 = ~w22537 & ~w22538;
assign w22540 = ~pi0737 & ~pi1088;
assign w22541 = ~pi0847 & ~pi0894;
assign w22542 = ~w22540 & ~w22541;
assign w22543 = w22539 & w22542;
assign w22544 = w22536 & w22543;
assign w22545 = w22529 & w22544;
assign w22546 = ~pi0617 & ~pi0896;
assign w22547 = pi0748 & pi0931;
assign w22548 = ~w22546 & ~w22547;
assign w22549 = pi0617 & pi0896;
assign w22550 = ~pi0869 & ~pi1085;
assign w22551 = ~w22549 & ~w22550;
assign w22552 = w22548 & w22551;
assign w22553 = ~pi0745 & pi1068;
assign w22554 = pi0745 & ~pi1068;
assign w22555 = ~w22553 & ~w22554;
assign w22556 = ~pi0600 & pi0895;
assign w22557 = pi0600 & ~pi0895;
assign w22558 = ~w22556 & ~w22557;
assign w22559 = ~w22555 & ~w22558;
assign w22560 = w22552 & w22559;
assign w22561 = ~pi0870 & ~pi1087;
assign w22562 = pi0742 & pi0940;
assign w22563 = ~w22561 & ~w22562;
assign w22564 = ~pi0727 & ~pi0897;
assign w22565 = pi0746 & pi1069;
assign w22566 = ~w22564 & ~w22565;
assign w22567 = w22563 & w22566;
assign w22568 = ~pi0748 & ~pi0931;
assign w22569 = pi0727 & pi0897;
assign w22570 = ~w22568 & ~w22569;
assign w22571 = pi0869 & pi1085;
assign w22572 = pi0744 & pi1083;
assign w22573 = ~w22571 & ~w22572;
assign w22574 = w22570 & w22573;
assign w22575 = w22567 & w22574;
assign w22576 = w22560 & w22575;
assign w22577 = w22545 & w22576;
assign w22578 = ~w22514 & ~w22577;
assign w22579 = pi1931 & pi3647;
assign w22580 = ~w22578 & w22579;
assign w22581 = ~w22495 & ~w22580;
assign w22582 = ~w22513 & w22581;
assign w22583 = ~w22512 & w22582;
assign w22584 = ~w22496 & ~w22583;
assign w22585 = pi3576 & pi3635;
assign w22586 = pi0969 & w22585;
assign w22587 = ~pi0933 & pi3635;
assign w22588 = ~pi1071 & w22587;
assign w22589 = ~pi1040 & w22588;
assign w22590 = ~pi1072 & w22589;
assign w22591 = ~pi1027 & w22590;
assign w22592 = ~pi1026 & w22591;
assign w22593 = ~pi0934 & w22592;
assign w22594 = ~pi0935 & w22593;
assign w22595 = ~pi0848 & w22594;
assign w22596 = ~pi1091 & w22595;
assign w22597 = ~pi0690 & w22596;
assign w22598 = ~pi0652 & w22597;
assign w22599 = ~pi0698 & w22598;
assign w22600 = ~pi1070 & w22599;
assign w22601 = ~pi0618 & w22600;
assign w22602 = ~pi0601 & w22601;
assign w22603 = pi0601 & ~w22601;
assign w22604 = ~pi0792 & ~pi0941;
assign w22605 = pi0698 & pi0972;
assign w22606 = ~pi0846 & ~pi1040;
assign w22607 = ~w22605 & ~w22606;
assign w22608 = pi0801 & pi0934;
assign w22609 = ~pi0690 & ~pi0978;
assign w22610 = ~w22608 & ~w22609;
assign w22611 = w22607 & w22610;
assign w22612 = ~pi0848 & ~pi0968;
assign w22613 = pi0618 & pi0970;
assign w22614 = ~w22612 & ~w22613;
assign w22615 = ~pi0981 & ~pi1070;
assign w22616 = pi0848 & pi0968;
assign w22617 = ~w22615 & ~w22616;
assign w22618 = w22614 & w22617;
assign w22619 = w22611 & w22618;
assign w22620 = ~pi0800 & ~pi0935;
assign w22621 = ~pi0698 & ~pi0972;
assign w22622 = ~w22620 & ~w22621;
assign w22623 = ~pi0850 & ~pi1027;
assign w22624 = pi0601 & pi0969;
assign w22625 = ~w22623 & ~w22624;
assign w22626 = w22622 & w22625;
assign w22627 = pi0800 & pi0935;
assign w22628 = pi0802 & pi1026;
assign w22629 = ~w22627 & ~w22628;
assign w22630 = pi0846 & pi1040;
assign w22631 = ~pi0977 & ~pi1091;
assign w22632 = ~w22630 & ~w22631;
assign w22633 = w22629 & w22632;
assign w22634 = w22626 & w22633;
assign w22635 = w22619 & w22634;
assign w22636 = ~pi0803 & pi1072;
assign w22637 = pi0803 & ~pi1072;
assign w22638 = ~w22636 & ~w22637;
assign w22639 = ~pi0618 & ~pi0970;
assign w22640 = pi0805 & pi0933;
assign w22641 = ~w22639 & ~w22640;
assign w22642 = ~w22638 & w22641;
assign w22643 = ~pi0652 & pi0971;
assign w22644 = pi0652 & ~pi0971;
assign w22645 = ~w22643 & ~w22644;
assign w22646 = ~pi0804 & pi1071;
assign w22647 = pi0804 & ~pi1071;
assign w22648 = ~w22646 & ~w22647;
assign w22649 = ~w22645 & ~w22648;
assign w22650 = w22642 & w22649;
assign w22651 = pi0850 & pi1027;
assign w22652 = ~pi0805 & ~pi0933;
assign w22653 = ~w22651 & ~w22652;
assign w22654 = pi0981 & pi1070;
assign w22655 = pi0690 & pi0978;
assign w22656 = ~w22654 & ~w22655;
assign w22657 = w22653 & w22656;
assign w22658 = ~pi0601 & ~pi0969;
assign w22659 = ~pi0802 & ~pi1026;
assign w22660 = ~w22658 & ~w22659;
assign w22661 = pi0977 & pi1091;
assign w22662 = ~pi0801 & ~pi0934;
assign w22663 = ~w22661 & ~w22662;
assign w22664 = w22660 & w22663;
assign w22665 = w22657 & w22664;
assign w22666 = w22650 & w22665;
assign w22667 = w22635 & w22666;
assign w22668 = ~w22604 & ~w22667;
assign w22669 = pi2111 & pi3635;
assign w22670 = ~w22668 & w22669;
assign w22671 = ~w22585 & ~w22670;
assign w22672 = ~w22603 & w22671;
assign w22673 = ~w22602 & w22672;
assign w22674 = ~w22586 & ~w22673;
assign w22675 = w21040 & ~w21192;
assign w22676 = pi0602 & ~w21040;
assign w22677 = ~w22675 & ~w22676;
assign w22678 = w21040 & ~w21259;
assign w22679 = pi0603 & ~w21040;
assign w22680 = ~w22678 & ~w22679;
assign w22681 = pi3100 & w22058;
assign w22682 = pi0789 & pi3540;
assign w22683 = ~w22681 & w22682;
assign w22684 = ~pi0625 & w18003;
assign w22685 = w8240 & w18008;
assign w22686 = ~w22684 & ~w22685;
assign w22687 = ~w18368 & w22686;
assign w22688 = ~w18012 & ~w22687;
assign w22689 = pi0605 & ~w18375;
assign w22690 = ~w22688 & ~w22689;
assign w22691 = ~pi0623 & w18003;
assign w22692 = w1639 & w18008;
assign w22693 = ~w22691 & ~w22692;
assign w22694 = ~w18368 & w22693;
assign w22695 = ~w18012 & ~w22694;
assign w22696 = pi0606 & ~w18375;
assign w22697 = ~w22695 & ~w22696;
assign w22698 = w8081 & w18008;
assign w22699 = ~pi0624 & w18003;
assign w22700 = ~w22698 & ~w22699;
assign w22701 = ~w18368 & w22700;
assign w22702 = ~w18012 & ~w22701;
assign w22703 = pi0607 & ~w18375;
assign w22704 = ~w22702 & ~w22703;
assign w22705 = w21870 & w21879;
assign w22706 = ~w21429 & ~w22705;
assign w22707 = pi0608 & ~w22706;
assign w22708 = ~pi0955 & ~pi1017;
assign w22709 = ~pi0562 & ~pi0693;
assign w22710 = ~w22708 & w22709;
assign w22711 = pi0562 & ~pi0631;
assign w22712 = ~w22710 & ~w22711;
assign w22713 = w22706 & w22712;
assign w22714 = ~w22707 & ~w22713;
assign w22715 = w6506 & w22184;
assign w22716 = ~w6520 & w22182;
assign w22717 = w6177 & w22188;
assign w22718 = w6413 & w22190;
assign w22719 = ~w22178 & ~w22718;
assign w22720 = ~w22717 & w22719;
assign w22721 = ~w22716 & ~w22720;
assign w22722 = ~w22715 & w22721;
assign w22723 = w6421 & w22196;
assign w22724 = w22205 & ~w22723;
assign w22725 = ~w8824 & w22724;
assign w22726 = w22176 & w22181;
assign w22727 = w6473 & w22726;
assign w22728 = ~w6538 & w22179;
assign w22729 = ~w6561 & ~w22728;
assign w22730 = ~w22181 & w22729;
assign w22731 = w22187 & ~w22730;
assign w22732 = ~w22723 & w22731;
assign w22733 = ~w22727 & w22732;
assign w22734 = ~w22725 & ~w22733;
assign w22735 = ~w22722 & w22734;
assign w22736 = w22210 & ~w22735;
assign w22737 = w5053 & w22726;
assign w22738 = w22181 & ~w22187;
assign w22739 = ~w5320 & w22738;
assign w22740 = ~w22188 & ~w22739;
assign w22741 = ~w22737 & ~w22740;
assign w22742 = w5341 & w22178;
assign w22743 = ~w22741 & ~w22742;
assign w22744 = w5377 & w22182;
assign w22745 = ~w22743 & ~w22744;
assign w22746 = w4812 & ~w22176;
assign w22747 = ~w4835 & w22176;
assign w22748 = w22181 & ~w22747;
assign w22749 = ~w4826 & w22179;
assign w22750 = ~w5062 & ~w22749;
assign w22751 = w22182 & w22750;
assign w22752 = ~w22748 & ~w22751;
assign w22753 = ~w22746 & w22752;
assign w22754 = ~w5349 & w22196;
assign w22755 = w22187 & ~w22754;
assign w22756 = ~w22753 & w22755;
assign w22757 = ~w22745 & ~w22756;
assign w22758 = w4502 & w22182;
assign w22759 = ~w4464 & w22184;
assign w22760 = w1308 & w22188;
assign w22761 = w4749 & w22190;
assign w22762 = ~w22178 & ~w22761;
assign w22763 = ~w22760 & w22762;
assign w22764 = ~w22759 & ~w22763;
assign w22765 = ~w22758 & w22764;
assign w22766 = ~w819 & w22184;
assign w22767 = ~w4471 & w22196;
assign w22768 = ~w4757 & w22726;
assign w22769 = ~w883 & w22179;
assign w22770 = ~w4778 & ~w22769;
assign w22771 = ~w22768 & w22770;
assign w22772 = ~w22767 & w22771;
assign w22773 = ~w22766 & w22772;
assign w22774 = w22187 & ~w22773;
assign w22775 = ~w22765 & ~w22774;
assign w22776 = w22757 & ~w22775;
assign w22777 = w22736 & w22776;
assign w22778 = w3831 & ~w22176;
assign w22779 = ~w3878 & w22179;
assign w22780 = ~w3881 & w22187;
assign w22781 = ~w22779 & w22780;
assign w22782 = ~w22778 & w22781;
assign w22783 = ~w3934 & w22188;
assign w22784 = w9004 & w22190;
assign w22785 = ~w22181 & ~w22784;
assign w22786 = ~w22783 & w22785;
assign w22787 = ~w22782 & w22786;
assign w22788 = w22181 & ~w22188;
assign w22789 = w3851 & w22176;
assign w22790 = w22788 & ~w22789;
assign w22791 = w4141 & w22738;
assign w22792 = ~w22790 & ~w22791;
assign w22793 = ~w4380 & w22190;
assign w22794 = w3899 & w22205;
assign w22795 = ~w22793 & ~w22794;
assign w22796 = ~w22792 & w22795;
assign w22797 = ~w22787 & ~w22796;
assign w22798 = w6514 & w22178;
assign w22799 = w6518 & w22178;
assign w22800 = ~w2826 & w22799;
assign w22801 = ~w6177 & w22738;
assign w22802 = ~w22188 & ~w22801;
assign w22803 = ~w22800 & w22802;
assign w22804 = ~w22798 & w22803;
assign w22805 = w6505 & w22182;
assign w22806 = ~w6496 & w22182;
assign w22807 = ~w2826 & w22806;
assign w22808 = w6413 & w22726;
assign w22809 = ~w22807 & ~w22808;
assign w22810 = ~w22805 & w22809;
assign w22811 = ~w22804 & w22810;
assign w22812 = ~w6473 & w22196;
assign w22813 = w22205 & ~w22812;
assign w22814 = ~w5969 & w22813;
assign w22815 = ~w6421 & w22726;
assign w22816 = ~w6446 & w22179;
assign w22817 = ~w6454 & w22187;
assign w22818 = ~w22816 & w22817;
assign w22819 = ~w22184 & w22818;
assign w22820 = ~w22812 & w22819;
assign w22821 = ~w22815 & w22820;
assign w22822 = ~w22814 & ~w22821;
assign w22823 = ~w22811 & w22822;
assign w22824 = w2406 & w22184;
assign w22825 = ~w2413 & w22184;
assign w22826 = ~w798 & w22825;
assign w22827 = ~w2873 & w22726;
assign w22828 = ~w2923 & w22196;
assign w22829 = ~w2863 & w22179;
assign w22830 = ~w2902 & w22187;
assign w22831 = ~w22829 & w22830;
assign w22832 = ~w22828 & w22831;
assign w22833 = ~w22827 & w22832;
assign w22834 = ~w22826 & w22833;
assign w22835 = ~w22824 & w22834;
assign w22836 = ~w40134 & w22726;
assign w22837 = ~w3195 & w22196;
assign w22838 = ~w22836 & ~w22837;
assign w22839 = w2836 & w22184;
assign w22840 = w2834 & w22839;
assign w22841 = w22838 & ~w22840;
assign w22842 = w2829 & w22184;
assign w22843 = ~w2834 & w22842;
assign w22844 = ~w2948 & w22182;
assign w22845 = ~w22843 & ~w22844;
assign w22846 = w22841 & w22845;
assign w22847 = ~w2826 & w22846;
assign w22848 = w2843 & w22184;
assign w22849 = ~w2955 & w22182;
assign w22850 = w22838 & ~w22849;
assign w22851 = ~w22848 & w22850;
assign w22852 = w2826 & w22851;
assign w22853 = ~w22187 & ~w22852;
assign w22854 = ~w22847 & w22853;
assign w22855 = ~w22835 & ~w22854;
assign w22856 = ~w343 & ~w22170;
assign w22857 = w2838 & w22176;
assign w22858 = ~w40134 & w22190;
assign w22859 = ~w3195 & w22188;
assign w22860 = w22181 & ~w22859;
assign w22861 = ~w22858 & w22860;
assign w22862 = ~w22187 & ~w22861;
assign w22863 = w2948 & ~w22176;
assign w22864 = w22862 & ~w22863;
assign w22865 = ~w2826 & w22864;
assign w22866 = ~w22857 & w22865;
assign w22867 = ~w2843 & w22176;
assign w22868 = w2955 & ~w22176;
assign w22869 = w22862 & ~w22868;
assign w22870 = ~w22867 & w22869;
assign w22871 = w2826 & w22870;
assign w22872 = ~w22866 & ~w22871;
assign w22873 = w22856 & w22872;
assign w22874 = w22855 & w22873;
assign w22875 = w22823 & w22874;
assign w22876 = ~w4408 & w22184;
assign w22877 = ~w4423 & w22179;
assign w22878 = ~w4426 & w22187;
assign w22879 = ~w22877 & w22878;
assign w22880 = ~w22181 & ~w22879;
assign w22881 = ~w2873 & ~w22176;
assign w22882 = ~w2923 & w22176;
assign w22883 = w22187 & ~w22882;
assign w22884 = ~w22881 & w22883;
assign w22885 = w22861 & ~w22884;
assign w22886 = ~w22880 & ~w22885;
assign w22887 = ~w22876 & w22886;
assign w22888 = w22176 & w22178;
assign w22889 = ~w5397 & w22888;
assign w22890 = ~w5939 & w22196;
assign w22891 = w22205 & ~w22890;
assign w22892 = ~w5415 & w22891;
assign w22893 = ~w22176 & w22178;
assign w22894 = w5429 & w22893;
assign w22895 = ~w2826 & w22894;
assign w22896 = w5422 & w22893;
assign w22897 = w2826 & w22896;
assign w22898 = w5914 & ~w22176;
assign w22899 = w5635 & w22176;
assign w22900 = w22738 & ~w22899;
assign w22901 = ~w22898 & w22900;
assign w22902 = ~w5659 & w22726;
assign w22903 = ~w5650 & w22179;
assign w22904 = ~w5924 & w22187;
assign w22905 = ~w22903 & w22904;
assign w22906 = ~w22184 & w22905;
assign w22907 = ~w22890 & w22906;
assign w22908 = ~w22902 & w22907;
assign w22909 = ~w22901 & ~w22908;
assign w22910 = ~w22897 & w22909;
assign w22911 = ~w22895 & w22910;
assign w22912 = ~w22892 & w22911;
assign w22913 = ~w22889 & w22912;
assign w22914 = ~w22887 & w22913;
assign w22915 = w22875 & w22914;
assign w22916 = ~w22797 & w22915;
assign w22917 = w22777 & w22916;
assign w22918 = pi0609 & w343;
assign w22919 = ~w22917 & ~w22918;
assign w22920 = pi0610 & ~w22706;
assign w22921 = pi0562 & ~pi0622;
assign w22922 = ~w22710 & ~w22921;
assign w22923 = w22706 & w22922;
assign w22924 = ~w22920 & ~w22923;
assign w22925 = pi0611 & ~w22706;
assign w22926 = pi0562 & ~pi0628;
assign w22927 = ~w22710 & ~w22926;
assign w22928 = w22706 & w22927;
assign w22929 = ~w22925 & ~w22928;
assign w22930 = ~pi0612 & w21497;
assign w22931 = w833 & w926;
assign w22932 = ~w354 & w416;
assign w22933 = w22931 & ~w22932;
assign w22934 = ~pi3367 & ~w926;
assign w22935 = ~w22933 & ~w22934;
assign w22936 = w839 & w926;
assign w22937 = ~w354 & w408;
assign w22938 = w22936 & ~w22937;
assign w22939 = ~pi3391 & ~w926;
assign w22940 = ~w22938 & ~w22939;
assign w22941 = ~w22935 & ~w22940;
assign w22942 = ~pi1010 & w22941;
assign w22943 = w22935 & w22940;
assign w22944 = ~pi0987 & w22943;
assign w22945 = ~w22942 & ~w22944;
assign w22946 = w22935 & ~w22940;
assign w22947 = ~pi0989 & w22946;
assign w22948 = ~w22935 & w22940;
assign w22949 = ~pi0988 & w22948;
assign w22950 = ~w22947 & ~w22949;
assign w22951 = w22945 & w22950;
assign w22952 = w6668 & ~w22951;
assign w22953 = w4141 & w22952;
assign w22954 = ~pi1010 & w6668;
assign w22955 = pi2602 & ~w22954;
assign w22956 = w22941 & w22955;
assign w22957 = ~pi0989 & w6668;
assign w22958 = w22946 & ~w22957;
assign w22959 = pi2675 & w22958;
assign w22960 = ~w22956 & ~w22959;
assign w22961 = ~pi0987 & w6668;
assign w22962 = pi2550 & ~w22961;
assign w22963 = w22943 & w22962;
assign w22964 = ~pi0988 & w6668;
assign w22965 = pi2661 & ~w22964;
assign w22966 = w22948 & w22965;
assign w22967 = ~w22963 & ~w22966;
assign w22968 = w22960 & w22967;
assign w22969 = ~w21497 & w22968;
assign w22970 = ~w22953 & w22969;
assign w22971 = ~w22930 & ~w22970;
assign w22972 = ~pi0613 & w21497;
assign w22973 = w1308 & w22952;
assign w22974 = pi2657 & ~w22961;
assign w22975 = w22943 & w22974;
assign w22976 = pi2685 & w22958;
assign w22977 = ~w22975 & ~w22976;
assign w22978 = pi2671 & ~w22964;
assign w22979 = w22948 & w22978;
assign w22980 = pi2695 & ~w22954;
assign w22981 = w22941 & w22980;
assign w22982 = ~w22979 & ~w22981;
assign w22983 = w22977 & w22982;
assign w22984 = ~w21497 & w22983;
assign w22985 = ~w22973 & w22984;
assign w22986 = ~w22972 & ~w22985;
assign w22987 = ~pi0614 & w21497;
assign w22988 = w5635 & w22952;
assign w22989 = pi2672 & ~w22964;
assign w22990 = w22948 & w22989;
assign w22991 = pi2615 & w22958;
assign w22992 = ~w22990 & ~w22991;
assign w22993 = pi2658 & ~w22961;
assign w22994 = w22943 & w22993;
assign w22995 = pi2696 & ~w22954;
assign w22996 = w22941 & w22995;
assign w22997 = ~w22994 & ~w22996;
assign w22998 = w22992 & w22997;
assign w22999 = ~w21497 & w22998;
assign w23000 = ~w22988 & w22999;
assign w23001 = ~w22987 & ~w23000;
assign w23002 = ~pi0686 & ~pi0921;
assign w23003 = ~w370 & w23002;
assign w23004 = ~pi0616 & w23003;
assign w23005 = ~pi0647 & w23004;
assign w23006 = ~pi0615 & ~w23005;
assign w23007 = ~w370 & ~w21046;
assign w23008 = w21060 & ~w23003;
assign w23009 = w23007 & w23008;
assign w23010 = ~w23006 & ~w23009;
assign w23011 = pi0616 & ~w23003;
assign w23012 = ~w370 & w21047;
assign w23013 = w23011 & ~w23012;
assign w23014 = ~w23003 & ~w23012;
assign w23015 = pi0615 & ~pi0647;
assign w23016 = ~w23007 & w23015;
assign w23017 = ~pi0616 & ~w23016;
assign w23018 = ~w23014 & w23017;
assign w23019 = ~w23013 & ~w23018;
assign w23020 = pi0896 & w22495;
assign w23021 = pi0617 & ~w22510;
assign w23022 = ~w22511 & w22581;
assign w23023 = ~w23021 & w23022;
assign w23024 = ~w23020 & ~w23023;
assign w23025 = pi0970 & w22585;
assign w23026 = pi0618 & ~w22600;
assign w23027 = ~w22601 & w22671;
assign w23028 = ~w23026 & w23027;
assign w23029 = ~w23025 & ~w23028;
assign w23030 = w18318 & w18323;
assign w23031 = pi3439 & ~pi3469;
assign w23032 = pi0827 & ~w23031;
assign w23033 = ~w23030 & w23032;
assign w23034 = ~pi3681 & ~w23033;
assign w23035 = ~pi1428 & w23034;
assign w23036 = pi1370 & ~w18320;
assign w23037 = pi0691 & w23036;
assign w23038 = pi0619 & w23037;
assign w23039 = ~pi0619 & ~w23037;
assign w23040 = ~w23034 & ~w23039;
assign w23041 = ~w23038 & w23040;
assign w23042 = ~w23035 & ~w23041;
assign w23043 = ~pi1427 & w23034;
assign w23044 = ~pi0620 & ~w23038;
assign w23045 = ~w18324 & ~w23034;
assign w23046 = ~w23044 & w23045;
assign w23047 = ~w23043 & ~w23046;
assign w23048 = pi0621 & ~w22706;
assign w23049 = pi0562 & ~pi0608;
assign w23050 = ~w22710 & ~w23049;
assign w23051 = w22706 & w23050;
assign w23052 = ~w23048 & ~w23051;
assign w23053 = pi0622 & ~w22706;
assign w23054 = pi0562 & ~pi0621;
assign w23055 = ~w22710 & ~w23054;
assign w23056 = w22706 & w23055;
assign w23057 = ~w23053 & ~w23056;
assign w23058 = pi0623 & ~w22706;
assign w23059 = pi0562 & ~pi0610;
assign w23060 = ~w22710 & ~w23059;
assign w23061 = w22706 & w23060;
assign w23062 = ~w23058 & ~w23061;
assign w23063 = pi0624 & ~w22706;
assign w23064 = pi0562 & ~pi0623;
assign w23065 = ~w22710 & ~w23064;
assign w23066 = w22706 & w23065;
assign w23067 = ~w23063 & ~w23066;
assign w23068 = pi0625 & ~w22706;
assign w23069 = pi0562 & ~pi0624;
assign w23070 = ~w22710 & ~w23069;
assign w23071 = w22706 & w23070;
assign w23072 = ~w23068 & ~w23071;
assign w23073 = pi0626 & ~w22706;
assign w23074 = pi0562 & ~pi0694;
assign w23075 = ~w22710 & ~w23074;
assign w23076 = w22706 & w23075;
assign w23077 = ~w23073 & ~w23076;
assign w23078 = pi0627 & ~w22706;
assign w23079 = pi0562 & ~pi0626;
assign w23080 = ~w22710 & ~w23079;
assign w23081 = w22706 & w23080;
assign w23082 = ~w23078 & ~w23081;
assign w23083 = pi0628 & ~w22706;
assign w23084 = pi0562 & ~pi0627;
assign w23085 = ~w22710 & ~w23084;
assign w23086 = w22706 & w23085;
assign w23087 = ~w23083 & ~w23086;
assign w23088 = pi0629 & ~w22706;
assign w23089 = pi0562 & ~pi0611;
assign w23090 = ~w22710 & ~w23089;
assign w23091 = w22706 & w23090;
assign w23092 = ~w23088 & ~w23091;
assign w23093 = pi0630 & ~w22706;
assign w23094 = pi0562 & ~pi0629;
assign w23095 = ~w22710 & ~w23094;
assign w23096 = w22706 & w23095;
assign w23097 = ~w23093 & ~w23096;
assign w23098 = pi0631 & ~w22706;
assign w23099 = pi0562 & ~pi0630;
assign w23100 = ~w22710 & ~w23099;
assign w23101 = w22706 & w23100;
assign w23102 = ~w23098 & ~w23101;
assign w23103 = pi0632 & ~w21040;
assign w23104 = w21040 & w21140;
assign w23105 = ~w23103 & ~w23104;
assign w23106 = ~pi0700 & ~w21452;
assign w23107 = ~pi0634 & w21497;
assign w23108 = w5320 & w22952;
assign w23109 = pi2653 & ~w22961;
assign w23110 = w22943 & w23109;
assign w23111 = pi2691 & ~w22954;
assign w23112 = w22941 & w23111;
assign w23113 = ~w23110 & ~w23112;
assign w23114 = pi2681 & ~w22957;
assign w23115 = w22946 & w23114;
assign w23116 = pi2667 & ~w22964;
assign w23117 = w22948 & w23116;
assign w23118 = ~w23115 & ~w23117;
assign w23119 = w23113 & w23118;
assign w23120 = ~w21497 & w23119;
assign w23121 = ~w23108 & w23120;
assign w23122 = ~w23107 & ~w23121;
assign w23123 = ~pi0729 & ~w21366;
assign w23124 = ~pi0636 & w21497;
assign w23125 = w3195 & w22952;
assign w23126 = pi2649 & ~w22961;
assign w23127 = w22943 & w23126;
assign w23128 = pi2688 & ~w22954;
assign w23129 = w22941 & w23128;
assign w23130 = ~w23127 & ~w23129;
assign w23131 = pi2677 & ~w22957;
assign w23132 = w22946 & w23131;
assign w23133 = pi2663 & ~w22964;
assign w23134 = w22948 & w23133;
assign w23135 = ~w23132 & ~w23134;
assign w23136 = w23130 & w23135;
assign w23137 = ~w21497 & w23136;
assign w23138 = ~w23125 & w23137;
assign w23139 = ~w23124 & ~w23138;
assign w23140 = ~pi0637 & w21497;
assign w23141 = w40134 & w22952;
assign w23142 = pi2650 & ~w22961;
assign w23143 = w22943 & w23142;
assign w23144 = pi2678 & w22958;
assign w23145 = ~w23143 & ~w23144;
assign w23146 = pi2563 & ~w22954;
assign w23147 = w22941 & w23146;
assign w23148 = pi2664 & ~w22964;
assign w23149 = w22948 & w23148;
assign w23150 = ~w23147 & ~w23149;
assign w23151 = w23145 & w23150;
assign w23152 = ~w21497 & w23151;
assign w23153 = ~w23141 & w23152;
assign w23154 = ~w23140 & ~w23153;
assign w23155 = ~pi0638 & w21497;
assign w23156 = w4380 & w22952;
assign w23157 = pi2666 & ~w22964;
assign w23158 = w22948 & w23157;
assign w23159 = pi2680 & w22958;
assign w23160 = ~w23158 & ~w23159;
assign w23161 = pi2652 & ~w22961;
assign w23162 = w22943 & w23161;
assign w23163 = pi2690 & ~w22954;
assign w23164 = w22941 & w23163;
assign w23165 = ~w23162 & ~w23164;
assign w23166 = w23160 & w23165;
assign w23167 = ~w21497 & w23166;
assign w23168 = ~w23156 & w23167;
assign w23169 = ~w23155 & ~w23168;
assign w23170 = ~pi0639 & w21497;
assign w23171 = w5914 & w22952;
assign w23172 = pi2654 & ~w22961;
assign w23173 = w22943 & w23172;
assign w23174 = pi2682 & w22958;
assign w23175 = ~w23173 & ~w23174;
assign w23176 = pi2668 & ~w22964;
assign w23177 = w22948 & w23176;
assign w23178 = pi2692 & ~w22954;
assign w23179 = w22941 & w23178;
assign w23180 = ~w23177 & ~w23179;
assign w23181 = w23175 & w23180;
assign w23182 = ~w21497 & w23181;
assign w23183 = ~w23171 & w23182;
assign w23184 = ~w23170 & ~w23183;
assign w23185 = ~pi0640 & w21497;
assign w23186 = w4749 & w22952;
assign w23187 = pi2669 & ~w22964;
assign w23188 = w22948 & w23187;
assign w23189 = pi2683 & w22958;
assign w23190 = ~w23188 & ~w23189;
assign w23191 = pi2655 & ~w22961;
assign w23192 = w22943 & w23191;
assign w23193 = pi2693 & ~w22954;
assign w23194 = w22941 & w23193;
assign w23195 = ~w23192 & ~w23194;
assign w23196 = w23190 & w23195;
assign w23197 = ~w21497 & w23196;
assign w23198 = ~w23186 & w23197;
assign w23199 = ~w23185 & ~w23198;
assign w23200 = ~pi0641 & w21497;
assign w23201 = w3711 & w22952;
assign w23202 = pi2660 & ~w22961;
assign w23203 = w22943 & w23202;
assign w23204 = pi2603 & w22958;
assign w23205 = ~w23203 & ~w23204;
assign w23206 = pi2562 & ~w22954;
assign w23207 = w22941 & w23206;
assign w23208 = pi2674 & ~w22964;
assign w23209 = w22948 & w23208;
assign w23210 = ~w23207 & ~w23209;
assign w23211 = w23205 & w23210;
assign w23212 = ~w21497 & w23211;
assign w23213 = ~w23201 & w23212;
assign w23214 = ~w23200 & ~w23213;
assign w23215 = ~pi0642 & w21497;
assign w23216 = ~w414 & ~w417;
assign w23217 = w22943 & w23216;
assign w23218 = ~w844 & w22948;
assign w23219 = ~w23217 & ~w23218;
assign w23220 = ~w849 & w22941;
assign w23221 = ~w856 & w22946;
assign w23222 = ~w23220 & ~w23221;
assign w23223 = w23219 & w23222;
assign w23224 = ~w8802 & w23223;
assign w23225 = pi2272 & ~w856;
assign w23226 = w22946 & w23225;
assign w23227 = pi2258 & w23217;
assign w23228 = ~w23226 & ~w23227;
assign w23229 = pi2262 & w23218;
assign w23230 = pi1977 & w23220;
assign w23231 = ~w23229 & ~w23230;
assign w23232 = w23228 & w23231;
assign w23233 = ~w21497 & w23232;
assign w23234 = ~w23224 & w23233;
assign w23235 = ~w23215 & ~w23234;
assign w23236 = ~pi0643 & w21497;
assign w23237 = ~w22222 & w23223;
assign w23238 = pi2446 & w23221;
assign w23239 = pi1984 & ~w849;
assign w23240 = w22941 & w23239;
assign w23241 = ~w23238 & ~w23240;
assign w23242 = pi2436 & w23217;
assign w23243 = pi2269 & w23218;
assign w23244 = ~w23242 & ~w23243;
assign w23245 = w23241 & w23244;
assign w23246 = ~w21497 & w23245;
assign w23247 = ~w23237 & w23246;
assign w23248 = ~w23236 & ~w23247;
assign w23249 = ~pi0644 & w21621;
assign w23250 = pi0415 & ~w354;
assign w23251 = w22931 & ~w23250;
assign w23252 = ~pi3392 & ~w926;
assign w23253 = ~w23251 & ~w23252;
assign w23254 = pi0414 & ~w354;
assign w23255 = w22936 & ~w23254;
assign w23256 = ~pi3398 & ~w926;
assign w23257 = ~w23255 & ~w23256;
assign w23258 = w23253 & ~w23257;
assign w23259 = ~pi0920 & w6668;
assign w23260 = w23258 & ~w23259;
assign w23261 = ~w23253 & ~w23257;
assign w23262 = ~pi0991 & w6668;
assign w23263 = w23261 & ~w23262;
assign w23264 = w23253 & w23257;
assign w23265 = pi1051 & w23264;
assign w23266 = ~w23253 & w23257;
assign w23267 = pi0990 & w23266;
assign w23268 = w6668 & ~w23267;
assign w23269 = ~w23265 & w23268;
assign w23270 = ~w23263 & w23269;
assign w23271 = ~w23260 & w23270;
assign w23272 = w6177 & w23271;
assign w23273 = ~pi1051 & w6668;
assign w23274 = pi2709 & ~w23273;
assign w23275 = w23264 & w23274;
assign w23276 = pi2739 & w23263;
assign w23277 = ~w23275 & ~w23276;
assign w23278 = pi2566 & ~w23259;
assign w23279 = w23258 & w23278;
assign w23280 = ~pi0990 & w6668;
assign w23281 = pi2720 & ~w23280;
assign w23282 = w23266 & w23281;
assign w23283 = ~w23279 & ~w23282;
assign w23284 = w23277 & w23283;
assign w23285 = ~w21621 & w23284;
assign w23286 = ~w23272 & w23285;
assign w23287 = ~w23249 & ~w23286;
assign w23288 = ~pi0645 & w21621;
assign w23289 = w1639 & w23271;
assign w23290 = pi2744 & w23263;
assign w23291 = pi2774 & ~w23280;
assign w23292 = w23266 & w23291;
assign w23293 = ~w23290 & ~w23292;
assign w23294 = pi2561 & ~w23259;
assign w23295 = w23258 & w23294;
assign w23296 = pi2716 & ~w23273;
assign w23297 = w23264 & w23296;
assign w23298 = ~w23295 & ~w23297;
assign w23299 = w23293 & w23298;
assign w23300 = ~w21621 & w23299;
assign w23301 = ~w23289 & w23300;
assign w23302 = ~w23288 & ~w23301;
assign w23303 = ~pi0646 & w21621;
assign w23304 = w1308 & w23271;
assign w23305 = pi2543 & w23263;
assign w23306 = pi2725 & ~w23280;
assign w23307 = w23266 & w23306;
assign w23308 = ~w23305 & ~w23307;
assign w23309 = pi2735 & ~w23259;
assign w23310 = w23258 & w23309;
assign w23311 = pi2717 & ~w23273;
assign w23312 = w23264 & w23311;
assign w23313 = ~w23310 & ~w23312;
assign w23314 = w23308 & w23313;
assign w23315 = ~w21621 & w23314;
assign w23316 = ~w23304 & w23315;
assign w23317 = ~w23303 & ~w23316;
assign w23318 = w23011 & w23012;
assign w23319 = ~pi0647 & w23318;
assign w23320 = pi0647 & ~w23004;
assign w23321 = ~w23318 & w23320;
assign w23322 = ~pi0615 & w23005;
assign w23323 = ~w23321 & ~w23322;
assign w23324 = ~w23319 & w23323;
assign w23325 = pi1330 & ~w6682;
assign w23326 = pi1096 & ~pi1641;
assign w23327 = ~pi3681 & w23326;
assign w23328 = pi0648 & pi3238;
assign w23329 = ~w23327 & w23328;
assign w23330 = pi3227 & ~w23329;
assign w23331 = ~w23325 & w23330;
assign w23332 = ~w22333 & w22474;
assign w23333 = ~pi0649 & w6684;
assign w23334 = ~pi0419 & pi0420;
assign w23335 = w22336 & w23334;
assign w23336 = ~w23333 & ~w23335;
assign w23337 = ~w23332 & w23336;
assign w23338 = ~pi0650 & w343;
assign w23339 = ~pi0416 & ~w2232;
assign w23340 = pi0417 & ~w23339;
assign w23341 = ~w343 & ~w23340;
assign w23342 = ~pi0414 & ~w22362;
assign w23343 = ~w22306 & w23342;
assign w23344 = w21800 & w23343;
assign w23345 = pi0427 & w21800;
assign w23346 = w2343 & ~w10683;
assign w23347 = ~w23345 & w23346;
assign w23348 = ~w23344 & ~w23347;
assign w23349 = ~w21950 & ~w23348;
assign w23350 = ~w21973 & ~w23349;
assign w23351 = w23341 & w23350;
assign w23352 = ~w23338 & ~w23351;
assign w23353 = pi0872 & w22495;
assign w23354 = pi0651 & ~w22507;
assign w23355 = ~w22508 & w22581;
assign w23356 = ~w23354 & w23355;
assign w23357 = ~w23353 & ~w23356;
assign w23358 = pi0971 & w22585;
assign w23359 = pi0652 & ~w22597;
assign w23360 = ~w22598 & w22671;
assign w23361 = ~w23359 & w23360;
assign w23362 = ~w23358 & ~w23361;
assign w23363 = ~pi2393 & w18313;
assign w23364 = pi0653 & ~w18332;
assign w23365 = ~w18333 & ~w18359;
assign w23366 = ~w23364 & w23365;
assign w23367 = ~pi1717 & w18359;
assign w23368 = ~w18313 & ~w23367;
assign w23369 = ~w23366 & w23368;
assign w23370 = ~w23363 & ~w23369;
assign w23371 = ~pi0656 & w21621;
assign w23372 = w3711 & w23271;
assign w23373 = pi2532 & ~w23273;
assign w23374 = w23264 & w23373;
assign w23375 = pi2542 & w23263;
assign w23376 = ~w23374 & ~w23375;
assign w23377 = pi2552 & ~w23259;
assign w23378 = w23258 & w23377;
assign w23379 = pi2727 & ~w23280;
assign w23380 = w23266 & w23379;
assign w23381 = ~w23378 & ~w23380;
assign w23382 = w23376 & w23381;
assign w23383 = ~w21621 & w23382;
assign w23384 = ~w23372 & w23383;
assign w23385 = ~w23371 & ~w23384;
assign w23386 = ~pi0657 & w21621;
assign w23387 = w5320 & w23271;
assign w23388 = pi2713 & ~w23273;
assign w23389 = w23264 & w23388;
assign w23390 = pi2742 & w23263;
assign w23391 = ~w23389 & ~w23390;
assign w23392 = pi2733 & w23260;
assign w23393 = pi2723 & ~w23280;
assign w23394 = w23266 & w23393;
assign w23395 = ~w23392 & ~w23394;
assign w23396 = w23391 & w23395;
assign w23397 = ~w21621 & w23396;
assign w23398 = ~w23387 & w23397;
assign w23399 = ~w23386 & ~w23398;
assign w23400 = ~pi0658 & w21497;
assign w23401 = w6177 & w22952;
assign w23402 = pi2662 & ~w22964;
assign w23403 = w22948 & w23402;
assign w23404 = pi2648 & ~w22961;
assign w23405 = w22943 & w23404;
assign w23406 = ~w23403 & ~w23405;
assign w23407 = pi2676 & ~w22957;
assign w23408 = w22946 & w23407;
assign w23409 = pi2687 & ~w22954;
assign w23410 = w22941 & w23409;
assign w23411 = ~w23408 & ~w23410;
assign w23412 = w23406 & w23411;
assign w23413 = ~w21497 & w23412;
assign w23414 = ~w23401 & w23413;
assign w23415 = ~w23400 & ~w23414;
assign w23416 = ~w10711 & w17481;
assign w23417 = ~pi0660 & w21497;
assign w23418 = w874 & ~w4141;
assign w23419 = ~w874 & ~w3831;
assign w23420 = ~w23418 & ~w23419;
assign w23421 = w23223 & w23420;
assign w23422 = pi2257 & w23216;
assign w23423 = w22943 & w23422;
assign w23424 = pi2261 & ~w844;
assign w23425 = w22948 & w23424;
assign w23426 = ~w23423 & ~w23425;
assign w23427 = pi1976 & w23220;
assign w23428 = pi2271 & w23221;
assign w23429 = ~w23427 & ~w23428;
assign w23430 = w23426 & w23429;
assign w23431 = ~w21497 & w23430;
assign w23432 = ~w23421 & w23431;
assign w23433 = ~w23417 & ~w23432;
assign w23434 = ~pi0661 & w21497;
assign w23435 = w874 & ~w6413;
assign w23436 = ~w874 & ~w5969;
assign w23437 = ~w23435 & ~w23436;
assign w23438 = w23223 & w23437;
assign w23439 = pi2442 & ~w856;
assign w23440 = w22946 & w23439;
assign w23441 = pi1978 & w23220;
assign w23442 = ~w23440 & ~w23441;
assign w23443 = pi2432 & w23216;
assign w23444 = w22943 & w23443;
assign w23445 = pi2263 & w23218;
assign w23446 = ~w23444 & ~w23445;
assign w23447 = w23442 & w23446;
assign w23448 = ~w21497 & w23447;
assign w23449 = ~w23438 & w23448;
assign w23450 = ~w23434 & ~w23449;
assign w23451 = ~pi0662 & w21497;
assign w23452 = w8745 & w23223;
assign w23453 = pi2264 & w23218;
assign w23454 = pi2259 & w23217;
assign w23455 = pi2273 & ~w856;
assign w23456 = w22946 & w23455;
assign w23457 = pi1979 & ~w849;
assign w23458 = w22941 & w23457;
assign w23459 = ~w23456 & ~w23458;
assign w23460 = ~w23454 & w23459;
assign w23461 = ~w23453 & w23460;
assign w23462 = ~w21497 & w23461;
assign w23463 = ~w23452 & w23462;
assign w23464 = ~w23451 & ~w23463;
assign w23465 = ~pi0663 & w21497;
assign w23466 = w8699 & w23223;
assign w23467 = pi2443 & ~w856;
assign w23468 = w22946 & w23467;
assign w23469 = pi2260 & w23216;
assign w23470 = w22943 & w23469;
assign w23471 = ~w23468 & ~w23470;
assign w23472 = pi2265 & w23218;
assign w23473 = pi1980 & w23220;
assign w23474 = ~w23472 & ~w23473;
assign w23475 = w23471 & w23474;
assign w23476 = ~w21497 & w23475;
assign w23477 = ~w23466 & w23476;
assign w23478 = ~w23465 & ~w23477;
assign w23479 = ~pi0664 & w21497;
assign w23480 = ~w8667 & w23223;
assign w23481 = pi2266 & ~w844;
assign w23482 = w22948 & w23481;
assign w23483 = pi2274 & w23221;
assign w23484 = ~w23482 & ~w23483;
assign w23485 = pi1981 & w23220;
assign w23486 = pi2433 & w23216;
assign w23487 = w22943 & w23486;
assign w23488 = ~w23485 & ~w23487;
assign w23489 = w23484 & w23488;
assign w23490 = ~w21497 & w23489;
assign w23491 = ~w23480 & w23490;
assign w23492 = ~w23479 & ~w23491;
assign w23493 = ~pi0665 & w21497;
assign w23494 = ~w874 & w8602;
assign w23495 = w874 & w4749;
assign w23496 = ~w23494 & ~w23495;
assign w23497 = w23223 & ~w23496;
assign w23498 = pi2267 & ~w844;
assign w23499 = w22948 & w23498;
assign w23500 = pi1982 & w23220;
assign w23501 = ~w23499 & ~w23500;
assign w23502 = pi2444 & w23221;
assign w23503 = pi2434 & w23216;
assign w23504 = w22943 & w23503;
assign w23505 = ~w23502 & ~w23504;
assign w23506 = w23501 & w23505;
assign w23507 = ~w21497 & w23506;
assign w23508 = ~w23497 & w23507;
assign w23509 = ~w23493 & ~w23508;
assign w23510 = ~pi0666 & w21497;
assign w23511 = w22214 & w23223;
assign w23512 = pi2435 & w23216;
assign w23513 = w22943 & w23512;
assign w23514 = pi2268 & ~w844;
assign w23515 = w22948 & w23514;
assign w23516 = ~w23513 & ~w23515;
assign w23517 = pi1983 & w23220;
assign w23518 = pi2445 & w23221;
assign w23519 = ~w23517 & ~w23518;
assign w23520 = w23516 & w23519;
assign w23521 = ~w21497 & w23520;
assign w23522 = ~w23511 & w23521;
assign w23523 = ~w23510 & ~w23522;
assign w23524 = ~pi0667 & w21497;
assign w23525 = w8560 & w23223;
assign w23526 = pi2437 & w23216;
assign w23527 = w22943 & w23526;
assign w23528 = pi1985 & w23220;
assign w23529 = ~w23527 & ~w23528;
assign w23530 = pi2447 & w23221;
assign w23531 = pi2270 & w23218;
assign w23532 = ~w23530 & ~w23531;
assign w23533 = w23529 & w23532;
assign w23534 = ~w21497 & w23533;
assign w23535 = ~w23525 & w23534;
assign w23536 = ~w23524 & ~w23535;
assign w23537 = ~pi0668 & w21621;
assign w23538 = w4141 & w23271;
assign w23539 = pi2738 & w23263;
assign w23540 = pi2719 & ~w23280;
assign w23541 = w23266 & w23540;
assign w23542 = ~w23539 & ~w23541;
assign w23543 = pi2728 & ~w23259;
assign w23544 = w23258 & w23543;
assign w23545 = pi2708 & ~w23273;
assign w23546 = w23264 & w23545;
assign w23547 = ~w23544 & ~w23546;
assign w23548 = w23542 & w23547;
assign w23549 = ~w21621 & w23548;
assign w23550 = ~w23538 & w23549;
assign w23551 = ~w23537 & ~w23550;
assign w23552 = ~pi0669 & w21621;
assign w23553 = w3195 & w23271;
assign w23554 = pi2729 & w23260;
assign w23555 = pi2531 & ~w23280;
assign w23556 = w23266 & w23555;
assign w23557 = ~w23554 & ~w23556;
assign w23558 = pi2548 & ~w23262;
assign w23559 = w23261 & w23558;
assign w23560 = pi2710 & ~w23273;
assign w23561 = w23264 & w23560;
assign w23562 = ~w23559 & ~w23561;
assign w23563 = w23557 & w23562;
assign w23564 = ~w21621 & w23563;
assign w23565 = ~w23553 & w23564;
assign w23566 = ~w23552 & ~w23565;
assign w23567 = ~pi0670 & w21621;
assign w23568 = w40134 & w23271;
assign w23569 = pi2740 & w23263;
assign w23570 = pi2528 & ~w23280;
assign w23571 = w23266 & w23570;
assign w23572 = ~w23569 & ~w23571;
assign w23573 = pi2730 & ~w23259;
assign w23574 = w23258 & w23573;
assign w23575 = pi2711 & ~w23273;
assign w23576 = w23264 & w23575;
assign w23577 = ~w23574 & ~w23576;
assign w23578 = w23572 & w23577;
assign w23579 = ~w21621 & w23578;
assign w23580 = ~w23568 & w23579;
assign w23581 = ~w23567 & ~w23580;
assign w23582 = ~pi0671 & w21621;
assign w23583 = w6413 & w23271;
assign w23584 = pi2721 & ~w23280;
assign w23585 = w23266 & w23584;
assign w23586 = pi2741 & w23263;
assign w23587 = ~w23585 & ~w23586;
assign w23588 = pi2731 & ~w23259;
assign w23589 = w23258 & w23588;
assign w23590 = pi2536 & ~w23273;
assign w23591 = w23264 & w23590;
assign w23592 = ~w23589 & ~w23591;
assign w23593 = w23587 & w23592;
assign w23594 = ~w21621 & w23593;
assign w23595 = ~w23583 & w23594;
assign w23596 = ~w23582 & ~w23595;
assign w23597 = ~pi0672 & w21621;
assign w23598 = w4380 & w23271;
assign w23599 = pi2722 & ~w23280;
assign w23600 = w23266 & w23599;
assign w23601 = pi2732 & w23260;
assign w23602 = ~w23600 & ~w23601;
assign w23603 = pi2546 & ~w23262;
assign w23604 = w23261 & w23603;
assign w23605 = pi2712 & ~w23273;
assign w23606 = w23264 & w23605;
assign w23607 = ~w23604 & ~w23606;
assign w23608 = w23602 & w23607;
assign w23609 = ~w21621 & w23608;
assign w23610 = ~w23598 & w23609;
assign w23611 = ~w23597 & ~w23610;
assign w23612 = ~pi0673 & w21621;
assign w23613 = w4749 & w23271;
assign w23614 = pi2773 & ~w23280;
assign w23615 = w23266 & w23614;
assign w23616 = pi2743 & w23263;
assign w23617 = ~w23615 & ~w23616;
assign w23618 = pi2734 & ~w23259;
assign w23619 = w23258 & w23618;
assign w23620 = pi2715 & ~w23273;
assign w23621 = w23264 & w23620;
assign w23622 = ~w23619 & ~w23621;
assign w23623 = w23617 & w23622;
assign w23624 = ~w21621 & w23623;
assign w23625 = ~w23613 & w23624;
assign w23626 = ~w23612 & ~w23625;
assign w23627 = ~pi0674 & w21621;
assign w23628 = w5914 & w23271;
assign w23629 = pi2547 & w23263;
assign w23630 = pi2724 & ~w23280;
assign w23631 = w23266 & w23630;
assign w23632 = ~w23629 & ~w23631;
assign w23633 = pi2560 & ~w23259;
assign w23634 = w23258 & w23633;
assign w23635 = pi2714 & ~w23273;
assign w23636 = w23264 & w23635;
assign w23637 = ~w23634 & ~w23636;
assign w23638 = w23632 & w23637;
assign w23639 = ~w21621 & w23638;
assign w23640 = ~w23628 & w23639;
assign w23641 = ~w23627 & ~w23640;
assign w23642 = ~pi0675 & w21621;
assign w23643 = w5635 & w23271;
assign w23644 = pi2565 & ~w23280;
assign w23645 = w23266 & w23644;
assign w23646 = pi2545 & w23263;
assign w23647 = ~w23645 & ~w23646;
assign w23648 = pi2736 & ~w23259;
assign w23649 = w23258 & w23648;
assign w23650 = pi2534 & ~w23273;
assign w23651 = w23264 & w23650;
assign w23652 = ~w23649 & ~w23651;
assign w23653 = w23647 & w23652;
assign w23654 = ~w21621 & w23653;
assign w23655 = ~w23643 & w23654;
assign w23656 = ~w23642 & ~w23655;
assign w23657 = ~pi0676 & w21621;
assign w23658 = w5053 & w23271;
assign w23659 = pi2737 & w23260;
assign w23660 = pi2718 & ~w23273;
assign w23661 = w23264 & w23660;
assign w23662 = ~w23659 & ~w23661;
assign w23663 = pi2745 & ~w23262;
assign w23664 = w23261 & w23663;
assign w23665 = pi2726 & ~w23280;
assign w23666 = w23266 & w23665;
assign w23667 = ~w23664 & ~w23666;
assign w23668 = w23662 & w23667;
assign w23669 = ~w21621 & w23668;
assign w23670 = ~w23658 & w23669;
assign w23671 = ~w23657 & ~w23670;
assign w23672 = ~pi0677 & w21621;
assign w23673 = w2875 & w23261;
assign w23674 = ~w2294 & w23266;
assign w23675 = ~w2315 & w23264;
assign w23676 = ~w2323 & w23258;
assign w23677 = ~w23675 & ~w23676;
assign w23678 = ~w23674 & w23677;
assign w23679 = ~w23673 & w23678;
assign w23680 = ~w2382 & ~w6520;
assign w23681 = w2382 & ~w6177;
assign w23682 = ~w23680 & ~w23681;
assign w23683 = w23679 & w23682;
assign w23684 = w6475 & w23261;
assign w23685 = pi2520 & w23674;
assign w23686 = pi2752 & ~w2323;
assign w23687 = w23258 & w23686;
assign w23688 = pi2535 & w23675;
assign w23689 = ~w23687 & ~w23688;
assign w23690 = ~w23685 & w23689;
assign w23691 = ~w23684 & w23690;
assign w23692 = ~w21621 & w23691;
assign w23693 = ~w23683 & w23692;
assign w23694 = ~w23672 & ~w23693;
assign w23695 = ~pi0678 & w21621;
assign w23696 = ~w2382 & w6506;
assign w23697 = w2382 & ~w6413;
assign w23698 = ~w23696 & ~w23697;
assign w23699 = w23679 & w23698;
assign w23700 = w6423 & w23261;
assign w23701 = pi2527 & w23674;
assign w23702 = pi2753 & ~w2323;
assign w23703 = w23258 & w23702;
assign w23704 = pi2746 & w23675;
assign w23705 = ~w23703 & ~w23704;
assign w23706 = ~w23701 & w23705;
assign w23707 = ~w23700 & w23706;
assign w23708 = ~w21621 & w23707;
assign w23709 = ~w23699 & w23708;
assign w23710 = ~w23695 & ~w23709;
assign w23711 = ~pi0679 & w21621;
assign w23712 = ~w2382 & ~w4464;
assign w23713 = w2382 & ~w4749;
assign w23714 = ~w23712 & ~w23713;
assign w23715 = w23679 & w23714;
assign w23716 = pi2466 & w23673;
assign w23717 = pi2457 & w23674;
assign w23718 = pi2747 & ~w2315;
assign w23719 = w23264 & w23718;
assign w23720 = pi2754 & ~w2323;
assign w23721 = w23258 & w23720;
assign w23722 = ~w23719 & ~w23721;
assign w23723 = ~w23717 & w23722;
assign w23724 = ~w23716 & w23723;
assign w23725 = ~w21621 & w23724;
assign w23726 = ~w23715 & w23725;
assign w23727 = ~w23711 & ~w23726;
assign w23728 = ~pi0680 & w21621;
assign w23729 = ~w1639 & w2382;
assign w23730 = ~w2382 & w3465;
assign w23731 = ~w23729 & ~w23730;
assign w23732 = w23679 & w23731;
assign w23733 = pi2410 & w2875;
assign w23734 = w23261 & w23733;
assign w23735 = pi2530 & ~w2323;
assign w23736 = w23258 & w23735;
assign w23737 = pi2458 & w23674;
assign w23738 = pi2748 & w23675;
assign w23739 = ~w23737 & ~w23738;
assign w23740 = ~w23736 & w23739;
assign w23741 = ~w23734 & w23740;
assign w23742 = ~w21621 & w23741;
assign w23743 = ~w23732 & w23742;
assign w23744 = ~w23728 & ~w23743;
assign w23745 = ~pi0681 & w21621;
assign w23746 = ~w2382 & ~w4502;
assign w23747 = w1308 & w2382;
assign w23748 = ~w23746 & ~w23747;
assign w23749 = w23679 & ~w23748;
assign w23750 = w4759 & w23261;
assign w23751 = w4764 & w23258;
assign w23752 = w4761 & w23264;
assign w23753 = w4766 & w23266;
assign w23754 = ~w23752 & ~w23753;
assign w23755 = ~w23751 & w23754;
assign w23756 = ~w23750 & w23755;
assign w23757 = ~w21621 & w23756;
assign w23758 = ~w23749 & w23757;
assign w23759 = ~w23745 & ~w23758;
assign w23760 = ~pi0682 & w21621;
assign w23761 = ~w2382 & w5397;
assign w23762 = w2382 & w5635;
assign w23763 = ~w23761 & ~w23762;
assign w23764 = w23679 & ~w23763;
assign w23765 = w5661 & w23261;
assign w23766 = pi2459 & w23674;
assign w23767 = pi2749 & w23675;
assign w23768 = pi2544 & ~w2323;
assign w23769 = w23258 & w23768;
assign w23770 = ~w23767 & ~w23769;
assign w23771 = ~w23766 & w23770;
assign w23772 = ~w23765 & w23771;
assign w23773 = ~w21621 & w23772;
assign w23774 = ~w23764 & w23773;
assign w23775 = ~w23760 & ~w23774;
assign w23776 = ~pi0683 & w21621;
assign w23777 = ~w2382 & w5377;
assign w23778 = w2382 & w5053;
assign w23779 = ~w23777 & ~w23778;
assign w23780 = w23679 & ~w23779;
assign w23781 = pi2469 & w23673;
assign w23782 = pi2460 & w23674;
assign w23783 = pi2756 & ~w2323;
assign w23784 = w23258 & w23783;
assign w23785 = pi2750 & w23675;
assign w23786 = ~w23784 & ~w23785;
assign w23787 = ~w23782 & w23786;
assign w23788 = ~w23781 & w23787;
assign w23789 = ~w21621 & w23788;
assign w23790 = ~w23780 & w23789;
assign w23791 = ~w23776 & ~w23790;
assign w23792 = ~pi3203 & ~w342;
assign w23793 = pi0684 & ~w23792;
assign w23794 = ~pi0648 & pi0708;
assign w23795 = ~pi0544 & pi0917;
assign w23796 = pi0916 & ~pi1822;
assign w23797 = pi0912 & pi3538;
assign w23798 = pi2402 & ~w23797;
assign w23799 = pi0913 & ~pi2381;
assign w23800 = w23798 & ~w23799;
assign w23801 = ~pi0522 & pi0914;
assign w23802 = w23800 & ~w23801;
assign w23803 = pi0915 & pi3539;
assign w23804 = w23802 & ~w23803;
assign w23805 = ~w23796 & w23804;
assign w23806 = ~w23795 & w23805;
assign w23807 = pi3641 & ~w23806;
assign w23808 = ~w23794 & ~w23807;
assign w23809 = pi0570 & pi1931;
assign w23810 = ~pi1931 & pi2403;
assign w23811 = pi0918 & pi3641;
assign w23812 = ~w23810 & w23811;
assign w23813 = ~w23809 & w23812;
assign w23814 = w23808 & ~w23813;
assign w23815 = pi0546 & pi1931;
assign w23816 = ~pi1931 & pi2401;
assign w23817 = pi0919 & ~w23816;
assign w23818 = ~w23815 & w23817;
assign w23819 = w23814 & ~w23818;
assign w23820 = ~pi0545 & pi0980;
assign w23821 = w23819 & ~w23820;
assign w23822 = pi3641 & ~w23821;
assign w23823 = ~pi3481 & ~w23822;
assign w23824 = ~pi1046 & pi3481;
assign w23825 = w23792 & ~w23824;
assign w23826 = ~w23823 & w23825;
assign w23827 = w2230 & w23826;
assign w23828 = ~w23793 & ~w23827;
assign w23829 = pi0685 & ~w23003;
assign w23830 = ~w23007 & ~w23829;
assign w23831 = ~w21060 & w23012;
assign w23832 = ~w23830 & ~w23831;
assign w23833 = ~w370 & ~w21035;
assign w23834 = pi0686 & ~w23833;
assign w23835 = ~pi0615 & w21035;
assign w23836 = w23007 & w23835;
assign w23837 = ~w23834 & ~w23836;
assign w23838 = pi2789 & w6668;
assign w23839 = w1213 & w23838;
assign w23840 = w1222 & w1265;
assign w23841 = w23839 & w23840;
assign w23842 = w1639 & w23841;
assign w23843 = ~pi0787 & w22043;
assign w23844 = ~pi0733 & w23843;
assign w23845 = ~pi0786 & w23844;
assign w23846 = ~pi0772 & w23845;
assign w23847 = ~pi0782 & w23846;
assign w23848 = ~pi0771 & w23847;
assign w23849 = ~pi0770 & w23848;
assign w23850 = ~pi0769 & w23849;
assign w23851 = ~pi0732 & w23850;
assign w23852 = ~pi0723 & w23851;
assign w23853 = ~pi0726 & w23852;
assign w23854 = ~pi0725 & w23853;
assign w23855 = ~pi0724 & w23854;
assign w23856 = pi0687 & w23855;
assign w23857 = ~pi0687 & ~w23855;
assign w23858 = ~w23841 & ~w23857;
assign w23859 = ~w23856 & w23858;
assign w23860 = ~w23842 & ~w23859;
assign w23861 = w1204 & w23839;
assign w23862 = w1215 & w23861;
assign w23863 = w1308 & w23862;
assign w23864 = ~pi2059 & ~w903;
assign w23865 = w22040 & ~w23864;
assign w23866 = pi2061 & w23865;
assign w23867 = pi2058 & w23866;
assign w23868 = pi1841 & w23867;
assign w23869 = pi1467 & w23868;
assign w23870 = pi1603 & w23869;
assign w23871 = pi1474 & w23870;
assign w23872 = pi1602 & w23871;
assign w23873 = pi0928 & w23872;
assign w23874 = pi1066 & w23873;
assign w23875 = pi1090 & w23874;
assign w23876 = pi0930 & w23875;
assign w23877 = pi0688 & w23876;
assign w23878 = ~pi0688 & ~w23876;
assign w23879 = ~w23862 & ~w23878;
assign w23880 = ~w23877 & w23879;
assign w23881 = ~w23863 & ~w23880;
assign w23882 = pi0871 & w22495;
assign w23883 = pi0689 & ~w22506;
assign w23884 = ~w22507 & w22581;
assign w23885 = ~w23883 & w23884;
assign w23886 = ~w23882 & ~w23885;
assign w23887 = pi0978 & w22585;
assign w23888 = pi0690 & ~w22596;
assign w23889 = ~w22597 & w22671;
assign w23890 = ~w23888 & w23889;
assign w23891 = ~w23887 & ~w23890;
assign w23892 = ~pi1429 & w23034;
assign w23893 = ~pi0691 & ~w23036;
assign w23894 = ~w23034 & ~w23037;
assign w23895 = ~w23893 & w23894;
assign w23896 = ~w23892 & ~w23895;
assign w23897 = ~w343 & w22227;
assign w23898 = ~pi0692 & w343;
assign w23899 = ~w23897 & ~w23898;
assign w23900 = pi0693 & ~w22706;
assign w23901 = ~pi0958 & pi3664;
assign w23902 = pi0958 & ~w248;
assign w23903 = ~w23901 & ~w23902;
assign w23904 = w22706 & w23903;
assign w23905 = ~w23900 & ~w23904;
assign w23906 = pi0694 & ~w22706;
assign w23907 = pi0693 & w22706;
assign w23908 = ~w23906 & ~w23907;
assign w23909 = ~pi0695 & w6684;
assign w23910 = w21968 & ~w22327;
assign w23911 = w22473 & w23910;
assign w23912 = ~w22356 & w23911;
assign w23913 = ~w23909 & ~w23912;
assign w23914 = pi0696 & ~w20935;
assign w23915 = pi0886 & ~w293;
assign w23916 = ~pi0886 & ~pi3665;
assign w23917 = ~w23915 & ~w23916;
assign w23918 = w20935 & ~w23917;
assign w23919 = ~w23914 & ~w23918;
assign w23920 = ~pi0697 & ~w20935;
assign w23921 = ~w20936 & ~w23920;
assign w23922 = pi0972 & w22585;
assign w23923 = pi0698 & ~w22598;
assign w23924 = ~w22599 & w22671;
assign w23925 = ~w23923 & w23924;
assign w23926 = ~w23922 & ~w23925;
assign w23927 = ~pi2396 & w18313;
assign w23928 = pi0699 & ~w18327;
assign w23929 = ~w18328 & ~w18359;
assign w23930 = ~w23928 & w23929;
assign w23931 = ~pi1721 & w18359;
assign w23932 = ~w18313 & ~w23931;
assign w23933 = ~w23930 & w23932;
assign w23934 = ~w23927 & ~w23933;
assign w23935 = ~pi0701 & w21621;
assign w23936 = w2382 & ~w4141;
assign w23937 = ~w2382 & ~w3934;
assign w23938 = ~w23936 & ~w23937;
assign w23939 = w23679 & w23938;
assign w23940 = w3853 & w23261;
assign w23941 = pi2452 & w23674;
assign w23942 = pi2960 & w23675;
assign w23943 = pi2965 & ~w2323;
assign w23944 = w23258 & w23943;
assign w23945 = ~w23942 & ~w23944;
assign w23946 = ~w23941 & w23945;
assign w23947 = ~w23940 & w23946;
assign w23948 = ~w21621 & w23947;
assign w23949 = ~w23939 & w23948;
assign w23950 = ~w23935 & ~w23949;
assign w23951 = ~pi0702 & w21621;
assign w23952 = ~w2382 & w2845;
assign w23953 = w2382 & ~w3195;
assign w23954 = ~w23952 & ~w23953;
assign w23955 = w23679 & w23954;
assign w23956 = pi2461 & w2875;
assign w23957 = w23261 & w23956;
assign w23958 = pi3096 & ~w2323;
assign w23959 = w23258 & w23958;
assign w23960 = w2930 & w23266;
assign w23961 = pi2961 & w23675;
assign w23962 = ~w23960 & ~w23961;
assign w23963 = ~w23959 & w23962;
assign w23964 = ~w23957 & w23963;
assign w23965 = ~w21621 & w23964;
assign w23966 = ~w23955 & w23965;
assign w23967 = ~w23951 & ~w23966;
assign w23968 = ~pi0703 & w21621;
assign w23969 = w2382 & ~w40134;
assign w23970 = ~w2382 & ~w2957;
assign w23971 = ~w23969 & ~w23970;
assign w23972 = w23679 & w23971;
assign w23973 = pi2462 & w2875;
assign w23974 = w23261 & w23973;
assign w23975 = pi3093 & ~w2323;
assign w23976 = w23258 & w23975;
assign w23977 = pi2962 & w23675;
assign w23978 = pi2454 & w23674;
assign w23979 = ~w23977 & ~w23978;
assign w23980 = ~w23976 & w23979;
assign w23981 = ~w23974 & w23980;
assign w23982 = ~w21621 & w23981;
assign w23983 = ~w23972 & w23982;
assign w23984 = ~w23968 & ~w23983;
assign w23985 = ~pi0704 & w21621;
assign w23986 = ~w2382 & w9004;
assign w23987 = w2382 & ~w4380;
assign w23988 = ~w23986 & ~w23987;
assign w23989 = w23679 & w23988;
assign w23990 = w3901 & w23261;
assign w23991 = pi2455 & w23674;
assign w23992 = pi2963 & ~w2315;
assign w23993 = w23264 & w23992;
assign w23994 = pi2966 & w23676;
assign w23995 = ~w23993 & ~w23994;
assign w23996 = ~w23991 & w23995;
assign w23997 = ~w23990 & w23996;
assign w23998 = ~w21621 & w23997;
assign w23999 = ~w23989 & w23998;
assign w24000 = ~w23985 & ~w23999;
assign w24001 = ~pi0705 & w21621;
assign w24002 = ~w2382 & w5341;
assign w24003 = w2382 & ~w5320;
assign w24004 = ~w24002 & ~w24003;
assign w24005 = w23679 & w24004;
assign w24006 = w5351 & w23261;
assign w24007 = pi2456 & w23674;
assign w24008 = pi2810 & ~w2323;
assign w24009 = w23258 & w24008;
assign w24010 = pi2780 & w23675;
assign w24011 = ~w24009 & ~w24010;
assign w24012 = ~w24007 & w24011;
assign w24013 = ~w24006 & w24012;
assign w24014 = ~w21621 & w24013;
assign w24015 = ~w24005 & w24014;
assign w24016 = ~w24001 & ~w24015;
assign w24017 = ~pi0706 & w21621;
assign w24018 = ~w2382 & ~w8963;
assign w24019 = w2382 & w5914;
assign w24020 = ~w24018 & ~w24019;
assign w24021 = w23679 & ~w24020;
assign w24022 = w5941 & w23261;
assign w24023 = pi2776 & ~w2315;
assign w24024 = w23264 & w24023;
assign w24025 = pi2967 & ~w2323;
assign w24026 = w23258 & w24025;
assign w24027 = pi2526 & w23674;
assign w24028 = ~w24026 & ~w24027;
assign w24029 = ~w24024 & w24028;
assign w24030 = ~w24022 & w24029;
assign w24031 = ~w21621 & w24030;
assign w24032 = ~w24021 & w24031;
assign w24033 = ~w24017 & ~w24032;
assign w24034 = ~pi0707 & w21621;
assign w24035 = ~w2382 & w3814;
assign w24036 = w2382 & ~w3711;
assign w24037 = ~w24035 & ~w24036;
assign w24038 = w23679 & w24037;
assign w24039 = w3763 & w23261;
assign w24040 = pi2524 & w23674;
assign w24041 = w3768 & w23258;
assign w24042 = pi2964 & w23675;
assign w24043 = ~w24041 & ~w24042;
assign w24044 = ~w24040 & w24043;
assign w24045 = ~w24039 & w24044;
assign w24046 = ~w21621 & w24045;
assign w24047 = ~w24038 & w24046;
assign w24048 = ~w24034 & ~w24047;
assign w24049 = pi3641 & ~w6681;
assign w24050 = pi1007 & ~w370;
assign w24051 = ~w10688 & ~w24050;
assign w24052 = ~w24049 & ~w24051;
assign w24053 = pi3293 & ~w9334;
assign w24054 = w24049 & ~w24053;
assign w24055 = pi1048 & pi3293;
assign w24056 = w24054 & ~w24055;
assign w24057 = pi0708 & ~w24056;
assign w24058 = ~w24052 & w24057;
assign w24059 = pi1007 & ~w5320;
assign w24060 = ~pi1041 & ~pi1486;
assign w24061 = pi1041 & ~pi1558;
assign w24062 = ~pi1093 & ~w24061;
assign w24063 = ~w24060 & w24062;
assign w24064 = pi1041 & pi1093;
assign w24065 = pi1590 & w24064;
assign w24066 = ~pi1041 & pi1093;
assign w24067 = pi1523 & w24066;
assign w24068 = pi1042 & ~w24067;
assign w24069 = ~w24065 & w24068;
assign w24070 = ~w24063 & w24069;
assign w24071 = pi1619 & w24064;
assign w24072 = ~pi1041 & pi1624;
assign w24073 = ~pi1042 & ~w24072;
assign w24074 = ~pi1041 & ~pi1093;
assign w24075 = ~pi1093 & pi1415;
assign w24076 = ~w24074 & ~w24075;
assign w24077 = w24073 & w24076;
assign w24078 = ~w24071 & w24077;
assign w24079 = ~pi1007 & ~w24078;
assign w24080 = ~w24070 & w24079;
assign w24081 = w24052 & ~w24080;
assign w24082 = ~w24059 & w24081;
assign w24083 = ~w24058 & ~w24082;
assign w24084 = pi0709 & w6684;
assign w24085 = ~w22365 & w23911;
assign w24086 = ~w24084 & ~w24085;
assign w24087 = pi0710 & w6684;
assign w24088 = w22324 & w23910;
assign w24089 = ~w22365 & w24088;
assign w24090 = ~w24087 & ~w24089;
assign w24091 = ~pi0711 & w6684;
assign w24092 = ~w22333 & w24088;
assign w24093 = ~w24091 & ~w24092;
assign w24094 = ~pi0712 & w6684;
assign w24095 = ~w22333 & w23911;
assign w24096 = ~w24094 & ~w24095;
assign w24097 = ~pi0713 & w6684;
assign w24098 = ~w22489 & w23911;
assign w24099 = ~w24097 & ~w24098;
assign w24100 = ~pi0714 & w6684;
assign w24101 = ~w22489 & w24088;
assign w24102 = ~w24100 & ~w24101;
assign w24103 = pi0715 & w6684;
assign w24104 = ~w22356 & w24088;
assign w24105 = ~w24103 & ~w24104;
assign w24106 = pi0716 & w343;
assign w24107 = ~w21823 & ~w22362;
assign w24108 = w21823 & ~w21944;
assign w24109 = ~w24107 & ~w24108;
assign w24110 = ~w343 & w24109;
assign w24111 = w21831 & w24110;
assign w24112 = ~w24106 & ~w24111;
assign w24113 = pi0717 & w343;
assign w24114 = ~w343 & ~w21844;
assign w24115 = w21841 & w24114;
assign w24116 = w22303 & w24115;
assign w24117 = ~w24113 & ~w24116;
assign w24118 = pi0718 & w343;
assign w24119 = w21831 & w24115;
assign w24120 = ~w24118 & ~w24119;
assign w24121 = pi0719 & w343;
assign w24122 = ~w343 & ~w21841;
assign w24123 = w21831 & w24122;
assign w24124 = ~w24121 & ~w24123;
assign w24125 = pi0720 & w343;
assign w24126 = w22303 & w24122;
assign w24127 = ~w24125 & ~w24126;
assign w24128 = pi0721 & w343;
assign w24129 = ~w343 & w21836;
assign w24130 = ~w24128 & ~w24129;
assign w24131 = pi0722 & w343;
assign w24132 = ~w343 & w21801;
assign w24133 = ~w2343 & w24132;
assign w24134 = ~w24131 & ~w24133;
assign w24135 = ~w4141 & w23841;
assign w24136 = pi0723 & ~w23851;
assign w24137 = ~w23841 & ~w23852;
assign w24138 = ~w24136 & w24137;
assign w24139 = ~w24135 & ~w24138;
assign w24140 = ~w1308 & w23841;
assign w24141 = pi0724 & ~w23854;
assign w24142 = ~w23841 & ~w23855;
assign w24143 = ~w24141 & w24142;
assign w24144 = ~w24140 & ~w24143;
assign w24145 = ~w5635 & w23841;
assign w24146 = pi0725 & ~w23853;
assign w24147 = ~w23841 & ~w23854;
assign w24148 = ~w24146 & w24147;
assign w24149 = ~w24145 & ~w24148;
assign w24150 = ~w5053 & w23841;
assign w24151 = pi0726 & ~w23852;
assign w24152 = ~w23841 & ~w23853;
assign w24153 = ~w24151 & w24152;
assign w24154 = ~w24150 & ~w24153;
assign w24155 = pi0897 & w22495;
assign w24156 = pi0727 & ~w22508;
assign w24157 = ~w22509 & w22581;
assign w24158 = ~w24156 & w24157;
assign w24159 = ~w24155 & ~w24158;
assign w24160 = ~pi2094 & w18313;
assign w24161 = pi0728 & ~w18328;
assign w24162 = ~w18329 & ~w18359;
assign w24163 = ~w24161 & w24162;
assign w24164 = ~pi1720 & w18359;
assign w24165 = ~w18313 & ~w24164;
assign w24166 = ~w24163 & w24165;
assign w24167 = ~w24160 & ~w24166;
assign w24168 = pi3502 & pi3506;
assign w24169 = pi3677 & ~w24168;
assign w24170 = ~pi3502 & ~pi3506;
assign w24171 = ~pi3425 & ~w24170;
assign w24172 = w24169 & ~w24171;
assign w24173 = ~pi3425 & ~w24169;
assign w24174 = ~w24172 & ~w24173;
assign w24175 = pi3502 & w24174;
assign w24176 = pi3502 & ~pi3677;
assign w24177 = ~w24175 & ~w24176;
assign w24178 = pi0730 & w24177;
assign w24179 = pi3677 & w24175;
assign w24180 = ~pi3266 & ~pi3271;
assign w24181 = w19515 & w24180;
assign w24182 = w24179 & ~w24181;
assign w24183 = pi3266 & pi3271;
assign w24184 = pi3246 & pi3255;
assign w24185 = w24183 & w24184;
assign w24186 = ~pi3090 & w24185;
assign w24187 = pi0406 & w19957;
assign w24188 = ~w24186 & ~w24187;
assign w24189 = w19956 & w24183;
assign w24190 = ~pi1386 & w24189;
assign w24191 = pi0381 & w19516;
assign w24192 = ~w24190 & ~w24191;
assign w24193 = ~pi3246 & pi3255;
assign w24194 = w19514 & w24193;
assign w24195 = ~pi3004 & w24194;
assign w24196 = w24180 & w24193;
assign w24197 = ~pi3018 & w24196;
assign w24198 = ~w24195 & ~w24197;
assign w24199 = w24192 & w24198;
assign w24200 = w24188 & w24199;
assign w24201 = ~pi3266 & pi3271;
assign w24202 = ~pi3049 & w24193;
assign w24203 = ~pi2898 & w24184;
assign w24204 = ~w24202 & ~w24203;
assign w24205 = ~pi2761 & w19515;
assign w24206 = pi0812 & w19956;
assign w24207 = ~w24205 & ~w24206;
assign w24208 = w24204 & w24207;
assign w24209 = w24201 & ~w24208;
assign w24210 = w24180 & w24184;
assign w24211 = ~pi3011 & w24210;
assign w24212 = w19514 & w24184;
assign w24213 = ~pi2995 & w24212;
assign w24214 = ~w24211 & ~w24213;
assign w24215 = w19515 & w24183;
assign w24216 = ~pi1361 & w24215;
assign w24217 = w24183 & w24193;
assign w24218 = ~pi2881 & w24217;
assign w24219 = ~w24216 & ~w24218;
assign w24220 = w24214 & w24219;
assign w24221 = ~w24209 & w24220;
assign w24222 = w24200 & w24221;
assign w24223 = w24182 & w24222;
assign w24224 = ~pi0859 & ~w24175;
assign w24225 = pi3425 & w24176;
assign w24226 = ~pi0731 & w24225;
assign w24227 = ~w24177 & ~w24226;
assign w24228 = ~w24224 & w24227;
assign w24229 = ~w24223 & w24228;
assign w24230 = ~w24178 & ~w24229;
assign w24231 = pi0731 & w24177;
assign w24232 = ~pi2956 & w24196;
assign w24233 = w24193 & w24201;
assign w24234 = ~pi3050 & w24233;
assign w24235 = ~w24232 & ~w24234;
assign w24236 = w24184 & w24201;
assign w24237 = ~pi3092 & w24236;
assign w24238 = ~pi1363 & w24189;
assign w24239 = ~w24237 & ~w24238;
assign w24240 = w24235 & w24239;
assign w24241 = pi0425 & w19957;
assign w24242 = ~pi3056 & w24210;
assign w24243 = ~w24241 & ~w24242;
assign w24244 = ~pi2900 & w24212;
assign w24245 = ~pi3027 & w24185;
assign w24246 = ~w24244 & ~w24245;
assign w24247 = w24243 & w24246;
assign w24248 = w24240 & w24247;
assign w24249 = w19956 & w24201;
assign w24250 = w19515 & w24201;
assign w24251 = ~pi2643 & w24250;
assign w24252 = ~w24249 & ~w24251;
assign w24253 = ~pi0813 & pi3246;
assign w24254 = ~w24252 & ~w24253;
assign w24255 = ~pi1701 & w24215;
assign w24256 = pi0391 & w19516;
assign w24257 = ~w24255 & ~w24256;
assign w24258 = ~pi2884 & w24194;
assign w24259 = ~pi3035 & w24217;
assign w24260 = ~w24258 & ~w24259;
assign w24261 = w24257 & w24260;
assign w24262 = ~w24254 & w24261;
assign w24263 = w24248 & w24262;
assign w24264 = w24182 & w24263;
assign w24265 = ~pi0730 & ~w24175;
assign w24266 = ~pi0938 & w24225;
assign w24267 = ~w24177 & ~w24266;
assign w24268 = ~w24265 & w24267;
assign w24269 = ~w24264 & w24268;
assign w24270 = ~w24231 & ~w24269;
assign w24271 = ~w6177 & w23841;
assign w24272 = pi0732 & ~w23850;
assign w24273 = ~w23841 & ~w23851;
assign w24274 = ~w24272 & w24273;
assign w24275 = ~w24271 & ~w24274;
assign w24276 = ~w4749 & w23841;
assign w24277 = pi0733 & ~w23843;
assign w24278 = ~w23844 & ~w24277;
assign w24279 = ~w23841 & w24278;
assign w24280 = ~w24276 & ~w24279;
assign w24281 = ~pi0734 & w6684;
assign w24282 = ~w343 & w21991;
assign w24283 = w21994 & w24282;
assign w24284 = w6682 & ~w21975;
assign w24285 = ~w21980 & w24284;
assign w24286 = w24283 & w24285;
assign w24287 = ~pi0413 & w21983;
assign w24288 = ~w22330 & ~w24287;
assign w24289 = w24286 & ~w24288;
assign w24290 = ~w24281 & ~w24289;
assign w24291 = ~pi0735 & w21497;
assign w24292 = w5053 & w22952;
assign w24293 = pi2697 & ~w22954;
assign w24294 = w22941 & w24293;
assign w24295 = pi2686 & w22958;
assign w24296 = ~w24294 & ~w24295;
assign w24297 = pi2673 & ~w22964;
assign w24298 = w22948 & w24297;
assign w24299 = pi2659 & ~w22961;
assign w24300 = w22943 & w24299;
assign w24301 = ~w24298 & ~w24300;
assign w24302 = w24296 & w24301;
assign w24303 = ~w21497 & w24302;
assign w24304 = ~w24292 & w24303;
assign w24305 = ~w24291 & ~w24304;
assign w24306 = ~pi0736 & w21497;
assign w24307 = w6413 & w22952;
assign w24308 = pi2665 & ~w22964;
assign w24309 = w22948 & w24308;
assign w24310 = pi2679 & w22958;
assign w24311 = ~w24309 & ~w24310;
assign w24312 = pi2689 & ~w22954;
assign w24313 = w22941 & w24312;
assign w24314 = pi2651 & ~w22961;
assign w24315 = w22943 & w24314;
assign w24316 = ~w24313 & ~w24315;
assign w24317 = w24311 & w24316;
assign w24318 = ~w21497 & w24317;
assign w24319 = ~w24307 & w24318;
assign w24320 = ~w24306 & ~w24319;
assign w24321 = w1231 & w23839;
assign w24322 = pi0609 & w24321;
assign w24323 = w1204 & w24322;
assign w24324 = ~pi1033 & w24323;
assign w24325 = ~w5914 & w24324;
assign w24326 = pi1033 & ~w8081;
assign w24327 = w24323 & ~w24326;
assign w24328 = ~pi0737 & ~w24327;
assign w24329 = ~w24325 & ~w24328;
assign w24330 = pi0609 & pi1032;
assign w24331 = w23861 & w24330;
assign w24332 = w1214 & w24331;
assign w24333 = ~w4141 & w24332;
assign w24334 = pi1033 & w24331;
assign w24335 = ~pi1012 & w24334;
assign w24336 = w8081 & w24335;
assign w24337 = ~w24332 & ~w24336;
assign w24338 = ~pi0738 & w24337;
assign w24339 = ~w24333 & ~w24338;
assign w24340 = w1241 & w23861;
assign w24341 = w8081 & w24340;
assign w24342 = ~w4749 & ~w24341;
assign w24343 = ~w24337 & w24342;
assign w24344 = ~pi0739 & w24337;
assign w24345 = ~w24343 & ~w24344;
assign w24346 = ~w5053 & w24332;
assign w24347 = ~pi0740 & w24337;
assign w24348 = ~w24346 & ~w24347;
assign w24349 = ~w3711 & ~w24341;
assign w24350 = ~w24337 & w24349;
assign w24351 = ~pi0741 & w24337;
assign w24352 = ~w24350 & ~w24351;
assign w24353 = ~w3195 & w24324;
assign w24354 = ~pi0742 & ~w24327;
assign w24355 = ~w24353 & ~w24354;
assign w24356 = ~w40134 & w24324;
assign w24357 = ~pi0743 & ~w24327;
assign w24358 = ~w24356 & ~w24357;
assign w24359 = ~w6413 & w24324;
assign w24360 = ~pi0744 & ~w24327;
assign w24361 = ~w24359 & ~w24360;
assign w24362 = ~w4380 & w24324;
assign w24363 = ~pi0745 & ~w24327;
assign w24364 = ~w24362 & ~w24363;
assign w24365 = ~w5320 & w24324;
assign w24366 = ~pi0746 & ~w24327;
assign w24367 = ~w24365 & ~w24366;
assign w24368 = w24327 & ~w24342;
assign w24369 = pi0747 & ~w24327;
assign w24370 = ~w24368 & ~w24369;
assign w24371 = w24327 & ~w24349;
assign w24372 = pi0748 & ~w24327;
assign w24373 = ~w24371 & ~w24372;
assign w24374 = w1225 & w23839;
assign w24375 = w1265 & w24374;
assign w24376 = w3711 & w24375;
assign w24377 = pi0749 & w22043;
assign w24378 = ~pi0749 & ~w22043;
assign w24379 = ~w24377 & ~w24378;
assign w24380 = ~w24375 & w24379;
assign w24381 = ~w24376 & ~w24380;
assign w24382 = w10752 & w16068;
assign w24383 = ~w40171 & w18039;
assign w24384 = ~pi0750 & ~w18039;
assign w24385 = ~w10753 & ~w24384;
assign w24386 = ~w24383 & w24385;
assign w24387 = w15173 & ~w24386;
assign w24388 = ~w24382 & ~w24387;
assign w24389 = w13923 & w16068;
assign w24390 = ~w40171 & w18046;
assign w24391 = ~pi0751 & ~w18046;
assign w24392 = ~w13925 & ~w24391;
assign w24393 = ~w24390 & w24392;
assign w24394 = w14336 & ~w24393;
assign w24395 = ~w24389 & ~w24394;
assign w24396 = w1639 & w24375;
assign w24397 = pi0778 & w24377;
assign w24398 = pi0777 & w24397;
assign w24399 = pi0776 & w24398;
assign w24400 = pi0775 & w24399;
assign w24401 = pi0774 & w24400;
assign w24402 = pi0773 & w24401;
assign w24403 = pi0861 & w24402;
assign w24404 = pi0862 & w24403;
assign w24405 = pi0845 & w24404;
assign w24406 = pi0781 & w24405;
assign w24407 = pi0780 & w24406;
assign w24408 = pi0779 & w24407;
assign w24409 = pi0752 & w24408;
assign w24410 = ~pi0752 & ~w24408;
assign w24411 = ~w24375 & ~w24410;
assign w24412 = ~w24409 & w24411;
assign w24413 = ~w24396 & ~w24412;
assign w24414 = ~pi0753 & w21497;
assign w24415 = w1639 & w22952;
assign w24416 = pi2670 & ~w22964;
assign w24417 = w22948 & w24416;
assign w24418 = pi2684 & w22958;
assign w24419 = ~w24417 & ~w24418;
assign w24420 = pi2694 & ~w22954;
assign w24421 = w22941 & w24420;
assign w24422 = pi2656 & ~w22961;
assign w24423 = w22943 & w24422;
assign w24424 = ~w24421 & ~w24423;
assign w24425 = w24419 & w24424;
assign w24426 = ~w21497 & w24425;
assign w24427 = ~w24415 & w24426;
assign w24428 = ~w24414 & ~w24427;
assign w24429 = ~pi0754 & w21497;
assign w24430 = w8826 & w23223;
assign w24431 = pi2275 & ~w849;
assign w24432 = w22941 & w24431;
assign w24433 = pi2701 & w23221;
assign w24434 = ~w24432 & ~w24433;
assign w24435 = pi2438 & w23218;
assign w24436 = pi2698 & w23217;
assign w24437 = ~w24435 & ~w24436;
assign w24438 = w24434 & w24437;
assign w24439 = ~w21497 & w24438;
assign w24440 = ~w24430 & w24439;
assign w24441 = ~w24429 & ~w24440;
assign w24442 = ~pi0755 & w21497;
assign w24443 = ~w874 & w4408;
assign w24444 = w874 & ~w3195;
assign w24445 = ~w24443 & ~w24444;
assign w24446 = w23223 & w24445;
assign w24447 = pi2699 & w23216;
assign w24448 = w22943 & w24447;
assign w24449 = pi2702 & ~w856;
assign w24450 = w22946 & w24449;
assign w24451 = ~w24448 & ~w24450;
assign w24452 = pi2439 & w23218;
assign w24453 = pi2276 & w23220;
assign w24454 = ~w24452 & ~w24453;
assign w24455 = w24451 & w24454;
assign w24456 = ~w21497 & w24455;
assign w24457 = ~w24446 & w24456;
assign w24458 = ~w24442 & ~w24457;
assign w24459 = ~pi0756 & w21497;
assign w24460 = w874 & ~w5635;
assign w24461 = ~w874 & ~w5415;
assign w24462 = ~w24460 & ~w24461;
assign w24463 = w23223 & w24462;
assign w24464 = pi2277 & w23220;
assign w24465 = pi2539 & w23217;
assign w24466 = pi2440 & ~w844;
assign w24467 = w22948 & w24466;
assign w24468 = pi2703 & ~w856;
assign w24469 = w22946 & w24468;
assign w24470 = ~w24467 & ~w24469;
assign w24471 = ~w24465 & w24470;
assign w24472 = ~w24464 & w24471;
assign w24473 = ~w21497 & w24472;
assign w24474 = ~w24463 & w24473;
assign w24475 = ~w24459 & ~w24474;
assign w24476 = ~pi0757 & w21497;
assign w24477 = ~w874 & ~w4812;
assign w24478 = w874 & w5053;
assign w24479 = ~w24477 & ~w24478;
assign w24480 = w23223 & ~w24479;
assign w24481 = pi2751 & ~w856;
assign w24482 = w22946 & w24481;
assign w24483 = pi2278 & w23220;
assign w24484 = ~w24482 & ~w24483;
assign w24485 = pi2441 & w23218;
assign w24486 = pi2700 & w23216;
assign w24487 = w22943 & w24486;
assign w24488 = ~w24485 & ~w24487;
assign w24489 = w24484 & w24488;
assign w24490 = ~w21497 & w24489;
assign w24491 = ~w24480 & w24490;
assign w24492 = ~w24476 & ~w24491;
assign w24493 = ~pi0758 & w6684;
assign w24494 = ~w21984 & w21987;
assign w24495 = w24286 & w24494;
assign w24496 = ~w24493 & ~w24495;
assign w24497 = pi0759 & w6684;
assign w24498 = w21988 & w24286;
assign w24499 = w2230 & w24498;
assign w24500 = ~w24497 & ~w24499;
assign w24501 = ~pi0760 & w6684;
assign w24502 = w6682 & w21994;
assign w24503 = ~w343 & ~w21991;
assign w24504 = w22000 & w24503;
assign w24505 = w24502 & w24504;
assign w24506 = w21984 & ~w21987;
assign w24507 = w24505 & w24506;
assign w24508 = ~w24501 & ~w24507;
assign w24509 = pi0761 & w343;
assign w24510 = w22303 & w24110;
assign w24511 = ~w24509 & ~w24510;
assign w24512 = pi0762 & w343;
assign w24513 = ~w343 & w21951;
assign w24514 = w385 & w24513;
assign w24515 = ~w24512 & ~w24514;
assign w24516 = pi0763 & w343;
assign w24517 = w21830 & w21843;
assign w24518 = w24110 & w24517;
assign w24519 = ~w24516 & ~w24518;
assign w24520 = pi0764 & w343;
assign w24521 = ~w21830 & w21843;
assign w24522 = w24110 & w24521;
assign w24523 = ~w24520 & ~w24522;
assign w24524 = pi0765 & w343;
assign w24525 = ~w343 & w21835;
assign w24526 = w24517 & w24525;
assign w24527 = ~w24524 & ~w24526;
assign w24528 = pi0766 & w343;
assign w24529 = w24521 & w24525;
assign w24530 = ~w24528 & ~w24529;
assign w24531 = pi0767 & w343;
assign w24532 = w24122 & w24517;
assign w24533 = ~w24531 & ~w24532;
assign w24534 = pi0768 & w343;
assign w24535 = w24122 & w24521;
assign w24536 = ~w24534 & ~w24535;
assign w24537 = ~w3195 & w23841;
assign w24538 = pi0769 & ~w23849;
assign w24539 = ~w23841 & ~w23850;
assign w24540 = ~w24538 & w24539;
assign w24541 = ~w24537 & ~w24540;
assign w24542 = ~w40134 & w23841;
assign w24543 = pi0770 & ~w23848;
assign w24544 = ~w23841 & ~w23849;
assign w24545 = ~w24543 & w24544;
assign w24546 = ~w24542 & ~w24545;
assign w24547 = ~pi3651 & ~pi3652;
assign w24548 = ~pi3525 & ~w24547;
assign w24549 = ~pi3525 & w24547;
assign w24550 = ~w6413 & w23841;
assign w24551 = pi0771 & ~w23847;
assign w24552 = ~w23841 & ~w23848;
assign w24553 = ~w24551 & w24552;
assign w24554 = ~w24550 & ~w24553;
assign w24555 = ~w5320 & w23841;
assign w24556 = pi0772 & ~w23845;
assign w24557 = ~w23846 & ~w24556;
assign w24558 = ~w23841 & w24557;
assign w24559 = ~w24555 & ~w24558;
assign w24560 = w40134 & w24375;
assign w24561 = ~pi0773 & ~w24401;
assign w24562 = ~w24375 & ~w24402;
assign w24563 = ~w24561 & w24562;
assign w24564 = ~w24560 & ~w24563;
assign w24565 = w6413 & w24375;
assign w24566 = ~pi0774 & ~w24400;
assign w24567 = ~w24375 & ~w24401;
assign w24568 = ~w24566 & w24567;
assign w24569 = ~w24565 & ~w24568;
assign w24570 = w4380 & w24375;
assign w24571 = ~pi0775 & ~w24399;
assign w24572 = ~w24400 & ~w24571;
assign w24573 = ~w24375 & w24572;
assign w24574 = ~w24570 & ~w24573;
assign w24575 = w5320 & w24375;
assign w24576 = ~pi0776 & ~w24398;
assign w24577 = ~w24399 & ~w24576;
assign w24578 = ~w24375 & w24577;
assign w24579 = ~w24575 & ~w24578;
assign w24580 = w5914 & w24375;
assign w24581 = ~pi0777 & ~w24397;
assign w24582 = ~w24398 & ~w24581;
assign w24583 = ~w24375 & w24582;
assign w24584 = ~w24580 & ~w24583;
assign w24585 = w4749 & w24375;
assign w24586 = ~pi0778 & ~w24377;
assign w24587 = ~w24397 & ~w24586;
assign w24588 = ~w24375 & w24587;
assign w24589 = ~w24585 & ~w24588;
assign w24590 = w1308 & w24375;
assign w24591 = ~pi0779 & ~w24407;
assign w24592 = ~w24375 & ~w24408;
assign w24593 = ~w24591 & w24592;
assign w24594 = ~w24590 & ~w24593;
assign w24595 = w5635 & w24375;
assign w24596 = ~pi0780 & ~w24406;
assign w24597 = ~w24375 & ~w24407;
assign w24598 = ~w24596 & w24597;
assign w24599 = ~w24595 & ~w24598;
assign w24600 = w5053 & w24375;
assign w24601 = ~pi0781 & ~w24405;
assign w24602 = ~w24375 & ~w24406;
assign w24603 = ~w24601 & w24602;
assign w24604 = ~w24600 & ~w24603;
assign w24605 = ~w4380 & w23841;
assign w24606 = pi0782 & ~w23846;
assign w24607 = ~w23841 & ~w23847;
assign w24608 = ~w24606 & w24607;
assign w24609 = ~w24605 & ~w24608;
assign w24610 = pi0784 & ~w22058;
assign w24611 = pi0785 & w24177;
assign w24612 = w24179 & ~w24250;
assign w24613 = ~pi3014 & w24210;
assign w24614 = ~pi3089 & w24217;
assign w24615 = ~w24613 & ~w24614;
assign w24616 = pi0403 & w19957;
assign w24617 = ~pi3006 & w24194;
assign w24618 = ~w24616 & ~w24617;
assign w24619 = ~pi1086 & w24189;
assign w24620 = ~pi2997 & w24212;
assign w24621 = ~w24619 & ~w24620;
assign w24622 = w24618 & w24621;
assign w24623 = w24615 & w24622;
assign w24624 = w19956 & w24180;
assign w24625 = ~pi3205 & w24624;
assign w24626 = pi0816 & w24249;
assign w24627 = ~w24625 & ~w24626;
assign w24628 = ~pi2806 & w24236;
assign w24629 = ~pi3057 & w24185;
assign w24630 = ~w24628 & ~w24629;
assign w24631 = w24627 & w24630;
assign w24632 = ~pi1674 & w24215;
assign w24633 = ~pi2837 & w24196;
assign w24634 = ~w24632 & ~w24633;
assign w24635 = pi0369 & w19516;
assign w24636 = ~pi3053 & w24233;
assign w24637 = ~w24635 & ~w24636;
assign w24638 = w24634 & w24637;
assign w24639 = w24631 & w24638;
assign w24640 = w24623 & w24639;
assign w24641 = w24612 & w24640;
assign w24642 = ~pi0854 & ~w24175;
assign w24643 = ~pi0825 & w24225;
assign w24644 = ~w24177 & ~w24643;
assign w24645 = ~w24642 & w24644;
assign w24646 = ~w24641 & w24645;
assign w24647 = ~w24611 & ~w24646;
assign w24648 = ~w5914 & w23841;
assign w24649 = pi0786 & ~w23844;
assign w24650 = ~w23845 & ~w24649;
assign w24651 = ~w23841 & w24650;
assign w24652 = ~w24648 & ~w24651;
assign w24653 = ~w3711 & w23841;
assign w24654 = ~w22044 & ~w23843;
assign w24655 = ~w23841 & w24654;
assign w24656 = ~w24653 & ~w24655;
assign w24657 = pi3420 & ~w341;
assign w24658 = w19517 & w24249;
assign w24659 = ~pi0788 & ~w24658;
assign w24660 = ~pi0855 & w24658;
assign w24661 = ~w24659 & ~w24660;
assign w24662 = w341 & w24661;
assign w24663 = ~w24657 & ~w24662;
assign w24664 = ~w6177 & w24332;
assign w24665 = ~pi0790 & w24337;
assign w24666 = ~w24664 & ~w24665;
assign w24667 = ~w5635 & w24332;
assign w24668 = ~pi0791 & w24337;
assign w24669 = ~w24667 & ~w24668;
assign w24670 = pi1012 & w24330;
assign w24671 = w23839 & w24670;
assign w24672 = w1223 & w24671;
assign w24673 = ~w4141 & w24672;
assign w24674 = ~pi1033 & w1236;
assign w24675 = w24671 & w24674;
assign w24676 = w8081 & w24675;
assign w24677 = ~w24672 & ~w24676;
assign w24678 = ~pi0792 & w24677;
assign w24679 = ~w24673 & ~w24678;
assign w24680 = ~pi0793 & w24677;
assign w24681 = w1236 & w23839;
assign w24682 = w1244 & w24681;
assign w24683 = w8081 & w24682;
assign w24684 = ~w4749 & ~w24683;
assign w24685 = w24672 & w24684;
assign w24686 = ~w24680 & ~w24685;
assign w24687 = ~w5053 & w24672;
assign w24688 = ~pi0794 & w24677;
assign w24689 = ~w24687 & ~w24688;
assign w24690 = ~pi0795 & w24677;
assign w24691 = ~w3711 & ~w24683;
assign w24692 = w24672 & w24691;
assign w24693 = ~w24690 & ~w24692;
assign w24694 = ~w8081 & w24675;
assign w24695 = ~pi0796 & ~w24675;
assign w24696 = ~w24694 & ~w24695;
assign w24697 = ~w5320 & w24694;
assign w24698 = ~pi0797 & ~w24675;
assign w24699 = ~w24697 & ~w24698;
assign w24700 = ~w5914 & w24694;
assign w24701 = ~pi0798 & ~w24675;
assign w24702 = ~w24700 & ~w24701;
assign w24703 = ~w8240 & w24694;
assign w24704 = ~pi0799 & ~w24675;
assign w24705 = ~w24703 & ~w24704;
assign w24706 = w1223 & w24322;
assign w24707 = ~w3195 & w24706;
assign w24708 = ~w24676 & ~w24706;
assign w24709 = ~pi0800 & w24708;
assign w24710 = ~w24707 & ~w24709;
assign w24711 = ~w40134 & w24706;
assign w24712 = ~pi0801 & w24708;
assign w24713 = ~w24711 & ~w24712;
assign w24714 = ~w6413 & w24706;
assign w24715 = ~pi0802 & w24708;
assign w24716 = ~w24714 & ~w24715;
assign w24717 = ~w5320 & w24706;
assign w24718 = ~pi0803 & w24708;
assign w24719 = ~w24717 & ~w24718;
assign w24720 = ~pi0804 & w24708;
assign w24721 = w24684 & w24706;
assign w24722 = ~w24720 & ~w24721;
assign w24723 = ~pi0805 & w24708;
assign w24724 = w24691 & w24706;
assign w24725 = ~w24723 & ~w24724;
assign w24726 = pi3411 & ~w341;
assign w24727 = ~pi0806 & ~w24658;
assign w24728 = ~pi0856 & w24658;
assign w24729 = ~w24727 & ~w24728;
assign w24730 = w341 & w24729;
assign w24731 = ~w24726 & ~w24730;
assign w24732 = pi3406 & ~w341;
assign w24733 = ~pi0807 & ~w24658;
assign w24734 = ~pi0857 & w24658;
assign w24735 = ~w24733 & ~w24734;
assign w24736 = w341 & w24735;
assign w24737 = ~w24732 & ~w24736;
assign w24738 = pi3413 & ~w341;
assign w24739 = ~pi0808 & ~w24658;
assign w24740 = ~pi0858 & w24658;
assign w24741 = ~w24739 & ~w24740;
assign w24742 = w341 & w24741;
assign w24743 = ~w24738 & ~w24742;
assign w24744 = pi3405 & ~w341;
assign w24745 = ~pi0809 & ~w24658;
assign w24746 = ~pi0824 & w24658;
assign w24747 = ~w24745 & ~w24746;
assign w24748 = w341 & w24747;
assign w24749 = ~w24744 & ~w24748;
assign w24750 = pi3414 & ~w341;
assign w24751 = ~pi0810 & ~w24658;
assign w24752 = ~pi0823 & w24658;
assign w24753 = ~w24751 & ~w24752;
assign w24754 = w341 & w24753;
assign w24755 = ~w24750 & ~w24754;
assign w24756 = pi3404 & ~w341;
assign w24757 = ~pi0811 & ~w24658;
assign w24758 = ~pi0859 & w24658;
assign w24759 = ~w24757 & ~w24758;
assign w24760 = w341 & w24759;
assign w24761 = ~w24756 & ~w24760;
assign w24762 = pi3402 & ~w341;
assign w24763 = ~pi0812 & ~w24658;
assign w24764 = ~pi0730 & w24658;
assign w24765 = ~w24763 & ~w24764;
assign w24766 = w341 & w24765;
assign w24767 = ~w24762 & ~w24766;
assign w24768 = pi3403 & ~w341;
assign w24769 = ~pi0813 & ~w24658;
assign w24770 = ~pi0731 & w24658;
assign w24771 = ~w24769 & ~w24770;
assign w24772 = w341 & w24771;
assign w24773 = ~w24768 & ~w24772;
assign w24774 = pi3430 & ~w341;
assign w24775 = ~pi0814 & ~w24658;
assign w24776 = ~pi0853 & w24658;
assign w24777 = ~w24775 & ~w24776;
assign w24778 = w341 & w24777;
assign w24779 = ~w24774 & ~w24778;
assign w24780 = pi3421 & ~w341;
assign w24781 = ~pi0815 & ~w24658;
assign w24782 = ~pi0854 & w24658;
assign w24783 = ~w24781 & ~w24782;
assign w24784 = w341 & w24783;
assign w24785 = ~w24780 & ~w24784;
assign w24786 = pi3422 & ~w341;
assign w24787 = ~pi0816 & ~w24658;
assign w24788 = ~pi0785 & w24658;
assign w24789 = ~w24787 & ~w24788;
assign w24790 = w341 & w24789;
assign w24791 = ~w24786 & ~w24790;
assign w24792 = pi3401 & ~w341;
assign w24793 = ~pi0817 & ~w24658;
assign w24794 = ~pi0825 & w24658;
assign w24795 = ~w24793 & ~w24794;
assign w24796 = w341 & w24795;
assign w24797 = ~w24792 & ~w24796;
assign w24798 = pi3400 & ~w341;
assign w24799 = ~pi0818 & ~w24658;
assign w24800 = ~pi0938 & w24658;
assign w24801 = ~w24799 & ~w24800;
assign w24802 = w341 & w24801;
assign w24803 = ~w24798 & ~w24802;
assign w24804 = pi1935 & pi2056;
assign w24805 = pi1936 & w24804;
assign w24806 = w20669 & ~w24805;
assign w24807 = pi3428 & ~w20669;
assign w24808 = ~w24806 & ~w24807;
assign w24809 = pi2769 & w24808;
assign w24810 = ~w19039 & ~w24809;
assign w24811 = ~pi0609 & ~pi1771;
assign w24812 = ~pi3579 & w24811;
assign w24813 = ~w20669 & ~w24812;
assign w24814 = ~w24810 & w24813;
assign w24815 = pi0873 & w24814;
assign w24816 = pi0908 & w24815;
assign w24817 = pi0907 & w24816;
assign w24818 = pi0874 & w24817;
assign w24819 = pi0906 & w24818;
assign w24820 = pi0905 & w24819;
assign w24821 = pi0904 & w24820;
assign w24822 = pi0876 & w24821;
assign w24823 = pi0903 & w24822;
assign w24824 = pi0902 & w24823;
assign w24825 = pi0910 & w24824;
assign w24826 = pi0820 & w24825;
assign w24827 = pi0819 & w24826;
assign w24828 = pi3578 & pi3579;
assign w24829 = pi3467 & w24828;
assign w24830 = w1204 & w1265;
assign w24831 = w1225 & w1241;
assign w24832 = ~w24830 & ~w24831;
assign w24833 = w23839 & ~w24832;
assign w24834 = ~pi1033 & ~w24812;
assign w24835 = w24833 & w24834;
assign w24836 = ~w24829 & ~w24835;
assign w24837 = ~pi0819 & ~w24826;
assign w24838 = w24836 & ~w24837;
assign w24839 = ~w24827 & w24838;
assign w24840 = ~pi3579 & ~w1308;
assign w24841 = pi3447 & pi3579;
assign w24842 = ~w24836 & ~w24841;
assign w24843 = ~w24840 & w24842;
assign w24844 = ~w24839 & ~w24843;
assign w24845 = ~pi3579 & ~w5635;
assign w24846 = pi3463 & pi3579;
assign w24847 = ~w24845 & ~w24846;
assign w24848 = ~w24836 & w24847;
assign w24849 = ~pi0820 & ~w24825;
assign w24850 = ~w24826 & w24836;
assign w24851 = ~w24849 & w24850;
assign w24852 = ~w24848 & ~w24851;
assign w24853 = ~pi3008 & w24194;
assign w24854 = ~pi2973 & w24217;
assign w24855 = ~w24853 & ~w24854;
assign w24856 = pi0385 & w19516;
assign w24857 = ~pi3025 & w24196;
assign w24858 = ~w24856 & ~w24857;
assign w24859 = w24855 & w24858;
assign w24860 = ~pi3042 & w24236;
assign w24861 = ~pi1368 & w24189;
assign w24862 = ~w24860 & ~w24861;
assign w24863 = ~pi3001 & w24212;
assign w24864 = ~pi1678 & w24215;
assign w24865 = ~w24863 & ~w24864;
assign w24866 = w24862 & w24865;
assign w24867 = ~pi2818 & w24233;
assign w24868 = ~pi3032 & w24185;
assign w24869 = ~w24867 & ~w24868;
assign w24870 = pi0412 & w19957;
assign w24871 = ~pi3016 & w24210;
assign w24872 = ~w24870 & ~w24871;
assign w24873 = w24869 & w24872;
assign w24874 = w24866 & w24873;
assign w24875 = w24859 & w24874;
assign w24876 = w24179 & w24875;
assign w24877 = ~pi0821 & ~w24175;
assign w24878 = ~w24176 & w24877;
assign w24879 = pi0937 & w24225;
assign w24880 = ~pi0852 & w24176;
assign w24881 = ~w24174 & w24880;
assign w24882 = ~w24879 & ~w24881;
assign w24883 = ~w24878 & w24882;
assign w24884 = ~w24876 & w24883;
assign w24885 = ~pi2397 & w18313;
assign w24886 = pi0822 & ~w18329;
assign w24887 = ~w18330 & ~w18359;
assign w24888 = ~w24886 & w24887;
assign w24889 = ~pi1719 & w18359;
assign w24890 = ~w18313 & ~w24889;
assign w24891 = ~w24888 & w24890;
assign w24892 = ~w24885 & ~w24891;
assign w24893 = pi0823 & w24177;
assign w24894 = ~pi3266 & w19515;
assign w24895 = w24179 & ~w24894;
assign w24896 = pi0810 & w24249;
assign w24897 = pi0423 & w19957;
assign w24898 = ~w24896 & ~w24897;
assign w24899 = ~pi2792 & w24217;
assign w24900 = ~pi3081 & w24185;
assign w24901 = ~w24899 & ~w24900;
assign w24902 = ~pi3040 & w24236;
assign w24903 = ~pi3017 & w24196;
assign w24904 = ~w24902 & ~w24903;
assign w24905 = w24901 & w24904;
assign w24906 = w24898 & w24905;
assign w24907 = ~pi1700 & w24215;
assign w24908 = ~pi2899 & w24233;
assign w24909 = ~pi1364 & w24189;
assign w24910 = ~w24908 & ~w24909;
assign w24911 = ~w24907 & w24910;
assign w24912 = ~pi3002 & w24194;
assign w24913 = ~pi2994 & w24212;
assign w24914 = ~w24912 & ~w24913;
assign w24915 = ~pi3010 & w24210;
assign w24916 = pi0377 & w19516;
assign w24917 = ~w24915 & ~w24916;
assign w24918 = w24914 & w24917;
assign w24919 = w24911 & w24918;
assign w24920 = w24906 & w24919;
assign w24921 = w24895 & w24920;
assign w24922 = ~pi0824 & ~w24175;
assign w24923 = ~pi0859 & w24225;
assign w24924 = ~w24177 & ~w24923;
assign w24925 = ~w24922 & w24924;
assign w24926 = ~w24921 & w24925;
assign w24927 = ~w24893 & ~w24926;
assign w24928 = pi0376 & w19516;
assign w24929 = ~pi2815 & w24196;
assign w24930 = ~w24928 & ~w24929;
assign w24931 = ~pi3033 & w24217;
assign w24932 = ~pi1385 & w24189;
assign w24933 = ~w24931 & ~w24932;
assign w24934 = ~pi3026 & w24185;
assign w24935 = pi0422 & w19957;
assign w24936 = ~w24934 & ~w24935;
assign w24937 = w24933 & w24936;
assign w24938 = w24930 & w24937;
assign w24939 = ~pi3061 & w24236;
assign w24940 = ~pi3009 & w24210;
assign w24941 = pi0809 & w24249;
assign w24942 = ~w24940 & ~w24941;
assign w24943 = ~w24939 & w24942;
assign w24944 = ~pi2954 & w24212;
assign w24945 = ~pi1387 & w24215;
assign w24946 = ~w24944 & ~w24945;
assign w24947 = ~pi2880 & w24194;
assign w24948 = ~pi2775 & w24233;
assign w24949 = ~w24947 & ~w24948;
assign w24950 = w24946 & w24949;
assign w24951 = w24943 & w24950;
assign w24952 = w24938 & w24951;
assign w24953 = w24895 & w24952;
assign w24954 = pi0823 & pi3425;
assign w24955 = pi0858 & ~pi3425;
assign w24956 = w24176 & ~w24955;
assign w24957 = ~w24954 & w24956;
assign w24958 = ~pi0824 & w24177;
assign w24959 = ~w24957 & ~w24958;
assign w24960 = ~w24953 & w24959;
assign w24961 = pi0825 & w24177;
assign w24962 = pi0817 & w24249;
assign w24963 = ~pi3058 & w24185;
assign w24964 = ~w24962 & ~w24963;
assign w24965 = ~pi2972 & w24210;
assign w24966 = pi0418 & w19957;
assign w24967 = ~w24965 & ~w24966;
assign w24968 = w24964 & w24967;
assign w24969 = ~pi2857 & w24194;
assign w24970 = ~pi2887 & w24212;
assign w24971 = ~w24969 & ~w24970;
assign w24972 = ~pi3044 & w24236;
assign w24973 = ~pi2930 & w24233;
assign w24974 = ~w24972 & ~w24973;
assign w24975 = w24971 & w24974;
assign w24976 = w24968 & w24975;
assign w24977 = pi0565 & w24181;
assign w24978 = pi3551 & w24624;
assign w24979 = ~pi1005 & w24189;
assign w24980 = ~w24978 & ~w24979;
assign w24981 = ~w24977 & w24980;
assign w24982 = ~pi1073 & w24215;
assign w24983 = pi0371 & w19516;
assign w24984 = ~w24982 & ~w24983;
assign w24985 = ~pi2910 & w24196;
assign w24986 = ~pi3039 & w24217;
assign w24987 = ~w24985 & ~w24986;
assign w24988 = w24984 & w24987;
assign w24989 = w24981 & w24988;
assign w24990 = w24976 & w24989;
assign w24991 = w24612 & w24990;
assign w24992 = ~pi0785 & ~w24175;
assign w24993 = ~pi0855 & w24225;
assign w24994 = ~w24177 & ~w24993;
assign w24995 = ~w24992 & w24994;
assign w24996 = ~w24991 & w24995;
assign w24997 = ~w24961 & ~w24996;
assign w24998 = ~pi0866 & ~pi3120;
assign w24999 = ~w370 & ~w24998;
assign w25000 = ~w10688 & ~w24999;
assign w25001 = ~pi0826 & w25000;
assign w25002 = pi0866 & w40134;
assign w25003 = ~pi0866 & pi3120;
assign w25004 = pi0826 & ~pi3398;
assign w25005 = ~w2307 & ~w25004;
assign w25006 = w25003 & ~w25005;
assign w25007 = ~pi1411 & w10561;
assign w25008 = ~pi1593 & w10559;
assign w25009 = ~pi1621 & w10566;
assign w25010 = ~w25008 & ~w25009;
assign w25011 = ~w25007 & w25010;
assign w25012 = pi1041 & ~w25011;
assign w25013 = ~pi1042 & pi1507;
assign w25014 = pi1042 & pi1526;
assign w25015 = w24066 & ~w25014;
assign w25016 = ~w25013 & w25015;
assign w25017 = ~pi1041 & pi1489;
assign w25018 = pi1041 & pi1561;
assign w25019 = w10564 & ~w25018;
assign w25020 = ~w25017 & w25019;
assign w25021 = ~w25016 & ~w25020;
assign w25022 = ~w25012 & w25021;
assign w25023 = w24998 & ~w25022;
assign w25024 = ~w25006 & ~w25023;
assign w25025 = ~w25000 & w25024;
assign w25026 = ~w25002 & w25025;
assign w25027 = ~w25001 & ~w25026;
assign w25028 = ~pi0827 & w25000;
assign w25029 = pi0866 & w6413;
assign w25030 = ~pi3504 & pi3513;
assign w25031 = ~pi0827 & ~pi3513;
assign w25032 = w25003 & ~w25031;
assign w25033 = ~w25030 & w25032;
assign w25034 = ~pi1423 & w10559;
assign w25035 = pi1041 & ~w25034;
assign w25036 = ~pi1577 & w10566;
assign w25037 = ~pi1391 & w10564;
assign w25038 = ~pi1545 & w10561;
assign w25039 = ~w25037 & ~w25038;
assign w25040 = ~w25036 & w25039;
assign w25041 = w25035 & w25040;
assign w25042 = ~pi1421 & w10559;
assign w25043 = ~pi1041 & ~w25042;
assign w25044 = ~pi1508 & w10566;
assign w25045 = ~pi1490 & w10564;
assign w25046 = ~w25044 & ~w25045;
assign w25047 = w25043 & w25046;
assign w25048 = w24998 & ~w25047;
assign w25049 = ~w25041 & w25048;
assign w25050 = ~w25033 & ~w25049;
assign w25051 = ~w25000 & w25050;
assign w25052 = ~w25029 & w25051;
assign w25053 = ~w25028 & ~w25052;
assign w25054 = ~pi0828 & w25000;
assign w25055 = pi0866 & w5320;
assign w25056 = pi3514 & ~pi3517;
assign w25057 = ~pi0828 & ~pi3514;
assign w25058 = w25003 & ~w25057;
assign w25059 = ~w25056 & w25058;
assign w25060 = ~pi1578 & w10566;
assign w25061 = pi1041 & ~w25060;
assign w25062 = ~pi1546 & w10561;
assign w25063 = ~pi1399 & w10564;
assign w25064 = ~pi1401 & w10559;
assign w25065 = ~w25063 & ~w25064;
assign w25066 = ~w25062 & w25065;
assign w25067 = w25061 & w25066;
assign w25068 = ~pi1509 & w10566;
assign w25069 = ~pi1041 & ~w25068;
assign w25070 = ~pi1390 & w10564;
assign w25071 = ~pi1528 & w10559;
assign w25072 = ~w25070 & ~w25071;
assign w25073 = w25069 & w25072;
assign w25074 = w24998 & ~w25073;
assign w25075 = ~w25067 & w25074;
assign w25076 = ~w25059 & ~w25075;
assign w25077 = ~w25000 & w25076;
assign w25078 = ~w25055 & w25077;
assign w25079 = ~w25054 & ~w25078;
assign w25080 = ~pi0829 & w25000;
assign w25081 = pi0866 & w5914;
assign w25082 = ~pi1595 & w10559;
assign w25083 = pi1041 & ~w25082;
assign w25084 = ~pi1412 & w10561;
assign w25085 = ~pi1579 & w10566;
assign w25086 = ~pi1563 & w10564;
assign w25087 = ~w25085 & ~w25086;
assign w25088 = ~w25084 & w25087;
assign w25089 = w25083 & w25088;
assign w25090 = ~pi1510 & w10566;
assign w25091 = ~pi1041 & ~w25090;
assign w25092 = ~pi1492 & w10564;
assign w25093 = ~pi1529 & w10559;
assign w25094 = ~w25092 & ~w25093;
assign w25095 = w25091 & w25094;
assign w25096 = w24998 & ~w25095;
assign w25097 = ~w25089 & w25096;
assign w25098 = pi3508 & ~pi3509;
assign w25099 = ~pi0829 & ~pi3508;
assign w25100 = w25003 & ~w25099;
assign w25101 = ~w25098 & w25100;
assign w25102 = ~w25097 & ~w25101;
assign w25103 = ~w25000 & w25102;
assign w25104 = ~w25081 & w25103;
assign w25105 = ~w25080 & ~w25104;
assign w25106 = ~pi0830 & w25000;
assign w25107 = pi0866 & w4749;
assign w25108 = pi3510 & pi3511;
assign w25109 = pi0830 & ~pi3511;
assign w25110 = ~w25108 & ~w25109;
assign w25111 = w25003 & ~w25110;
assign w25112 = ~pi1611 & w10559;
assign w25113 = pi1041 & ~w25112;
assign w25114 = ~pi1565 & w10566;
assign w25115 = ~pi1548 & w10564;
assign w25116 = ~pi1530 & w10561;
assign w25117 = ~w25115 & ~w25116;
assign w25118 = ~w25114 & w25117;
assign w25119 = w25113 & w25118;
assign w25120 = ~pi1476 & w10564;
assign w25121 = ~pi1041 & ~w25120;
assign w25122 = ~pi1615 & w10559;
assign w25123 = ~pi1494 & w10566;
assign w25124 = ~w25122 & ~w25123;
assign w25125 = w25121 & w25124;
assign w25126 = w24998 & ~w25125;
assign w25127 = ~w25119 & w25126;
assign w25128 = ~w25111 & ~w25127;
assign w25129 = ~w25000 & w25128;
assign w25130 = ~w25107 & w25129;
assign w25131 = ~w25106 & ~w25130;
assign w25132 = ~pi0831 & w6684;
assign w25133 = ~w21994 & w24282;
assign w25134 = w24285 & w25133;
assign w25135 = ~w24288 & w25134;
assign w25136 = ~w25132 & ~w25135;
assign w25137 = ~pi0832 & w6684;
assign w25138 = w2230 & w24506;
assign w25139 = w24286 & w25138;
assign w25140 = ~w25137 & ~w25139;
assign w25141 = ~pi0833 & w6684;
assign w25142 = w25134 & w25138;
assign w25143 = ~w25141 & ~w25142;
assign w25144 = ~pi0834 & w6684;
assign w25145 = ~w21999 & w24284;
assign w25146 = w25133 & w25145;
assign w25147 = w25138 & w25146;
assign w25148 = ~w25144 & ~w25147;
assign w25149 = ~pi0835 & w6684;
assign w25150 = ~w24288 & w25146;
assign w25151 = ~w25149 & ~w25150;
assign w25152 = pi0836 & w343;
assign w25153 = w24115 & w24517;
assign w25154 = ~w25152 & ~w25153;
assign w25155 = pi0837 & w343;
assign w25156 = w24115 & w24521;
assign w25157 = ~w25155 & ~w25156;
assign w25158 = pi0838 & w343;
assign w25159 = ~w343 & w22304;
assign w25160 = ~w25158 & ~w25159;
assign w25161 = pi2986 & ~pi2990;
assign w25162 = ~w2893 & ~w25161;
assign w25163 = ~w902 & w25162;
assign w25164 = w156 & ~w25163;
assign w25165 = pi2990 & ~w2889;
assign w25166 = ~w7233 & ~w25165;
assign w25167 = w156 & ~w25166;
assign w25168 = ~w25161 & ~w25167;
assign w25169 = ~w25164 & ~w25168;
assign w25170 = pi0839 & ~w25169;
assign w25171 = pi3690 & w25167;
assign w25172 = ~w25170 & ~w25171;
assign w25173 = pi0840 & ~w25169;
assign w25174 = pi3689 & w25167;
assign w25175 = ~w25173 & ~w25174;
assign w25176 = pi0841 & ~w25169;
assign w25177 = pi3687 & w25167;
assign w25178 = ~w25176 & ~w25177;
assign w25179 = pi0842 & ~w25169;
assign w25180 = pi3685 & w25167;
assign w25181 = ~w25179 & ~w25180;
assign w25182 = pi0843 & ~w25169;
assign w25183 = pi3684 & w25167;
assign w25184 = ~w25182 & ~w25183;
assign w25185 = pi0844 & ~w25169;
assign w25186 = pi3683 & w25167;
assign w25187 = ~w25185 & ~w25186;
assign w25188 = w4141 & w24375;
assign w25189 = ~pi0845 & ~w24404;
assign w25190 = ~w24375 & ~w24405;
assign w25191 = ~w25189 & w25190;
assign w25192 = ~w25188 & ~w25191;
assign w25193 = ~w5914 & w24706;
assign w25194 = ~pi0846 & w24708;
assign w25195 = ~w25193 & ~w25194;
assign w25196 = pi0894 & w22495;
assign w25197 = pi0847 & ~w22504;
assign w25198 = ~w22505 & ~w25197;
assign w25199 = w22581 & w25198;
assign w25200 = ~w25196 & ~w25199;
assign w25201 = pi0968 & w22585;
assign w25202 = pi0848 & ~w22594;
assign w25203 = ~w22595 & w22671;
assign w25204 = ~w25202 & w25203;
assign w25205 = ~w25201 & ~w25204;
assign w25206 = ~pi2098 & w18313;
assign w25207 = pi0849 & w18326;
assign w25208 = ~w18327 & ~w18359;
assign w25209 = ~w25207 & w25208;
assign w25210 = ~pi1726 & w18359;
assign w25211 = ~w18313 & ~w25210;
assign w25212 = ~w25209 & w25211;
assign w25213 = ~w25206 & ~w25212;
assign w25214 = ~w4380 & w24706;
assign w25215 = ~pi0850 & w24708;
assign w25216 = ~w25214 & ~w25215;
assign w25217 = ~pi1698 & w24215;
assign w25218 = pi0409 & w19957;
assign w25219 = ~w25217 & ~w25218;
assign w25220 = ~pi1381 & w24189;
assign w25221 = ~pi3060 & w24185;
assign w25222 = ~w25220 & ~w25221;
assign w25223 = w25219 & w25222;
assign w25224 = ~pi3036 & w24217;
assign w25225 = ~pi2971 & w24233;
assign w25226 = ~w25224 & ~w25225;
assign w25227 = ~pi2790 & w24196;
assign w25228 = ~pi2991 & w24210;
assign w25229 = ~w25227 & ~w25228;
assign w25230 = w25226 & w25229;
assign w25231 = ~pi2970 & w24236;
assign w25232 = ~pi2822 & w24194;
assign w25233 = ~w25231 & ~w25232;
assign w25234 = ~pi3067 & w24212;
assign w25235 = pi0382 & w19516;
assign w25236 = ~w25234 & ~w25235;
assign w25237 = w25233 & w25236;
assign w25238 = w25230 & w25237;
assign w25239 = w25223 & w25238;
assign w25240 = w24179 & w25239;
assign w25241 = pi0851 & ~w24176;
assign w25242 = ~pi0938 & ~pi3425;
assign w25243 = ~pi0860 & pi3425;
assign w25244 = w24176 & ~w25243;
assign w25245 = ~w25242 & w25244;
assign w25246 = ~w25241 & ~w25245;
assign w25247 = ~w24179 & w25246;
assign w25248 = ~w25240 & ~w25247;
assign w25249 = pi0411 & w19957;
assign w25250 = ~pi1679 & w24215;
assign w25251 = ~w25249 & ~w25250;
assign w25252 = ~pi2977 & w24210;
assign w25253 = ~pi2907 & w24212;
assign w25254 = ~w25252 & ~w25253;
assign w25255 = w25251 & w25254;
assign w25256 = ~pi3021 & w24196;
assign w25257 = ~pi2958 & w24233;
assign w25258 = ~w25256 & ~w25257;
assign w25259 = ~pi1105 & w24189;
assign w25260 = ~pi2838 & w24194;
assign w25261 = ~w25259 & ~w25260;
assign w25262 = w25258 & w25261;
assign w25263 = ~pi2811 & w24236;
assign w25264 = ~pi3028 & w24185;
assign w25265 = ~w25263 & ~w25264;
assign w25266 = pi0384 & w19516;
assign w25267 = ~pi3037 & w24217;
assign w25268 = ~w25266 & ~w25267;
assign w25269 = w25265 & w25268;
assign w25270 = w25262 & w25269;
assign w25271 = w25255 & w25270;
assign w25272 = w24179 & w25271;
assign w25273 = pi0821 & pi3425;
assign w25274 = pi0860 & ~pi3425;
assign w25275 = w24176 & ~w25274;
assign w25276 = ~w25273 & w25275;
assign w25277 = ~pi0852 & w24177;
assign w25278 = ~w25276 & ~w25277;
assign w25279 = ~w25272 & w25278;
assign w25280 = ~pi0854 & pi3425;
assign w25281 = ~pi3425 & ~pi3678;
assign w25282 = w24176 & ~w25281;
assign w25283 = ~w25280 & w25282;
assign w25284 = pi0853 & ~w24176;
assign w25285 = ~w25283 & ~w25284;
assign w25286 = ~w24179 & w25285;
assign w25287 = ~pi1074 & w24215;
assign w25288 = ~pi2902 & w24236;
assign w25289 = ~w25287 & ~w25288;
assign w25290 = ~pi1084 & w24189;
assign w25291 = pi0416 & w19957;
assign w25292 = ~w25290 & ~w25291;
assign w25293 = pi0379 & w19516;
assign w25294 = ~pi3013 & w24210;
assign w25295 = ~w25293 & ~w25294;
assign w25296 = w25292 & w25295;
assign w25297 = w25289 & w25296;
assign w25298 = ~pi3083 & w24185;
assign w25299 = ~pi3022 & w24196;
assign w25300 = ~w25298 & ~w25299;
assign w25301 = ~pi3255 & w24180;
assign w25302 = ~pi2813 & ~pi3246;
assign w25303 = ~pi3055 & pi3246;
assign w25304 = ~w25302 & ~w25303;
assign w25305 = w25301 & w25304;
assign w25306 = ~pi3082 & w24217;
assign w25307 = ~w25305 & ~w25306;
assign w25308 = w25300 & w25307;
assign w25309 = ~pi2996 & w24212;
assign w25310 = ~pi3005 & w24194;
assign w25311 = ~w25309 & ~w25310;
assign w25312 = pi0814 & w24249;
assign w25313 = ~pi3051 & w24233;
assign w25314 = ~w25312 & ~w25313;
assign w25315 = w25311 & w25314;
assign w25316 = w25308 & w25315;
assign w25317 = w25297 & w25316;
assign w25318 = w24612 & w25317;
assign w25319 = ~w25286 & ~w25318;
assign w25320 = ~pi1078 & w24189;
assign w25321 = ~pi2984 & w24210;
assign w25322 = ~w25320 & ~w25321;
assign w25323 = ~pi3029 & w24185;
assign w25324 = ~pi3052 & w24233;
assign w25325 = ~w25323 & ~w25324;
assign w25326 = w25322 & w25325;
assign w25327 = ~pi3038 & w24217;
assign w25328 = pi0417 & w19957;
assign w25329 = ~w25327 & ~w25328;
assign w25330 = ~pi1610 & w24215;
assign w25331 = pi0815 & w24249;
assign w25332 = ~w25330 & ~w25331;
assign w25333 = w25329 & w25332;
assign w25334 = w25326 & w25333;
assign w25335 = pi0380 & w19516;
assign w25336 = ~pi3188 & w24624;
assign w25337 = ~pi3145 & w24181;
assign w25338 = ~w25336 & ~w25337;
assign w25339 = ~w25335 & w25338;
assign w25340 = ~pi2858 & w24194;
assign w25341 = ~pi3043 & w24236;
assign w25342 = ~w25340 & ~w25341;
assign w25343 = ~pi2908 & w24212;
assign w25344 = ~pi2909 & w24196;
assign w25345 = ~w25343 & ~w25344;
assign w25346 = w25342 & w25345;
assign w25347 = w25339 & w25346;
assign w25348 = w25334 & w25347;
assign w25349 = w24612 & w25348;
assign w25350 = pi0785 & pi3425;
assign w25351 = pi0853 & ~pi3425;
assign w25352 = w24176 & ~w25351;
assign w25353 = ~w25350 & w25352;
assign w25354 = ~pi0854 & w24177;
assign w25355 = ~w25353 & ~w25354;
assign w25356 = ~w25349 & w25355;
assign w25357 = pi0855 & w24177;
assign w25358 = ~pi3007 & w24194;
assign w25359 = ~pi1604 & w24215;
assign w25360 = ~w25358 & ~w25359;
assign w25361 = pi0419 & w19957;
assign w25362 = ~pi3070 & w24185;
assign w25363 = ~w25361 & ~w25362;
assign w25364 = w25360 & w25363;
assign w25365 = ~pi2998 & w24212;
assign w25366 = ~pi3064 & w24217;
assign w25367 = ~w25365 & ~w25366;
assign w25368 = pi0372 & w19516;
assign w25369 = ~pi3015 & w24210;
assign w25370 = ~w25368 & ~w25369;
assign w25371 = w25367 & w25370;
assign w25372 = w25364 & w25371;
assign w25373 = pi2860 & ~pi3573;
assign w25374 = w24624 & ~w25373;
assign w25375 = pi3452 & w24181;
assign w25376 = ~pi3054 & w24233;
assign w25377 = ~w25375 & ~w25376;
assign w25378 = ~w25374 & w25377;
assign w25379 = ~pi2906 & w24196;
assign w25380 = ~pi2904 & w24236;
assign w25381 = ~w25379 & ~w25380;
assign w25382 = ~pi1077 & w24189;
assign w25383 = pi0788 & w24249;
assign w25384 = ~w25382 & ~w25383;
assign w25385 = w25381 & w25384;
assign w25386 = w25378 & w25385;
assign w25387 = w25372 & w25386;
assign w25388 = w24612 & w25387;
assign w25389 = ~pi0825 & ~w24175;
assign w25390 = ~pi0856 & w24225;
assign w25391 = ~w24177 & ~w25390;
assign w25392 = ~w25389 & w25391;
assign w25393 = ~w25388 & w25392;
assign w25394 = ~w25357 & ~w25393;
assign w25395 = pi0856 & w24177;
assign w25396 = ~pi3080 & w24233;
assign w25397 = ~pi2886 & w24210;
assign w25398 = ~w25396 & ~w25397;
assign w25399 = ~pi3071 & w24217;
assign w25400 = pi0806 & w24249;
assign w25401 = ~w25399 & ~w25400;
assign w25402 = w25398 & w25401;
assign w25403 = ~pi2885 & w24196;
assign w25404 = ~pi3030 & w24185;
assign w25405 = ~w25403 & ~w25404;
assign w25406 = pi0420 & w19957;
assign w25407 = ~pi1672 & w24215;
assign w25408 = ~w25406 & ~w25407;
assign w25409 = w25405 & w25408;
assign w25410 = w25402 & w25409;
assign w25411 = ~pi3200 & w24624;
assign w25412 = ~pi3641 & w24181;
assign w25413 = pi0373 & w19516;
assign w25414 = ~w25412 & ~w25413;
assign w25415 = ~w25411 & w25414;
assign w25416 = ~pi3094 & w24194;
assign w25417 = ~pi3045 & w24236;
assign w25418 = ~w25416 & ~w25417;
assign w25419 = ~pi1076 & w24189;
assign w25420 = ~pi2901 & w24212;
assign w25421 = ~w25419 & ~w25420;
assign w25422 = w25418 & w25421;
assign w25423 = w25415 & w25422;
assign w25424 = w25410 & w25423;
assign w25425 = w24612 & w25424;
assign w25426 = ~pi0855 & ~w24175;
assign w25427 = ~pi0857 & w24225;
assign w25428 = ~w24177 & ~w25427;
assign w25429 = ~w25426 & w25428;
assign w25430 = ~w25425 & w25429;
assign w25431 = ~w25395 & ~w25430;
assign w25432 = pi0857 & w24177;
assign w25433 = ~pi3078 & w24185;
assign w25434 = ~pi2959 & w24210;
assign w25435 = ~w25433 & ~w25434;
assign w25436 = ~pi1673 & w24215;
assign w25437 = ~pi2915 & w24233;
assign w25438 = ~w25436 & ~w25437;
assign w25439 = ~pi3023 & w24196;
assign w25440 = pi0374 & w19516;
assign w25441 = ~w25439 & ~w25440;
assign w25442 = w25438 & w25441;
assign w25443 = w25435 & w25442;
assign w25444 = ~pi2823 & w24217;
assign w25445 = ~pi3088 & w24236;
assign w25446 = ~pi1366 & w24189;
assign w25447 = ~w25445 & ~w25446;
assign w25448 = ~w25444 & w25447;
assign w25449 = ~pi3077 & w24194;
assign w25450 = pi0807 & w24249;
assign w25451 = ~w25449 & ~w25450;
assign w25452 = pi0421 & w19957;
assign w25453 = ~pi2999 & w24212;
assign w25454 = ~w25452 & ~w25453;
assign w25455 = w25451 & w25454;
assign w25456 = w25448 & w25455;
assign w25457 = w25443 & w25456;
assign w25458 = w24895 & w25457;
assign w25459 = ~pi0856 & ~w24175;
assign w25460 = ~pi0858 & w24225;
assign w25461 = ~w24177 & ~w25460;
assign w25462 = ~w25459 & w25461;
assign w25463 = ~w25458 & w25462;
assign w25464 = ~w25432 & ~w25463;
assign w25465 = ~pi0824 & pi3425;
assign w25466 = ~pi0857 & ~pi3425;
assign w25467 = w24176 & ~w25466;
assign w25468 = ~w25465 & w25467;
assign w25469 = pi0858 & ~w24176;
assign w25470 = ~w25468 & ~w25469;
assign w25471 = ~w24179 & w25470;
assign w25472 = ~pi2883 & w24217;
assign w25473 = ~pi3069 & w24233;
assign w25474 = ~w25472 & ~w25473;
assign w25475 = ~pi1004 & w24189;
assign w25476 = ~pi3085 & w24194;
assign w25477 = ~w25475 & ~w25476;
assign w25478 = ~pi2786 & w24210;
assign w25479 = ~pi3031 & w24185;
assign w25480 = ~w25478 & ~w25479;
assign w25481 = w25477 & w25480;
assign w25482 = w25474 & w25481;
assign w25483 = pi0405 & w19957;
assign w25484 = pi0375 & w19516;
assign w25485 = ~pi1003 & w24215;
assign w25486 = ~w25484 & ~w25485;
assign w25487 = ~w25483 & w25486;
assign w25488 = ~pi3000 & w24212;
assign w25489 = ~pi3046 & w24236;
assign w25490 = ~w25488 & ~w25489;
assign w25491 = pi0808 & w24249;
assign w25492 = ~pi3024 & w24196;
assign w25493 = ~w25491 & ~w25492;
assign w25494 = w25490 & w25493;
assign w25495 = w25487 & w25494;
assign w25496 = w25482 & w25495;
assign w25497 = w24895 & w25496;
assign w25498 = ~w25471 & ~w25497;
assign w25499 = ~w24176 & ~w24224;
assign w25500 = ~pi0823 & ~pi3425;
assign w25501 = ~pi0730 & pi3425;
assign w25502 = w24176 & ~w25501;
assign w25503 = ~w25500 & w25502;
assign w25504 = ~w25499 & ~w25503;
assign w25505 = ~pi2955 & w24212;
assign w25506 = ~pi3095 & w24210;
assign w25507 = ~w25505 & ~w25506;
assign w25508 = ~pi3048 & w24233;
assign w25509 = pi0424 & w19957;
assign w25510 = ~w25508 & ~w25509;
assign w25511 = ~pi1671 & w24215;
assign w25512 = ~pi3103 & w24236;
assign w25513 = ~w25511 & ~w25512;
assign w25514 = w25510 & w25513;
assign w25515 = w25507 & w25514;
assign w25516 = ~pi1365 & w24189;
assign w25517 = pi0378 & w19516;
assign w25518 = ~pi3066 & w24196;
assign w25519 = ~w25517 & ~w25518;
assign w25520 = ~w25516 & w25519;
assign w25521 = ~pi3087 & w24185;
assign w25522 = pi0811 & w24249;
assign w25523 = ~w25521 & ~w25522;
assign w25524 = ~pi3034 & w24217;
assign w25525 = ~pi3003 & w24194;
assign w25526 = ~w25524 & ~w25525;
assign w25527 = w25523 & w25526;
assign w25528 = w25520 & w25527;
assign w25529 = w25515 & w25528;
assign w25530 = w24895 & w25529;
assign w25531 = ~w25504 & ~w25530;
assign w25532 = pi0860 & w24177;
assign w25533 = ~pi2905 & w24217;
assign w25534 = ~pi1369 & w24189;
assign w25535 = ~w25533 & ~w25534;
assign w25536 = pi0383 & w19516;
assign w25537 = ~pi3073 & w24212;
assign w25538 = ~w25536 & ~w25537;
assign w25539 = w25535 & w25538;
assign w25540 = pi0410 & w19957;
assign w25541 = ~pi3041 & w24236;
assign w25542 = ~w25540 & ~w25541;
assign w25543 = ~pi2957 & w24233;
assign w25544 = ~pi1680 & w24215;
assign w25545 = ~w25543 & ~w25544;
assign w25546 = w25542 & w25545;
assign w25547 = ~pi2859 & w24185;
assign w25548 = ~pi3012 & w24210;
assign w25549 = ~w25547 & ~w25548;
assign w25550 = ~pi3020 & w24196;
assign w25551 = ~pi2839 & w24194;
assign w25552 = ~w25550 & ~w25551;
assign w25553 = w25549 & w25552;
assign w25554 = w25546 & w25553;
assign w25555 = w25539 & w25554;
assign w25556 = w24179 & w25555;
assign w25557 = ~pi0851 & ~w24175;
assign w25558 = ~pi0852 & w24225;
assign w25559 = ~w24177 & ~w25558;
assign w25560 = ~w25557 & w25559;
assign w25561 = ~w25556 & w25560;
assign w25562 = ~w25532 & ~w25561;
assign w25563 = w3195 & w24375;
assign w25564 = ~pi0861 & ~w24402;
assign w25565 = ~w24375 & ~w24403;
assign w25566 = ~w25564 & w25565;
assign w25567 = ~w25563 & ~w25566;
assign w25568 = w6177 & w24375;
assign w25569 = ~pi0862 & ~w24403;
assign w25570 = ~w24375 & ~w24404;
assign w25571 = ~w25569 & w25570;
assign w25572 = ~w25568 & ~w25571;
assign w25573 = ~pi2093 & w18313;
assign w25574 = pi0863 & w18331;
assign w25575 = ~w18332 & ~w18359;
assign w25576 = ~w25574 & w25575;
assign w25577 = ~pi1718 & w18359;
assign w25578 = ~w18313 & ~w25577;
assign w25579 = ~w25576 & w25578;
assign w25580 = ~w25573 & ~w25579;
assign w25581 = pi0864 & ~w25169;
assign w25582 = pi3686 & w25167;
assign w25583 = ~w25581 & ~w25582;
assign w25584 = pi0865 & ~w25169;
assign w25585 = pi3688 & w25167;
assign w25586 = ~w25584 & ~w25585;
assign w25587 = pi0866 & w6684;
assign w25588 = w24283 & w25145;
assign w25589 = w2230 & w25588;
assign w25590 = ~w24288 & w25589;
assign w25591 = ~w25587 & ~w25590;
assign w25592 = pi0867 & w6684;
assign w25593 = w21988 & w25146;
assign w25594 = ~w25592 & ~w25593;
assign w25595 = pi0868 & w25000;
assign w25596 = pi0866 & ~w4380;
assign w25597 = ~pi1616 & w10566;
assign w25598 = pi1041 & ~w25597;
assign w25599 = ~pi1413 & w10561;
assign w25600 = ~pi1562 & w10564;
assign w25601 = ~pi1594 & w10559;
assign w25602 = ~w25600 & ~w25601;
assign w25603 = ~w25599 & w25602;
assign w25604 = w25598 & w25603;
assign w25605 = ~pi1617 & w10566;
assign w25606 = ~pi1041 & ~w25605;
assign w25607 = ~pi1527 & w10559;
assign w25608 = ~pi1491 & w10564;
assign w25609 = ~w25607 & ~w25608;
assign w25610 = w25606 & w25609;
assign w25611 = ~pi3120 & ~w25610;
assign w25612 = ~w25604 & w25611;
assign w25613 = ~pi0868 & ~pi3516;
assign w25614 = pi3120 & ~w10005;
assign w25615 = ~w25613 & w25614;
assign w25616 = ~pi0866 & ~w25615;
assign w25617 = ~w25612 & w25616;
assign w25618 = ~w25000 & ~w25617;
assign w25619 = ~w25596 & w25618;
assign w25620 = ~w25595 & ~w25619;
assign w25621 = w4141 & w24324;
assign w25622 = pi0869 & ~w24327;
assign w25623 = ~w25621 & ~w25622;
assign w25624 = pi0870 & ~w24327;
assign w25625 = w1639 & ~w24341;
assign w25626 = w24327 & w25625;
assign w25627 = ~w25624 & ~w25626;
assign w25628 = w5053 & w24324;
assign w25629 = pi0871 & ~w24327;
assign w25630 = ~w25628 & ~w25629;
assign w25631 = w5635 & w24324;
assign w25632 = pi0872 & ~w24327;
assign w25633 = ~w25631 & ~w25632;
assign w25634 = ~pi3579 & ~w3711;
assign w25635 = pi3464 & pi3579;
assign w25636 = ~w25634 & ~w25635;
assign w25637 = ~w24836 & w25636;
assign w25638 = ~pi0873 & ~w24814;
assign w25639 = ~w24815 & ~w25638;
assign w25640 = w24836 & w25639;
assign w25641 = ~w25637 & ~w25640;
assign w25642 = ~pi3579 & ~w5320;
assign w25643 = pi3446 & pi3579;
assign w25644 = ~w25642 & ~w25643;
assign w25645 = ~w24836 & w25644;
assign w25646 = ~pi0874 & ~w24817;
assign w25647 = ~w24818 & ~w25646;
assign w25648 = w24836 & w25647;
assign w25649 = ~w25645 & ~w25648;
assign w25650 = pi3451 & ~w437;
assign w25651 = w798 & w25650;
assign w25652 = ~pi3451 & ~w2555;
assign w25653 = ~w2826 & w25652;
assign w25654 = ~w25651 & ~w25653;
assign w25655 = pi3427 & ~w25654;
assign w25656 = ~pi3579 & ~w3195;
assign w25657 = pi3477 & pi3579;
assign w25658 = ~w25656 & ~w25657;
assign w25659 = ~w24836 & w25658;
assign w25660 = ~pi0876 & ~w24821;
assign w25661 = ~w24822 & ~w25660;
assign w25662 = w24836 & w25661;
assign w25663 = ~w25659 & ~w25662;
assign w25664 = pi3395 & ~w25654;
assign w25665 = pi3424 & ~w25654;
assign w25666 = pi3429 & ~w25654;
assign w25667 = w3195 & w24332;
assign w25668 = pi0880 & w24337;
assign w25669 = ~w25667 & ~w25668;
assign w25670 = w40134 & w24332;
assign w25671 = pi0881 & w24337;
assign w25672 = ~w25670 & ~w25671;
assign w25673 = w6413 & w24332;
assign w25674 = pi0882 & w24337;
assign w25675 = ~w25673 & ~w25674;
assign w25676 = w4380 & w24332;
assign w25677 = pi0883 & w24337;
assign w25678 = ~w25676 & ~w25677;
assign w25679 = w5320 & w24332;
assign w25680 = pi0884 & w24337;
assign w25681 = ~w25679 & ~w25680;
assign w25682 = w5914 & w24332;
assign w25683 = pi0885 & w24337;
assign w25684 = ~w25682 & ~w25683;
assign w25685 = w8240 & ~w24341;
assign w25686 = ~w24337 & w25685;
assign w25687 = pi0886 & w24337;
assign w25688 = ~w25686 & ~w25687;
assign w25689 = w8081 & w24332;
assign w25690 = pi0887 & w24337;
assign w25691 = ~w25689 & ~w25690;
assign w25692 = ~w24337 & w25625;
assign w25693 = pi0888 & w24337;
assign w25694 = ~w25692 & ~w25693;
assign w25695 = w1308 & ~w24341;
assign w25696 = ~w24337 & w25695;
assign w25697 = pi0889 & w24337;
assign w25698 = ~w25696 & ~w25697;
assign w25699 = ~w8081 & w24335;
assign w25700 = ~pi0890 & ~w24335;
assign w25701 = ~w25699 & ~w25700;
assign w25702 = ~w5320 & w25699;
assign w25703 = ~pi0891 & ~w24335;
assign w25704 = ~w25702 & ~w25703;
assign w25705 = ~w5914 & w25699;
assign w25706 = ~pi0892 & ~w24335;
assign w25707 = ~w25705 & ~w25706;
assign w25708 = ~w8240 & w25699;
assign w25709 = ~pi0893 & ~w24335;
assign w25710 = ~w25708 & ~w25709;
assign w25711 = w6177 & w24324;
assign w25712 = pi0894 & ~w24327;
assign w25713 = ~w25711 & ~w25712;
assign w25714 = pi0895 & ~w24327;
assign w25715 = w24327 & w25685;
assign w25716 = ~w25714 & ~w25715;
assign w25717 = w8081 & w24324;
assign w25718 = pi0896 & ~w24327;
assign w25719 = ~w25717 & ~w25718;
assign w25720 = pi0897 & ~w24327;
assign w25721 = w24327 & w25695;
assign w25722 = ~w25720 & ~w25721;
assign w25723 = ~pi1868 & ~pi1896;
assign w25724 = ~pi1895 & w25723;
assign w25725 = ~pi1871 & w25724;
assign w25726 = ~pi1894 & w25725;
assign w25727 = ~pi1870 & w25726;
assign w25728 = ~pi1893 & w25727;
assign w25729 = ~pi1740 & w25728;
assign w25730 = ~pi1435 & w25729;
assign w25731 = ~pi1872 & w25730;
assign w25732 = ~pi1016 & w25731;
assign w25733 = ~pi1094 & w25732;
assign w25734 = ~pi1097 & w25733;
assign w25735 = ~pi1715 & w25734;
assign w25736 = ~pi0946 & w25735;
assign w25737 = pi0898 & ~w25736;
assign w25738 = pi1886 & pi1894;
assign w25739 = ~pi1094 & ~pi1892;
assign w25740 = ~w25738 & ~w25739;
assign w25741 = ~pi1871 & ~pi1887;
assign w25742 = pi0946 & pi1869;
assign w25743 = ~w25741 & ~w25742;
assign w25744 = w25740 & w25743;
assign w25745 = pi1740 & pi1884;
assign w25746 = pi1872 & pi1952;
assign w25747 = ~w25745 & ~w25746;
assign w25748 = ~pi1872 & ~pi1952;
assign w25749 = pi1871 & pi1887;
assign w25750 = ~w25748 & ~w25749;
assign w25751 = w25747 & w25750;
assign w25752 = w25744 & w25751;
assign w25753 = pi1885 & pi1893;
assign w25754 = ~pi1888 & ~pi1895;
assign w25755 = ~w25753 & ~w25754;
assign w25756 = pi0898 & pi1889;
assign w25757 = pi1016 & pi1891;
assign w25758 = ~w25756 & ~w25757;
assign w25759 = w25755 & w25758;
assign w25760 = pi1862 & pi1868;
assign w25761 = pi1873 & pi1896;
assign w25762 = ~w25760 & ~w25761;
assign w25763 = ~pi1740 & ~pi1884;
assign w25764 = ~pi1715 & ~pi1890;
assign w25765 = ~w25763 & ~w25764;
assign w25766 = w25762 & w25765;
assign w25767 = w25759 & w25766;
assign w25768 = w25752 & w25767;
assign w25769 = pi1870 & pi1920;
assign w25770 = ~pi1873 & ~pi1896;
assign w25771 = ~w25769 & ~w25770;
assign w25772 = ~pi1435 & ~pi1883;
assign w25773 = pi1888 & pi1895;
assign w25774 = ~w25772 & ~w25773;
assign w25775 = w25771 & w25774;
assign w25776 = ~pi1097 & pi1874;
assign w25777 = pi1097 & ~pi1874;
assign w25778 = ~w25776 & ~w25777;
assign w25779 = pi1435 & pi1883;
assign w25780 = ~pi0946 & ~pi1869;
assign w25781 = ~w25779 & ~w25780;
assign w25782 = ~w25778 & w25781;
assign w25783 = w25775 & w25782;
assign w25784 = ~pi1886 & ~pi1894;
assign w25785 = pi1715 & pi1890;
assign w25786 = ~w25784 & ~w25785;
assign w25787 = ~pi1870 & ~pi1920;
assign w25788 = ~pi0898 & ~pi1889;
assign w25789 = ~w25787 & ~w25788;
assign w25790 = w25786 & w25789;
assign w25791 = ~pi1016 & ~pi1891;
assign w25792 = ~pi1862 & ~pi1868;
assign w25793 = ~w25791 & ~w25792;
assign w25794 = pi1094 & pi1892;
assign w25795 = ~pi1885 & ~pi1893;
assign w25796 = ~w25794 & ~w25795;
assign w25797 = w25793 & w25796;
assign w25798 = w25790 & w25797;
assign w25799 = w25783 & w25798;
assign w25800 = w25768 & w25799;
assign w25801 = pi3647 & ~w25800;
assign w25802 = ~pi0898 & w25736;
assign w25803 = w25801 & ~w25802;
assign w25804 = ~w25737 & w25803;
assign w25805 = ~w5635 & w24672;
assign w25806 = ~pi0899 & w24677;
assign w25807 = ~w25805 & ~w25806;
assign w25808 = pi0900 & ~w24675;
assign w25809 = w4380 & w24694;
assign w25810 = ~w25808 & ~w25809;
assign w25811 = ~pi1876 & ~pi1912;
assign w25812 = ~pi1913 & w25811;
assign w25813 = ~pi1914 & w25812;
assign w25814 = ~pi1911 & w25813;
assign w25815 = ~pi1916 & w25814;
assign w25816 = ~pi1910 & w25815;
assign w25817 = ~pi1748 & w25816;
assign w25818 = ~pi1448 & w25817;
assign w25819 = ~pi1915 & w25818;
assign w25820 = ~pi1018 & w25819;
assign w25821 = ~pi1095 & w25820;
assign w25822 = ~pi1098 & w25821;
assign w25823 = ~pi1747 & w25822;
assign w25824 = ~pi0973 & w25823;
assign w25825 = pi0901 & ~w25824;
assign w25826 = pi1901 & pi1914;
assign w25827 = pi1900 & pi1911;
assign w25828 = ~w25826 & ~w25827;
assign w25829 = pi1018 & pi2051;
assign w25830 = ~pi1748 & ~pi2055;
assign w25831 = ~w25829 & ~w25830;
assign w25832 = w25828 & w25831;
assign w25833 = ~pi1902 & ~pi1913;
assign w25834 = pi1902 & pi1913;
assign w25835 = ~w25833 & ~w25834;
assign w25836 = ~pi0901 & ~pi1903;
assign w25837 = ~pi1747 & ~pi1905;
assign w25838 = ~w25836 & ~w25837;
assign w25839 = w25835 & w25838;
assign w25840 = w25832 & w25839;
assign w25841 = pi1916 & pi2054;
assign w25842 = pi1747 & pi1905;
assign w25843 = ~w25841 & ~w25842;
assign w25844 = pi1915 & pi2057;
assign w25845 = ~pi1900 & ~pi1911;
assign w25846 = ~w25844 & ~w25845;
assign w25847 = w25843 & w25846;
assign w25848 = ~pi0973 & ~pi1904;
assign w25849 = ~pi1876 & ~pi1907;
assign w25850 = ~w25848 & ~w25849;
assign w25851 = pi1448 & pi1898;
assign w25852 = ~pi1018 & ~pi2051;
assign w25853 = ~w25851 & ~w25852;
assign w25854 = w25850 & w25853;
assign w25855 = w25847 & w25854;
assign w25856 = w25840 & w25855;
assign w25857 = ~pi1912 & ~pi2052;
assign w25858 = pi1876 & pi1907;
assign w25859 = ~w25857 & ~w25858;
assign w25860 = ~pi1901 & ~pi1914;
assign w25861 = ~pi1916 & ~pi2054;
assign w25862 = ~w25860 & ~w25861;
assign w25863 = w25859 & w25862;
assign w25864 = ~pi1899 & pi1910;
assign w25865 = pi1899 & ~pi1910;
assign w25866 = ~w25864 & ~w25865;
assign w25867 = ~pi1098 & pi2053;
assign w25868 = pi1098 & ~pi2053;
assign w25869 = ~w25867 & ~w25868;
assign w25870 = ~w25866 & ~w25869;
assign w25871 = w25863 & w25870;
assign w25872 = ~pi1095 & ~pi1906;
assign w25873 = ~pi1448 & ~pi1898;
assign w25874 = ~w25872 & ~w25873;
assign w25875 = pi1748 & pi2055;
assign w25876 = pi1095 & pi1906;
assign w25877 = ~w25875 & ~w25876;
assign w25878 = w25874 & w25877;
assign w25879 = pi1912 & pi2052;
assign w25880 = pi0973 & pi1904;
assign w25881 = ~w25879 & ~w25880;
assign w25882 = ~pi1915 & ~pi2057;
assign w25883 = pi0901 & pi1903;
assign w25884 = ~w25882 & ~w25883;
assign w25885 = w25881 & w25884;
assign w25886 = w25878 & w25885;
assign w25887 = w25871 & w25886;
assign w25888 = w25856 & w25887;
assign w25889 = pi3635 & ~w25888;
assign w25890 = ~pi0901 & w25824;
assign w25891 = w25889 & ~w25890;
assign w25892 = ~w25825 & w25891;
assign w25893 = ~pi3579 & ~w4141;
assign w25894 = pi3445 & pi3579;
assign w25895 = ~w25893 & ~w25894;
assign w25896 = ~w24836 & w25895;
assign w25897 = ~pi0902 & ~w24823;
assign w25898 = ~w24824 & w24836;
assign w25899 = ~w25897 & w25898;
assign w25900 = ~w25896 & ~w25899;
assign w25901 = ~pi3579 & ~w6177;
assign w25902 = pi3474 & pi3579;
assign w25903 = ~w25901 & ~w25902;
assign w25904 = ~w24836 & w25903;
assign w25905 = ~pi0903 & ~w24822;
assign w25906 = ~w24823 & w24836;
assign w25907 = ~w25905 & w25906;
assign w25908 = ~w25904 & ~w25907;
assign w25909 = ~pi3579 & ~w40134;
assign w25910 = pi3476 & pi3579;
assign w25911 = ~w25909 & ~w25910;
assign w25912 = ~w24836 & w25911;
assign w25913 = ~pi0904 & ~w24820;
assign w25914 = ~w24821 & ~w25913;
assign w25915 = w24836 & w25914;
assign w25916 = ~w25912 & ~w25915;
assign w25917 = ~pi3579 & ~w6413;
assign w25918 = pi3475 & pi3579;
assign w25919 = ~w25917 & ~w25918;
assign w25920 = ~w24836 & w25919;
assign w25921 = ~pi0905 & ~w24819;
assign w25922 = ~w24820 & ~w25921;
assign w25923 = w24836 & w25922;
assign w25924 = ~w25920 & ~w25923;
assign w25925 = ~pi3579 & ~w4380;
assign w25926 = pi3470 & pi3579;
assign w25927 = ~w25925 & ~w25926;
assign w25928 = ~w24836 & w25927;
assign w25929 = ~pi0906 & ~w24818;
assign w25930 = ~w24819 & ~w25929;
assign w25931 = w24836 & w25930;
assign w25932 = ~w25928 & ~w25931;
assign w25933 = ~pi3579 & ~w5914;
assign w25934 = pi3462 & pi3579;
assign w25935 = ~w25933 & ~w25934;
assign w25936 = ~w24836 & w25935;
assign w25937 = ~pi0907 & ~w24816;
assign w25938 = ~w24817 & ~w25937;
assign w25939 = w24836 & w25938;
assign w25940 = ~w25936 & ~w25939;
assign w25941 = ~pi3579 & ~w4749;
assign w25942 = pi3468 & pi3579;
assign w25943 = ~w25941 & ~w25942;
assign w25944 = ~w24836 & w25943;
assign w25945 = ~pi0908 & ~w24815;
assign w25946 = ~w24816 & ~w25945;
assign w25947 = w24836 & w25946;
assign w25948 = ~w25944 & ~w25947;
assign w25949 = ~pi3579 & ~w1639;
assign w25950 = pi3466 & pi3579;
assign w25951 = ~w24836 & ~w25950;
assign w25952 = ~w25949 & w25951;
assign w25953 = ~pi0909 & ~w24827;
assign w25954 = pi0909 & w24827;
assign w25955 = w24836 & ~w25954;
assign w25956 = ~w25953 & w25955;
assign w25957 = ~w25952 & ~w25956;
assign w25958 = ~pi3579 & ~w5053;
assign w25959 = pi3448 & pi3579;
assign w25960 = ~w25958 & ~w25959;
assign w25961 = ~w24836 & w25960;
assign w25962 = ~pi0910 & ~w24824;
assign w25963 = ~w24825 & w24836;
assign w25964 = ~w25962 & w25963;
assign w25965 = ~w25961 & ~w25964;
assign w25966 = ~pi1075 & w24189;
assign w25967 = ~pi0427 & w19957;
assign w25968 = ~w25966 & ~w25967;
assign w25969 = pi0393 & w19516;
assign w25970 = ~pi1670 & w24215;
assign w25971 = ~w25969 & ~w25970;
assign w25972 = w25968 & w25971;
assign w25973 = w24179 & ~w25972;
assign w25974 = pi0911 & ~w24176;
assign w25975 = pi1052 & w24176;
assign w25976 = ~w25974 & ~w25975;
assign w25977 = ~w24175 & w25976;
assign w25978 = ~w25973 & ~w25977;
assign w25979 = pi1598 & pi3293;
assign w25980 = w24056 & ~w25979;
assign w25981 = pi3293 & ~w9286;
assign w25982 = w25980 & ~w25981;
assign w25983 = pi1597 & pi3293;
assign w25984 = w25982 & ~w25983;
assign w25985 = pi2017 & pi3293;
assign w25986 = w25984 & ~w25985;
assign w25987 = pi2474 & pi3293;
assign w25988 = w25986 & ~w25987;
assign w25989 = pi0912 & ~w25988;
assign w25990 = ~w24052 & ~w25989;
assign w25991 = pi1007 & w4141;
assign w25992 = ~pi1482 & w10564;
assign w25993 = ~pi1500 & w10566;
assign w25994 = ~pi1463 & w10559;
assign w25995 = ~w25993 & ~w25994;
assign w25996 = ~w25992 & w25995;
assign w25997 = ~pi1041 & ~w25996;
assign w25998 = pi1536 & w10561;
assign w25999 = pi1041 & ~w25998;
assign w26000 = pi1571 & w10566;
assign w26001 = pi1464 & w10559;
assign w26002 = pi1408 & w10564;
assign w26003 = ~w26001 & ~w26002;
assign w26004 = ~w26000 & w26003;
assign w26005 = w25999 & w26004;
assign w26006 = ~w25997 & ~w26005;
assign w26007 = ~pi1007 & ~w26006;
assign w26008 = w24052 & ~w26007;
assign w26009 = ~w25991 & w26008;
assign w26010 = ~w25990 & ~w26009;
assign w26011 = pi0913 & ~w25986;
assign w26012 = ~w24052 & w26011;
assign w26013 = pi1007 & ~w6177;
assign w26014 = ~pi1554 & w10564;
assign w26015 = ~pi1537 & w10561;
assign w26016 = ~pi1586 & w10559;
assign w26017 = ~w26015 & ~w26016;
assign w26018 = ~w26014 & w26017;
assign w26019 = pi1041 & ~w26018;
assign w26020 = pi1041 & pi1618;
assign w26021 = ~pi1041 & pi1627;
assign w26022 = w10566 & ~w26021;
assign w26023 = ~w26020 & w26022;
assign w26024 = ~pi1093 & pi1483;
assign w26025 = pi1093 & pi1518;
assign w26026 = w17569 & ~w26025;
assign w26027 = ~w26024 & w26026;
assign w26028 = ~pi1007 & ~w26027;
assign w26029 = ~w26023 & w26028;
assign w26030 = ~w26019 & w26029;
assign w26031 = w24052 & ~w26030;
assign w26032 = ~w26013 & w26031;
assign w26033 = ~w26012 & ~w26032;
assign w26034 = pi0914 & ~w25984;
assign w26035 = ~w24052 & w26034;
assign w26036 = pi1007 & ~w3195;
assign w26037 = pi1404 & w10564;
assign w26038 = pi1475 & w10559;
assign w26039 = ~w26037 & ~w26038;
assign w26040 = pi1572 & w10566;
assign w26041 = pi1538 & w10561;
assign w26042 = ~w26040 & ~w26041;
assign w26043 = w26039 & w26042;
assign w26044 = pi1041 & ~w26043;
assign w26045 = ~pi1400 & w10564;
assign w26046 = ~pi1041 & ~w26045;
assign w26047 = ~pi1519 & w10559;
assign w26048 = ~pi1501 & w10566;
assign w26049 = ~w26047 & ~w26048;
assign w26050 = w26046 & w26049;
assign w26051 = ~w26044 & ~w26050;
assign w26052 = ~pi1007 & ~w26051;
assign w26053 = w24052 & ~w26052;
assign w26054 = ~w26036 & w26053;
assign w26055 = ~w26035 & ~w26054;
assign w26056 = pi0915 & ~w25982;
assign w26057 = ~w24052 & w26056;
assign w26058 = pi1007 & ~w40134;
assign w26059 = ~pi1520 & w10559;
assign w26060 = ~pi1502 & w10566;
assign w26061 = ~pi1484 & w10564;
assign w26062 = ~w26060 & ~w26061;
assign w26063 = ~w26059 & w26062;
assign w26064 = ~pi1041 & ~w26063;
assign w26065 = pi1555 & w10564;
assign w26066 = pi1041 & ~w26065;
assign w26067 = pi1628 & w10566;
assign w26068 = pi1587 & w10559;
assign w26069 = pi1416 & w10561;
assign w26070 = ~w26068 & ~w26069;
assign w26071 = ~w26067 & w26070;
assign w26072 = w26066 & w26071;
assign w26073 = ~pi1007 & ~w26072;
assign w26074 = ~w26064 & w26073;
assign w26075 = w24052 & ~w26074;
assign w26076 = ~w26058 & w26075;
assign w26077 = ~w26057 & ~w26076;
assign w26078 = pi2019 & pi3293;
assign w26079 = w25980 & ~w26078;
assign w26080 = pi0916 & ~w26079;
assign w26081 = ~w24052 & w26080;
assign w26082 = pi1007 & ~w6413;
assign w26083 = ~pi1395 & w24066;
assign w26084 = ~pi1093 & pi1556;
assign w26085 = pi1093 & pi1466;
assign w26086 = pi1041 & ~w26085;
assign w26087 = ~w26084 & w26086;
assign w26088 = ~w26083 & ~w26087;
assign w26089 = pi1042 & ~w26088;
assign w26090 = ~pi1503 & w10566;
assign w26091 = ~pi1398 & w10564;
assign w26092 = ~w26090 & ~w26091;
assign w26093 = ~pi1041 & ~w26092;
assign w26094 = pi1093 & pi1573;
assign w26095 = pi1041 & ~pi1042;
assign w26096 = ~pi1093 & pi1539;
assign w26097 = w26095 & ~w26096;
assign w26098 = ~w26094 & w26097;
assign w26099 = ~pi1007 & ~w26098;
assign w26100 = ~w26093 & w26099;
assign w26101 = ~w26089 & w26100;
assign w26102 = w24052 & ~w26101;
assign w26103 = ~w26082 & w26102;
assign w26104 = ~w26081 & ~w26103;
assign w26105 = pi0917 & ~w25980;
assign w26106 = ~w24052 & ~w26105;
assign w26107 = pi1007 & w4380;
assign w26108 = ~pi1397 & w10564;
assign w26109 = ~pi1504 & w10566;
assign w26110 = ~pi1522 & w10559;
assign w26111 = ~w26109 & ~w26110;
assign w26112 = ~w26108 & w26111;
assign w26113 = ~pi1041 & ~w26112;
assign w26114 = pi1541 & w10561;
assign w26115 = pi1041 & ~w26114;
assign w26116 = pi1589 & w10559;
assign w26117 = pi1574 & w10566;
assign w26118 = pi1405 & w10564;
assign w26119 = ~w26117 & ~w26118;
assign w26120 = ~w26116 & w26119;
assign w26121 = w26115 & w26120;
assign w26122 = ~w26113 & ~w26121;
assign w26123 = ~pi1007 & ~w26122;
assign w26124 = w24052 & ~w26123;
assign w26125 = ~w26107 & w26124;
assign w26126 = ~w26106 & ~w26125;
assign w26127 = pi0918 & ~w24054;
assign w26128 = ~w24052 & w26127;
assign w26129 = pi1007 & ~w5914;
assign w26130 = ~pi1393 & w10559;
assign w26131 = ~pi1542 & w10561;
assign w26132 = ~pi1559 & w10564;
assign w26133 = ~w26131 & ~w26132;
assign w26134 = ~w26130 & w26133;
assign w26135 = pi1041 & ~w26134;
assign w26136 = ~pi1041 & pi1505;
assign w26137 = pi1041 & pi1575;
assign w26138 = w10566 & ~w26137;
assign w26139 = ~w26136 & w26138;
assign w26140 = pi1093 & pi1419;
assign w26141 = ~pi1093 & pi1487;
assign w26142 = w17569 & ~w26141;
assign w26143 = ~w26140 & w26142;
assign w26144 = ~pi1007 & ~w26143;
assign w26145 = ~w26139 & w26144;
assign w26146 = ~w26135 & w26145;
assign w26147 = w24052 & ~w26146;
assign w26148 = ~w26129 & w26147;
assign w26149 = ~w26128 & ~w26148;
assign w26150 = pi0919 & pi1330;
assign w26151 = pi3293 & w26150;
assign w26152 = w24049 & w26151;
assign w26153 = pi1007 & w4749;
assign w26154 = ~pi1591 & w10559;
assign w26155 = pi1041 & ~w26154;
assign w26156 = ~pi1560 & w10564;
assign w26157 = ~pi1543 & w10561;
assign w26158 = ~pi1623 & w10566;
assign w26159 = ~w26157 & ~w26158;
assign w26160 = ~w26156 & w26159;
assign w26161 = w26155 & w26160;
assign w26162 = ~pi1488 & w10564;
assign w26163 = ~pi1041 & ~w26162;
assign w26164 = ~pi1524 & w10559;
assign w26165 = ~pi1622 & w10566;
assign w26166 = ~w26164 & ~w26165;
assign w26167 = w26163 & w26166;
assign w26168 = ~pi1007 & ~w26167;
assign w26169 = ~w26161 & w26168;
assign w26170 = ~w24051 & ~w26169;
assign w26171 = ~w26153 & w26170;
assign w26172 = ~pi0919 & w24051;
assign w26173 = ~w24049 & ~w26172;
assign w26174 = ~w26171 & w26173;
assign w26175 = ~w26152 & ~w26174;
assign w26176 = ~pi0920 & w6684;
assign w26177 = w21981 & w24503;
assign w26178 = ~w24288 & w24502;
assign w26179 = w26177 & w26178;
assign w26180 = ~w26176 & ~w26179;
assign w26181 = ~pi0921 & w6684;
assign w26182 = w24506 & w25589;
assign w26183 = ~w26181 & ~w26182;
assign w26184 = ~pi3252 & w896;
assign w26185 = pi0445 & w26184;
assign w26186 = ~pi3252 & ~w25166;
assign w26187 = pi0440 & w26186;
assign w26188 = ~pi0922 & ~w26186;
assign w26189 = ~pi3252 & ~w25163;
assign w26190 = ~w26188 & ~w26189;
assign w26191 = ~w26187 & w26190;
assign w26192 = ~pi0453 & w26189;
assign w26193 = ~w26184 & ~w26192;
assign w26194 = ~w26191 & w26193;
assign w26195 = ~w26185 & ~w26194;
assign w26196 = ~pi0446 & w26184;
assign w26197 = pi0923 & ~w26186;
assign w26198 = ~pi0441 & w26186;
assign w26199 = ~w26189 & ~w26198;
assign w26200 = ~w26197 & w26199;
assign w26201 = pi0454 & w26189;
assign w26202 = ~w26184 & ~w26201;
assign w26203 = ~w26200 & w26202;
assign w26204 = ~w26196 & ~w26203;
assign w26205 = ~pi0447 & w26184;
assign w26206 = pi0924 & ~w26186;
assign w26207 = ~pi0442 & w26186;
assign w26208 = ~w26189 & ~w26207;
assign w26209 = ~w26206 & w26208;
assign w26210 = pi0461 & w26189;
assign w26211 = ~w26184 & ~w26210;
assign w26212 = ~w26209 & w26211;
assign w26213 = ~w26205 & ~w26212;
assign w26214 = ~pi0450 & w26184;
assign w26215 = pi0925 & ~w26186;
assign w26216 = ~pi0444 & w26186;
assign w26217 = ~w26189 & ~w26216;
assign w26218 = ~w26215 & w26217;
assign w26219 = pi0456 & w26189;
assign w26220 = ~w26184 & ~w26219;
assign w26221 = ~w26218 & w26220;
assign w26222 = ~w26214 & ~w26221;
assign w26223 = pi0451 & w26184;
assign w26224 = pi0459 & w26186;
assign w26225 = ~pi0926 & ~w26186;
assign w26226 = ~w26189 & ~w26225;
assign w26227 = ~w26224 & w26226;
assign w26228 = ~pi0457 & w26189;
assign w26229 = ~w26184 & ~w26228;
assign w26230 = ~w26227 & w26229;
assign w26231 = ~w26223 & ~w26230;
assign w26232 = ~pi0462 & w26184;
assign w26233 = pi0927 & ~w26186;
assign w26234 = ~pi0449 & w26186;
assign w26235 = ~w26189 & ~w26234;
assign w26236 = ~w26233 & w26235;
assign w26237 = pi0438 & w26189;
assign w26238 = ~w26184 & ~w26237;
assign w26239 = ~w26236 & w26238;
assign w26240 = ~w26232 & ~w26239;
assign w26241 = w6177 & w23862;
assign w26242 = ~pi0928 & ~w23872;
assign w26243 = ~w23862 & ~w23873;
assign w26244 = ~w26242 & w26243;
assign w26245 = ~w26241 & ~w26244;
assign w26246 = w1639 & w23862;
assign w26247 = pi0929 & w23877;
assign w26248 = ~pi0929 & ~w23877;
assign w26249 = ~w23862 & ~w26248;
assign w26250 = ~w26247 & w26249;
assign w26251 = ~w26246 & ~w26250;
assign w26252 = w5635 & w23862;
assign w26253 = ~pi0930 & ~w23875;
assign w26254 = ~w23862 & ~w23876;
assign w26255 = ~w26253 & w26254;
assign w26256 = ~w26252 & ~w26255;
assign w26257 = pi0748 & w22495;
assign w26258 = pi0931 & ~pi3647;
assign w26259 = ~w22497 & ~w26258;
assign w26260 = w22581 & w26259;
assign w26261 = ~w26257 & ~w26260;
assign w26262 = pi0743 & w22495;
assign w26263 = pi0932 & ~w22502;
assign w26264 = ~w22503 & ~w26263;
assign w26265 = w22581 & w26264;
assign w26266 = ~w26262 & ~w26265;
assign w26267 = pi0805 & w22585;
assign w26268 = pi0933 & ~pi3635;
assign w26269 = ~w22587 & ~w26268;
assign w26270 = w22671 & w26269;
assign w26271 = ~w26267 & ~w26270;
assign w26272 = pi0801 & w22585;
assign w26273 = pi0934 & ~w22592;
assign w26274 = ~w22593 & ~w26273;
assign w26275 = w22671 & w26274;
assign w26276 = ~w26272 & ~w26275;
assign w26277 = pi0800 & w22585;
assign w26278 = pi0935 & ~w22593;
assign w26279 = ~w22594 & ~w26278;
assign w26280 = w22671 & w26279;
assign w26281 = ~w26277 & ~w26280;
assign w26282 = pi3568 & w0;
assign w26283 = pi1380 & pi1668;
assign w26284 = pi1788 & w26283;
assign w26285 = pi1695 & pi2416;
assign w26286 = pi1081 & pi1379;
assign w26287 = w26285 & w26286;
assign w26288 = w26284 & w26287;
assign w26289 = pi3681 & w26288;
assign w26290 = ~pi1695 & ~pi2416;
assign w26291 = ~pi3681 & w26290;
assign w26292 = ~pi1081 & ~pi1379;
assign w26293 = ~pi1380 & ~pi1668;
assign w26294 = ~pi1788 & w26293;
assign w26295 = w26292 & w26294;
assign w26296 = w26291 & w26295;
assign w26297 = ~w26289 & ~w26296;
assign w26298 = ~pi2510 & ~pi2824;
assign w26299 = ~pi3247 & w26298;
assign w26300 = ~pi3290 & w26299;
assign w26301 = pi1908 & pi1917;
assign w26302 = ~pi1851 & w26301;
assign w26303 = w26300 & w26302;
assign w26304 = ~w26297 & w26303;
assign w26305 = ~pi1006 & ~w26301;
assign w26306 = ~pi0936 & ~w26305;
assign w26307 = ~w26304 & w26306;
assign w26308 = ~pi3583 & ~w26307;
assign w26309 = ~pi0937 & w24177;
assign w26310 = ~pi3502 & pi3506;
assign w26311 = ~w24174 & w26310;
assign w26312 = ~pi3677 & ~w26311;
assign w26313 = pi0386 & w19516;
assign w26314 = ~pi1699 & w24215;
assign w26315 = ~w26313 & ~w26314;
assign w26316 = ~pi2882 & w24233;
assign w26317 = ~pi1079 & w24189;
assign w26318 = ~w26316 & ~w26317;
assign w26319 = pi0413 & w19957;
assign w26320 = ~pi3047 & w24236;
assign w26321 = ~w26319 & ~w26320;
assign w26322 = w26318 & w26321;
assign w26323 = w26315 & w26322;
assign w26324 = ~w26312 & w26323;
assign w26325 = pi1045 & w24225;
assign w26326 = ~w24177 & ~w26325;
assign w26327 = ~w24877 & w26326;
assign w26328 = ~w26324 & w26327;
assign w26329 = ~w26309 & ~w26328;
assign w26330 = ~pi1669 & w24215;
assign w26331 = ~pi3019 & w24196;
assign w26332 = ~w26330 & ~w26331;
assign w26333 = ~pi2903 & w24217;
assign w26334 = ~pi2791 & w24236;
assign w26335 = ~w26333 & ~w26334;
assign w26336 = ~pi3062 & w24185;
assign w26337 = ~pi3072 & w24212;
assign w26338 = ~w26336 & ~w26337;
assign w26339 = w26335 & w26338;
assign w26340 = w26332 & w26339;
assign w26341 = ~pi2762 & w24250;
assign w26342 = pi0818 & w24249;
assign w26343 = ~w26341 & ~w26342;
assign w26344 = pi0392 & w19516;
assign w26345 = ~pi3108 & w24210;
assign w26346 = ~w26344 & ~w26345;
assign w26347 = w26343 & w26346;
assign w26348 = ~pi1362 & w24189;
assign w26349 = ~pi2821 & w24194;
assign w26350 = ~w26348 & ~w26349;
assign w26351 = pi0426 & w19957;
assign w26352 = ~pi3110 & w24233;
assign w26353 = ~w26351 & ~w26352;
assign w26354 = w26350 & w26353;
assign w26355 = w26347 & w26354;
assign w26356 = w26340 & w26355;
assign w26357 = w24182 & w26356;
assign w26358 = pi0851 & pi3425;
assign w26359 = pi0731 & ~pi3425;
assign w26360 = w24176 & ~w26359;
assign w26361 = ~w26358 & w26360;
assign w26362 = ~pi0938 & w24177;
assign w26363 = ~w26361 & ~w26362;
assign w26364 = ~w26357 & w26363;
assign w26365 = pi3410 & ~pi3416;
assign w26366 = w7 & ~w26365;
assign w26367 = pi3330 & ~pi3392;
assign w26368 = pi3394 & w26367;
assign w26369 = ~pi3382 & pi3410;
assign w26370 = ~w26368 & w26369;
assign w26371 = ~pi3416 & w26370;
assign w26372 = ~pi0939 & ~w26370;
assign w26373 = w25373 & ~w26372;
assign w26374 = ~w26371 & w26373;
assign w26375 = ~w23822 & w26374;
assign w26376 = pi0742 & w22495;
assign w26377 = pi0940 & ~w22503;
assign w26378 = ~w22504 & ~w26377;
assign w26379 = w22581 & w26378;
assign w26380 = ~w26376 & ~w26379;
assign w26381 = ~w6177 & w24672;
assign w26382 = ~pi0941 & w24677;
assign w26383 = ~w26381 & ~w26382;
assign w26384 = ~pi0452 & w26184;
assign w26385 = pi0942 & ~w26186;
assign w26386 = ~pi0460 & w26186;
assign w26387 = ~w26189 & ~w26386;
assign w26388 = ~w26385 & w26387;
assign w26389 = pi0439 & w26189;
assign w26390 = ~w26184 & ~w26389;
assign w26391 = ~w26388 & w26390;
assign w26392 = ~w26384 & ~w26391;
assign w26393 = ~pi0448 & w26184;
assign w26394 = pi0943 & ~w26186;
assign w26395 = ~pi0443 & w26186;
assign w26396 = ~w26189 & ~w26395;
assign w26397 = ~w26394 & w26396;
assign w26398 = pi0455 & w26189;
assign w26399 = ~w26184 & ~w26398;
assign w26400 = ~w26397 & w26399;
assign w26401 = ~w26393 & ~w26400;
assign w26402 = ~pi0944 & w6684;
assign w26403 = w6682 & ~w21994;
assign w26404 = w26177 & w26403;
assign w26405 = w21988 & w26404;
assign w26406 = ~w26402 & ~w26405;
assign w26407 = ~pi0945 & w6684;
assign w26408 = w24504 & w26403;
assign w26409 = w24506 & w26408;
assign w26410 = ~w26407 & ~w26409;
assign w26411 = pi0946 & ~w25735;
assign w26412 = ~w25736 & w25801;
assign w26413 = ~w26411 & w26412;
assign w26414 = pi0947 & ~w24335;
assign w26415 = w1639 & w24335;
assign w26416 = ~w26414 & ~w26415;
assign w26417 = pi0948 & ~w24335;
assign w26418 = w3195 & w25699;
assign w26419 = ~w26417 & ~w26418;
assign w26420 = pi0949 & ~w24335;
assign w26421 = w40134 & w25699;
assign w26422 = ~w26420 & ~w26421;
assign w26423 = pi0950 & ~w24335;
assign w26424 = w6413 & w25699;
assign w26425 = ~w26423 & ~w26424;
assign w26426 = pi0951 & ~w24335;
assign w26427 = w4380 & w25699;
assign w26428 = ~w26426 & ~w26427;
assign w26429 = pi0952 & ~w24335;
assign w26430 = w4749 & w25699;
assign w26431 = ~w26429 & ~w26430;
assign w26432 = pi0953 & ~w24335;
assign w26433 = w3711 & w25699;
assign w26434 = ~w26432 & ~w26433;
assign w26435 = w40134 & w24672;
assign w26436 = pi0954 & w24677;
assign w26437 = ~w26435 & ~w26436;
assign w26438 = w6413 & w24672;
assign w26439 = pi0955 & w24677;
assign w26440 = ~w26438 & ~w26439;
assign w26441 = w3195 & w24672;
assign w26442 = pi0956 & w24677;
assign w26443 = ~w26441 & ~w26442;
assign w26444 = w5320 & w24672;
assign w26445 = pi0957 & w24677;
assign w26446 = ~w26444 & ~w26445;
assign w26447 = w8240 & w24672;
assign w26448 = pi0958 & w24677;
assign w26449 = ~w26447 & ~w26448;
assign w26450 = w8081 & w24672;
assign w26451 = pi0959 & w24677;
assign w26452 = ~w26450 & ~w26451;
assign w26453 = w1639 & w24672;
assign w26454 = pi0960 & w24677;
assign w26455 = ~w26453 & ~w26454;
assign w26456 = w1308 & w24672;
assign w26457 = pi0961 & w24677;
assign w26458 = ~w26456 & ~w26457;
assign w26459 = pi0962 & ~w24675;
assign w26460 = w1639 & w24675;
assign w26461 = ~w26459 & ~w26460;
assign w26462 = pi0963 & ~w24675;
assign w26463 = w3195 & w24694;
assign w26464 = ~w26462 & ~w26463;
assign w26465 = pi0964 & ~w24675;
assign w26466 = w40134 & w24694;
assign w26467 = ~w26465 & ~w26466;
assign w26468 = pi0965 & ~w24675;
assign w26469 = w6413 & w24694;
assign w26470 = ~w26468 & ~w26469;
assign w26471 = pi0966 & ~w24675;
assign w26472 = w4749 & w24694;
assign w26473 = ~w26471 & ~w26472;
assign w26474 = pi0967 & ~w24675;
assign w26475 = w3711 & w24694;
assign w26476 = ~w26474 & ~w26475;
assign w26477 = w6177 & w24706;
assign w26478 = pi0968 & w24708;
assign w26479 = ~w26477 & ~w26478;
assign w26480 = w8240 & w24706;
assign w26481 = pi0969 & w24708;
assign w26482 = ~w26480 & ~w26481;
assign w26483 = w8081 & w24706;
assign w26484 = pi0970 & w24708;
assign w26485 = ~w26483 & ~w26484;
assign w26486 = w5635 & w24706;
assign w26487 = pi0971 & w24708;
assign w26488 = ~w26486 & ~w26487;
assign w26489 = w1308 & w24706;
assign w26490 = pi0972 & w24708;
assign w26491 = ~w26489 & ~w26490;
assign w26492 = pi0973 & ~w25823;
assign w26493 = ~w25824 & w25889;
assign w26494 = ~w26492 & w26493;
assign w26495 = ~pi1761 & pi3243;
assign w26496 = ~pi0609 & pi1761;
assign w26497 = pi1762 & w26496;
assign w26498 = w1265 & w24681;
assign w26499 = ~w26497 & w26498;
assign w26500 = w1639 & w26499;
assign w26501 = pi0974 & ~w26499;
assign w26502 = pi1761 & ~w26501;
assign w26503 = ~w26500 & w26502;
assign w26504 = ~w26495 & ~w26503;
assign w26505 = ~w24828 & ~w24833;
assign w26506 = w19033 & ~w24810;
assign w26507 = ~pi1422 & ~w24810;
assign w26508 = ~pi0975 & ~w26507;
assign w26509 = ~w26506 & ~w26508;
assign w26510 = w26505 & w26509;
assign w26511 = ~pi3211 & ~w2214;
assign w26512 = ~pi2487 & pi3520;
assign w26513 = ~pi1331 & ~w26512;
assign w26514 = ~w26511 & w26513;
assign w26515 = ~w7009 & w26514;
assign w26516 = ~w370 & ~w26515;
assign w26517 = pi1015 & w26516;
assign w26518 = pi0684 & ~w6681;
assign w26519 = ~pi2491 & ~w2214;
assign w26520 = ~pi0759 & pi3191;
assign w26521 = ~w26519 & w26520;
assign w26522 = ~w370 & ~w26521;
assign w26523 = ~w26518 & ~w26522;
assign w26524 = pi1015 & w1661;
assign w26525 = ~w26523 & ~w26524;
assign w26526 = pi0976 & ~w26525;
assign w26527 = ~w26517 & w26526;
assign w26528 = ~pi0976 & w26517;
assign w26529 = ~pi0976 & ~w26523;
assign w26530 = ~w26528 & ~w26529;
assign w26531 = ~w26527 & w26530;
assign w26532 = w4141 & w24706;
assign w26533 = pi0977 & w24708;
assign w26534 = ~w26532 & ~w26533;
assign w26535 = w5053 & w24706;
assign w26536 = pi0978 & w24708;
assign w26537 = ~w26535 & ~w26536;
assign w26538 = pi0866 & ~w3711;
assign w26539 = pi0979 & ~pi3521;
assign w26540 = pi3520 & pi3521;
assign w26541 = w25003 & ~w26540;
assign w26542 = ~w26539 & w26541;
assign w26543 = ~pi1512 & w10559;
assign w26544 = ~pi1041 & ~w26543;
assign w26545 = ~pi1477 & w10564;
assign w26546 = ~pi1465 & w10566;
assign w26547 = ~w26545 & ~w26546;
assign w26548 = w26544 & w26547;
assign w26549 = ~pi1581 & w10559;
assign w26550 = pi1041 & ~w26549;
assign w26551 = ~pi1531 & w10561;
assign w26552 = ~pi1392 & w10566;
assign w26553 = ~pi1549 & w10564;
assign w26554 = ~w26552 & ~w26553;
assign w26555 = ~w26551 & w26554;
assign w26556 = w26550 & w26555;
assign w26557 = ~w26548 & ~w26556;
assign w26558 = w24998 & ~w26557;
assign w26559 = ~w26542 & ~w26558;
assign w26560 = ~w26538 & w26559;
assign w26561 = pi0980 & ~w24049;
assign w26562 = ~w24052 & ~w26561;
assign w26563 = pi1007 & w3711;
assign w26564 = ~pi1042 & pi1544;
assign w26565 = pi1042 & pi1403;
assign w26566 = pi1041 & ~w26565;
assign w26567 = ~w26564 & w26566;
assign w26568 = ~pi1396 & w17569;
assign w26569 = ~pi1093 & ~w26568;
assign w26570 = ~w26567 & w26569;
assign w26571 = ~pi1042 & ~pi1576;
assign w26572 = pi1042 & ~pi1592;
assign w26573 = w24064 & ~w26572;
assign w26574 = ~w26571 & w26573;
assign w26575 = pi1042 & ~pi1525;
assign w26576 = ~pi1042 & ~pi1506;
assign w26577 = w24066 & ~w26576;
assign w26578 = ~w26575 & w26577;
assign w26579 = ~pi1007 & ~w26578;
assign w26580 = ~w26574 & w26579;
assign w26581 = ~w26570 & w26580;
assign w26582 = ~w24051 & ~w26581;
assign w26583 = ~w26563 & w26582;
assign w26584 = ~w26562 & ~w26583;
assign w26585 = w1639 & w24706;
assign w26586 = pi0981 & w24708;
assign w26587 = ~w26585 & ~w26586;
assign w26588 = ~pi0982 & w6684;
assign w26589 = w24494 & w25134;
assign w26590 = ~w26588 & ~w26589;
assign w26591 = ~pi0983 & w6684;
assign w26592 = pi0414 & ~pi0420;
assign w26593 = pi0411 & ~pi0426;
assign w26594 = w21795 & w26593;
assign w26595 = ~w26592 & ~w26594;
assign w26596 = ~w21976 & ~w21978;
assign w26597 = w26595 & w26596;
assign w26598 = w24284 & w26597;
assign w26599 = w25133 & w26598;
assign w26600 = w21988 & w26599;
assign w26601 = ~w26591 & ~w26600;
assign w26602 = ~pi0984 & w6684;
assign w26603 = w24506 & w26599;
assign w26604 = ~w26602 & ~w26603;
assign w26605 = ~pi0985 & w6684;
assign w26606 = w21988 & w26408;
assign w26607 = ~w26605 & ~w26606;
assign w26608 = ~pi0986 & w6684;
assign w26609 = w21988 & w24505;
assign w26610 = ~w26608 & ~w26609;
assign w26611 = ~pi0987 & w6684;
assign w26612 = w24284 & ~w26595;
assign w26613 = w24494 & w26612;
assign w26614 = w24283 & w26613;
assign w26615 = ~w26611 & ~w26614;
assign w26616 = ~pi0988 & w6684;
assign w26617 = w25133 & w26613;
assign w26618 = ~w26616 & ~w26617;
assign w26619 = ~pi0989 & w6684;
assign w26620 = ~w24288 & w26612;
assign w26621 = w24283 & w26620;
assign w26622 = ~w26619 & ~w26621;
assign w26623 = ~pi0990 & w6684;
assign w26624 = w24494 & w26404;
assign w26625 = ~w26623 & ~w26624;
assign w26626 = ~pi0991 & w6684;
assign w26627 = ~w24288 & w26404;
assign w26628 = ~w26626 & ~w26627;
assign w26629 = pi0992 & w6684;
assign w26630 = w24283 & w26598;
assign w26631 = w24494 & w26630;
assign w26632 = ~w26629 & ~w26631;
assign w26633 = pi0993 & w6684;
assign w26634 = w24494 & w26599;
assign w26635 = ~w26633 & ~w26634;
assign w26636 = pi0994 & w6684;
assign w26637 = ~w24288 & w26630;
assign w26638 = ~w26636 & ~w26637;
assign w26639 = pi0995 & w6684;
assign w26640 = ~w24288 & w26599;
assign w26641 = ~w26639 & ~w26640;
assign w26642 = pi0996 & w6684;
assign w26643 = w24494 & w24505;
assign w26644 = ~w26642 & ~w26643;
assign w26645 = pi0997 & w6684;
assign w26646 = w24494 & w26408;
assign w26647 = ~w26645 & ~w26646;
assign w26648 = pi0998 & w6684;
assign w26649 = w24504 & w26178;
assign w26650 = ~w26648 & ~w26649;
assign w26651 = pi0999 & w6684;
assign w26652 = ~w24288 & w26408;
assign w26653 = ~w26651 & ~w26652;
assign w26654 = ~pi1000 & w6684;
assign w26655 = w21989 & w24502;
assign w26656 = w24503 & w26655;
assign w26657 = ~w26654 & ~w26656;
assign w26658 = ~pi1001 & w22580;
assign w26659 = ~pi0884 & ~pi1069;
assign w26660 = ~pi0741 & ~pi0931;
assign w26661 = ~w26659 & ~w26660;
assign w26662 = pi0741 & pi0931;
assign w26663 = pi0884 & pi1069;
assign w26664 = ~w26662 & ~w26663;
assign w26665 = w26661 & w26664;
assign w26666 = ~pi0739 & pi1067;
assign w26667 = pi0739 & ~pi1067;
assign w26668 = ~w26666 & ~w26667;
assign w26669 = ~pi0885 & pi1088;
assign w26670 = pi0885 & ~pi1088;
assign w26671 = ~w26669 & ~w26670;
assign w26672 = ~pi0893 & pi1068;
assign w26673 = pi0893 & ~pi1068;
assign w26674 = ~w26672 & ~w26673;
assign w26675 = ~w26671 & ~w26674;
assign w26676 = ~w26668 & w26675;
assign w26677 = w26665 & w26676;
assign w26678 = pi0890 & ~pi0931;
assign w26679 = ~pi1067 & pi1068;
assign w26680 = w26678 & w26679;
assign w26681 = w22499 & w26680;
assign w26682 = pi0740 & pi1001;
assign w26683 = pi3647 & w26682;
assign w26684 = ~w26681 & w26683;
assign w26685 = ~w26677 & w26684;
assign w26686 = ~w26658 & ~w26685;
assign w26687 = ~pi1002 & w22670;
assign w26688 = ~pi0957 & pi1072;
assign w26689 = pi0957 & ~pi1072;
assign w26690 = ~w26688 & ~w26689;
assign w26691 = ~pi1009 & ~pi1040;
assign w26692 = pi1009 & pi1040;
assign w26693 = ~w26691 & ~w26692;
assign w26694 = ~w26690 & w26693;
assign w26695 = ~pi0793 & pi1071;
assign w26696 = pi0793 & ~pi1071;
assign w26697 = ~w26695 & ~w26696;
assign w26698 = ~pi0795 & pi0933;
assign w26699 = pi0795 & ~pi0933;
assign w26700 = ~w26698 & ~w26699;
assign w26701 = ~pi0799 & pi1027;
assign w26702 = pi0799 & ~pi1027;
assign w26703 = ~w26701 & ~w26702;
assign w26704 = ~w26700 & ~w26703;
assign w26705 = ~w26697 & w26704;
assign w26706 = w26694 & w26705;
assign w26707 = pi0796 & ~pi0933;
assign w26708 = pi1027 & ~pi1040;
assign w26709 = ~pi1071 & ~pi1072;
assign w26710 = w26708 & w26709;
assign w26711 = w26707 & w26710;
assign w26712 = pi0794 & pi1002;
assign w26713 = pi3635 & w26712;
assign w26714 = ~w26711 & w26713;
assign w26715 = ~w26706 & w26714;
assign w26716 = ~w26687 & ~w26715;
assign w26717 = pi3086 & w10741;
assign w26718 = ~pi3559 & w10;
assign w26719 = ~pi1676 & ~pi1677;
assign w26720 = ~pi1387 & ~pi1604;
assign w26721 = ~pi1645 & ~pi1669;
assign w26722 = w26720 & w26721;
assign w26723 = ~pi1003 & ~pi1361;
assign w26724 = w26719 & w26723;
assign w26725 = w26722 & w26724;
assign w26726 = ~pi1698 & ~pi1699;
assign w26727 = ~pi1700 & ~pi1701;
assign w26728 = w26726 & w26727;
assign w26729 = ~pi1675 & ~pi1678;
assign w26730 = ~pi1679 & ~pi1680;
assign w26731 = w26729 & w26730;
assign w26732 = ~pi1670 & ~pi1671;
assign w26733 = ~pi1672 & ~pi1673;
assign w26734 = w26732 & w26733;
assign w26735 = w26731 & w26734;
assign w26736 = w26728 & w26735;
assign w26737 = w26725 & w26736;
assign w26738 = ~pi1074 & ~pi1610;
assign w26739 = ~pi1674 & w26738;
assign w26740 = ~pi1073 & w26739;
assign w26741 = w26736 & w40062;
assign w26742 = pi3641 & ~w26741;
assign w26743 = ~pi1670 & w26742;
assign w26744 = ~pi1645 & w26743;
assign w26745 = ~pi1675 & w26744;
assign w26746 = w26719 & w26745;
assign w26747 = ~pi1699 & w26746;
assign w26748 = ~pi1678 & w26747;
assign w26749 = ~pi1679 & w26748;
assign w26750 = ~pi1680 & w26749;
assign w26751 = ~pi1698 & w26750;
assign w26752 = ~pi1669 & w26751;
assign w26753 = ~pi1701 & w26752;
assign w26754 = ~pi1361 & w26753;
assign w26755 = ~pi1671 & w26754;
assign w26756 = ~pi1700 & w26755;
assign w26757 = ~pi1387 & w26756;
assign w26758 = pi1003 & ~w26757;
assign w26759 = ~pi1003 & w26757;
assign w26760 = ~w26758 & ~w26759;
assign w26761 = ~pi3426 & w26742;
assign w26762 = ~w341 & w26761;
assign w26763 = ~pi1075 & w26762;
assign w26764 = ~pi1382 & w26763;
assign w26765 = ~pi1367 & w26764;
assign w26766 = ~pi1384 & w26765;
assign w26767 = ~pi1383 & w26766;
assign w26768 = ~pi1079 & w26767;
assign w26769 = ~pi1368 & w26768;
assign w26770 = ~pi1105 & w26769;
assign w26771 = ~pi1369 & w26770;
assign w26772 = ~pi1381 & w26771;
assign w26773 = ~pi1362 & w26772;
assign w26774 = ~pi1363 & w26773;
assign w26775 = ~pi1386 & w26774;
assign w26776 = ~pi1365 & w26775;
assign w26777 = ~pi1364 & w26776;
assign w26778 = ~pi1385 & w26777;
assign w26779 = pi1004 & ~w26778;
assign w26780 = ~pi1004 & w26778;
assign w26781 = ~w26779 & ~w26780;
assign w26782 = ~pi1366 & w26780;
assign w26783 = ~pi1076 & w26782;
assign w26784 = ~pi1077 & w26783;
assign w26785 = pi1005 & ~w26784;
assign w26786 = ~pi1005 & w26784;
assign w26787 = ~w26785 & ~w26786;
assign w26788 = ~pi1851 & ~w26291;
assign w26789 = pi3681 & w26285;
assign w26790 = pi1851 & ~w26789;
assign w26791 = w26300 & ~w26790;
assign w26792 = ~w26788 & w26791;
assign w26793 = pi1908 & ~w26792;
assign w26794 = pi1851 & pi2510;
assign w26795 = pi2824 & pi3247;
assign w26796 = pi3290 & w26795;
assign w26797 = w26794 & w26796;
assign w26798 = w26288 & w26797;
assign w26799 = ~w26793 & ~w26798;
assign w26800 = pi1006 & ~w26799;
assign w26801 = ~pi3583 & ~w26800;
assign w26802 = pi1007 & w6684;
assign w26803 = w24494 & w25589;
assign w26804 = ~w26802 & ~w26803;
assign w26805 = ~pi1008 & w6684;
assign w26806 = w24506 & w26404;
assign w26807 = ~w26805 & ~w26806;
assign w26808 = w5914 & w24672;
assign w26809 = pi1009 & w24677;
assign w26810 = ~w26808 & ~w26809;
assign w26811 = ~pi1010 & w6684;
assign w26812 = w25133 & w26620;
assign w26813 = ~w26811 & ~w26812;
assign w26814 = ~pi1011 & w6684;
assign w26815 = w24506 & w26630;
assign w26816 = ~w26814 & ~w26815;
assign w26817 = ~w343 & ~w22171;
assign w26818 = pi1012 & ~w26817;
assign w26819 = ~w4502 & w22184;
assign w26820 = ~w4749 & w22188;
assign w26821 = ~w1308 & w22190;
assign w26822 = ~w22178 & ~w26821;
assign w26823 = ~w26820 & w26822;
assign w26824 = w4464 & w22182;
assign w26825 = ~w26823 & ~w26824;
assign w26826 = ~w26819 & w26825;
assign w26827 = w8602 & w22184;
assign w26828 = ~w4471 & w22726;
assign w26829 = ~w4757 & w22196;
assign w26830 = ~w8609 & w22179;
assign w26831 = ~w8924 & w22187;
assign w26832 = ~w26830 & w26831;
assign w26833 = ~w26829 & w26832;
assign w26834 = ~w26828 & w26833;
assign w26835 = ~w26827 & w26834;
assign w26836 = w26817 & ~w26835;
assign w26837 = ~w26826 & w26836;
assign w26838 = ~w26818 & ~w26837;
assign w26839 = pi1013 & ~w26817;
assign w26840 = w22823 & w26817;
assign w26841 = ~w26839 & ~w26840;
assign w26842 = w26517 & w26523;
assign w26843 = w1045 & w26842;
assign w26844 = ~w1030 & ~w1045;
assign w26845 = w26525 & w26844;
assign w26846 = ~pi1014 & w26523;
assign w26847 = ~w26528 & w26846;
assign w26848 = ~w26845 & ~w26847;
assign w26849 = ~w26843 & w26848;
assign w26850 = w1661 & w26525;
assign w26851 = pi1015 & ~w1040;
assign w26852 = w26516 & ~w26851;
assign w26853 = ~w26525 & w26852;
assign w26854 = pi1015 & ~w26853;
assign w26855 = ~w26850 & ~w26854;
assign w26856 = pi1016 & ~w25731;
assign w26857 = ~w25732 & w25801;
assign w26858 = ~w26856 & w26857;
assign w26859 = w4380 & w24672;
assign w26860 = pi1017 & w24677;
assign w26861 = ~w26859 & ~w26860;
assign w26862 = pi1018 & ~w25819;
assign w26863 = ~w25820 & w25889;
assign w26864 = ~w26862 & w26863;
assign w26865 = ~pi1762 & pi3219;
assign w26866 = w1308 & w26499;
assign w26867 = pi1019 & ~w26499;
assign w26868 = pi1762 & ~w26867;
assign w26869 = ~w26866 & w26868;
assign w26870 = ~w26865 & ~w26869;
assign w26871 = ~pi1857 & pi3241;
assign w26872 = ~pi0609 & pi1763;
assign w26873 = pi1857 & w26872;
assign w26874 = w26498 & ~w26873;
assign w26875 = w3195 & w26874;
assign w26876 = pi1020 & ~w26874;
assign w26877 = pi1857 & ~w26876;
assign w26878 = ~w26875 & w26877;
assign w26879 = ~w26871 & ~w26878;
assign w26880 = ~pi1764 & pi3242;
assign w26881 = ~pi0609 & pi1764;
assign w26882 = pi1765 & w26881;
assign w26883 = w26498 & ~w26882;
assign w26884 = w6413 & w26883;
assign w26885 = pi1021 & ~w26883;
assign w26886 = pi1764 & ~w26885;
assign w26887 = ~w26884 & w26886;
assign w26888 = ~w26880 & ~w26887;
assign w26889 = ~pi1858 & pi3218;
assign w26890 = ~pi0609 & pi1766;
assign w26891 = pi1858 & w26890;
assign w26892 = w26498 & ~w26891;
assign w26893 = w5320 & w26892;
assign w26894 = pi1022 & ~w26892;
assign w26895 = pi1858 & ~w26894;
assign w26896 = ~w26893 & w26895;
assign w26897 = ~w26889 & ~w26896;
assign w26898 = ~pi1767 & pi3223;
assign w26899 = ~pi0609 & pi1767;
assign w26900 = pi1769 & w26899;
assign w26901 = w26498 & ~w26900;
assign w26902 = w4749 & w26901;
assign w26903 = pi1023 & ~w26901;
assign w26904 = pi1767 & ~w26903;
assign w26905 = ~w26902 & w26904;
assign w26906 = ~w26898 & ~w26905;
assign w26907 = ~pi1768 & pi3224;
assign w26908 = ~pi0609 & pi1768;
assign w26909 = pi1854 & w26908;
assign w26910 = w26498 & ~w26909;
assign w26911 = pi1024 & ~w26910;
assign w26912 = w8240 & w26910;
assign w26913 = pi1768 & ~w26912;
assign w26914 = ~w26911 & w26913;
assign w26915 = ~w26907 & ~w26914;
assign w26916 = ~pi1025 & w370;
assign w26917 = ~pi0835 & w40134;
assign w26918 = ~pi1496 & w10566;
assign w26919 = ~pi1514 & w10559;
assign w26920 = ~pi1478 & w10564;
assign w26921 = ~w26919 & ~w26920;
assign w26922 = ~w26918 & w26921;
assign w26923 = ~pi1041 & ~w26922;
assign w26924 = ~pi1582 & w10559;
assign w26925 = ~pi1550 & w10564;
assign w26926 = ~w26924 & ~w26925;
assign w26927 = pi1041 & ~w26926;
assign w26928 = pi1093 & pi1567;
assign w26929 = ~pi1093 & pi1407;
assign w26930 = w26095 & ~w26929;
assign w26931 = ~w26928 & w26930;
assign w26932 = ~w26927 & ~w26931;
assign w26933 = ~w26923 & w26932;
assign w26934 = w10627 & ~w26933;
assign w26935 = ~w370 & ~w26934;
assign w26936 = ~w26917 & w26935;
assign w26937 = ~w26916 & ~w26936;
assign w26938 = pi0802 & w22585;
assign w26939 = pi1026 & ~w22591;
assign w26940 = ~w22592 & ~w26939;
assign w26941 = w22671 & w26940;
assign w26942 = ~w26938 & ~w26941;
assign w26943 = pi0850 & w22585;
assign w26944 = pi1027 & ~w22590;
assign w26945 = ~w22591 & ~w26944;
assign w26946 = w22671 & w26945;
assign w26947 = ~w26943 & ~w26946;
assign w26948 = ~w22797 & w26817;
assign w26949 = pi1028 & ~w26817;
assign w26950 = ~w26948 & ~w26949;
assign w26951 = ~w22735 & w26817;
assign w26952 = pi1029 & ~w26817;
assign w26953 = ~w26951 & ~w26952;
assign w26954 = pi1030 & ~w26817;
assign w26955 = w22872 & w26817;
assign w26956 = ~w22887 & w26955;
assign w26957 = ~w26954 & ~w26956;
assign w26958 = pi1031 & ~w26817;
assign w26959 = w22855 & w26817;
assign w26960 = ~w26958 & ~w26959;
assign w26961 = pi1032 & ~w26817;
assign w26962 = w3934 & w22184;
assign w26963 = ~w4380 & w22188;
assign w26964 = ~w4141 & w22190;
assign w26965 = ~w22178 & ~w26964;
assign w26966 = ~w26963 & w26965;
assign w26967 = ~w9004 & w22182;
assign w26968 = ~w26966 & ~w26967;
assign w26969 = ~w26962 & w26968;
assign w26970 = ~w8743 & w22184;
assign w26971 = ~w3899 & w22726;
assign w26972 = ~w3851 & w22196;
assign w26973 = ~w8752 & w22179;
assign w26974 = ~w9016 & w22187;
assign w26975 = ~w26973 & w26974;
assign w26976 = ~w26972 & w26975;
assign w26977 = ~w26971 & w26976;
assign w26978 = ~w26970 & w26977;
assign w26979 = w26817 & ~w26978;
assign w26980 = ~w26969 & w26979;
assign w26981 = ~w26961 & ~w26980;
assign w26982 = pi1033 & ~w26817;
assign w26983 = ~w8697 & w22205;
assign w26984 = w5377 & w22190;
assign w26985 = ~w5341 & w22188;
assign w26986 = ~w8707 & w22179;
assign w26987 = ~w8975 & ~w26986;
assign w26988 = ~w22181 & w26987;
assign w26989 = ~w26985 & w26988;
assign w26990 = ~w26984 & w26989;
assign w26991 = ~w26983 & w26990;
assign w26992 = ~w5349 & w22176;
assign w26993 = w22788 & ~w26992;
assign w26994 = ~w22739 & ~w26993;
assign w26995 = ~w4835 & w22205;
assign w26996 = w5053 & w22190;
assign w26997 = ~w26995 & ~w26996;
assign w26998 = ~w26994 & w26997;
assign w26999 = w26817 & ~w26998;
assign w27000 = ~w26991 & w26999;
assign w27001 = ~w26982 & ~w27000;
assign w27002 = pi1034 & ~w26817;
assign w27003 = w8665 & ~w22176;
assign w27004 = ~w8674 & w22179;
assign w27005 = ~w8950 & ~w27004;
assign w27006 = ~w22181 & w27005;
assign w27007 = ~w27003 & w27006;
assign w27008 = ~w22178 & ~w27007;
assign w27009 = ~w8963 & w22188;
assign w27010 = w5397 & w22190;
assign w27011 = ~w27009 & ~w27010;
assign w27012 = ~w27008 & w27011;
assign w27013 = w5659 & w22196;
assign w27014 = w5939 & w22726;
assign w27015 = ~w22738 & ~w27014;
assign w27016 = ~w27013 & w27015;
assign w27017 = w5914 & w22188;
assign w27018 = w5635 & w22190;
assign w27019 = ~w27017 & ~w27018;
assign w27020 = ~w27016 & w27019;
assign w27021 = w26817 & ~w27020;
assign w27022 = ~w27012 & w27021;
assign w27023 = ~w27002 & ~w27022;
assign w27024 = pi1035 & ~w26817;
assign w27025 = w22210 & w26817;
assign w27026 = ~w27024 & ~w27025;
assign w27027 = ~w22775 & w26817;
assign w27028 = pi1036 & ~w26817;
assign w27029 = ~w27027 & ~w27028;
assign w27030 = pi1037 & ~w26817;
assign w27031 = w22913 & w26817;
assign w27032 = ~w27030 & ~w27031;
assign w27033 = pi1038 & ~w26817;
assign w27034 = w22757 & w26817;
assign w27035 = ~w27033 & ~w27034;
assign w27036 = ~pi1039 & ~w26817;
assign w27037 = ~w8558 & w22184;
assign w27038 = w22176 & w22206;
assign w27039 = ~w22176 & w22198;
assign w27040 = ~w8567 & w22179;
assign w27041 = ~w8896 & ~w27040;
assign w27042 = ~w27039 & w27041;
assign w27043 = ~w27038 & w27042;
assign w27044 = ~w27037 & w27043;
assign w27045 = w22187 & ~w27044;
assign w27046 = w3465 & w22184;
assign w27047 = w3814 & w22182;
assign w27048 = w3711 & w22188;
assign w27049 = w1639 & w22190;
assign w27050 = ~w22178 & ~w27049;
assign w27051 = ~w27048 & w27050;
assign w27052 = ~w27047 & ~w27051;
assign w27053 = ~w27046 & w27052;
assign w27054 = w26817 & ~w27053;
assign w27055 = ~w27045 & w27054;
assign w27056 = ~w27036 & ~w27055;
assign w27057 = pi0846 & w22585;
assign w27058 = pi1040 & ~w22588;
assign w27059 = ~w22589 & ~w27058;
assign w27060 = w22671 & w27059;
assign w27061 = ~w27057 & ~w27060;
assign w27062 = ~pi2487 & ~w370;
assign w27063 = w21032 & w27062;
assign w27064 = ~w26518 & ~w27063;
assign w27065 = ~w10561 & ~w27064;
assign w27066 = w10559 & w10687;
assign w27067 = w27064 & ~w27066;
assign w27068 = ~w27065 & ~w27067;
assign w27069 = ~pi1041 & w27068;
assign w27070 = pi1041 & ~w27068;
assign w27071 = ~w27069 & ~w27070;
assign w27072 = ~w370 & ~w10556;
assign w27073 = ~w26518 & ~w27072;
assign w27074 = ~pi1042 & w27073;
assign w27075 = w24074 & w27064;
assign w27076 = ~pi1042 & ~w27075;
assign w27077 = ~w24074 & ~w27064;
assign w27078 = ~w10687 & ~w27077;
assign w27079 = ~w27076 & ~w27078;
assign w27080 = ~w27074 & ~w27079;
assign w27081 = pi1014 & w26525;
assign w27082 = w26517 & w26846;
assign w27083 = ~w27081 & ~w27082;
assign w27084 = ~w26529 & ~w27083;
assign w27085 = pi1043 & ~w27084;
assign w27086 = ~pi1043 & w1036;
assign w27087 = w26842 & w27086;
assign w27088 = pi0976 & pi1043;
assign w27089 = w26523 & w27088;
assign w27090 = w1754 & ~w26523;
assign w27091 = ~w27089 & ~w27090;
assign w27092 = ~w27087 & w27091;
assign w27093 = ~w27085 & w27092;
assign w27094 = w1381 & ~w26523;
assign w27095 = ~w27087 & ~w27094;
assign w27096 = pi1044 & ~w27083;
assign w27097 = ~w27095 & ~w27096;
assign w27098 = pi1044 & w27095;
assign w27099 = ~w27097 & ~w27098;
assign w27100 = ~pi1045 & w24177;
assign w27101 = ~w24177 & ~w24225;
assign w27102 = ~pi1082 & w24176;
assign w27103 = ~w27101 & ~w27102;
assign w27104 = pi0937 & ~w24175;
assign w27105 = pi0387 & w19516;
assign w27106 = ~pi1383 & w24189;
assign w27107 = ~w27105 & ~w27106;
assign w27108 = pi0408 & w19957;
assign w27109 = ~pi1677 & w24215;
assign w27110 = ~w27108 & ~w27109;
assign w27111 = w27107 & w27110;
assign w27112 = w24179 & w27111;
assign w27113 = ~w27104 & ~w27112;
assign w27114 = ~w27103 & w27113;
assign w27115 = ~w27100 & ~w27114;
assign w27116 = ~pi0939 & pi3484;
assign w27117 = pi3571 & w27116;
assign w27118 = w23822 & w27117;
assign w27119 = pi1047 & w26523;
assign w27120 = ~w26516 & w27119;
assign w27121 = ~w26852 & ~w27120;
assign w27122 = pi1048 & ~w23792;
assign w27123 = w23808 & w23813;
assign w27124 = w23792 & w27123;
assign w27125 = ~w27122 & ~w27124;
assign w27126 = pi1049 & ~w23792;
assign w27127 = pi3641 & w23792;
assign w27128 = w23814 & w23818;
assign w27129 = w27127 & w27128;
assign w27130 = ~w27126 & ~w27129;
assign w27131 = ~pi1050 & w6684;
assign w27132 = w21988 & w26630;
assign w27133 = ~w27131 & ~w27132;
assign w27134 = ~pi1051 & w6684;
assign w27135 = w24494 & w24502;
assign w27136 = w26177 & w27135;
assign w27137 = ~w27134 & ~w27136;
assign w27138 = ~pi1052 & w24177;
assign w27139 = pi0390 & w19516;
assign w27140 = ~pi1645 & w24215;
assign w27141 = ~w27139 & ~w27140;
assign w27142 = ~pi1382 & w24189;
assign w27143 = ~pi0407 & w19957;
assign w27144 = ~w27142 & ~w27143;
assign w27145 = w27141 & w27144;
assign w27146 = w24179 & w27145;
assign w27147 = pi0911 & w24225;
assign w27148 = ~pi1080 & w24176;
assign w27149 = ~w24175 & ~w27148;
assign w27150 = ~w27147 & ~w27149;
assign w27151 = ~w27146 & w27150;
assign w27152 = ~w27138 & ~w27151;
assign w27153 = pi1053 & w343;
assign w27154 = ~w21800 & w21965;
assign w27155 = w2343 & w27154;
assign w27156 = w21952 & w27155;
assign w27157 = ~w27153 & ~w27156;
assign w27158 = pi1054 & w343;
assign w27159 = w385 & w10685;
assign w27160 = w27154 & w27159;
assign w27161 = ~w27158 & ~w27160;
assign w27162 = pi1055 & w343;
assign w27163 = w385 & w27154;
assign w27164 = w21952 & w27163;
assign w27165 = ~w27162 & ~w27164;
assign w27166 = pi1056 & w343;
assign w27167 = w10653 & w27163;
assign w27168 = ~w27166 & ~w27167;
assign w27169 = pi1057 & w343;
assign w27170 = w10653 & w27155;
assign w27171 = ~w27169 & ~w27170;
assign w27172 = pi1058 & w343;
assign w27173 = w397 & w10653;
assign w27174 = w24513 & w27173;
assign w27175 = ~w27172 & ~w27174;
assign w27176 = pi1059 & w343;
assign w27177 = w10685 & w27155;
assign w27178 = ~w27176 & ~w27177;
assign w27179 = pi3684 & w25164;
assign w27180 = pi2986 & pi2990;
assign w27181 = ~w156 & w27180;
assign w27182 = ~w25164 & ~w27181;
assign w27183 = pi1060 & w27182;
assign w27184 = ~w27179 & ~w27183;
assign w27185 = pi3690 & w25164;
assign w27186 = pi1061 & w27182;
assign w27187 = ~w27185 & ~w27186;
assign w27188 = pi3689 & w25164;
assign w27189 = pi1062 & w27182;
assign w27190 = ~w27188 & ~w27189;
assign w27191 = pi3688 & w25164;
assign w27192 = pi1063 & w27182;
assign w27193 = ~w27191 & ~w27192;
assign w27194 = pi3687 & w25164;
assign w27195 = pi1064 & w27182;
assign w27196 = ~w27194 & ~w27195;
assign w27197 = pi3686 & w25164;
assign w27198 = pi1065 & w27182;
assign w27199 = ~w27197 & ~w27198;
assign w27200 = w4141 & w23862;
assign w27201 = ~pi1066 & ~w23873;
assign w27202 = ~w23862 & ~w23874;
assign w27203 = ~w27201 & w27202;
assign w27204 = ~w27200 & ~w27203;
assign w27205 = pi0747 & w22495;
assign w27206 = pi1067 & ~w22497;
assign w27207 = ~w22498 & ~w27206;
assign w27208 = w22581 & w27207;
assign w27209 = ~w27205 & ~w27208;
assign w27210 = pi0745 & w22495;
assign w27211 = pi1068 & ~w22500;
assign w27212 = ~w22501 & ~w27211;
assign w27213 = w22581 & w27212;
assign w27214 = ~w27210 & ~w27213;
assign w27215 = pi0746 & w22495;
assign w27216 = ~pi1088 & w22498;
assign w27217 = pi1069 & ~w27216;
assign w27218 = ~w22500 & ~w27217;
assign w27219 = w22581 & w27218;
assign w27220 = ~w27215 & ~w27219;
assign w27221 = pi0981 & w22585;
assign w27222 = pi1070 & ~w22599;
assign w27223 = ~w22600 & w22671;
assign w27224 = ~w27222 & w27223;
assign w27225 = ~w27221 & ~w27224;
assign w27226 = pi0804 & w22585;
assign w27227 = pi1071 & ~w22587;
assign w27228 = ~w22588 & ~w27227;
assign w27229 = w22671 & w27228;
assign w27230 = ~w27226 & ~w27229;
assign w27231 = pi0803 & w22585;
assign w27232 = pi1072 & ~w22589;
assign w27233 = ~w22590 & ~w27232;
assign w27234 = w22671 & w27233;
assign w27235 = ~w27231 & ~w27234;
assign w27236 = pi3641 & w26737;
assign w27237 = ~pi1073 & w27236;
assign w27238 = pi1073 & ~w27236;
assign w27239 = ~w27237 & ~w27238;
assign w27240 = ~w26740 & ~w27239;
assign w27241 = ~pi1674 & w27237;
assign w27242 = ~pi1610 & w27241;
assign w27243 = pi1074 & ~w27242;
assign w27244 = pi1075 & ~w26762;
assign w27245 = ~w26763 & ~w27244;
assign w27246 = pi1076 & ~w26782;
assign w27247 = ~w26783 & ~w27246;
assign w27248 = pi1077 & ~w26783;
assign w27249 = ~w26784 & ~w27248;
assign w27250 = ~pi1086 & w26786;
assign w27251 = pi1078 & ~w27250;
assign w27252 = ~pi1078 & w27250;
assign w27253 = ~w27251 & ~w27252;
assign w27254 = pi1079 & ~w26767;
assign w27255 = ~w26768 & ~w27254;
assign w27256 = ~pi1080 & w24177;
assign w27257 = pi0389 & w19516;
assign w27258 = ~pi1367 & w24189;
assign w27259 = ~w27257 & ~w27258;
assign w27260 = pi0415 & w19957;
assign w27261 = ~pi1675 & w24215;
assign w27262 = ~w27260 & ~w27261;
assign w27263 = w27259 & w27262;
assign w27264 = w24179 & w27263;
assign w27265 = ~w24175 & ~w27102;
assign w27266 = pi1052 & w24225;
assign w27267 = ~w27265 & ~w27266;
assign w27268 = ~w27264 & w27267;
assign w27269 = ~w27256 & ~w27268;
assign w27270 = ~pi3583 & w26282;
assign w27271 = pi3397 & pi3481;
assign w27272 = ~pi2492 & w27271;
assign w27273 = ~pi3290 & w27272;
assign w27274 = w26299 & w27273;
assign w27275 = ~pi1851 & w27274;
assign w27276 = ~pi2416 & w27275;
assign w27277 = ~pi1695 & w27276;
assign w27278 = ~pi1668 & w27277;
assign w27279 = ~pi1380 & w27278;
assign w27280 = ~pi1788 & w27279;
assign w27281 = w26292 & w27280;
assign w27282 = ~pi1379 & w27280;
assign w27283 = pi1081 & ~w27282;
assign w27284 = ~w27281 & ~w27283;
assign w27285 = ~pi1082 & w24177;
assign w27286 = ~w27101 & ~w27148;
assign w27287 = pi1045 & ~w24175;
assign w27288 = ~pi1676 & w24215;
assign w27289 = ~pi1384 & w24189;
assign w27290 = ~w27288 & ~w27289;
assign w27291 = pi0388 & w19516;
assign w27292 = pi0414 & w19957;
assign w27293 = ~w27291 & ~w27292;
assign w27294 = w27290 & w27293;
assign w27295 = w24179 & w27294;
assign w27296 = ~w27287 & ~w27295;
assign w27297 = ~w27286 & w27296;
assign w27298 = ~w27285 & ~w27297;
assign w27299 = pi0744 & w22495;
assign w27300 = pi1083 & ~w22501;
assign w27301 = ~w22502 & ~w27300;
assign w27302 = w22581 & w27301;
assign w27303 = ~w27299 & ~w27302;
assign w27304 = ~pi1084 & w27252;
assign w27305 = pi1084 & ~w27252;
assign w27306 = ~w27304 & ~w27305;
assign w27307 = pi0869 & w22495;
assign w27308 = pi1085 & ~w22505;
assign w27309 = ~w22506 & w22581;
assign w27310 = ~w27308 & w27309;
assign w27311 = ~w27307 & ~w27310;
assign w27312 = pi1086 & ~w26786;
assign w27313 = ~w27250 & ~w27312;
assign w27314 = pi0870 & w22495;
assign w27315 = pi1087 & ~w22509;
assign w27316 = ~w22510 & w22581;
assign w27317 = ~w27315 & w27316;
assign w27318 = ~w27314 & ~w27317;
assign w27319 = pi0737 & w22495;
assign w27320 = pi1088 & ~w22498;
assign w27321 = ~w27216 & ~w27320;
assign w27322 = w22581 & w27321;
assign w27323 = ~w27319 & ~w27322;
assign w27324 = pi3685 & w25164;
assign w27325 = pi1089 & w27182;
assign w27326 = ~w27324 & ~w27325;
assign w27327 = w5053 & w23862;
assign w27328 = ~pi1090 & ~w23874;
assign w27329 = ~w23862 & ~w23875;
assign w27330 = ~w27328 & w27329;
assign w27331 = ~w27327 & ~w27330;
assign w27332 = pi0977 & w22585;
assign w27333 = pi1091 & ~w22595;
assign w27334 = ~w22596 & w22671;
assign w27335 = ~w27333 & w27334;
assign w27336 = ~w27332 & ~w27335;
assign w27337 = pi3683 & w25164;
assign w27338 = pi1092 & w27182;
assign w27339 = ~w27337 & ~w27338;
assign w27340 = ~w10561 & ~w27066;
assign w27341 = w27064 & ~w27340;
assign w27342 = ~w10559 & ~w24074;
assign w27343 = w27065 & w27342;
assign w27344 = w10564 & ~w10687;
assign w27345 = ~w27343 & ~w27344;
assign w27346 = ~w27341 & w27345;
assign w27347 = pi1094 & ~w25732;
assign w27348 = ~w25733 & w25801;
assign w27349 = ~w27347 & w27348;
assign w27350 = pi1095 & ~w25820;
assign w27351 = ~w25821 & w25889;
assign w27352 = ~w27350 & w27351;
assign w27353 = pi1097 & ~w25733;
assign w27354 = ~w25734 & w25801;
assign w27355 = ~w27353 & w27354;
assign w27356 = pi1098 & ~w25821;
assign w27357 = ~w25822 & w25889;
assign w27358 = ~w27356 & w27357;
assign w27359 = ~pi1763 & pi3220;
assign w27360 = w40134 & w26874;
assign w27361 = pi1099 & ~w26874;
assign w27362 = pi1763 & ~w27361;
assign w27363 = ~w27360 & w27362;
assign w27364 = ~w27359 & ~w27363;
assign w27365 = ~pi1765 & pi3221;
assign w27366 = w4380 & w26883;
assign w27367 = pi1100 & ~w26883;
assign w27368 = pi1765 & ~w27367;
assign w27369 = ~w27366 & w27368;
assign w27370 = ~w27365 & ~w27369;
assign w27371 = ~pi1766 & pi3222;
assign w27372 = w5914 & w26892;
assign w27373 = pi1101 & ~w26892;
assign w27374 = pi1766 & ~w27373;
assign w27375 = ~w27372 & w27374;
assign w27376 = ~w27371 & ~w27375;
assign w27377 = ~pi1854 & pi3240;
assign w27378 = pi1102 & ~w26910;
assign w27379 = w8081 & w26910;
assign w27380 = pi1854 & ~w27379;
assign w27381 = ~w27378 & w27380;
assign w27382 = ~w27377 & ~w27381;
assign w27383 = ~pi1769 & pi3225;
assign w27384 = w3711 & w26901;
assign w27385 = pi1103 & ~w26901;
assign w27386 = pi1769 & ~w27385;
assign w27387 = ~w27384 & w27386;
assign w27388 = ~w27383 & ~w27387;
assign w27389 = ~pi1104 & ~pi1373;
assign w27390 = ~pi1372 & w27389;
assign w27391 = ~pi1388 & w27390;
assign w27392 = ~pi1371 & w27391;
assign w27393 = pi1683 & ~pi1702;
assign w27394 = ~pi1846 & ~pi1847;
assign w27395 = w27393 & w27394;
assign w27396 = ~pi1684 & pi1703;
assign w27397 = pi1607 & pi1682;
assign w27398 = w27396 & w27397;
assign w27399 = w27395 & w27398;
assign w27400 = w27392 & w27399;
assign w27401 = ~pi2992 & ~w27400;
assign w27402 = pi3588 & ~w27401;
assign w27403 = ~pi2992 & ~pi3588;
assign w27404 = ~pi2508 & ~w27403;
assign w27405 = ~w27402 & w27404;
assign w27406 = pi0738 & ~w318;
assign w27407 = ~pi0738 & pi3671;
assign w27408 = ~w27406 & ~w27407;
assign w27409 = ~pi0880 & w27408;
assign w27410 = pi0880 & ~w27408;
assign w27411 = ~w27409 & ~w27410;
assign w27412 = pi3646 & pi3647;
assign w27413 = w27411 & w27412;
assign w27414 = ~pi0889 & w27413;
assign w27415 = pi0889 & pi3637;
assign w27416 = ~pi0791 & ~w27415;
assign w27417 = ~w27414 & w27416;
assign w27418 = pi0889 & pi3634;
assign w27419 = ~pi0889 & pi3640;
assign w27420 = pi0791 & ~w27419;
assign w27421 = ~w27418 & w27420;
assign w27422 = pi2508 & w27403;
assign w27423 = ~w27421 & w27422;
assign w27424 = ~w27417 & w27423;
assign w27425 = ~w27405 & ~w27424;
assign w27426 = ~pi2508 & ~pi2992;
assign w27427 = pi3588 & w27426;
assign w27428 = ~w27399 & w27427;
assign w27429 = w27392 & w27428;
assign w27430 = ~w27425 & ~w27429;
assign w27431 = pi1104 & pi1373;
assign w27432 = ~w27389 & ~w27431;
assign w27433 = w27430 & ~w27432;
assign w27434 = pi0739 & ~w27430;
assign w27435 = pi1685 & ~w27434;
assign w27436 = ~w27433 & w27435;
assign w27437 = pi1105 & ~w26769;
assign w27438 = ~w26770 & ~w27437;
assign w27439 = w1037 & ~w26523;
assign w27440 = pi1106 & ~w27439;
assign w27441 = ~pi0759 & ~w7086;
assign w27442 = ~pi0684 & ~w27441;
assign w27443 = pi0759 & w4141;
assign w27444 = w27442 & ~w27443;
assign w27445 = ~pi0759 & ~w7085;
assign w27446 = ~pi0684 & ~w27445;
assign w27447 = ~pi3420 & ~w27446;
assign w27448 = ~w27444 & ~w27447;
assign w27449 = w27439 & w27448;
assign w27450 = ~w27440 & ~w27449;
assign w27451 = pi1107 & ~w27439;
assign w27452 = pi0759 & w6177;
assign w27453 = w27446 & ~w27452;
assign w27454 = ~pi0759 & ~w7084;
assign w27455 = ~pi0684 & ~w27454;
assign w27456 = ~pi3411 & ~w27455;
assign w27457 = ~w27453 & ~w27456;
assign w27458 = w27439 & w27457;
assign w27459 = ~w27451 & ~w27458;
assign w27460 = pi1108 & ~w27439;
assign w27461 = pi0759 & w3195;
assign w27462 = w27455 & ~w27461;
assign w27463 = ~pi0759 & ~w7083;
assign w27464 = ~pi0684 & ~w27463;
assign w27465 = ~pi3406 & ~w27464;
assign w27466 = ~w27462 & ~w27465;
assign w27467 = w27439 & w27466;
assign w27468 = ~w27460 & ~w27467;
assign w27469 = pi1109 & ~w27439;
assign w27470 = pi0759 & w40134;
assign w27471 = w27464 & ~w27470;
assign w27472 = ~pi0759 & ~w7082;
assign w27473 = ~pi0684 & ~w27472;
assign w27474 = ~pi3413 & ~w27473;
assign w27475 = ~w27471 & ~w27474;
assign w27476 = w27439 & w27475;
assign w27477 = ~w27469 & ~w27476;
assign w27478 = pi1110 & ~w27439;
assign w27479 = pi0759 & w6413;
assign w27480 = w27473 & ~w27479;
assign w27481 = ~pi0759 & ~w7081;
assign w27482 = ~pi0684 & ~w27481;
assign w27483 = ~pi3405 & ~w27482;
assign w27484 = ~w27480 & ~w27483;
assign w27485 = w27439 & w27484;
assign w27486 = ~w27478 & ~w27485;
assign w27487 = pi1111 & ~w27439;
assign w27488 = pi0759 & w4380;
assign w27489 = w27482 & ~w27488;
assign w27490 = ~pi0759 & ~w7080;
assign w27491 = ~pi0684 & ~w27490;
assign w27492 = ~pi3414 & ~w27491;
assign w27493 = ~w27489 & ~w27492;
assign w27494 = w27439 & w27493;
assign w27495 = ~w27487 & ~w27494;
assign w27496 = pi1112 & ~w27439;
assign w27497 = pi0759 & w5320;
assign w27498 = w27491 & ~w27497;
assign w27499 = ~pi0759 & ~w7079;
assign w27500 = ~pi0684 & ~w27499;
assign w27501 = ~pi3404 & ~w27500;
assign w27502 = ~w27498 & ~w27501;
assign w27503 = w27439 & w27502;
assign w27504 = ~w27496 & ~w27503;
assign w27505 = pi1113 & ~w27439;
assign w27506 = pi0759 & w5914;
assign w27507 = w27500 & ~w27506;
assign w27508 = ~pi0759 & ~w7078;
assign w27509 = ~pi0684 & ~w27508;
assign w27510 = ~pi3402 & ~w27509;
assign w27511 = ~w27507 & ~w27510;
assign w27512 = w27439 & w27511;
assign w27513 = ~w27505 & ~w27512;
assign w27514 = pi1114 & ~w27439;
assign w27515 = pi0759 & w4749;
assign w27516 = w27509 & ~w27515;
assign w27517 = ~pi0759 & ~pi3400;
assign w27518 = ~pi0684 & ~w27517;
assign w27519 = ~pi3403 & ~w27518;
assign w27520 = ~w27516 & ~w27519;
assign w27521 = w27439 & w27520;
assign w27522 = ~w27514 & ~w27521;
assign w27523 = pi1115 & ~w27439;
assign w27524 = ~pi0759 & ~w7089;
assign w27525 = ~pi0684 & ~w27524;
assign w27526 = ~pi3430 & ~w27525;
assign w27527 = pi0759 & w1639;
assign w27528 = ~pi0759 & ~w7150;
assign w27529 = ~pi0684 & ~w27528;
assign w27530 = ~w27527 & w27529;
assign w27531 = ~w27526 & ~w27530;
assign w27532 = w27439 & w27531;
assign w27533 = ~w27523 & ~w27532;
assign w27534 = pi1116 & ~w27439;
assign w27535 = pi0759 & w1308;
assign w27536 = w27525 & ~w27535;
assign w27537 = ~pi0759 & ~w7088;
assign w27538 = ~pi0684 & ~w27537;
assign w27539 = ~pi3421 & ~w27538;
assign w27540 = ~w27536 & ~w27539;
assign w27541 = w27439 & w27540;
assign w27542 = ~w27534 & ~w27541;
assign w27543 = pi1117 & ~w27439;
assign w27544 = pi0759 & w5635;
assign w27545 = w27538 & ~w27544;
assign w27546 = ~pi0759 & ~w7087;
assign w27547 = ~pi0684 & ~w27546;
assign w27548 = ~pi3422 & ~w27547;
assign w27549 = ~w27545 & ~w27548;
assign w27550 = w27439 & w27549;
assign w27551 = ~w27543 & ~w27550;
assign w27552 = pi1118 & ~w27439;
assign w27553 = pi0759 & w5053;
assign w27554 = w27547 & ~w27553;
assign w27555 = ~pi3401 & ~w27442;
assign w27556 = ~w27554 & ~w27555;
assign w27557 = w27439 & w27556;
assign w27558 = ~w27552 & ~w27557;
assign w27559 = pi1119 & ~w27439;
assign w27560 = pi0759 & w3711;
assign w27561 = w27518 & ~w27560;
assign w27562 = pi0684 & ~pi3400;
assign w27563 = ~w27561 & ~w27562;
assign w27564 = w27439 & w27563;
assign w27565 = ~w27559 & ~w27564;
assign w27566 = w1382 & ~w26523;
assign w27567 = pi1120 & ~w27566;
assign w27568 = w27448 & w27566;
assign w27569 = ~w27567 & ~w27568;
assign w27570 = pi1121 & ~w27566;
assign w27571 = w27457 & w27566;
assign w27572 = ~w27570 & ~w27571;
assign w27573 = pi1122 & ~w27566;
assign w27574 = w27466 & w27566;
assign w27575 = ~w27573 & ~w27574;
assign w27576 = pi1123 & ~w27566;
assign w27577 = w27475 & w27566;
assign w27578 = ~w27576 & ~w27577;
assign w27579 = pi1124 & ~w27566;
assign w27580 = w27484 & w27566;
assign w27581 = ~w27579 & ~w27580;
assign w27582 = pi1125 & ~w27566;
assign w27583 = w27493 & w27566;
assign w27584 = ~w27582 & ~w27583;
assign w27585 = pi1126 & ~w27566;
assign w27586 = w27502 & w27566;
assign w27587 = ~w27585 & ~w27586;
assign w27588 = pi1127 & ~w27566;
assign w27589 = w27511 & w27566;
assign w27590 = ~w27588 & ~w27589;
assign w27591 = pi1128 & ~w27566;
assign w27592 = w27520 & w27566;
assign w27593 = ~w27591 & ~w27592;
assign w27594 = pi1129 & ~w27566;
assign w27595 = w27531 & w27566;
assign w27596 = ~w27594 & ~w27595;
assign w27597 = pi1130 & ~w27566;
assign w27598 = w27540 & w27566;
assign w27599 = ~w27597 & ~w27598;
assign w27600 = pi1131 & ~w27566;
assign w27601 = w27549 & w27566;
assign w27602 = ~w27600 & ~w27601;
assign w27603 = pi1132 & ~w27566;
assign w27604 = w27556 & w27566;
assign w27605 = ~w27603 & ~w27604;
assign w27606 = pi1133 & ~w27566;
assign w27607 = w27563 & w27566;
assign w27608 = ~w27606 & ~w27607;
assign w27609 = w1388 & ~w26523;
assign w27610 = pi1134 & ~w27609;
assign w27611 = w27448 & w27609;
assign w27612 = ~w27610 & ~w27611;
assign w27613 = pi1135 & ~w27609;
assign w27614 = w27457 & w27609;
assign w27615 = ~w27613 & ~w27614;
assign w27616 = pi1136 & ~w27609;
assign w27617 = w27466 & w27609;
assign w27618 = ~w27616 & ~w27617;
assign w27619 = pi1137 & ~w27609;
assign w27620 = w27475 & w27609;
assign w27621 = ~w27619 & ~w27620;
assign w27622 = pi1138 & ~w27609;
assign w27623 = w27484 & w27609;
assign w27624 = ~w27622 & ~w27623;
assign w27625 = pi1139 & ~w27609;
assign w27626 = w27493 & w27609;
assign w27627 = ~w27625 & ~w27626;
assign w27628 = pi1140 & ~w27609;
assign w27629 = w27502 & w27609;
assign w27630 = ~w27628 & ~w27629;
assign w27631 = pi1141 & ~w27609;
assign w27632 = w27511 & w27609;
assign w27633 = ~w27631 & ~w27632;
assign w27634 = pi1142 & ~w27609;
assign w27635 = w27520 & w27609;
assign w27636 = ~w27634 & ~w27635;
assign w27637 = pi1143 & ~w27609;
assign w27638 = w27531 & w27609;
assign w27639 = ~w27637 & ~w27638;
assign w27640 = pi1144 & ~w27609;
assign w27641 = w27540 & w27609;
assign w27642 = ~w27640 & ~w27641;
assign w27643 = pi1145 & ~w27609;
assign w27644 = w27549 & w27609;
assign w27645 = ~w27643 & ~w27644;
assign w27646 = pi1146 & ~w27609;
assign w27647 = w27556 & w27609;
assign w27648 = ~w27646 & ~w27647;
assign w27649 = pi1147 & ~w27609;
assign w27650 = w27563 & w27609;
assign w27651 = ~w27649 & ~w27650;
assign w27652 = w1411 & ~w26523;
assign w27653 = pi1148 & ~w27652;
assign w27654 = w27448 & w27652;
assign w27655 = ~w27653 & ~w27654;
assign w27656 = pi1149 & ~w27652;
assign w27657 = w27457 & w27652;
assign w27658 = ~w27656 & ~w27657;
assign w27659 = pi1150 & ~w27652;
assign w27660 = w27466 & w27652;
assign w27661 = ~w27659 & ~w27660;
assign w27662 = pi1151 & ~w27652;
assign w27663 = w27475 & w27652;
assign w27664 = ~w27662 & ~w27663;
assign w27665 = pi1152 & ~w27652;
assign w27666 = w27484 & w27652;
assign w27667 = ~w27665 & ~w27666;
assign w27668 = pi1153 & ~w27652;
assign w27669 = w27493 & w27652;
assign w27670 = ~w27668 & ~w27669;
assign w27671 = pi1154 & ~w27652;
assign w27672 = w27502 & w27652;
assign w27673 = ~w27671 & ~w27672;
assign w27674 = pi1155 & ~w27652;
assign w27675 = w27511 & w27652;
assign w27676 = ~w27674 & ~w27675;
assign w27677 = pi1156 & ~w27652;
assign w27678 = w27520 & w27652;
assign w27679 = ~w27677 & ~w27678;
assign w27680 = pi1157 & ~w27652;
assign w27681 = w27531 & w27652;
assign w27682 = ~w27680 & ~w27681;
assign w27683 = pi1158 & ~w27652;
assign w27684 = w27540 & w27652;
assign w27685 = ~w27683 & ~w27684;
assign w27686 = pi1159 & ~w27652;
assign w27687 = w27549 & w27652;
assign w27688 = ~w27686 & ~w27687;
assign w27689 = pi1160 & ~w27652;
assign w27690 = w27556 & w27652;
assign w27691 = ~w27689 & ~w27690;
assign w27692 = pi1161 & ~w27652;
assign w27693 = w27563 & w27652;
assign w27694 = ~w27692 & ~w27693;
assign w27695 = w1385 & ~w26523;
assign w27696 = pi1162 & ~w27695;
assign w27697 = w27448 & w27695;
assign w27698 = ~w27696 & ~w27697;
assign w27699 = pi1163 & ~w27695;
assign w27700 = w27457 & w27695;
assign w27701 = ~w27699 & ~w27700;
assign w27702 = pi1164 & ~w27695;
assign w27703 = w27466 & w27695;
assign w27704 = ~w27702 & ~w27703;
assign w27705 = pi1165 & ~w27695;
assign w27706 = w27475 & w27695;
assign w27707 = ~w27705 & ~w27706;
assign w27708 = pi1166 & ~w27695;
assign w27709 = w27484 & w27695;
assign w27710 = ~w27708 & ~w27709;
assign w27711 = pi1167 & ~w27695;
assign w27712 = w27493 & w27695;
assign w27713 = ~w27711 & ~w27712;
assign w27714 = pi1168 & ~w27695;
assign w27715 = w27502 & w27695;
assign w27716 = ~w27714 & ~w27715;
assign w27717 = pi1169 & ~w27695;
assign w27718 = w27511 & w27695;
assign w27719 = ~w27717 & ~w27718;
assign w27720 = pi1170 & ~w27695;
assign w27721 = w27520 & w27695;
assign w27722 = ~w27720 & ~w27721;
assign w27723 = pi1171 & ~w27695;
assign w27724 = w27531 & w27695;
assign w27725 = ~w27723 & ~w27724;
assign w27726 = pi1172 & ~w27695;
assign w27727 = w27540 & w27695;
assign w27728 = ~w27726 & ~w27727;
assign w27729 = pi1173 & ~w27695;
assign w27730 = w27549 & w27695;
assign w27731 = ~w27729 & ~w27730;
assign w27732 = pi1174 & ~w27695;
assign w27733 = w27556 & w27695;
assign w27734 = ~w27732 & ~w27733;
assign w27735 = pi1175 & ~w27695;
assign w27736 = w27563 & w27695;
assign w27737 = ~w27735 & ~w27736;
assign w27738 = w1687 & ~w26523;
assign w27739 = pi1176 & ~w27738;
assign w27740 = w27448 & w27738;
assign w27741 = ~w27739 & ~w27740;
assign w27742 = pi1177 & ~w27738;
assign w27743 = w27457 & w27738;
assign w27744 = ~w27742 & ~w27743;
assign w27745 = pi1178 & ~w27738;
assign w27746 = w27466 & w27738;
assign w27747 = ~w27745 & ~w27746;
assign w27748 = pi1179 & ~w27738;
assign w27749 = w27475 & w27738;
assign w27750 = ~w27748 & ~w27749;
assign w27751 = pi1180 & ~w27738;
assign w27752 = w27484 & w27738;
assign w27753 = ~w27751 & ~w27752;
assign w27754 = pi1181 & ~w27738;
assign w27755 = w27493 & w27738;
assign w27756 = ~w27754 & ~w27755;
assign w27757 = pi1182 & ~w27738;
assign w27758 = w27502 & w27738;
assign w27759 = ~w27757 & ~w27758;
assign w27760 = pi1183 & ~w27738;
assign w27761 = w27511 & w27738;
assign w27762 = ~w27760 & ~w27761;
assign w27763 = pi1184 & ~w27738;
assign w27764 = w27520 & w27738;
assign w27765 = ~w27763 & ~w27764;
assign w27766 = pi1185 & ~w27738;
assign w27767 = w27531 & w27738;
assign w27768 = ~w27766 & ~w27767;
assign w27769 = pi1186 & ~w27738;
assign w27770 = w27540 & w27738;
assign w27771 = ~w27769 & ~w27770;
assign w27772 = pi1187 & ~w27738;
assign w27773 = w27549 & w27738;
assign w27774 = ~w27772 & ~w27773;
assign w27775 = pi1188 & ~w27738;
assign w27776 = w27556 & w27738;
assign w27777 = ~w27775 & ~w27776;
assign w27778 = pi1189 & ~w27738;
assign w27779 = w27563 & w27738;
assign w27780 = ~w27778 & ~w27779;
assign w27781 = w1046 & ~w26523;
assign w27782 = pi1190 & ~w27781;
assign w27783 = w27448 & w27781;
assign w27784 = ~w27782 & ~w27783;
assign w27785 = pi1191 & ~w27781;
assign w27786 = w27457 & w27781;
assign w27787 = ~w27785 & ~w27786;
assign w27788 = pi1192 & ~w27781;
assign w27789 = w27466 & w27781;
assign w27790 = ~w27788 & ~w27789;
assign w27791 = pi1193 & ~w27781;
assign w27792 = w27475 & w27781;
assign w27793 = ~w27791 & ~w27792;
assign w27794 = pi1194 & ~w27781;
assign w27795 = w27484 & w27781;
assign w27796 = ~w27794 & ~w27795;
assign w27797 = pi1195 & ~w27781;
assign w27798 = w27493 & w27781;
assign w27799 = ~w27797 & ~w27798;
assign w27800 = pi1196 & ~w27781;
assign w27801 = w27502 & w27781;
assign w27802 = ~w27800 & ~w27801;
assign w27803 = pi1197 & ~w27781;
assign w27804 = w27511 & w27781;
assign w27805 = ~w27803 & ~w27804;
assign w27806 = pi1198 & ~w27781;
assign w27807 = w27520 & w27781;
assign w27808 = ~w27806 & ~w27807;
assign w27809 = pi1199 & ~w27781;
assign w27810 = w27531 & w27781;
assign w27811 = ~w27809 & ~w27810;
assign w27812 = pi1200 & ~w27781;
assign w27813 = w27540 & w27781;
assign w27814 = ~w27812 & ~w27813;
assign w27815 = pi1201 & ~w27781;
assign w27816 = w27549 & w27781;
assign w27817 = ~w27815 & ~w27816;
assign w27818 = pi1202 & ~w27781;
assign w27819 = w27556 & w27781;
assign w27820 = ~w27818 & ~w27819;
assign w27821 = pi1203 & ~w27781;
assign w27822 = w27563 & w27781;
assign w27823 = ~w27821 & ~w27822;
assign w27824 = w1043 & ~w26523;
assign w27825 = pi1204 & ~w27824;
assign w27826 = w27448 & w27824;
assign w27827 = ~w27825 & ~w27826;
assign w27828 = pi1205 & ~w27824;
assign w27829 = w27457 & w27824;
assign w27830 = ~w27828 & ~w27829;
assign w27831 = pi1206 & ~w27824;
assign w27832 = w27466 & w27824;
assign w27833 = ~w27831 & ~w27832;
assign w27834 = pi1207 & ~w27824;
assign w27835 = w27475 & w27824;
assign w27836 = ~w27834 & ~w27835;
assign w27837 = pi1208 & ~w27824;
assign w27838 = w27484 & w27824;
assign w27839 = ~w27837 & ~w27838;
assign w27840 = pi1209 & ~w27824;
assign w27841 = w27493 & w27824;
assign w27842 = ~w27840 & ~w27841;
assign w27843 = pi1210 & ~w27824;
assign w27844 = w27502 & w27824;
assign w27845 = ~w27843 & ~w27844;
assign w27846 = pi1211 & ~w27824;
assign w27847 = w27511 & w27824;
assign w27848 = ~w27846 & ~w27847;
assign w27849 = pi1212 & ~w27824;
assign w27850 = w27520 & w27824;
assign w27851 = ~w27849 & ~w27850;
assign w27852 = pi1213 & ~w27824;
assign w27853 = w27531 & w27824;
assign w27854 = ~w27852 & ~w27853;
assign w27855 = pi1214 & ~w27824;
assign w27856 = w27540 & w27824;
assign w27857 = ~w27855 & ~w27856;
assign w27858 = pi1215 & ~w27824;
assign w27859 = w27549 & w27824;
assign w27860 = ~w27858 & ~w27859;
assign w27861 = pi1216 & ~w27824;
assign w27862 = w27556 & w27824;
assign w27863 = ~w27861 & ~w27862;
assign w27864 = pi1217 & ~w27824;
assign w27865 = w27563 & w27824;
assign w27866 = ~w27864 & ~w27865;
assign w27867 = w1040 & ~w26523;
assign w27868 = pi1218 & ~w27867;
assign w27869 = w27448 & w27867;
assign w27870 = ~w27868 & ~w27869;
assign w27871 = pi1219 & ~w27867;
assign w27872 = w27457 & w27867;
assign w27873 = ~w27871 & ~w27872;
assign w27874 = pi1220 & ~w27867;
assign w27875 = w27466 & w27867;
assign w27876 = ~w27874 & ~w27875;
assign w27877 = pi1221 & ~w27867;
assign w27878 = w27475 & w27867;
assign w27879 = ~w27877 & ~w27878;
assign w27880 = pi1222 & ~w27867;
assign w27881 = w27484 & w27867;
assign w27882 = ~w27880 & ~w27881;
assign w27883 = pi1223 & ~w27867;
assign w27884 = w27493 & w27867;
assign w27885 = ~w27883 & ~w27884;
assign w27886 = pi1224 & ~w27867;
assign w27887 = w27502 & w27867;
assign w27888 = ~w27886 & ~w27887;
assign w27889 = pi1225 & ~w27867;
assign w27890 = w27511 & w27867;
assign w27891 = ~w27889 & ~w27890;
assign w27892 = pi1226 & ~w27867;
assign w27893 = w27520 & w27867;
assign w27894 = ~w27892 & ~w27893;
assign w27895 = pi1227 & ~w27867;
assign w27896 = w27531 & w27867;
assign w27897 = ~w27895 & ~w27896;
assign w27898 = pi1228 & ~w27867;
assign w27899 = w27540 & w27867;
assign w27900 = ~w27898 & ~w27899;
assign w27901 = pi1229 & ~w27867;
assign w27902 = w27549 & w27867;
assign w27903 = ~w27901 & ~w27902;
assign w27904 = pi1230 & ~w27867;
assign w27905 = w27556 & w27867;
assign w27906 = ~w27904 & ~w27905;
assign w27907 = pi1231 & ~w27867;
assign w27908 = w27563 & w27867;
assign w27909 = ~w27907 & ~w27908;
assign w27910 = w1414 & ~w26523;
assign w27911 = pi1232 & ~w27910;
assign w27912 = w27448 & w27910;
assign w27913 = ~w27911 & ~w27912;
assign w27914 = pi1233 & ~w27910;
assign w27915 = w27457 & w27910;
assign w27916 = ~w27914 & ~w27915;
assign w27917 = pi1234 & ~w27910;
assign w27918 = w27466 & w27910;
assign w27919 = ~w27917 & ~w27918;
assign w27920 = pi1235 & ~w27910;
assign w27921 = w27475 & w27910;
assign w27922 = ~w27920 & ~w27921;
assign w27923 = pi1236 & ~w27910;
assign w27924 = w27484 & w27910;
assign w27925 = ~w27923 & ~w27924;
assign w27926 = pi1237 & ~w27910;
assign w27927 = w27493 & w27910;
assign w27928 = ~w27926 & ~w27927;
assign w27929 = pi1238 & ~w27910;
assign w27930 = w27502 & w27910;
assign w27931 = ~w27929 & ~w27930;
assign w27932 = pi1239 & ~w27910;
assign w27933 = w27511 & w27910;
assign w27934 = ~w27932 & ~w27933;
assign w27935 = pi1240 & ~w27910;
assign w27936 = w27520 & w27910;
assign w27937 = ~w27935 & ~w27936;
assign w27938 = pi1241 & ~w27910;
assign w27939 = w27531 & w27910;
assign w27940 = ~w27938 & ~w27939;
assign w27941 = pi1242 & ~w27910;
assign w27942 = w27540 & w27910;
assign w27943 = ~w27941 & ~w27942;
assign w27944 = pi1243 & ~w27910;
assign w27945 = w27549 & w27910;
assign w27946 = ~w27944 & ~w27945;
assign w27947 = pi1244 & ~w27910;
assign w27948 = w27556 & w27910;
assign w27949 = ~w27947 & ~w27948;
assign w27950 = pi1245 & ~w27910;
assign w27951 = w27563 & w27910;
assign w27952 = ~w27950 & ~w27951;
assign w27953 = w1390 & ~w26523;
assign w27954 = pi1246 & ~w27953;
assign w27955 = w27448 & w27953;
assign w27956 = ~w27954 & ~w27955;
assign w27957 = pi1247 & ~w27953;
assign w27958 = w27457 & w27953;
assign w27959 = ~w27957 & ~w27958;
assign w27960 = pi1248 & ~w27953;
assign w27961 = w27466 & w27953;
assign w27962 = ~w27960 & ~w27961;
assign w27963 = pi1249 & ~w27953;
assign w27964 = w27475 & w27953;
assign w27965 = ~w27963 & ~w27964;
assign w27966 = pi1250 & ~w27953;
assign w27967 = w27484 & w27953;
assign w27968 = ~w27966 & ~w27967;
assign w27969 = pi1251 & ~w27953;
assign w27970 = w27493 & w27953;
assign w27971 = ~w27969 & ~w27970;
assign w27972 = pi1252 & ~w27953;
assign w27973 = w27502 & w27953;
assign w27974 = ~w27972 & ~w27973;
assign w27975 = pi1253 & ~w27953;
assign w27976 = w27511 & w27953;
assign w27977 = ~w27975 & ~w27976;
assign w27978 = pi1254 & ~w27953;
assign w27979 = w27520 & w27953;
assign w27980 = ~w27978 & ~w27979;
assign w27981 = pi1255 & ~w27953;
assign w27982 = w27531 & w27953;
assign w27983 = ~w27981 & ~w27982;
assign w27984 = pi1256 & ~w27953;
assign w27985 = w27540 & w27953;
assign w27986 = ~w27984 & ~w27985;
assign w27987 = pi1257 & ~w27953;
assign w27988 = w27549 & w27953;
assign w27989 = ~w27987 & ~w27988;
assign w27990 = pi1258 & ~w27953;
assign w27991 = w27556 & w27953;
assign w27992 = ~w27990 & ~w27991;
assign w27993 = pi1259 & ~w27953;
assign w27994 = w27563 & w27953;
assign w27995 = ~w27993 & ~w27994;
assign w27996 = w1678 & ~w26523;
assign w27997 = pi1260 & ~w27996;
assign w27998 = w27448 & w27996;
assign w27999 = ~w27997 & ~w27998;
assign w28000 = pi1261 & ~w27996;
assign w28001 = w27457 & w27996;
assign w28002 = ~w28000 & ~w28001;
assign w28003 = pi1262 & ~w27996;
assign w28004 = w27466 & w27996;
assign w28005 = ~w28003 & ~w28004;
assign w28006 = pi1263 & ~w27996;
assign w28007 = w27475 & w27996;
assign w28008 = ~w28006 & ~w28007;
assign w28009 = pi1264 & ~w27996;
assign w28010 = w27484 & w27996;
assign w28011 = ~w28009 & ~w28010;
assign w28012 = pi1265 & ~w27996;
assign w28013 = w27493 & w27996;
assign w28014 = ~w28012 & ~w28013;
assign w28015 = pi1266 & ~w27996;
assign w28016 = w27502 & w27996;
assign w28017 = ~w28015 & ~w28016;
assign w28018 = pi1267 & ~w27996;
assign w28019 = w27511 & w27996;
assign w28020 = ~w28018 & ~w28019;
assign w28021 = pi1268 & ~w27996;
assign w28022 = w27520 & w27996;
assign w28023 = ~w28021 & ~w28022;
assign w28024 = pi1269 & ~w27996;
assign w28025 = w27531 & w27996;
assign w28026 = ~w28024 & ~w28025;
assign w28027 = pi1270 & ~w27996;
assign w28028 = w27540 & w27996;
assign w28029 = ~w28027 & ~w28028;
assign w28030 = pi1271 & ~w27996;
assign w28031 = w27549 & w27996;
assign w28032 = ~w28030 & ~w28031;
assign w28033 = pi1272 & ~w27996;
assign w28034 = w27556 & w27996;
assign w28035 = ~w28033 & ~w28034;
assign w28036 = pi1273 & ~w27996;
assign w28037 = w27563 & w27996;
assign w28038 = ~w28036 & ~w28037;
assign w28039 = w1659 & ~w26523;
assign w28040 = pi1274 & ~w28039;
assign w28041 = w27448 & w28039;
assign w28042 = ~w28040 & ~w28041;
assign w28043 = pi1275 & ~w28039;
assign w28044 = w27457 & w28039;
assign w28045 = ~w28043 & ~w28044;
assign w28046 = pi1276 & ~w28039;
assign w28047 = w27466 & w28039;
assign w28048 = ~w28046 & ~w28047;
assign w28049 = pi1277 & ~w28039;
assign w28050 = w27475 & w28039;
assign w28051 = ~w28049 & ~w28050;
assign w28052 = pi1278 & ~w28039;
assign w28053 = w27484 & w28039;
assign w28054 = ~w28052 & ~w28053;
assign w28055 = pi1279 & ~w28039;
assign w28056 = w27493 & w28039;
assign w28057 = ~w28055 & ~w28056;
assign w28058 = pi1280 & ~w28039;
assign w28059 = w27502 & w28039;
assign w28060 = ~w28058 & ~w28059;
assign w28061 = pi1281 & ~w28039;
assign w28062 = w27511 & w28039;
assign w28063 = ~w28061 & ~w28062;
assign w28064 = pi1282 & ~w28039;
assign w28065 = w27520 & w28039;
assign w28066 = ~w28064 & ~w28065;
assign w28067 = pi1283 & ~w28039;
assign w28068 = w27531 & w28039;
assign w28069 = ~w28067 & ~w28068;
assign w28070 = pi1284 & ~w28039;
assign w28071 = w27540 & w28039;
assign w28072 = ~w28070 & ~w28071;
assign w28073 = pi1285 & ~w28039;
assign w28074 = w27549 & w28039;
assign w28075 = ~w28073 & ~w28074;
assign w28076 = pi1286 & ~w28039;
assign w28077 = w27556 & w28039;
assign w28078 = ~w28076 & ~w28077;
assign w28079 = pi1287 & ~w28039;
assign w28080 = w27563 & w28039;
assign w28081 = ~w28079 & ~w28080;
assign w28082 = w1416 & ~w26523;
assign w28083 = pi1288 & ~w28082;
assign w28084 = w27448 & w28082;
assign w28085 = ~w28083 & ~w28084;
assign w28086 = pi1289 & ~w28082;
assign w28087 = w27457 & w28082;
assign w28088 = ~w28086 & ~w28087;
assign w28089 = pi1290 & ~w28082;
assign w28090 = w27466 & w28082;
assign w28091 = ~w28089 & ~w28090;
assign w28092 = pi1291 & ~w28082;
assign w28093 = w27475 & w28082;
assign w28094 = ~w28092 & ~w28093;
assign w28095 = pi1292 & ~w28082;
assign w28096 = w27484 & w28082;
assign w28097 = ~w28095 & ~w28096;
assign w28098 = pi1293 & ~w28082;
assign w28099 = w27493 & w28082;
assign w28100 = ~w28098 & ~w28099;
assign w28101 = pi1294 & ~w28082;
assign w28102 = w27502 & w28082;
assign w28103 = ~w28101 & ~w28102;
assign w28104 = pi1295 & ~w28082;
assign w28105 = w27511 & w28082;
assign w28106 = ~w28104 & ~w28105;
assign w28107 = pi1296 & ~w28082;
assign w28108 = w27520 & w28082;
assign w28109 = ~w28107 & ~w28108;
assign w28110 = pi1297 & ~w28082;
assign w28111 = w27531 & w28082;
assign w28112 = ~w28110 & ~w28111;
assign w28113 = pi1298 & ~w28082;
assign w28114 = w27540 & w28082;
assign w28115 = ~w28113 & ~w28114;
assign w28116 = pi1299 & ~w28082;
assign w28117 = w27549 & w28082;
assign w28118 = ~w28116 & ~w28117;
assign w28119 = pi1300 & ~w28082;
assign w28120 = w27556 & w28082;
assign w28121 = ~w28119 & ~w28120;
assign w28122 = pi1301 & ~w28082;
assign w28123 = w27563 & w28082;
assign w28124 = ~w28122 & ~w28123;
assign w28125 = w1409 & ~w26523;
assign w28126 = pi1302 & ~w28125;
assign w28127 = w27448 & w28125;
assign w28128 = ~w28126 & ~w28127;
assign w28129 = pi1303 & ~w28125;
assign w28130 = w27457 & w28125;
assign w28131 = ~w28129 & ~w28130;
assign w28132 = pi1304 & ~w28125;
assign w28133 = w27466 & w28125;
assign w28134 = ~w28132 & ~w28133;
assign w28135 = pi1305 & ~w28125;
assign w28136 = w27475 & w28125;
assign w28137 = ~w28135 & ~w28136;
assign w28138 = pi1306 & ~w28125;
assign w28139 = w27484 & w28125;
assign w28140 = ~w28138 & ~w28139;
assign w28141 = pi1307 & ~w28125;
assign w28142 = w27493 & w28125;
assign w28143 = ~w28141 & ~w28142;
assign w28144 = pi1308 & ~w28125;
assign w28145 = w27502 & w28125;
assign w28146 = ~w28144 & ~w28145;
assign w28147 = pi1309 & ~w28125;
assign w28148 = w27511 & w28125;
assign w28149 = ~w28147 & ~w28148;
assign w28150 = pi1310 & ~w28125;
assign w28151 = w27520 & w28125;
assign w28152 = ~w28150 & ~w28151;
assign w28153 = pi1311 & ~w28125;
assign w28154 = w27531 & w28125;
assign w28155 = ~w28153 & ~w28154;
assign w28156 = pi1312 & ~w28125;
assign w28157 = w27540 & w28125;
assign w28158 = ~w28156 & ~w28157;
assign w28159 = pi1313 & ~w28125;
assign w28160 = w27549 & w28125;
assign w28161 = ~w28159 & ~w28160;
assign w28162 = pi1314 & ~w28125;
assign w28163 = w27556 & w28125;
assign w28164 = ~w28162 & ~w28163;
assign w28165 = pi1315 & ~w28125;
assign w28166 = w27563 & w28125;
assign w28167 = ~w28165 & ~w28166;
assign w28168 = pi1316 & ~w26850;
assign w28169 = w26850 & w27448;
assign w28170 = ~w28168 & ~w28169;
assign w28171 = pi1317 & ~w26850;
assign w28172 = w26850 & w27457;
assign w28173 = ~w28171 & ~w28172;
assign w28174 = pi1318 & ~w26850;
assign w28175 = w26850 & w27466;
assign w28176 = ~w28174 & ~w28175;
assign w28177 = pi1319 & ~w26850;
assign w28178 = w26850 & w27475;
assign w28179 = ~w28177 & ~w28178;
assign w28180 = pi1320 & ~w26850;
assign w28181 = w26850 & w27484;
assign w28182 = ~w28180 & ~w28181;
assign w28183 = pi1321 & ~w26850;
assign w28184 = w26850 & w27493;
assign w28185 = ~w28183 & ~w28184;
assign w28186 = pi1322 & ~w26850;
assign w28187 = w26850 & w27502;
assign w28188 = ~w28186 & ~w28187;
assign w28189 = pi1323 & ~w26850;
assign w28190 = w26850 & w27511;
assign w28191 = ~w28189 & ~w28190;
assign w28192 = pi1324 & ~w26850;
assign w28193 = w26850 & w27520;
assign w28194 = ~w28192 & ~w28193;
assign w28195 = pi1325 & ~w26850;
assign w28196 = w26850 & w27531;
assign w28197 = ~w28195 & ~w28196;
assign w28198 = pi1326 & ~w26850;
assign w28199 = w26850 & w27540;
assign w28200 = ~w28198 & ~w28199;
assign w28201 = pi1327 & ~w26850;
assign w28202 = w26850 & w27549;
assign w28203 = ~w28201 & ~w28202;
assign w28204 = pi1328 & ~w26850;
assign w28205 = w26850 & w27556;
assign w28206 = ~w28204 & ~w28205;
assign w28207 = pi1329 & ~w26850;
assign w28208 = w26850 & w27563;
assign w28209 = ~w28207 & ~w28208;
assign w28210 = pi1330 & ~w23792;
assign w28211 = w23819 & w23820;
assign w28212 = w27127 & w28211;
assign w28213 = ~w28210 & ~w28212;
assign w28214 = pi1331 & w6684;
assign w28215 = ~w21972 & ~w28214;
assign w28216 = pi1332 & w343;
assign w28217 = w24513 & w27159;
assign w28218 = ~w28216 & ~w28217;
assign w28219 = pi1333 & w343;
assign w28220 = w10684 & w24513;
assign w28221 = ~w28219 & ~w28220;
assign w28222 = pi1334 & w343;
assign w28223 = w2332 & w21952;
assign w28224 = w24513 & w28223;
assign w28225 = ~w28222 & ~w28224;
assign w28226 = pi1335 & w343;
assign w28227 = w385 & w21952;
assign w28228 = w24513 & w28227;
assign w28229 = ~w28226 & ~w28228;
assign w28230 = pi1336 & w343;
assign w28231 = w10720 & w24513;
assign w28232 = ~w28230 & ~w28231;
assign w28233 = pi1337 & w343;
assign w28234 = w21953 & w24132;
assign w28235 = ~w28233 & ~w28234;
assign w28236 = pi1338 & w343;
assign w28237 = w397 & w10683;
assign w28238 = w24132 & w28237;
assign w28239 = ~w28236 & ~w28238;
assign w28240 = pi1339 & w343;
assign w28241 = w24132 & w27173;
assign w28242 = ~w28240 & ~w28241;
assign w28243 = pi1340 & w343;
assign w28244 = w21962 & w27154;
assign w28245 = ~w28243 & ~w28244;
assign w28246 = pi1341 & w343;
assign w28247 = w21953 & w27154;
assign w28248 = ~w28246 & ~w28247;
assign w28249 = pi1342 & w343;
assign w28250 = w27154 & w28237;
assign w28251 = ~w28249 & ~w28250;
assign w28252 = pi1343 & w343;
assign w28253 = w27154 & w27173;
assign w28254 = ~w28252 & ~w28253;
assign w28255 = pi1344 & w343;
assign w28256 = w2332 & w10683;
assign w28257 = w24513 & w28256;
assign w28258 = ~w28255 & ~w28257;
assign w28259 = pi1345 & w343;
assign w28260 = w24132 & w27159;
assign w28261 = ~w28259 & ~w28260;
assign w28262 = pi1346 & w343;
assign w28263 = w24132 & w28227;
assign w28264 = ~w28262 & ~w28263;
assign w28265 = pi1347 & w343;
assign w28266 = w10684 & w24132;
assign w28267 = ~w28265 & ~w28266;
assign w28268 = pi1348 & w343;
assign w28269 = w10720 & w24132;
assign w28270 = ~w28268 & ~w28269;
assign w28271 = pi1349 & w343;
assign w28272 = w10684 & w27154;
assign w28273 = ~w28271 & ~w28272;
assign w28274 = pi1350 & w343;
assign w28275 = w2332 & w10685;
assign w28276 = w24132 & w28275;
assign w28277 = ~w28274 & ~w28276;
assign w28278 = pi1351 & w343;
assign w28279 = w24132 & w28223;
assign w28280 = ~w28278 & ~w28279;
assign w28281 = pi1352 & w343;
assign w28282 = w24132 & w28256;
assign w28283 = ~w28281 & ~w28282;
assign w28284 = pi1353 & w343;
assign w28285 = w22306 & w24132;
assign w28286 = ~w28284 & ~w28285;
assign w28287 = pi1354 & w343;
assign w28288 = w27154 & w28275;
assign w28289 = ~w28287 & ~w28288;
assign w28290 = pi1355 & w343;
assign w28291 = w2332 & w27154;
assign w28292 = w21952 & w28291;
assign w28293 = ~w28290 & ~w28292;
assign w28294 = pi1356 & w343;
assign w28295 = w10683 & w28291;
assign w28296 = ~w28294 & ~w28295;
assign w28297 = pi1357 & w343;
assign w28298 = w10653 & w28291;
assign w28299 = ~w28297 & ~w28298;
assign w28300 = pi1358 & w343;
assign w28301 = w24513 & w28275;
assign w28302 = ~w28300 & ~w28301;
assign w28303 = pi1359 & w343;
assign w28304 = w24513 & w28237;
assign w28305 = ~w28303 & ~w28304;
assign w28306 = ~w343 & w22307;
assign w28307 = pi1360 & w343;
assign w28308 = ~w28306 & ~w28307;
assign w28309 = pi1361 & ~w26753;
assign w28310 = ~w26754 & ~w28309;
assign w28311 = pi1362 & ~w26772;
assign w28312 = ~w26773 & ~w28311;
assign w28313 = pi1363 & ~w26773;
assign w28314 = ~w26774 & ~w28313;
assign w28315 = pi1364 & ~w26776;
assign w28316 = ~w26777 & ~w28315;
assign w28317 = pi1365 & ~w26775;
assign w28318 = ~w26776 & ~w28317;
assign w28319 = pi1366 & ~w26780;
assign w28320 = ~w26782 & ~w28319;
assign w28321 = pi1367 & ~w26764;
assign w28322 = ~w26765 & ~w28321;
assign w28323 = pi1368 & ~w26768;
assign w28324 = ~w26769 & ~w28323;
assign w28325 = pi1369 & ~w26770;
assign w28326 = ~w26771 & ~w28325;
assign w28327 = ~pi1430 & w23034;
assign w28328 = ~pi1370 & w18320;
assign w28329 = ~w23034 & ~w23036;
assign w28330 = ~w28328 & w28329;
assign w28331 = ~w28327 & ~w28330;
assign w28332 = ~pi0893 & ~w27430;
assign w28333 = pi1371 & ~w27391;
assign w28334 = ~w27392 & ~w28333;
assign w28335 = ~w27425 & w28334;
assign w28336 = pi1685 & ~w28335;
assign w28337 = ~w28332 & w28336;
assign w28338 = pi1372 & ~w27389;
assign w28339 = ~w27390 & ~w28338;
assign w28340 = w27430 & ~w28339;
assign w28341 = pi0885 & ~w27430;
assign w28342 = pi1685 & ~w28341;
assign w28343 = ~w28340 & w28342;
assign w28344 = pi0741 & ~w27430;
assign w28345 = ~pi1373 & w27430;
assign w28346 = pi1685 & ~w28345;
assign w28347 = ~w28344 & w28346;
assign w28348 = pi1608 & pi1648;
assign w28349 = pi1686 & w28348;
assign w28350 = ~pi1629 & pi1644;
assign w28351 = ~pi1687 & ~pi1848;
assign w28352 = ~pi1849 & w28351;
assign w28353 = w28350 & w28352;
assign w28354 = w28349 & w28353;
assign w28355 = ~pi1377 & ~pi1389;
assign w28356 = ~pi1376 & w28355;
assign w28357 = ~pi1375 & w28356;
assign w28358 = ~pi1374 & w28357;
assign w28359 = w28354 & w28358;
assign w28360 = ~pi2993 & ~w28359;
assign w28361 = pi3554 & ~w28360;
assign w28362 = ~pi2993 & ~pi3554;
assign w28363 = ~pi2509 & ~w28362;
assign w28364 = ~w28361 & w28363;
assign w28365 = pi0792 & ~w309;
assign w28366 = ~pi0792 & pi3669;
assign w28367 = ~w28365 & ~w28366;
assign w28368 = ~pi0956 & w28367;
assign w28369 = pi0956 & ~w28367;
assign w28370 = ~w28368 & ~w28369;
assign w28371 = pi3635 & pi3636;
assign w28372 = w28370 & w28371;
assign w28373 = ~pi0961 & w28372;
assign w28374 = pi0961 & pi3629;
assign w28375 = ~pi0899 & ~w28374;
assign w28376 = ~w28373 & w28375;
assign w28377 = pi0961 & pi3628;
assign w28378 = ~pi0961 & pi3630;
assign w28379 = pi0899 & ~w28378;
assign w28380 = ~w28377 & w28379;
assign w28381 = pi2509 & w28362;
assign w28382 = ~w28380 & w28381;
assign w28383 = ~w28376 & w28382;
assign w28384 = ~w28364 & ~w28383;
assign w28385 = ~pi2509 & ~pi2993;
assign w28386 = pi3554 & w28385;
assign w28387 = w28358 & w28386;
assign w28388 = ~w28354 & w28387;
assign w28389 = ~w28384 & ~w28388;
assign w28390 = ~pi0799 & ~w28389;
assign w28391 = pi1374 & ~w28357;
assign w28392 = ~w28358 & ~w28391;
assign w28393 = ~w28384 & w28392;
assign w28394 = pi1688 & ~w28393;
assign w28395 = ~w28390 & w28394;
assign w28396 = pi1375 & ~w28356;
assign w28397 = ~w28357 & ~w28396;
assign w28398 = w28389 & ~w28397;
assign w28399 = pi0957 & ~w28389;
assign w28400 = pi1688 & ~w28399;
assign w28401 = ~w28398 & w28400;
assign w28402 = pi1376 & ~w28355;
assign w28403 = ~w28356 & ~w28402;
assign w28404 = w28389 & ~w28403;
assign w28405 = pi1009 & ~w28389;
assign w28406 = pi1688 & ~w28405;
assign w28407 = ~w28404 & w28406;
assign w28408 = pi0795 & ~w28389;
assign w28409 = ~pi1377 & w28389;
assign w28410 = pi1688 & ~w28409;
assign w28411 = ~w28408 & w28410;
assign w28412 = ~pi1646 & ~pi1850;
assign w28413 = ~pi1694 & w28412;
assign w28414 = ~pi1643 & w28413;
assign w28415 = ~pi1692 & w28414;
assign w28416 = ~pi1691 & w28415;
assign w28417 = ~pi1693 & w28416;
assign w28418 = ~pi1649 & w28417;
assign w28419 = ~pi1690 & w28418;
assign w28420 = ~pi1689 & w28419;
assign w28421 = ~pi1378 & w28420;
assign w28422 = ~pi1689 & ~pi1831;
assign w28423 = ~pi1643 & ~pi1839;
assign w28424 = ~w28422 & ~w28423;
assign w28425 = pi1689 & pi1831;
assign w28426 = ~pi1691 & ~pi1834;
assign w28427 = ~w28425 & ~w28426;
assign w28428 = w28424 & w28427;
assign w28429 = ~pi1649 & pi1833;
assign w28430 = pi1649 & ~pi1833;
assign w28431 = ~w28429 & ~w28430;
assign w28432 = pi1692 & pi1853;
assign w28433 = pi1643 & pi1839;
assign w28434 = ~w28432 & ~w28433;
assign w28435 = ~w28431 & w28434;
assign w28436 = w28428 & w28435;
assign w28437 = ~pi1692 & ~pi1853;
assign w28438 = pi1690 & pi1832;
assign w28439 = ~w28437 & ~w28438;
assign w28440 = pi1378 & pi1830;
assign w28441 = ~pi1690 & ~pi1832;
assign w28442 = ~w28440 & ~w28441;
assign w28443 = w28439 & w28442;
assign w28444 = ~pi1378 & ~pi1830;
assign w28445 = ~pi1693 & ~pi1852;
assign w28446 = ~w28444 & ~w28445;
assign w28447 = pi1693 & pi1852;
assign w28448 = pi1691 & pi1834;
assign w28449 = ~w28447 & ~w28448;
assign w28450 = w28446 & w28449;
assign w28451 = w28443 & w28450;
assign w28452 = w28436 & w28451;
assign w28453 = pi1378 & ~w28420;
assign w28454 = ~w28452 & ~w28453;
assign w28455 = ~w28421 & w28454;
assign w28456 = pi1379 & ~w27280;
assign w28457 = ~w27282 & ~w28456;
assign w28458 = pi1380 & ~w27278;
assign w28459 = ~w27279 & ~w28458;
assign w28460 = pi1381 & ~w26771;
assign w28461 = ~w26772 & ~w28460;
assign w28462 = pi1382 & ~w26763;
assign w28463 = ~w26764 & ~w28462;
assign w28464 = pi1383 & ~w26766;
assign w28465 = ~w26767 & ~w28464;
assign w28466 = pi1384 & ~w26765;
assign w28467 = ~w26766 & ~w28466;
assign w28468 = pi1385 & ~w26777;
assign w28469 = ~w26778 & ~w28468;
assign w28470 = pi1386 & ~w26774;
assign w28471 = ~w26775 & ~w28470;
assign w28472 = pi1387 & ~w26756;
assign w28473 = ~w26757 & ~w28472;
assign w28474 = pi1388 & ~w27390;
assign w28475 = ~w27391 & ~w28474;
assign w28476 = w27430 & ~w28475;
assign w28477 = pi0884 & ~w27430;
assign w28478 = pi1685 & ~w28477;
assign w28479 = ~w28476 & w28478;
assign w28480 = pi1377 & pi1389;
assign w28481 = ~w28355 & ~w28480;
assign w28482 = w28389 & ~w28481;
assign w28483 = pi0793 & ~w28389;
assign w28484 = pi1688 & ~w28483;
assign w28485 = ~w28482 & w28484;
assign w28486 = ~pi1041 & ~w27064;
assign w28487 = w10566 & w28486;
assign w28488 = pi1390 & ~w28487;
assign w28489 = ~pi0828 & w28487;
assign w28490 = ~w28488 & ~w28489;
assign w28491 = pi1041 & ~w27064;
assign w28492 = w10566 & w28491;
assign w28493 = pi1391 & ~w28492;
assign w28494 = ~pi0827 & w28492;
assign w28495 = ~w28493 & ~w28494;
assign w28496 = w10559 & w28491;
assign w28497 = pi1392 & ~w28496;
assign w28498 = ~pi0979 & w28496;
assign w28499 = ~w28497 & ~w28498;
assign w28500 = w10561 & w28486;
assign w28501 = pi1393 & ~w28500;
assign w28502 = ~pi0918 & w28500;
assign w28503 = ~w28501 & ~w28502;
assign w28504 = pi1394 & ~w28496;
assign w28505 = ~pi0659 & w28496;
assign w28506 = ~w28504 & ~w28505;
assign w28507 = w10561 & w28491;
assign w28508 = pi1395 & ~w28507;
assign w28509 = ~pi0916 & w28507;
assign w28510 = ~w28508 & ~w28509;
assign w28511 = pi1396 & ~w28487;
assign w28512 = ~pi0980 & w28487;
assign w28513 = ~w28511 & ~w28512;
assign w28514 = pi1397 & ~w28487;
assign w28515 = ~pi0917 & w28487;
assign w28516 = ~w28514 & ~w28515;
assign w28517 = pi1398 & ~w28487;
assign w28518 = ~pi0916 & w28487;
assign w28519 = ~w28517 & ~w28518;
assign w28520 = pi1399 & ~w28492;
assign w28521 = ~pi0828 & w28492;
assign w28522 = ~w28520 & ~w28521;
assign w28523 = pi1400 & ~w28487;
assign w28524 = ~pi0914 & w28487;
assign w28525 = ~w28523 & ~w28524;
assign w28526 = pi1401 & ~w28500;
assign w28527 = ~pi0828 & w28500;
assign w28528 = ~w28526 & ~w28527;
assign w28529 = pi1402 & ~w28487;
assign w28530 = ~pi0586 & w28487;
assign w28531 = ~w28529 & ~w28530;
assign w28532 = pi1403 & ~w28492;
assign w28533 = ~pi0980 & w28492;
assign w28534 = ~w28532 & ~w28533;
assign w28535 = pi1404 & ~w28492;
assign w28536 = ~pi0914 & w28492;
assign w28537 = ~w28535 & ~w28536;
assign w28538 = pi1405 & ~w28492;
assign w28539 = ~pi0917 & w28492;
assign w28540 = ~w28538 & ~w28539;
assign w28541 = pi1406 & ~w28487;
assign w28542 = ~pi0196 & w28487;
assign w28543 = ~w28541 & ~w28542;
assign w28544 = w10564 & w28491;
assign w28545 = pi1407 & ~w28544;
assign w28546 = pi3633 & w28544;
assign w28547 = ~w28545 & ~w28546;
assign w28548 = pi1408 & ~w28492;
assign w28549 = ~pi0912 & w28492;
assign w28550 = ~w28548 & ~w28549;
assign w28551 = pi1409 & ~w28492;
assign w28552 = ~pi0196 & w28492;
assign w28553 = ~w28551 & ~w28552;
assign w28554 = pi1410 & ~w28492;
assign w28555 = ~pi0586 & w28492;
assign w28556 = ~w28554 & ~w28555;
assign w28557 = pi1411 & ~w28544;
assign w28558 = ~pi0826 & w28544;
assign w28559 = ~w28557 & ~w28558;
assign w28560 = pi1412 & ~w28544;
assign w28561 = ~pi0829 & w28544;
assign w28562 = ~w28560 & ~w28561;
assign w28563 = pi1413 & ~w28544;
assign w28564 = ~pi0868 & w28544;
assign w28565 = ~w28563 & ~w28564;
assign w28566 = pi1414 & ~w28500;
assign w28567 = ~pi0149 & w28500;
assign w28568 = ~w28566 & ~w28567;
assign w28569 = pi1415 & ~w28544;
assign w28570 = ~pi0708 & w28544;
assign w28571 = ~w28569 & ~w28570;
assign w28572 = pi1416 & ~w28544;
assign w28573 = ~pi0915 & w28544;
assign w28574 = ~w28572 & ~w28573;
assign w28575 = pi1417 & ~w28544;
assign w28576 = ~pi0152 & w28544;
assign w28577 = ~w28575 & ~w28576;
assign w28578 = pi0423 & pi0424;
assign w28579 = w14366 & w28578;
assign w28580 = ~w21802 & ~w28579;
assign w28581 = w14887 & ~w28580;
assign w28582 = ~pi1418 & ~w14887;
assign w28583 = ~w28581 & ~w28582;
assign w28584 = pi1419 & ~w28507;
assign w28585 = ~pi0918 & w28507;
assign w28586 = ~w28584 & ~w28585;
assign w28587 = pi1420 & ~w28507;
assign w28588 = ~pi0149 & w28507;
assign w28589 = ~w28587 & ~w28588;
assign w28590 = pi1421 & ~w28507;
assign w28591 = ~pi0827 & w28507;
assign w28592 = ~w28590 & ~w28591;
assign w28593 = ~pi1422 & w24836;
assign w28594 = ~pi3579 & w8081;
assign w28595 = ~pi3465 & pi3579;
assign w28596 = ~w24836 & ~w28595;
assign w28597 = ~w28594 & w28596;
assign w28598 = ~w28593 & ~w28597;
assign w28599 = pi1423 & ~w28500;
assign w28600 = ~pi0827 & w28500;
assign w28601 = ~w28599 & ~w28600;
assign w28602 = ~pi1424 & ~w14887;
assign w28603 = ~w28581 & ~w28602;
assign w28604 = ~pi1425 & ~w14887;
assign w28605 = ~w28581 & ~w28604;
assign w28606 = w1256 & w24330;
assign w28607 = w24374 & w28606;
assign w28608 = pi1426 & ~w28607;
assign w28609 = w8240 & w28607;
assign w28610 = ~w28608 & ~w28609;
assign w28611 = pi1427 & ~w28607;
assign w28612 = w3195 & w28607;
assign w28613 = ~w28611 & ~w28612;
assign w28614 = pi1428 & ~w28607;
assign w28615 = w40134 & w28607;
assign w28616 = ~w28614 & ~w28615;
assign w28617 = pi1429 & ~w28607;
assign w28618 = w6413 & w28607;
assign w28619 = ~w28617 & ~w28618;
assign w28620 = pi1430 & ~w28607;
assign w28621 = w4380 & w28607;
assign w28622 = ~w28620 & ~w28621;
assign w28623 = pi1431 & ~w28607;
assign w28624 = w5320 & w28607;
assign w28625 = ~w28623 & ~w28624;
assign w28626 = pi1432 & ~w28607;
assign w28627 = w5914 & w28607;
assign w28628 = ~w28626 & ~w28627;
assign w28629 = pi1433 & ~w28607;
assign w28630 = w4749 & w28607;
assign w28631 = ~w28629 & ~w28630;
assign w28632 = pi1434 & ~w28607;
assign w28633 = w3711 & w28607;
assign w28634 = ~w28632 & ~w28633;
assign w28635 = pi1435 & ~w25729;
assign w28636 = ~w25730 & w25801;
assign w28637 = ~w28635 & w28636;
assign w28638 = w1286 & w24671;
assign w28639 = pi1436 & ~w28638;
assign w28640 = w4141 & w28638;
assign w28641 = ~w28639 & ~w28640;
assign w28642 = pi1437 & ~w28638;
assign w28643 = w6177 & w28638;
assign w28644 = ~w28642 & ~w28643;
assign w28645 = pi1438 & ~w28638;
assign w28646 = w3195 & w28638;
assign w28647 = ~w28645 & ~w28646;
assign w28648 = pi1439 & ~w28638;
assign w28649 = w40134 & w28638;
assign w28650 = ~w28648 & ~w28649;
assign w28651 = pi1440 & ~w28638;
assign w28652 = w6413 & w28638;
assign w28653 = ~w28651 & ~w28652;
assign w28654 = pi1441 & ~w28638;
assign w28655 = w4380 & w28638;
assign w28656 = ~w28654 & ~w28655;
assign w28657 = pi1442 & ~w28638;
assign w28658 = w5320 & w28638;
assign w28659 = ~w28657 & ~w28658;
assign w28660 = pi1443 & ~w28638;
assign w28661 = w5914 & w28638;
assign w28662 = ~w28660 & ~w28661;
assign w28663 = pi1444 & ~w28638;
assign w28664 = w4749 & w28638;
assign w28665 = ~w28663 & ~w28664;
assign w28666 = pi1445 & ~w28638;
assign w28667 = w5635 & w28638;
assign w28668 = ~w28666 & ~w28667;
assign w28669 = pi1446 & ~w28638;
assign w28670 = w5053 & w28638;
assign w28671 = ~w28669 & ~w28670;
assign w28672 = pi1447 & ~w28638;
assign w28673 = w3711 & w28638;
assign w28674 = ~w28672 & ~w28673;
assign w28675 = pi1448 & ~w25817;
assign w28676 = ~w25818 & w25889;
assign w28677 = ~w28675 & w28676;
assign w28678 = pi3651 & ~pi3652;
assign w28679 = pi3529 & ~w28678;
assign w28680 = pi3529 & w28678;
assign w28681 = ~pi0873 & ~pi0874;
assign w28682 = ~pi0876 & ~pi0902;
assign w28683 = w28681 & w28682;
assign w28684 = ~pi0819 & ~pi0820;
assign w28685 = w19033 & w28684;
assign w28686 = w28683 & w28685;
assign w28687 = ~pi0907 & ~pi0908;
assign w28688 = ~pi0909 & ~pi0910;
assign w28689 = w28687 & w28688;
assign w28690 = ~pi0903 & ~pi0904;
assign w28691 = ~pi0905 & ~pi0906;
assign w28692 = w28690 & w28691;
assign w28693 = w28689 & w28692;
assign w28694 = w28686 & w28693;
assign w28695 = w24809 & w28694;
assign w28696 = pi1449 & ~w28695;
assign w28697 = ~pi3467 & w24828;
assign w28698 = ~w24812 & w24831;
assign w28699 = w23839 & w28698;
assign w28700 = ~w28697 & ~w28699;
assign w28701 = ~w25895 & ~w28700;
assign w28702 = ~pi1450 & w28700;
assign w28703 = ~w28701 & ~w28702;
assign w28704 = ~w25903 & ~w28700;
assign w28705 = ~pi1451 & w28700;
assign w28706 = ~w28704 & ~w28705;
assign w28707 = ~w25658 & ~w28700;
assign w28708 = ~pi1452 & w28700;
assign w28709 = ~w28707 & ~w28708;
assign w28710 = ~w25911 & ~w28700;
assign w28711 = ~pi1453 & w28700;
assign w28712 = ~w28710 & ~w28711;
assign w28713 = ~w25919 & ~w28700;
assign w28714 = ~pi1454 & w28700;
assign w28715 = ~w28713 & ~w28714;
assign w28716 = ~w25927 & ~w28700;
assign w28717 = ~pi1455 & w28700;
assign w28718 = ~w28716 & ~w28717;
assign w28719 = ~w25644 & ~w28700;
assign w28720 = ~pi1456 & w28700;
assign w28721 = ~w28719 & ~w28720;
assign w28722 = ~w25935 & ~w28700;
assign w28723 = ~pi1457 & w28700;
assign w28724 = ~w28722 & ~w28723;
assign w28725 = ~w25943 & ~w28700;
assign w28726 = ~pi1458 & w28700;
assign w28727 = ~w28725 & ~w28726;
assign w28728 = ~w24847 & ~w28700;
assign w28729 = ~pi1459 & w28700;
assign w28730 = ~w28728 & ~w28729;
assign w28731 = ~w25960 & ~w28700;
assign w28732 = ~pi1460 & w28700;
assign w28733 = ~w28731 & ~w28732;
assign w28734 = ~w25636 & ~w28700;
assign w28735 = ~pi1461 & w28700;
assign w28736 = ~w28734 & ~w28735;
assign w28737 = ~pi2529 & ~pi3680;
assign w28738 = pi2409 & pi2647;
assign w28739 = ~w28737 & w28738;
assign w28740 = pi3344 & w28739;
assign w28741 = ~w908 & ~w916;
assign w28742 = pi3641 & w28741;
assign w28743 = ~pi3631 & ~w28742;
assign w28744 = ~pi0565 & ~pi3641;
assign w28745 = ~pi0565 & pi3582;
assign w28746 = ~w28744 & ~w28745;
assign w28747 = w28743 & w28746;
assign w28748 = ~w28740 & w28747;
assign w28749 = pi3324 & ~w28745;
assign w28750 = w96 & w28749;
assign w28751 = pi3294 & w28740;
assign w28752 = w28750 & w28751;
assign w28753 = ~w28748 & ~w28752;
assign w28754 = ~pi2789 & ~pi3257;
assign w28755 = pi0565 & w117;
assign w28756 = ~w28754 & w28755;
assign w28757 = ~w28753 & w28756;
assign w28758 = w180 & w28749;
assign w28759 = pi1462 & ~w28758;
assign w28760 = w28753 & w28759;
assign w28761 = ~w28757 & ~w28760;
assign w28762 = pi1463 & ~w28507;
assign w28763 = ~pi0912 & w28507;
assign w28764 = ~w28762 & ~w28763;
assign w28765 = pi1464 & ~w28500;
assign w28766 = ~pi0912 & w28500;
assign w28767 = ~w28765 & ~w28766;
assign w28768 = w10559 & w28486;
assign w28769 = pi1465 & ~w28768;
assign w28770 = ~pi0979 & w28768;
assign w28771 = ~w28769 & ~w28770;
assign w28772 = pi1466 & ~w28500;
assign w28773 = ~pi0916 & w28500;
assign w28774 = ~w28772 & ~w28773;
assign w28775 = w4380 & w23862;
assign w28776 = ~pi1467 & ~w23868;
assign w28777 = ~w23869 & ~w28776;
assign w28778 = ~w23862 & w28777;
assign w28779 = ~w28775 & ~w28778;
assign w28780 = ~pi1468 & ~w14887;
assign w28781 = ~w28581 & ~w28780;
assign w28782 = ~pi1469 & ~w14887;
assign w28783 = ~w28581 & ~w28782;
assign w28784 = ~pi1470 & ~w14887;
assign w28785 = ~w28581 & ~w28784;
assign w28786 = ~pi1471 & ~w14887;
assign w28787 = ~w28581 & ~w28786;
assign w28788 = ~pi1472 & ~w14887;
assign w28789 = ~pi0423 & pi0424;
assign w28790 = ~pi0422 & ~w28789;
assign w28791 = ~pi0405 & ~w28790;
assign w28792 = w14887 & w28791;
assign w28793 = ~w28788 & ~w28792;
assign w28794 = ~pi1473 & ~w14887;
assign w28795 = ~w28581 & ~w28794;
assign w28796 = w40134 & w23862;
assign w28797 = ~pi1474 & ~w23870;
assign w28798 = ~w23862 & ~w23871;
assign w28799 = ~w28797 & w28798;
assign w28800 = ~w28796 & ~w28799;
assign w28801 = pi1475 & ~w28500;
assign w28802 = ~pi0914 & w28500;
assign w28803 = ~w28801 & ~w28802;
assign w28804 = pi1476 & ~w28487;
assign w28805 = ~pi0830 & w28487;
assign w28806 = ~w28804 & ~w28805;
assign w28807 = pi1477 & ~w28487;
assign w28808 = ~pi0979 & w28487;
assign w28809 = ~w28807 & ~w28808;
assign w28810 = pi1478 & ~w28487;
assign w28811 = pi3633 & w28487;
assign w28812 = ~w28810 & ~w28811;
assign w28813 = pi1479 & ~w28487;
assign w28814 = ~pi0143 & w28487;
assign w28815 = ~w28813 & ~w28814;
assign w28816 = pi1480 & ~w28487;
assign w28817 = ~pi0659 & w28487;
assign w28818 = ~w28816 & ~w28817;
assign w28819 = pi1481 & ~w28487;
assign w28820 = ~pi0152 & w28487;
assign w28821 = ~w28819 & ~w28820;
assign w28822 = pi1482 & ~w28487;
assign w28823 = ~pi0912 & w28487;
assign w28824 = ~w28822 & ~w28823;
assign w28825 = pi1483 & ~w28487;
assign w28826 = ~pi0913 & w28487;
assign w28827 = ~w28825 & ~w28826;
assign w28828 = pi1484 & ~w28487;
assign w28829 = ~pi0915 & w28487;
assign w28830 = ~w28828 & ~w28829;
assign w28831 = pi1485 & ~w28487;
assign w28832 = ~pi0134 & w28487;
assign w28833 = ~w28831 & ~w28832;
assign w28834 = pi1486 & ~w28487;
assign w28835 = ~pi0708 & w28487;
assign w28836 = ~w28834 & ~w28835;
assign w28837 = pi1487 & ~w28487;
assign w28838 = ~pi0918 & w28487;
assign w28839 = ~w28837 & ~w28838;
assign w28840 = pi1488 & ~w28487;
assign w28841 = ~pi0919 & w28487;
assign w28842 = ~w28840 & ~w28841;
assign w28843 = pi1489 & ~w28487;
assign w28844 = ~pi0826 & w28487;
assign w28845 = ~w28843 & ~w28844;
assign w28846 = pi1490 & ~w28487;
assign w28847 = ~pi0827 & w28487;
assign w28848 = ~w28846 & ~w28847;
assign w28849 = pi1491 & ~w28487;
assign w28850 = ~pi0868 & w28487;
assign w28851 = ~w28849 & ~w28850;
assign w28852 = pi1492 & ~w28487;
assign w28853 = ~pi0829 & w28487;
assign w28854 = ~w28852 & ~w28853;
assign w28855 = pi1493 & ~w28487;
assign w28856 = ~pi0149 & w28487;
assign w28857 = ~w28855 & ~w28856;
assign w28858 = pi1494 & ~w28768;
assign w28859 = ~pi0830 & w28768;
assign w28860 = ~w28858 & ~w28859;
assign w28861 = pi1495 & ~w28768;
assign w28862 = ~pi0586 & w28768;
assign w28863 = ~w28861 & ~w28862;
assign w28864 = pi1496 & ~w28768;
assign w28865 = pi3633 & w28768;
assign w28866 = ~w28864 & ~w28865;
assign w28867 = pi1497 & ~w28768;
assign w28868 = ~pi0143 & w28768;
assign w28869 = ~w28867 & ~w28868;
assign w28870 = pi1498 & ~w28768;
assign w28871 = ~pi0196 & w28768;
assign w28872 = ~w28870 & ~w28871;
assign w28873 = pi1499 & ~w28768;
assign w28874 = ~pi0152 & w28768;
assign w28875 = ~w28873 & ~w28874;
assign w28876 = pi1500 & ~w28768;
assign w28877 = ~pi0912 & w28768;
assign w28878 = ~w28876 & ~w28877;
assign w28879 = pi1501 & ~w28768;
assign w28880 = ~pi0914 & w28768;
assign w28881 = ~w28879 & ~w28880;
assign w28882 = pi1502 & ~w28768;
assign w28883 = ~pi0915 & w28768;
assign w28884 = ~w28882 & ~w28883;
assign w28885 = pi1503 & ~w28768;
assign w28886 = ~pi0916 & w28768;
assign w28887 = ~w28885 & ~w28886;
assign w28888 = pi1504 & ~w28768;
assign w28889 = ~pi0917 & w28768;
assign w28890 = ~w28888 & ~w28889;
assign w28891 = pi1505 & ~w28768;
assign w28892 = ~pi0918 & w28768;
assign w28893 = ~w28891 & ~w28892;
assign w28894 = pi1506 & ~w28768;
assign w28895 = ~pi0980 & w28768;
assign w28896 = ~w28894 & ~w28895;
assign w28897 = pi1507 & ~w28768;
assign w28898 = ~pi0826 & w28768;
assign w28899 = ~w28897 & ~w28898;
assign w28900 = pi1508 & ~w28768;
assign w28901 = ~pi0827 & w28768;
assign w28902 = ~w28900 & ~w28901;
assign w28903 = pi1509 & ~w28768;
assign w28904 = ~pi0828 & w28768;
assign w28905 = ~w28903 & ~w28904;
assign w28906 = pi1510 & ~w28768;
assign w28907 = ~pi0829 & w28768;
assign w28908 = ~w28906 & ~w28907;
assign w28909 = pi1511 & ~w28768;
assign w28910 = ~pi0149 & w28768;
assign w28911 = ~w28909 & ~w28910;
assign w28912 = pi1512 & ~w28507;
assign w28913 = ~pi0979 & w28507;
assign w28914 = ~w28912 & ~w28913;
assign w28915 = pi1513 & ~w28507;
assign w28916 = ~pi0586 & w28507;
assign w28917 = ~w28915 & ~w28916;
assign w28918 = pi1514 & ~w28507;
assign w28919 = pi3633 & w28507;
assign w28920 = ~w28918 & ~w28919;
assign w28921 = pi1515 & ~w28507;
assign w28922 = ~pi0659 & w28507;
assign w28923 = ~w28921 & ~w28922;
assign w28924 = pi1516 & ~w28507;
assign w28925 = ~pi0196 & w28507;
assign w28926 = ~w28924 & ~w28925;
assign w28927 = pi1517 & ~w28507;
assign w28928 = ~pi0152 & w28507;
assign w28929 = ~w28927 & ~w28928;
assign w28930 = pi1518 & ~w28507;
assign w28931 = ~pi0913 & w28507;
assign w28932 = ~w28930 & ~w28931;
assign w28933 = pi1519 & ~w28507;
assign w28934 = ~pi0914 & w28507;
assign w28935 = ~w28933 & ~w28934;
assign w28936 = pi1520 & ~w28507;
assign w28937 = ~pi0915 & w28507;
assign w28938 = ~w28936 & ~w28937;
assign w28939 = pi1521 & ~w28507;
assign w28940 = ~pi0134 & w28507;
assign w28941 = ~w28939 & ~w28940;
assign w28942 = pi1522 & ~w28507;
assign w28943 = ~pi0917 & w28507;
assign w28944 = ~w28942 & ~w28943;
assign w28945 = pi1523 & ~w28507;
assign w28946 = ~pi0708 & w28507;
assign w28947 = ~w28945 & ~w28946;
assign w28948 = pi1524 & ~w28507;
assign w28949 = ~pi0919 & w28507;
assign w28950 = ~w28948 & ~w28949;
assign w28951 = pi1525 & ~w28507;
assign w28952 = ~pi0980 & w28507;
assign w28953 = ~w28951 & ~w28952;
assign w28954 = pi1526 & ~w28507;
assign w28955 = ~pi0826 & w28507;
assign w28956 = ~w28954 & ~w28955;
assign w28957 = pi1527 & ~w28507;
assign w28958 = ~pi0868 & w28507;
assign w28959 = ~w28957 & ~w28958;
assign w28960 = pi1528 & ~w28507;
assign w28961 = ~pi0828 & w28507;
assign w28962 = ~w28960 & ~w28961;
assign w28963 = pi1529 & ~w28507;
assign w28964 = ~pi0829 & w28507;
assign w28965 = ~w28963 & ~w28964;
assign w28966 = pi1530 & ~w28544;
assign w28967 = ~pi0830 & w28544;
assign w28968 = ~w28966 & ~w28967;
assign w28969 = pi1531 & ~w28544;
assign w28970 = ~pi0979 & w28544;
assign w28971 = ~w28969 & ~w28970;
assign w28972 = pi1532 & ~w28544;
assign w28973 = ~pi0586 & w28544;
assign w28974 = ~w28972 & ~w28973;
assign w28975 = pi1533 & ~w28544;
assign w28976 = ~pi0143 & w28544;
assign w28977 = ~w28975 & ~w28976;
assign w28978 = pi1534 & ~w28544;
assign w28979 = ~pi0659 & w28544;
assign w28980 = ~w28978 & ~w28979;
assign w28981 = pi1535 & ~w28544;
assign w28982 = ~pi0196 & w28544;
assign w28983 = ~w28981 & ~w28982;
assign w28984 = pi1536 & ~w28544;
assign w28985 = ~pi0912 & w28544;
assign w28986 = ~w28984 & ~w28985;
assign w28987 = pi1537 & ~w28544;
assign w28988 = ~pi0913 & w28544;
assign w28989 = ~w28987 & ~w28988;
assign w28990 = pi1538 & ~w28544;
assign w28991 = ~pi0914 & w28544;
assign w28992 = ~w28990 & ~w28991;
assign w28993 = pi1539 & ~w28544;
assign w28994 = ~pi0916 & w28544;
assign w28995 = ~w28993 & ~w28994;
assign w28996 = pi1540 & ~w28544;
assign w28997 = ~pi0134 & w28544;
assign w28998 = ~w28996 & ~w28997;
assign w28999 = pi1541 & ~w28544;
assign w29000 = ~pi0917 & w28544;
assign w29001 = ~w28999 & ~w29000;
assign w29002 = pi1542 & ~w28544;
assign w29003 = ~pi0918 & w28544;
assign w29004 = ~w29002 & ~w29003;
assign w29005 = pi1543 & ~w28544;
assign w29006 = ~pi0919 & w28544;
assign w29007 = ~w29005 & ~w29006;
assign w29008 = pi1544 & ~w28544;
assign w29009 = ~pi0980 & w28544;
assign w29010 = ~w29008 & ~w29009;
assign w29011 = pi1545 & ~w28544;
assign w29012 = ~pi0827 & w28544;
assign w29013 = ~w29011 & ~w29012;
assign w29014 = pi1546 & ~w28544;
assign w29015 = ~pi0828 & w28544;
assign w29016 = ~w29014 & ~w29015;
assign w29017 = pi1547 & ~w28544;
assign w29018 = ~pi0149 & w28544;
assign w29019 = ~w29017 & ~w29018;
assign w29020 = pi1548 & ~w28492;
assign w29021 = ~pi0830 & w28492;
assign w29022 = ~w29020 & ~w29021;
assign w29023 = pi1549 & ~w28492;
assign w29024 = ~pi0979 & w28492;
assign w29025 = ~w29023 & ~w29024;
assign w29026 = pi1550 & ~w28492;
assign w29027 = pi3633 & w28492;
assign w29028 = ~w29026 & ~w29027;
assign w29029 = pi1551 & ~w28492;
assign w29030 = ~pi0143 & w28492;
assign w29031 = ~w29029 & ~w29030;
assign w29032 = pi1552 & ~w28492;
assign w29033 = ~pi0659 & w28492;
assign w29034 = ~w29032 & ~w29033;
assign w29035 = pi1553 & ~w28492;
assign w29036 = ~pi0152 & w28492;
assign w29037 = ~w29035 & ~w29036;
assign w29038 = pi1554 & ~w28492;
assign w29039 = ~pi0913 & w28492;
assign w29040 = ~w29038 & ~w29039;
assign w29041 = pi1555 & ~w28492;
assign w29042 = ~pi0915 & w28492;
assign w29043 = ~w29041 & ~w29042;
assign w29044 = pi1556 & ~w28492;
assign w29045 = ~pi0916 & w28492;
assign w29046 = ~w29044 & ~w29045;
assign w29047 = pi1557 & ~w28492;
assign w29048 = ~pi0134 & w28492;
assign w29049 = ~w29047 & ~w29048;
assign w29050 = pi1558 & ~w28492;
assign w29051 = ~pi0708 & w28492;
assign w29052 = ~w29050 & ~w29051;
assign w29053 = pi1559 & ~w28492;
assign w29054 = ~pi0918 & w28492;
assign w29055 = ~w29053 & ~w29054;
assign w29056 = pi1560 & ~w28492;
assign w29057 = ~pi0919 & w28492;
assign w29058 = ~w29056 & ~w29057;
assign w29059 = pi1561 & ~w28492;
assign w29060 = ~pi0826 & w28492;
assign w29061 = ~w29059 & ~w29060;
assign w29062 = pi1562 & ~w28492;
assign w29063 = ~pi0868 & w28492;
assign w29064 = ~w29062 & ~w29063;
assign w29065 = pi1563 & ~w28492;
assign w29066 = ~pi0829 & w28492;
assign w29067 = ~w29065 & ~w29066;
assign w29068 = pi1564 & ~w28492;
assign w29069 = ~pi0149 & w28492;
assign w29070 = ~w29068 & ~w29069;
assign w29071 = pi1565 & ~w28496;
assign w29072 = ~pi0830 & w28496;
assign w29073 = ~w29071 & ~w29072;
assign w29074 = pi1566 & ~w28496;
assign w29075 = ~pi0586 & w28496;
assign w29076 = ~w29074 & ~w29075;
assign w29077 = pi1567 & ~w28496;
assign w29078 = pi3633 & w28496;
assign w29079 = ~w29077 & ~w29078;
assign w29080 = pi1568 & ~w28496;
assign w29081 = ~pi0143 & w28496;
assign w29082 = ~w29080 & ~w29081;
assign w29083 = pi1569 & ~w28496;
assign w29084 = ~pi0196 & w28496;
assign w29085 = ~w29083 & ~w29084;
assign w29086 = pi1570 & ~w28496;
assign w29087 = ~pi0152 & w28496;
assign w29088 = ~w29086 & ~w29087;
assign w29089 = pi1571 & ~w28496;
assign w29090 = ~pi0912 & w28496;
assign w29091 = ~w29089 & ~w29090;
assign w29092 = pi1572 & ~w28496;
assign w29093 = ~pi0914 & w28496;
assign w29094 = ~w29092 & ~w29093;
assign w29095 = pi1573 & ~w28496;
assign w29096 = ~pi0916 & w28496;
assign w29097 = ~w29095 & ~w29096;
assign w29098 = pi1574 & ~w28496;
assign w29099 = ~pi0917 & w28496;
assign w29100 = ~w29098 & ~w29099;
assign w29101 = pi1575 & ~w28496;
assign w29102 = ~pi0918 & w28496;
assign w29103 = ~w29101 & ~w29102;
assign w29104 = pi1576 & ~w28496;
assign w29105 = ~pi0980 & w28496;
assign w29106 = ~w29104 & ~w29105;
assign w29107 = pi1577 & ~w28496;
assign w29108 = ~pi0827 & w28496;
assign w29109 = ~w29107 & ~w29108;
assign w29110 = pi1578 & ~w28496;
assign w29111 = ~pi0828 & w28496;
assign w29112 = ~w29110 & ~w29111;
assign w29113 = pi1579 & ~w28496;
assign w29114 = ~pi0829 & w28496;
assign w29115 = ~w29113 & ~w29114;
assign w29116 = pi1580 & ~w28496;
assign w29117 = ~pi0149 & w28496;
assign w29118 = ~w29116 & ~w29117;
assign w29119 = pi1581 & ~w28500;
assign w29120 = ~pi0979 & w28500;
assign w29121 = ~w29119 & ~w29120;
assign w29122 = pi1582 & ~w28500;
assign w29123 = pi3633 & w28500;
assign w29124 = ~w29122 & ~w29123;
assign w29125 = pi1583 & ~w28500;
assign w29126 = ~pi0659 & w28500;
assign w29127 = ~w29125 & ~w29126;
assign w29128 = pi1584 & ~w28500;
assign w29129 = ~pi0196 & w28500;
assign w29130 = ~w29128 & ~w29129;
assign w29131 = pi1585 & ~w28500;
assign w29132 = ~pi0152 & w28500;
assign w29133 = ~w29131 & ~w29132;
assign w29134 = pi1586 & ~w28500;
assign w29135 = ~pi0913 & w28500;
assign w29136 = ~w29134 & ~w29135;
assign w29137 = pi1587 & ~w28500;
assign w29138 = ~pi0915 & w28500;
assign w29139 = ~w29137 & ~w29138;
assign w29140 = pi1588 & ~w28500;
assign w29141 = ~pi0134 & w28500;
assign w29142 = ~w29140 & ~w29141;
assign w29143 = pi1589 & ~w28500;
assign w29144 = ~pi0917 & w28500;
assign w29145 = ~w29143 & ~w29144;
assign w29146 = pi1590 & ~w28500;
assign w29147 = ~pi0708 & w28500;
assign w29148 = ~w29146 & ~w29147;
assign w29149 = pi1591 & ~w28500;
assign w29150 = ~pi0919 & w28500;
assign w29151 = ~w29149 & ~w29150;
assign w29152 = pi1592 & ~w28500;
assign w29153 = ~pi0980 & w28500;
assign w29154 = ~w29152 & ~w29153;
assign w29155 = pi1593 & ~w28500;
assign w29156 = ~pi0826 & w28500;
assign w29157 = ~w29155 & ~w29156;
assign w29158 = pi1594 & ~w28500;
assign w29159 = ~pi0868 & w28500;
assign w29160 = ~w29158 & ~w29159;
assign w29161 = pi1595 & ~w28500;
assign w29162 = ~pi0829 & w28500;
assign w29163 = ~w29161 & ~w29162;
assign w29164 = pi1596 & pi2564;
assign w29165 = pi3137 & ~w29164;
assign w29166 = ~pi1596 & ~pi2564;
assign w29167 = ~w29165 & ~w29166;
assign w29168 = pi1597 & ~w23792;
assign w29169 = w23802 & w23803;
assign w29170 = w27127 & w29169;
assign w29171 = ~w29168 & ~w29170;
assign w29172 = pi1598 & ~w23792;
assign w29173 = w23794 & w23806;
assign w29174 = w27127 & w29173;
assign w29175 = ~w29172 & ~w29174;
assign w29176 = ~w343 & w21954;
assign w29177 = pi1599 & w343;
assign w29178 = ~w29176 & ~w29177;
assign w29179 = pi1600 & w343;
assign w29180 = w21962 & w24132;
assign w29181 = ~w29179 & ~w29180;
assign w29182 = pi1601 & pi3252;
assign w29183 = ~pi2505 & ~pi2522;
assign w29184 = ~w151 & w29183;
assign w29185 = ~w132 & ~w143;
assign w29186 = ~w126 & w150;
assign w29187 = ~w148 & ~w29186;
assign w29188 = ~w29185 & ~w29187;
assign w29189 = ~w29184 & w29188;
assign w29190 = ~w149 & ~w29183;
assign w29191 = ~pi2049 & ~w29190;
assign w29192 = w148 & ~w29191;
assign w29193 = w131 & ~w145;
assign w29194 = ~w29192 & w29193;
assign w29195 = w29189 & w29194;
assign w29196 = ~w29182 & ~w29195;
assign w29197 = w3195 & w23862;
assign w29198 = ~pi1602 & ~w23871;
assign w29199 = ~w23862 & ~w23872;
assign w29200 = ~w29198 & w29199;
assign w29201 = ~w29197 & ~w29200;
assign w29202 = w6413 & w23862;
assign w29203 = ~pi1603 & ~w23869;
assign w29204 = ~w23870 & ~w29203;
assign w29205 = ~w23862 & w29204;
assign w29206 = ~w29202 & ~w29205;
assign w29207 = ~pi1673 & w26759;
assign w29208 = ~pi1672 & w29207;
assign w29209 = ~pi1604 & w29208;
assign w29210 = pi1604 & ~w29208;
assign w29211 = ~w29209 & ~w29210;
assign w29212 = ~pi1434 & w23034;
assign w29213 = pi1605 & pi3641;
assign w29214 = ~pi1605 & ~pi3641;
assign w29215 = ~w29213 & ~w29214;
assign w29216 = ~w23034 & w29215;
assign w29217 = ~w29212 & ~w29216;
assign w29218 = ~pi1431 & w23034;
assign w29219 = pi1681 & w29213;
assign w29220 = pi1704 & w29219;
assign w29221 = ~pi1606 & ~w29220;
assign w29222 = ~w18319 & ~w29221;
assign w29223 = ~w23034 & w29222;
assign w29224 = ~w29218 & ~w29223;
assign w29225 = ~pi0950 & w27425;
assign w29226 = ~pi1847 & w27429;
assign w29227 = ~pi1846 & w29226;
assign w29228 = ~pi1702 & w29227;
assign w29229 = w27396 & w29228;
assign w29230 = ~pi1607 & ~w29229;
assign w29231 = pi1607 & w29229;
assign w29232 = ~w29230 & ~w29231;
assign w29233 = ~w27425 & w29232;
assign w29234 = ~w29225 & ~w29233;
assign w29235 = pi0965 & w28384;
assign w29236 = w28353 & w28387;
assign w29237 = pi1608 & w29236;
assign w29238 = ~pi1608 & ~w29236;
assign w29239 = ~w29237 & ~w29238;
assign w29240 = ~w28349 & ~w29239;
assign w29241 = ~w28384 & w29240;
assign w29242 = ~w29235 & ~w29241;
assign w29243 = ~pi1609 & w28452;
assign w29244 = pi1609 & ~w28452;
assign w29245 = ~w29243 & ~w29244;
assign w29246 = pi1610 & ~w27241;
assign w29247 = pi1074 & w27242;
assign w29248 = ~w29246 & ~w29247;
assign w29249 = pi1611 & ~w28500;
assign w29250 = ~pi0830 & w28500;
assign w29251 = ~w29249 & ~w29250;
assign w29252 = pi1612 & ~w28507;
assign w29253 = ~pi0143 & w28507;
assign w29254 = ~w29252 & ~w29253;
assign w29255 = pi1613 & ~w28500;
assign w29256 = ~pi0143 & w28500;
assign w29257 = ~w29255 & ~w29256;
assign w29258 = pi1614 & ~w28500;
assign w29259 = ~pi0586 & w28500;
assign w29260 = ~w29258 & ~w29259;
assign w29261 = pi1615 & ~w28507;
assign w29262 = ~pi0830 & w28507;
assign w29263 = ~w29261 & ~w29262;
assign w29264 = pi1616 & ~w28496;
assign w29265 = ~pi0868 & w28496;
assign w29266 = ~w29264 & ~w29265;
assign w29267 = pi1617 & ~w28768;
assign w29268 = ~pi0868 & w28768;
assign w29269 = ~w29267 & ~w29268;
assign w29270 = pi1618 & ~w28496;
assign w29271 = ~pi0913 & w28496;
assign w29272 = ~w29270 & ~w29271;
assign w29273 = pi1619 & ~w28496;
assign w29274 = ~pi0708 & w28496;
assign w29275 = ~w29273 & ~w29274;
assign w29276 = pi1620 & ~w28768;
assign w29277 = ~pi0134 & w28768;
assign w29278 = ~w29276 & ~w29277;
assign w29279 = pi1621 & ~w28496;
assign w29280 = ~pi0826 & w28496;
assign w29281 = ~w29279 & ~w29280;
assign w29282 = pi1622 & ~w28768;
assign w29283 = ~pi0919 & w28768;
assign w29284 = ~w29282 & ~w29283;
assign w29285 = pi1623 & ~w28496;
assign w29286 = ~pi0919 & w28496;
assign w29287 = ~w29285 & ~w29286;
assign w29288 = pi1624 & ~w28768;
assign w29289 = ~pi0708 & w28768;
assign w29290 = ~w29288 & ~w29289;
assign w29291 = pi1625 & ~w28496;
assign w29292 = ~pi0134 & w28496;
assign w29293 = ~w29291 & ~w29292;
assign w29294 = pi1626 & ~w28768;
assign w29295 = ~pi0659 & w28768;
assign w29296 = ~w29294 & ~w29295;
assign w29297 = pi1627 & ~w28768;
assign w29298 = ~pi0913 & w28768;
assign w29299 = ~w29297 & ~w29298;
assign w29300 = pi1628 & ~w28496;
assign w29301 = ~pi0915 & w28496;
assign w29302 = ~w29300 & ~w29301;
assign w29303 = ~pi0798 & w28384;
assign w29304 = ~pi1848 & w28388;
assign w29305 = ~pi1849 & w29304;
assign w29306 = ~pi1629 & w29305;
assign w29307 = pi1629 & ~w29305;
assign w29308 = ~w29306 & ~w29307;
assign w29309 = ~w28384 & w29308;
assign w29310 = ~w29303 & ~w29309;
assign w29311 = w21060 & w23003;
assign w29312 = pi1630 & ~w29311;
assign w29313 = ~pi0632 & w29311;
assign w29314 = ~w29312 & ~w29313;
assign w29315 = pi1631 & ~w29311;
assign w29316 = ~pi0593 & w29311;
assign w29317 = ~w29315 & ~w29316;
assign w29318 = pi1632 & ~w29311;
assign w29319 = ~pi0594 & w29311;
assign w29320 = ~w29318 & ~w29319;
assign w29321 = pi1633 & ~w29311;
assign w29322 = ~pi0571 & w29311;
assign w29323 = ~w29321 & ~w29322;
assign w29324 = pi0647 & w23004;
assign w29325 = pi1634 & ~w29324;
assign w29326 = ~pi0594 & w29324;
assign w29327 = ~w29325 & ~w29326;
assign w29328 = pi1635 & ~w29311;
assign w29329 = ~pi0590 & w29311;
assign w29330 = ~w29328 & ~w29329;
assign w29331 = pi1636 & ~w29324;
assign w29332 = ~pi0593 & w29324;
assign w29333 = ~w29331 & ~w29332;
assign w29334 = pi1637 & ~w29324;
assign w29335 = ~pi0603 & w29324;
assign w29336 = ~w29334 & ~w29335;
assign w29337 = pi1638 & ~w29324;
assign w29338 = ~pi0632 & w29324;
assign w29339 = ~w29337 & ~w29338;
assign w29340 = pi1639 & ~w29324;
assign w29341 = ~pi0571 & w29324;
assign w29342 = ~w29340 & ~w29341;
assign w29343 = ~pi1640 & ~w14887;
assign w29344 = ~w14366 & w14887;
assign w29345 = pi0423 & w29344;
assign w29346 = ~w29343 & ~w29345;
assign w29347 = ~pi3395 & ~pi3638;
assign w29348 = ~w18003 & ~w18007;
assign w29349 = ~pi0955 & ~w29348;
assign w29350 = ~w18366 & ~w29349;
assign w29351 = pi1447 & pi3635;
assign w29352 = ~w29350 & w29351;
assign w29353 = ~pi1642 & ~w29352;
assign w29354 = pi1643 & ~w28413;
assign w29355 = ~w28414 & ~w29354;
assign w29356 = ~w28452 & w29355;
assign w29357 = ~pi0900 & w28384;
assign w29358 = ~w28349 & w29236;
assign w29359 = ~pi1687 & w29306;
assign w29360 = ~pi1644 & ~w29359;
assign w29361 = ~w29358 & ~w29360;
assign w29362 = ~w28384 & w29361;
assign w29363 = ~w29357 & ~w29362;
assign w29364 = pi1645 & ~w26743;
assign w29365 = ~w26744 & ~w29364;
assign w29366 = pi1646 & ~w28452;
assign w29367 = ~pi1647 & ~w14887;
assign w29368 = pi0424 & w29344;
assign w29369 = ~w29367 & ~w29368;
assign w29370 = ~pi0964 & w28384;
assign w29371 = pi1648 & w29237;
assign w29372 = ~pi1686 & w29371;
assign w29373 = ~pi1648 & ~w29237;
assign w29374 = ~w29372 & ~w29373;
assign w29375 = ~w28384 & w29374;
assign w29376 = ~w29370 & ~w29375;
assign w29377 = pi1649 & ~w28417;
assign w29378 = ~w28418 & ~w28452;
assign w29379 = ~w29377 & w29378;
assign w29380 = pi1650 & ~w29324;
assign w29381 = ~pi0590 & w29324;
assign w29382 = ~w29380 & ~w29381;
assign w29383 = pi1651 & ~w29324;
assign w29384 = ~pi0602 & w29324;
assign w29385 = ~w29383 & ~w29384;
assign w29386 = pi1652 & ~w29324;
assign w29387 = ~pi0572 & w29324;
assign w29388 = ~w29386 & ~w29387;
assign w29389 = pi1653 & ~w29324;
assign w29390 = ~pi0591 & w29324;
assign w29391 = ~w29389 & ~w29390;
assign w29392 = pi1654 & ~w29324;
assign w29393 = ~pi0592 & w29324;
assign w29394 = ~w29392 & ~w29393;
assign w29395 = pi1655 & ~w29324;
assign w29396 = ~pi0573 & w29324;
assign w29397 = ~w29395 & ~w29396;
assign w29398 = pi1656 & ~w29324;
assign w29399 = ~pi0595 & w29324;
assign w29400 = ~w29398 & ~w29399;
assign w29401 = pi1657 & ~w29324;
assign w29402 = ~pi0585 & w29324;
assign w29403 = ~w29401 & ~w29402;
assign w29404 = pi1658 & ~w29311;
assign w29405 = ~pi0602 & w29311;
assign w29406 = ~w29404 & ~w29405;
assign w29407 = pi1659 & ~w29311;
assign w29408 = ~pi0572 & w29311;
assign w29409 = ~w29407 & ~w29408;
assign w29410 = pi1660 & ~w29311;
assign w29411 = ~pi0591 & w29311;
assign w29412 = ~w29410 & ~w29411;
assign w29413 = pi1661 & ~w29311;
assign w29414 = ~pi0603 & w29311;
assign w29415 = ~w29413 & ~w29414;
assign w29416 = pi1662 & ~w29311;
assign w29417 = ~pi0592 & w29311;
assign w29418 = ~w29416 & ~w29417;
assign w29419 = pi1663 & ~w29311;
assign w29420 = ~pi0573 & w29311;
assign w29421 = ~w29419 & ~w29420;
assign w29422 = pi1664 & ~w29311;
assign w29423 = ~pi0595 & w29311;
assign w29424 = ~w29422 & ~w29423;
assign w29425 = pi1665 & ~w29311;
assign w29426 = ~pi0585 & w29311;
assign w29427 = ~w29425 & ~w29426;
assign w29428 = ~pi1666 & w6684;
assign w29429 = pi0420 & ~w375;
assign w29430 = w22020 & ~w29429;
assign w29431 = ~w29428 & ~w29430;
assign w29432 = ~pi1667 & w6684;
assign w29433 = w22020 & w29429;
assign w29434 = ~w29432 & ~w29433;
assign w29435 = pi1668 & ~w27277;
assign w29436 = ~w27278 & ~w29435;
assign w29437 = pi1669 & ~w26751;
assign w29438 = ~w26752 & ~w29437;
assign w29439 = pi1670 & ~w26742;
assign w29440 = ~w26743 & ~w29439;
assign w29441 = pi1671 & ~w26754;
assign w29442 = ~w26755 & ~w29441;
assign w29443 = pi1672 & ~w29207;
assign w29444 = ~w29208 & ~w29443;
assign w29445 = pi1673 & ~w26759;
assign w29446 = ~w29207 & ~w29445;
assign w29447 = pi1674 & ~w27237;
assign w29448 = ~w27241 & ~w29447;
assign w29449 = ~w26739 & ~w29448;
assign w29450 = pi1675 & ~w26744;
assign w29451 = ~w26745 & ~w29450;
assign w29452 = ~pi1676 & w26745;
assign w29453 = pi1676 & ~w26745;
assign w29454 = ~w29452 & ~w29453;
assign w29455 = pi1677 & ~w29452;
assign w29456 = ~w26746 & ~w29455;
assign w29457 = pi1678 & ~w26747;
assign w29458 = ~w26748 & ~w29457;
assign w29459 = pi1679 & ~w26748;
assign w29460 = ~w26749 & ~w29459;
assign w29461 = pi1680 & ~w26749;
assign w29462 = ~w26750 & ~w29461;
assign w29463 = ~pi1433 & w23034;
assign w29464 = ~pi1681 & ~w29213;
assign w29465 = ~w29219 & ~w29464;
assign w29466 = ~w23034 & w29465;
assign w29467 = ~w29463 & ~w29466;
assign w29468 = pi0948 & w27425;
assign w29469 = pi1683 & w29231;
assign w29470 = ~w27425 & ~w29469;
assign w29471 = ~pi1682 & w29470;
assign w29472 = ~w29468 & ~w29471;
assign w29473 = ~pi1683 & ~w29231;
assign w29474 = w29470 & ~w29473;
assign w29475 = ~pi0949 & w27425;
assign w29476 = ~w29474 & ~w29475;
assign w29477 = ~pi0891 & w27425;
assign w29478 = ~pi1684 & w29228;
assign w29479 = pi1684 & ~w29228;
assign w29480 = ~w29478 & ~w29479;
assign w29481 = ~w27425 & w29480;
assign w29482 = ~w29477 & ~w29481;
assign w29483 = pi0890 & w22580;
assign w29484 = pi0963 & w28384;
assign w29485 = ~pi1686 & ~w29371;
assign w29486 = ~w28384 & w29485;
assign w29487 = ~w29484 & ~w29486;
assign w29488 = ~pi0797 & w28384;
assign w29489 = pi1687 & ~w29306;
assign w29490 = ~w29359 & ~w29489;
assign w29491 = ~w28384 & w29490;
assign w29492 = ~w29488 & ~w29491;
assign w29493 = pi0796 & w22670;
assign w29494 = pi1689 & ~w28419;
assign w29495 = ~w28420 & ~w28452;
assign w29496 = ~w29494 & w29495;
assign w29497 = pi1690 & ~w28418;
assign w29498 = ~w28419 & ~w28452;
assign w29499 = ~w29497 & w29498;
assign w29500 = pi1691 & ~w28415;
assign w29501 = ~w28416 & ~w28452;
assign w29502 = ~w29500 & w29501;
assign w29503 = pi1692 & ~w28414;
assign w29504 = ~w28415 & ~w29503;
assign w29505 = ~w28452 & w29504;
assign w29506 = pi1693 & ~w28416;
assign w29507 = ~w28417 & ~w28452;
assign w29508 = ~w29506 & w29507;
assign w29509 = pi1694 & ~w28412;
assign w29510 = ~w28413 & ~w29509;
assign w29511 = ~w28452 & w29510;
assign w29512 = pi1695 & ~w27276;
assign w29513 = ~w27277 & ~w29512;
assign w29514 = pi1698 & ~w26750;
assign w29515 = ~w26751 & ~w29514;
assign w29516 = pi1699 & ~w26746;
assign w29517 = ~w26747 & ~w29516;
assign w29518 = pi1700 & ~w26755;
assign w29519 = ~w26756 & ~w29518;
assign w29520 = pi1701 & ~w26752;
assign w29521 = ~w26753 & ~w29520;
assign w29522 = ~pi0892 & w27425;
assign w29523 = pi1702 & ~w29227;
assign w29524 = ~w29228 & ~w29523;
assign w29525 = ~w27425 & w29524;
assign w29526 = ~w29522 & ~w29525;
assign w29527 = ~pi0951 & w27425;
assign w29528 = ~pi1703 & ~w29478;
assign w29529 = ~w29229 & ~w29528;
assign w29530 = ~w27425 & w29529;
assign w29531 = ~w29527 & ~w29530;
assign w29532 = ~pi1432 & w23034;
assign w29533 = ~pi1704 & ~w29219;
assign w29534 = ~w29220 & ~w29533;
assign w29535 = ~w23034 & w29534;
assign w29536 = ~w29532 & ~w29535;
assign w29537 = pi1012 & w24334;
assign w29538 = pi1705 & ~w29537;
assign w29539 = w5053 & w29537;
assign w29540 = ~w29538 & ~w29539;
assign w29541 = pi1033 & w1236;
assign w29542 = w24322 & w29541;
assign w29543 = pi1706 & ~w29542;
assign w29544 = w3195 & w29542;
assign w29545 = ~w29543 & ~w29544;
assign w29546 = pi1707 & ~w23322;
assign w29547 = ~pi0603 & w23322;
assign w29548 = ~w29546 & ~w29547;
assign w29549 = pi1708 & ~w23322;
assign w29550 = ~pi0571 & w23322;
assign w29551 = ~w29549 & ~w29550;
assign w29552 = pi1709 & ~w29311;
assign w29553 = ~pi0578 & w29311;
assign w29554 = ~w29552 & ~w29553;
assign w29555 = w21062 & w23003;
assign w29556 = pi1710 & ~w29555;
assign w29557 = ~pi0594 & w29555;
assign w29558 = ~w29556 & ~w29557;
assign w29559 = pi1711 & ~w29555;
assign w29560 = ~pi0632 & w29555;
assign w29561 = ~w29559 & ~w29560;
assign w29562 = pi1712 & ~w29555;
assign w29563 = ~pi0590 & w29555;
assign w29564 = ~w29562 & ~w29563;
assign w29565 = pi2383 & ~w7009;
assign w29566 = ~w370 & ~w29565;
assign w29567 = ~pi1797 & w29566;
assign w29568 = pi3191 & w29567;
assign w29569 = ~pi1713 & ~w29568;
assign w29570 = pi1713 & ~pi1797;
assign w29571 = ~pi1798 & ~w29570;
assign w29572 = ~w29569 & w29571;
assign w29573 = ~pi3191 & ~w370;
assign w29574 = ~w29570 & w29573;
assign w29575 = ~w29567 & ~w29574;
assign w29576 = pi1713 & w29575;
assign w29577 = ~pi1798 & ~w29573;
assign w29578 = w29570 & ~w29577;
assign w29579 = w6760 & w29573;
assign w29580 = ~w29578 & ~w29579;
assign w29581 = ~w29576 & w29580;
assign w29582 = ~w29572 & w29581;
assign w29583 = ~pi1897 & pi2555;
assign w29584 = ~w5635 & ~w15388;
assign w29585 = ~pi1714 & w15388;
assign w29586 = ~pi2555 & ~w29585;
assign w29587 = ~w29584 & w29586;
assign w29588 = ~w29583 & ~w29587;
assign w29589 = pi1715 & ~w25734;
assign w29590 = ~w25735 & w25801;
assign w29591 = ~w29589 & w29590;
assign w29592 = pi1716 & ~w29542;
assign w29593 = w40134 & w29542;
assign w29594 = ~w29592 & ~w29593;
assign w29595 = pi1717 & ~w29542;
assign w29596 = w6413 & w29542;
assign w29597 = ~w29595 & ~w29596;
assign w29598 = pi1718 & ~w29542;
assign w29599 = w4380 & w29542;
assign w29600 = ~w29598 & ~w29599;
assign w29601 = pi1719 & ~w29542;
assign w29602 = w5320 & w29542;
assign w29603 = ~w29601 & ~w29602;
assign w29604 = pi1720 & ~w29542;
assign w29605 = w5914 & w29542;
assign w29606 = ~w29604 & ~w29605;
assign w29607 = pi1721 & ~w29542;
assign w29608 = w4749 & w29542;
assign w29609 = ~w29607 & ~w29608;
assign w29610 = pi1722 & ~w29542;
assign w29611 = w8240 & w29542;
assign w29612 = ~w29610 & ~w29611;
assign w29613 = pi1723 & ~w29542;
assign w29614 = w8081 & w29542;
assign w29615 = ~w29613 & ~w29614;
assign w29616 = pi1724 & ~w29542;
assign w29617 = w5635 & w29542;
assign w29618 = ~w29616 & ~w29617;
assign w29619 = pi1725 & ~w29542;
assign w29620 = w5053 & w29542;
assign w29621 = ~w29619 & ~w29620;
assign w29622 = pi1726 & ~w29542;
assign w29623 = w3711 & w29542;
assign w29624 = ~w29622 & ~w29623;
assign w29625 = pi0609 & w3144;
assign w29626 = w24681 & w29625;
assign w29627 = pi1727 & ~w29626;
assign w29628 = w4141 & w29626;
assign w29629 = ~w29627 & ~w29628;
assign w29630 = pi1728 & ~w29626;
assign w29631 = w6177 & w29626;
assign w29632 = ~w29630 & ~w29631;
assign w29633 = pi1729 & ~w29626;
assign w29634 = w3195 & w29626;
assign w29635 = ~w29633 & ~w29634;
assign w29636 = pi1730 & ~w29626;
assign w29637 = w40134 & w29626;
assign w29638 = ~w29636 & ~w29637;
assign w29639 = pi1731 & ~w29626;
assign w29640 = w6413 & w29626;
assign w29641 = ~w29639 & ~w29640;
assign w29642 = pi1732 & ~w29626;
assign w29643 = w4380 & w29626;
assign w29644 = ~w29642 & ~w29643;
assign w29645 = pi1733 & ~w29626;
assign w29646 = w5320 & w29626;
assign w29647 = ~w29645 & ~w29646;
assign w29648 = pi1734 & ~w29626;
assign w29649 = w5914 & w29626;
assign w29650 = ~w29648 & ~w29649;
assign w29651 = pi1735 & ~w29626;
assign w29652 = w4749 & w29626;
assign w29653 = ~w29651 & ~w29652;
assign w29654 = pi1736 & ~w29626;
assign w29655 = w5635 & w29626;
assign w29656 = ~w29654 & ~w29655;
assign w29657 = pi1737 & ~w29626;
assign w29658 = w5053 & w29626;
assign w29659 = ~w29657 & ~w29658;
assign w29660 = pi1738 & ~w29626;
assign w29661 = w3711 & w29626;
assign w29662 = ~w29660 & ~w29661;
assign w29663 = ~pi1739 & w25801;
assign w29664 = pi1739 & ~w25801;
assign w29665 = ~w29663 & ~w29664;
assign w29666 = pi1740 & ~w25728;
assign w29667 = ~w25729 & w25801;
assign w29668 = ~w29666 & w29667;
assign w29669 = ~w6177 & ~w15388;
assign w29670 = ~pi1741 & w15388;
assign w29671 = ~pi2555 & ~w29670;
assign w29672 = ~w29669 & w29671;
assign w29673 = ~w29583 & ~w29672;
assign w29674 = ~w4141 & ~w15388;
assign w29675 = ~pi1742 & w15388;
assign w29676 = ~pi2555 & ~w29675;
assign w29677 = ~w29674 & w29676;
assign w29678 = ~w29583 & ~w29677;
assign w29679 = ~w1639 & ~w15388;
assign w29680 = ~pi1743 & w15388;
assign w29681 = ~pi2555 & ~w29680;
assign w29682 = ~w29679 & w29681;
assign w29683 = ~w29583 & ~w29682;
assign w29684 = ~w1308 & ~w15388;
assign w29685 = ~pi1744 & w15388;
assign w29686 = ~pi2555 & ~w29685;
assign w29687 = ~w29684 & w29686;
assign w29688 = ~w29583 & ~w29687;
assign w29689 = ~w5053 & ~w15388;
assign w29690 = ~pi1745 & w15388;
assign w29691 = ~pi2555 & ~w29690;
assign w29692 = ~w29689 & w29691;
assign w29693 = ~w29583 & ~w29692;
assign w29694 = ~pi1746 & w25889;
assign w29695 = pi1746 & ~w25889;
assign w29696 = ~w29694 & ~w29695;
assign w29697 = pi1747 & ~w25822;
assign w29698 = ~w25823 & w25889;
assign w29699 = ~w29697 & w29698;
assign w29700 = pi1748 & ~w25816;
assign w29701 = ~w25817 & w25889;
assign w29702 = ~w29700 & w29701;
assign w29703 = pi0609 & w1216;
assign w29704 = w23838 & w29703;
assign w29705 = w1236 & w29704;
assign w29706 = pi1749 & ~w29705;
assign w29707 = w1639 & w29705;
assign w29708 = ~w29706 & ~w29707;
assign w29709 = pi1750 & ~w29705;
assign w29710 = w1308 & w29705;
assign w29711 = ~w29709 & ~w29710;
assign w29712 = pi1751 & ~w29705;
assign w29713 = w3195 & w29705;
assign w29714 = ~w29712 & ~w29713;
assign w29715 = pi1752 & ~w29705;
assign w29716 = w40134 & w29705;
assign w29717 = ~w29715 & ~w29716;
assign w29718 = pi1753 & ~w29705;
assign w29719 = w6413 & w29705;
assign w29720 = ~w29718 & ~w29719;
assign w29721 = pi1754 & ~w29705;
assign w29722 = w4380 & w29705;
assign w29723 = ~w29721 & ~w29722;
assign w29724 = pi1755 & ~w29705;
assign w29725 = w5320 & w29705;
assign w29726 = ~w29724 & ~w29725;
assign w29727 = pi1756 & ~w29705;
assign w29728 = w5914 & w29705;
assign w29729 = ~w29727 & ~w29728;
assign w29730 = pi1757 & ~w29705;
assign w29731 = w4749 & w29705;
assign w29732 = ~w29730 & ~w29731;
assign w29733 = pi1758 & ~w29705;
assign w29734 = w8240 & w29705;
assign w29735 = ~w29733 & ~w29734;
assign w29736 = pi1759 & ~w29705;
assign w29737 = w8081 & w29705;
assign w29738 = ~w29736 & ~w29737;
assign w29739 = pi1760 & ~w29705;
assign w29740 = w3711 & w29705;
assign w29741 = ~w29739 & ~w29740;
assign w29742 = w1222 & w29704;
assign w29743 = pi1761 & ~w29742;
assign w29744 = w1639 & w29742;
assign w29745 = ~w29743 & ~w29744;
assign w29746 = pi1762 & ~w29742;
assign w29747 = w1308 & w29742;
assign w29748 = ~w29746 & ~w29747;
assign w29749 = pi1763 & ~w29742;
assign w29750 = w40134 & w29742;
assign w29751 = ~w29749 & ~w29750;
assign w29752 = pi1764 & ~w29742;
assign w29753 = w6413 & w29742;
assign w29754 = ~w29752 & ~w29753;
assign w29755 = pi1765 & ~w29742;
assign w29756 = w4380 & w29742;
assign w29757 = ~w29755 & ~w29756;
assign w29758 = pi1766 & ~w29742;
assign w29759 = w5914 & w29742;
assign w29760 = ~w29758 & ~w29759;
assign w29761 = pi1767 & ~w29742;
assign w29762 = w4749 & w29742;
assign w29763 = ~w29761 & ~w29762;
assign w29764 = pi1768 & ~w29742;
assign w29765 = w8240 & w29742;
assign w29766 = ~w29764 & ~w29765;
assign w29767 = pi1769 & ~w29742;
assign w29768 = w3711 & w29742;
assign w29769 = ~w29767 & ~w29768;
assign w29770 = w19033 & ~w20671;
assign w29771 = pi3572 & pi3645;
assign w29772 = w29770 & w29771;
assign w29773 = ~pi1923 & w29772;
assign w29774 = pi2515 & w29770;
assign w29775 = pi1855 & w29774;
assign w29776 = pi1770 & w29775;
assign w29777 = ~pi1770 & ~w29775;
assign w29778 = ~w29772 & ~w29777;
assign w29779 = ~w29776 & w29778;
assign w29780 = ~w29773 & ~w29779;
assign w29781 = pi3440 & pi3507;
assign w29782 = ~pi1771 & ~w29771;
assign w29783 = ~w29781 & w29782;
assign w29784 = w24810 & ~w29783;
assign w29785 = pi1033 & w1222;
assign w29786 = w24671 & w29785;
assign w29787 = pi1772 & ~w29786;
assign w29788 = w4141 & w29786;
assign w29789 = ~w29787 & ~w29788;
assign w29790 = pi1773 & ~w29786;
assign w29791 = w6177 & w29786;
assign w29792 = ~w29790 & ~w29791;
assign w29793 = pi1774 & ~w29786;
assign w29794 = w3195 & w29786;
assign w29795 = ~w29793 & ~w29794;
assign w29796 = pi1775 & ~w29786;
assign w29797 = w40134 & w29786;
assign w29798 = ~w29796 & ~w29797;
assign w29799 = pi1776 & ~w29786;
assign w29800 = w6413 & w29786;
assign w29801 = ~w29799 & ~w29800;
assign w29802 = pi1777 & ~w29786;
assign w29803 = w4380 & w29786;
assign w29804 = ~w29802 & ~w29803;
assign w29805 = pi1778 & ~w29786;
assign w29806 = w5320 & w29786;
assign w29807 = ~w29805 & ~w29806;
assign w29808 = pi1779 & ~w29786;
assign w29809 = w5914 & w29786;
assign w29810 = ~w29808 & ~w29809;
assign w29811 = pi1780 & ~w29786;
assign w29812 = w4749 & w29786;
assign w29813 = ~w29811 & ~w29812;
assign w29814 = pi1781 & ~w29786;
assign w29815 = w8081 & w29786;
assign w29816 = ~w29814 & ~w29815;
assign w29817 = pi1782 & ~w29786;
assign w29818 = w1639 & w29786;
assign w29819 = ~w29817 & ~w29818;
assign w29820 = pi1783 & ~w29786;
assign w29821 = w1308 & w29786;
assign w29822 = ~w29820 & ~w29821;
assign w29823 = pi1784 & ~w29786;
assign w29824 = w5635 & w29786;
assign w29825 = ~w29823 & ~w29824;
assign w29826 = pi1785 & ~w29786;
assign w29827 = w5053 & w29786;
assign w29828 = ~w29826 & ~w29827;
assign w29829 = pi1786 & ~w29786;
assign w29830 = w3711 & w29786;
assign w29831 = ~w29829 & ~w29830;
assign w29832 = pi3257 & w117;
assign w29833 = ~pi2779 & ~w29832;
assign w29834 = ~w28753 & ~w29833;
assign w29835 = ~w343 & ~w28745;
assign w29836 = pi1787 & ~w29835;
assign w29837 = w28753 & w29836;
assign w29838 = ~w29834 & ~w29837;
assign w29839 = pi1788 & ~w27279;
assign w29840 = ~w27280 & ~w29839;
assign w29841 = pi1789 & ~w14887;
assign w29842 = ~w29344 & ~w29841;
assign w29843 = w4749 & w14856;
assign w29844 = ~w15116 & ~w29843;
assign w29845 = ~w17425 & w29844;
assign w29846 = w3593 & w17425;
assign w29847 = ~w29845 & ~w29846;
assign w29848 = w17421 & ~w29847;
assign w29849 = ~pi1790 & ~w17421;
assign w29850 = ~w29848 & ~w29849;
assign w29851 = w8081 & w14856;
assign w29852 = ~w16647 & ~w29851;
assign w29853 = ~w17425 & w29852;
assign w29854 = w1445 & w17425;
assign w29855 = ~w29853 & ~w29854;
assign w29856 = w17421 & ~w29855;
assign w29857 = ~pi1791 & ~w17421;
assign w29858 = ~w29856 & ~w29857;
assign w29859 = pi1792 & ~w29537;
assign w29860 = w8081 & w29537;
assign w29861 = ~w29859 & ~w29860;
assign w29862 = w7160 & w14360;
assign w29863 = pi0411 & pi0425;
assign w29864 = pi0406 & w29863;
assign w29865 = ~pi0413 & ~w29864;
assign w29866 = w29862 & ~w29865;
assign w29867 = ~w21945 & w29864;
assign w29868 = w29866 & ~w29867;
assign w29869 = ~pi0408 & ~pi0411;
assign w29870 = w21943 & w29869;
assign w29871 = w14359 & ~w29870;
assign w29872 = w7160 & w29871;
assign w29873 = ~pi1793 & ~w29872;
assign w29874 = ~w29868 & ~w29873;
assign w29875 = w21945 & w29864;
assign w29876 = w29866 & ~w29875;
assign w29877 = ~pi1794 & ~w29872;
assign w29878 = ~w29876 & ~w29877;
assign w29879 = ~pi0411 & pi0425;
assign w29880 = pi0406 & w29879;
assign w29881 = ~pi0413 & ~w29880;
assign w29882 = w29862 & ~w29881;
assign w29883 = ~w21945 & w29880;
assign w29884 = w29882 & ~w29883;
assign w29885 = ~pi1795 & ~w29872;
assign w29886 = ~w29884 & ~w29885;
assign w29887 = w21945 & w29880;
assign w29888 = w29882 & ~w29887;
assign w29889 = ~pi1796 & ~w29872;
assign w29890 = ~w29888 & ~w29889;
assign w29891 = pi1713 & w29573;
assign w29892 = pi1797 & ~w29891;
assign w29893 = ~w29572 & ~w29892;
assign w29894 = ~w29567 & w29577;
assign w29895 = pi1798 & ~w29575;
assign w29896 = ~w29894 & ~w29895;
assign w29897 = ~pi1798 & w29891;
assign w29898 = ~pi3330 & w29897;
assign w29899 = pi1799 & ~w29897;
assign w29900 = ~w29898 & ~w29899;
assign w29901 = w6758 & w29573;
assign w29902 = ~pi3330 & w29901;
assign w29903 = pi1800 & ~w29901;
assign w29904 = ~w29902 & ~w29903;
assign w29905 = pi1801 & ~w29555;
assign w29906 = ~pi0602 & w29555;
assign w29907 = ~w29905 & ~w29906;
assign w29908 = pi1802 & ~w29555;
assign w29909 = ~pi0571 & w29555;
assign w29910 = ~w29908 & ~w29909;
assign w29911 = pi1803 & ~w29555;
assign w29912 = ~pi0572 & w29555;
assign w29913 = ~w29911 & ~w29912;
assign w29914 = pi1804 & ~w29555;
assign w29915 = ~pi0591 & w29555;
assign w29916 = ~w29914 & ~w29915;
assign w29917 = pi1805 & ~w29555;
assign w29918 = ~pi0603 & w29555;
assign w29919 = ~w29917 & ~w29918;
assign w29920 = pi1806 & ~w29555;
assign w29921 = ~pi0592 & w29555;
assign w29922 = ~w29920 & ~w29921;
assign w29923 = pi1807 & ~w29555;
assign w29924 = ~pi0573 & w29555;
assign w29925 = ~w29923 & ~w29924;
assign w29926 = pi1808 & ~w29555;
assign w29927 = ~pi0593 & w29555;
assign w29928 = ~w29926 & ~w29927;
assign w29929 = pi1809 & ~w29555;
assign w29930 = ~pi0595 & w29555;
assign w29931 = ~w29929 & ~w29930;
assign w29932 = pi1810 & ~w29555;
assign w29933 = ~pi0585 & w29555;
assign w29934 = ~w29932 & ~w29933;
assign w29935 = pi1811 & ~w29324;
assign w29936 = ~pi0578 & w29324;
assign w29937 = ~w29935 & ~w29936;
assign w29938 = pi1812 & ~w23322;
assign w29939 = ~pi0590 & w23322;
assign w29940 = ~w29938 & ~w29939;
assign w29941 = pi1813 & ~w23322;
assign w29942 = ~pi0602 & w23322;
assign w29943 = ~w29941 & ~w29942;
assign w29944 = pi1814 & ~w23322;
assign w29945 = ~pi0572 & w23322;
assign w29946 = ~w29944 & ~w29945;
assign w29947 = pi1815 & ~w23322;
assign w29948 = ~pi0591 & w23322;
assign w29949 = ~w29947 & ~w29948;
assign w29950 = pi1816 & ~w23322;
assign w29951 = ~pi0592 & w23322;
assign w29952 = ~w29950 & ~w29951;
assign w29953 = pi1817 & ~w23322;
assign w29954 = ~pi0632 & w23322;
assign w29955 = ~w29953 & ~w29954;
assign w29956 = pi1818 & ~w23322;
assign w29957 = ~pi0573 & w23322;
assign w29958 = ~w29956 & ~w29957;
assign w29959 = pi1819 & ~w23322;
assign w29960 = ~pi0595 & w23322;
assign w29961 = ~w29959 & ~w29960;
assign w29962 = pi1820 & ~w23322;
assign w29963 = ~pi0594 & w23322;
assign w29964 = ~w29962 & ~w29963;
assign w29965 = pi1821 & ~w23322;
assign w29966 = ~pi0585 & w23322;
assign w29967 = ~w29965 & ~w29966;
assign w29968 = pi2019 & ~w6682;
assign w29969 = ~pi3443 & ~pi3536;
assign w29970 = pi1822 & pi3374;
assign w29971 = ~w29969 & w29970;
assign w29972 = pi3217 & ~w29971;
assign w29973 = ~w29968 & w29972;
assign w29974 = ~w6970 & ~w19954;
assign w29975 = pi1823 & w19954;
assign w29976 = w6682 & ~w29975;
assign w29977 = ~w29974 & w29976;
assign w29978 = ~w343 & ~w14359;
assign w29979 = w6974 & ~w23334;
assign w29980 = w2233 & w23334;
assign w29981 = ~w382 & ~w29980;
assign w29982 = ~w29979 & w29981;
assign w29983 = w29978 & w29982;
assign w29984 = pi1824 & w343;
assign w29985 = w6682 & ~w29984;
assign w29986 = ~w29983 & w29985;
assign w29987 = pi1930 & ~w19954;
assign w29988 = ~pi1825 & ~w29987;
assign w29989 = w6749 & ~w19954;
assign w29990 = w6729 & w29989;
assign w29991 = ~w29988 & ~w29990;
assign w29992 = w6682 & ~w29991;
assign w29993 = ~pi1826 & ~w29987;
assign w29994 = w7046 & w29989;
assign w29995 = ~w29993 & ~w29994;
assign w29996 = w6682 & ~w29995;
assign w29997 = ~w7050 & w29987;
assign w29998 = pi1827 & ~w29987;
assign w29999 = w6682 & ~w29998;
assign w30000 = ~w29997 & w29999;
assign w30001 = pi1828 & ~w29537;
assign w30002 = w4141 & w29537;
assign w30003 = ~w30001 & ~w30002;
assign w30004 = pi1829 & ~w29537;
assign w30005 = w6177 & w29537;
assign w30006 = ~w30004 & ~w30005;
assign w30007 = pi1830 & ~w29537;
assign w30008 = w3195 & w29537;
assign w30009 = ~w30007 & ~w30008;
assign w30010 = pi1831 & ~w29537;
assign w30011 = w40134 & w29537;
assign w30012 = ~w30010 & ~w30011;
assign w30013 = pi1832 & ~w29537;
assign w30014 = w6413 & w29537;
assign w30015 = ~w30013 & ~w30014;
assign w30016 = pi1833 & ~w29537;
assign w30017 = w4380 & w29537;
assign w30018 = ~w30016 & ~w30017;
assign w30019 = pi1834 & ~w29537;
assign w30020 = w5914 & w29537;
assign w30021 = ~w30019 & ~w30020;
assign w30022 = pi1835 & ~w29537;
assign w30023 = w8240 & w29537;
assign w30024 = ~w30022 & ~w30023;
assign w30025 = pi1836 & ~w29537;
assign w30026 = w1639 & w29537;
assign w30027 = ~w30025 & ~w30026;
assign w30028 = pi1837 & ~w29537;
assign w30029 = w1308 & w29537;
assign w30030 = ~w30028 & ~w30029;
assign w30031 = pi1838 & ~w29537;
assign w30032 = w5635 & w29537;
assign w30033 = ~w30031 & ~w30032;
assign w30034 = pi1839 & ~w29537;
assign w30035 = w3711 & w29537;
assign w30036 = ~w30034 & ~w30035;
assign w30037 = w894 & w22040;
assign w30038 = ~pi1861 & w891;
assign w30039 = w30037 & ~w30038;
assign w30040 = pi1840 & ~w30039;
assign w30041 = ~w903 & w22040;
assign w30042 = w902 & w30041;
assign w30043 = ~w30040 & ~w30042;
assign w30044 = w5320 & w23862;
assign w30045 = ~pi1841 & ~w23867;
assign w30046 = ~w23868 & ~w30045;
assign w30047 = ~w23862 & w30046;
assign w30048 = ~w30044 & ~w30047;
assign w30049 = pi0492 & pi0493;
assign w30050 = pi0497 & ~pi0552;
assign w30051 = ~pi0553 & ~pi0563;
assign w30052 = w30050 & w30051;
assign w30053 = w30049 & w30052;
assign w30054 = w21353 & w30053;
assign w30055 = pi0498 & ~pi0504;
assign w30056 = w30054 & w30055;
assign w30057 = pi1842 & ~w30056;
assign w30058 = w23917 & w30056;
assign w30059 = ~w30057 & ~w30058;
assign w30060 = w21482 & w30054;
assign w30061 = pi1843 & ~w30060;
assign w30062 = w23917 & w30060;
assign w30063 = ~w30061 & ~w30062;
assign w30064 = pi0501 & ~pi0502;
assign w30065 = ~pi0559 & ~pi0561;
assign w30066 = ~pi0564 & w30065;
assign w30067 = w30064 & w30066;
assign w30068 = w21440 & w30067;
assign w30069 = pi0503 & w30068;
assign w30070 = pi1844 & ~w30069;
assign w30071 = ~w23903 & w30069;
assign w30072 = ~w30070 & ~w30071;
assign w30073 = ~pi0503 & w30068;
assign w30074 = pi1845 & ~w30073;
assign w30075 = ~w23903 & w30073;
assign w30076 = ~w30074 & ~w30075;
assign w30077 = ~pi0952 & w27425;
assign w30078 = pi1846 & ~w29226;
assign w30079 = ~w29227 & ~w30078;
assign w30080 = ~w27425 & w30079;
assign w30081 = ~w30077 & ~w30080;
assign w30082 = ~pi0953 & w27425;
assign w30083 = pi1847 & ~w27429;
assign w30084 = ~w29226 & ~w30083;
assign w30085 = ~w27425 & w30084;
assign w30086 = ~w30082 & ~w30085;
assign w30087 = ~pi0967 & w28384;
assign w30088 = pi1848 & ~w28387;
assign w30089 = ~w29304 & ~w30088;
assign w30090 = ~w28384 & w30089;
assign w30091 = ~w30087 & ~w30090;
assign w30092 = ~pi0966 & w28384;
assign w30093 = pi1849 & ~w29304;
assign w30094 = ~w29305 & ~w30093;
assign w30095 = ~w28384 & w30094;
assign w30096 = ~w30092 & ~w30095;
assign w30097 = pi1646 & pi1850;
assign w30098 = ~w28412 & ~w30097;
assign w30099 = ~w28452 & w30098;
assign w30100 = pi1851 & ~w27274;
assign w30101 = ~w27275 & ~w30100;
assign w30102 = pi1852 & ~w29537;
assign w30103 = w5320 & w29537;
assign w30104 = ~w30102 & ~w30103;
assign w30105 = pi1853 & ~w29537;
assign w30106 = w4749 & w29537;
assign w30107 = ~w30105 & ~w30106;
assign w30108 = pi1854 & ~w29742;
assign w30109 = w8081 & w29742;
assign w30110 = ~w30108 & ~w30109;
assign w30111 = ~pi1924 & w29772;
assign w30112 = ~pi1855 & ~w29774;
assign w30113 = ~w29772 & ~w29775;
assign w30114 = ~w30112 & w30113;
assign w30115 = ~w30111 & ~w30114;
assign w30116 = ~pi1422 & ~pi3572;
assign w30117 = ~pi3645 & w30116;
assign w30118 = ~pi1856 & w30117;
assign w30119 = pi1856 & ~w30117;
assign w30120 = ~w30118 & ~w30119;
assign w30121 = w26505 & w30120;
assign w30122 = pi1857 & ~w29742;
assign w30123 = w3195 & w29742;
assign w30124 = ~w30122 & ~w30123;
assign w30125 = pi1858 & ~w29742;
assign w30126 = w5320 & w29742;
assign w30127 = ~w30125 & ~w30126;
assign w30128 = pi1859 & ~w23322;
assign w30129 = ~pi0593 & w23322;
assign w30130 = ~w30128 & ~w30129;
assign w30131 = ~pi3419 & pi3562;
assign w30132 = ~w897 & ~w2896;
assign w30133 = pi3590 & ~w30132;
assign w30134 = w156 & ~w22042;
assign w30135 = ~pi1860 & ~w30134;
assign w30136 = ~w30133 & w30135;
assign w30137 = pi1861 & ~w30037;
assign w30138 = w895 & ~w7232;
assign w30139 = w22040 & w30138;
assign w30140 = ~w30137 & ~w30139;
assign w30141 = w1286 & w24322;
assign w30142 = pi1862 & ~w30141;
assign w30143 = w4749 & w30141;
assign w30144 = ~w30142 & ~w30143;
assign w30145 = pi1863 & ~w29987;
assign w30146 = ~pi0036 & w29987;
assign w30147 = ~w30145 & ~w30146;
assign w30148 = pi1864 & ~w23322;
assign w30149 = ~pi0578 & w23322;
assign w30150 = ~w30148 & ~w30149;
assign w30151 = pi1865 & ~w29555;
assign w30152 = ~pi0578 & w29555;
assign w30153 = ~w30151 & ~w30152;
assign w30154 = ~w8081 & ~w15388;
assign w30155 = ~pi1866 & w15388;
assign w30156 = ~pi2555 & ~w30155;
assign w30157 = ~w30154 & w30156;
assign w30158 = ~w29583 & ~w30157;
assign w30159 = ~w3195 & ~w15388;
assign w30160 = ~pi1867 & w15388;
assign w30161 = ~pi2555 & ~w30160;
assign w30162 = ~w30159 & w30161;
assign w30163 = ~w29583 & ~w30162;
assign w30164 = pi1868 & pi1896;
assign w30165 = ~w25723 & ~w30164;
assign w30166 = w25801 & w30165;
assign w30167 = pi1869 & ~w30141;
assign w30168 = w8081 & w30141;
assign w30169 = ~w30167 & ~w30168;
assign w30170 = pi1870 & ~w25726;
assign w30171 = ~w25727 & ~w30170;
assign w30172 = w25801 & w30171;
assign w30173 = pi1871 & ~w25724;
assign w30174 = ~w25725 & ~w30173;
assign w30175 = w25801 & w30174;
assign w30176 = pi1872 & ~w25730;
assign w30177 = ~w25731 & w25801;
assign w30178 = ~w30176 & w30177;
assign w30179 = pi1873 & ~w30141;
assign w30180 = w3711 & w30141;
assign w30181 = ~w30179 & ~w30180;
assign w30182 = pi1874 & ~w30141;
assign w30183 = w1308 & w30141;
assign w30184 = ~w30182 & ~w30183;
assign w30185 = ~pi3681 & w23031;
assign w30186 = pi3444 & ~w18313;
assign w30187 = ~w30185 & w30186;
assign w30188 = w18357 & w30187;
assign w30189 = pi1876 & w25889;
assign w30190 = pi1877 & ~w29542;
assign w30191 = w4141 & w29542;
assign w30192 = ~w30190 & ~w30191;
assign w30193 = pi1878 & ~w29542;
assign w30194 = w6177 & w29542;
assign w30195 = ~w30193 & ~w30194;
assign w30196 = pi1879 & ~w29542;
assign w30197 = w1639 & w29542;
assign w30198 = ~w30196 & ~w30197;
assign w30199 = pi1880 & ~w29542;
assign w30200 = w1308 & w29542;
assign w30201 = ~w30199 & ~w30200;
assign w30202 = w24322 & w29785;
assign w30203 = ~w5635 & w30202;
assign w30204 = pi1881 & ~w30202;
assign w30205 = ~w30203 & ~w30204;
assign w30206 = w10741 & ~w30185;
assign w30207 = pi1882 & ~pi2814;
assign w30208 = pi1883 & ~w30141;
assign w30209 = w6177 & w30141;
assign w30210 = ~w30208 & ~w30209;
assign w30211 = pi1884 & ~w30141;
assign w30212 = w3195 & w30141;
assign w30213 = ~w30211 & ~w30212;
assign w30214 = pi1885 & ~w30141;
assign w30215 = w40134 & w30141;
assign w30216 = ~w30214 & ~w30215;
assign w30217 = pi1886 & ~w30141;
assign w30218 = w4380 & w30141;
assign w30219 = ~w30217 & ~w30218;
assign w30220 = pi1887 & ~w30141;
assign w30221 = w5320 & w30141;
assign w30222 = ~w30220 & ~w30221;
assign w30223 = pi1888 & ~w30141;
assign w30224 = w5914 & w30141;
assign w30225 = ~w30223 & ~w30224;
assign w30226 = pi1889 & ~w30141;
assign w30227 = w8240 & w30141;
assign w30228 = ~w30226 & ~w30227;
assign w30229 = pi1890 & ~w30141;
assign w30230 = w1639 & w30141;
assign w30231 = ~w30229 & ~w30230;
assign w30232 = pi1891 & ~w30141;
assign w30233 = w5053 & w30141;
assign w30234 = ~w30232 & ~w30233;
assign w30235 = pi1892 & ~w30141;
assign w30236 = w5635 & w30141;
assign w30237 = ~w30235 & ~w30236;
assign w30238 = pi1893 & ~w25727;
assign w30239 = ~w25728 & ~w30238;
assign w30240 = w25801 & w30239;
assign w30241 = pi1894 & ~w25725;
assign w30242 = ~w25726 & ~w30241;
assign w30243 = w25801 & w30242;
assign w30244 = pi1895 & ~w25723;
assign w30245 = ~w25724 & ~w30244;
assign w30246 = w25801 & w30245;
assign w30247 = pi1896 & w25801;
assign w30248 = ~w8240 & ~w15388;
assign w30249 = ~pi1897 & w15388;
assign w30250 = ~pi2555 & ~w30249;
assign w30251 = ~w30248 & w30250;
assign w30252 = ~w29583 & ~w30251;
assign w30253 = w24322 & w24674;
assign w30254 = pi1898 & ~w30253;
assign w30255 = w6177 & w30253;
assign w30256 = ~w30254 & ~w30255;
assign w30257 = pi1899 & ~w30253;
assign w30258 = w40134 & w30253;
assign w30259 = ~w30257 & ~w30258;
assign w30260 = pi1900 & ~w30253;
assign w30261 = w4380 & w30253;
assign w30262 = ~w30260 & ~w30261;
assign w30263 = pi1901 & ~w30253;
assign w30264 = w5320 & w30253;
assign w30265 = ~w30263 & ~w30264;
assign w30266 = pi1902 & ~w30253;
assign w30267 = w5914 & w30253;
assign w30268 = ~w30266 & ~w30267;
assign w30269 = pi1903 & ~w30253;
assign w30270 = w8240 & w30253;
assign w30271 = ~w30269 & ~w30270;
assign w30272 = pi1904 & ~w30253;
assign w30273 = w8081 & w30253;
assign w30274 = ~w30272 & ~w30273;
assign w30275 = pi1905 & ~w30253;
assign w30276 = w1639 & w30253;
assign w30277 = ~w30275 & ~w30276;
assign w30278 = pi1906 & ~w30253;
assign w30279 = w5635 & w30253;
assign w30280 = ~w30278 & ~w30279;
assign w30281 = pi1907 & ~w30253;
assign w30282 = w3711 & w30253;
assign w30283 = ~w30281 & ~w30282;
assign w30284 = w1244 & w24374;
assign w30285 = pi1908 & ~w30284;
assign w30286 = w8240 & w30284;
assign w30287 = ~w30285 & ~w30286;
assign w30288 = pi1909 & ~w30284;
assign w30289 = w1308 & w30284;
assign w30290 = ~w30288 & ~w30289;
assign w30291 = pi1910 & ~w25815;
assign w30292 = ~w25816 & ~w30291;
assign w30293 = w25889 & w30292;
assign w30294 = pi1911 & ~w25813;
assign w30295 = ~w25814 & ~w30294;
assign w30296 = w25889 & w30295;
assign w30297 = pi1876 & pi1912;
assign w30298 = ~w25811 & ~w30297;
assign w30299 = w25889 & w30298;
assign w30300 = pi1913 & ~w25811;
assign w30301 = ~w25812 & ~w30300;
assign w30302 = w25889 & w30301;
assign w30303 = pi1914 & ~w25812;
assign w30304 = ~w25813 & ~w30303;
assign w30305 = w25889 & w30304;
assign w30306 = pi1915 & ~w25818;
assign w30307 = ~w25819 & w25889;
assign w30308 = ~w30306 & w30307;
assign w30309 = pi1916 & ~w25814;
assign w30310 = ~w25815 & ~w30309;
assign w30311 = w25889 & w30310;
assign w30312 = pi1917 & ~w30284;
assign w30313 = w8081 & w30284;
assign w30314 = ~w30312 & ~w30313;
assign w30315 = w24681 & w28606;
assign w30316 = pi1918 & ~w30315;
assign w30317 = w4141 & w30315;
assign w30318 = ~w30316 & ~w30317;
assign w30319 = pi1919 & ~w30315;
assign w30320 = w6177 & w30315;
assign w30321 = ~w30319 & ~w30320;
assign w30322 = pi1920 & ~w30141;
assign w30323 = w6413 & w30141;
assign w30324 = ~w30322 & ~w30323;
assign w30325 = pi1921 & ~w30315;
assign w30326 = w3195 & w30315;
assign w30327 = ~w30325 & ~w30326;
assign w30328 = pi1922 & ~w30315;
assign w30329 = w40134 & w30315;
assign w30330 = ~w30328 & ~w30329;
assign w30331 = pi1923 & ~w30315;
assign w30332 = w6413 & w30315;
assign w30333 = ~w30331 & ~w30332;
assign w30334 = pi1924 & ~w30315;
assign w30335 = w4380 & w30315;
assign w30336 = ~w30334 & ~w30335;
assign w30337 = pi1925 & ~w30315;
assign w30338 = w5320 & w30315;
assign w30339 = ~w30337 & ~w30338;
assign w30340 = pi1926 & ~w30315;
assign w30341 = w5914 & w30315;
assign w30342 = ~w30340 & ~w30341;
assign w30343 = pi1927 & ~w30315;
assign w30344 = w4749 & w30315;
assign w30345 = ~w30343 & ~w30344;
assign w30346 = pi1928 & ~w30315;
assign w30347 = w8240 & w30315;
assign w30348 = ~w30346 & ~w30347;
assign w30349 = pi1929 & ~w30315;
assign w30350 = w8081 & w30315;
assign w30351 = ~w30349 & ~w30350;
assign w30352 = pi1930 & ~w30315;
assign w30353 = w1639 & w30315;
assign w30354 = ~w30352 & ~w30353;
assign w30355 = pi1931 & ~w30315;
assign w30356 = w5635 & w30315;
assign w30357 = ~w30355 & ~w30356;
assign w30358 = pi1932 & ~w30315;
assign w30359 = w5053 & w30315;
assign w30360 = ~w30358 & ~w30359;
assign w30361 = pi1933 & ~w30315;
assign w30362 = w3711 & w30315;
assign w30363 = ~w30361 & ~w30362;
assign w30364 = w343 & w928;
assign w30365 = ~w6612 & ~w30364;
assign w30366 = w6598 & w30365;
assign w30367 = w4797 & w30366;
assign w30368 = pi1934 & w30364;
assign w30369 = ~w30367 & ~w30368;
assign w30370 = pi1936 & ~pi3147;
assign w30371 = ~w29781 & ~w30370;
assign w30372 = ~w20671 & ~w30371;
assign w30373 = ~w29781 & w30370;
assign w30374 = ~pi2056 & w30373;
assign w30375 = w30372 & ~w30374;
assign w30376 = ~pi1935 & ~w30375;
assign w30377 = w24804 & w30373;
assign w30378 = pi1918 & w29781;
assign w30379 = ~w30377 & ~w30378;
assign w30380 = ~w20671 & ~w30379;
assign w30381 = ~w30376 & ~w30380;
assign w30382 = pi3147 & ~w29781;
assign w30383 = ~w20671 & ~w30382;
assign w30384 = ~pi1936 & ~w30383;
assign w30385 = ~pi1921 & w29781;
assign w30386 = w30372 & ~w30385;
assign w30387 = ~w30384 & ~w30386;
assign w30388 = ~pi1922 & w29772;
assign w30389 = ~pi1937 & ~w29776;
assign w30390 = w19035 & w29774;
assign w30391 = ~w29772 & ~w30390;
assign w30392 = ~w30389 & w30391;
assign w30393 = ~w30388 & ~w30392;
assign w30394 = w24374 & w29625;
assign w30395 = pi1938 & ~w30394;
assign w30396 = w3195 & w30394;
assign w30397 = ~w30395 & ~w30396;
assign w30398 = pi1939 & ~w30394;
assign w30399 = w40134 & w30394;
assign w30400 = ~w30398 & ~w30399;
assign w30401 = pi1940 & ~w30394;
assign w30402 = w6413 & w30394;
assign w30403 = ~w30401 & ~w30402;
assign w30404 = pi1941 & ~w30394;
assign w30405 = w4380 & w30394;
assign w30406 = ~w30404 & ~w30405;
assign w30407 = pi1942 & ~w30394;
assign w30408 = w5320 & w30394;
assign w30409 = ~w30407 & ~w30408;
assign w30410 = pi1943 & ~w30394;
assign w30411 = w5914 & w30394;
assign w30412 = ~w30410 & ~w30411;
assign w30413 = pi1944 & ~w30394;
assign w30414 = w4749 & w30394;
assign w30415 = ~w30413 & ~w30414;
assign w30416 = pi1945 & ~w30394;
assign w30417 = w3711 & w30394;
assign w30418 = ~w30416 & ~w30417;
assign w30419 = pi3256 & ~w28745;
assign w30420 = w116 & w30419;
assign w30421 = w85 & w30420;
assign w30422 = pi1946 & ~w30421;
assign w30423 = pi3698 & w30421;
assign w30424 = ~w30422 & ~w30423;
assign w30425 = pi1947 & ~w30421;
assign w30426 = pi3697 & w30421;
assign w30427 = ~w30425 & ~w30426;
assign w30428 = pi1948 & ~w30421;
assign w30429 = pi3696 & w30421;
assign w30430 = ~w30428 & ~w30429;
assign w30431 = pi1949 & ~w30421;
assign w30432 = pi3695 & w30421;
assign w30433 = ~w30431 & ~w30432;
assign w30434 = pi1950 & ~w30421;
assign w30435 = pi3694 & w30421;
assign w30436 = ~w30434 & ~w30435;
assign w30437 = pi1951 & ~w30421;
assign w30438 = pi3693 & w30421;
assign w30439 = ~w30437 & ~w30438;
assign w30440 = pi1952 & ~w30141;
assign w30441 = w4141 & w30141;
assign w30442 = ~w30440 & ~w30441;
assign w30443 = ~pi1953 & w6684;
assign w30444 = w7160 & ~w14373;
assign w30445 = w6682 & w30444;
assign w30446 = w29429 & w30445;
assign w30447 = ~w30443 & ~w30446;
assign w30448 = pi1954 & ~w29987;
assign w30449 = ~pi0007 & w29987;
assign w30450 = ~w30448 & ~w30449;
assign w30451 = w4141 & w14856;
assign w30452 = ~w16540 & ~w30451;
assign w30453 = ~w17425 & w30452;
assign w30454 = w6115 & w17425;
assign w30455 = ~w30453 & ~w30454;
assign w30456 = w17421 & ~w30455;
assign w30457 = ~pi1955 & ~w17421;
assign w30458 = ~w30456 & ~w30457;
assign w30459 = w6177 & w14856;
assign w30460 = ~w16243 & ~w30459;
assign w30461 = ~w17425 & w30460;
assign w30462 = w3088 & w17425;
assign w30463 = ~w30461 & ~w30462;
assign w30464 = w17421 & ~w30463;
assign w30465 = ~pi1956 & ~w17421;
assign w30466 = ~w30464 & ~w30465;
assign w30467 = w3195 & w14856;
assign w30468 = ~w16331 & ~w30467;
assign w30469 = ~w17425 & w30468;
assign w30470 = w3362 & w17425;
assign w30471 = ~w30469 & ~w30470;
assign w30472 = w17421 & ~w30471;
assign w30473 = ~pi1957 & ~w17421;
assign w30474 = ~w30472 & ~w30473;
assign w30475 = w40134 & w14856;
assign w30476 = ~w15549 & ~w30475;
assign w30477 = ~w17425 & w30476;
assign w30478 = w6275 & w17425;
assign w30479 = ~w30477 & ~w30478;
assign w30480 = w17421 & ~w30479;
assign w30481 = ~pi1958 & ~w17421;
assign w30482 = ~w30480 & ~w30481;
assign w30483 = w6413 & w14856;
assign w30484 = ~w15649 & ~w30483;
assign w30485 = ~w17425 & w30484;
assign w30486 = w4298 & w17425;
assign w30487 = ~w30485 & ~w30486;
assign w30488 = w17421 & ~w30487;
assign w30489 = ~pi1959 & ~w17421;
assign w30490 = ~w30488 & ~w30489;
assign w30491 = w4380 & w14856;
assign w30492 = ~w15754 & ~w30491;
assign w30493 = ~w17425 & w30492;
assign w30494 = w5183 & w17425;
assign w30495 = ~w30493 & ~w30494;
assign w30496 = w17421 & ~w30495;
assign w30497 = ~pi1960 & ~w17421;
assign w30498 = ~w30496 & ~w30497;
assign w30499 = w5320 & w14856;
assign w30500 = ~w16434 & ~w30499;
assign w30501 = ~w17425 & w30500;
assign w30502 = w5778 & w17425;
assign w30503 = ~w30501 & ~w30502;
assign w30504 = w17421 & ~w30503;
assign w30505 = ~pi1961 & ~w17421;
assign w30506 = ~w30504 & ~w30505;
assign w30507 = w5914 & w14856;
assign w30508 = ~w14857 & ~w30507;
assign w30509 = ~w17425 & w30508;
assign w30510 = w4716 & w17425;
assign w30511 = ~w30509 & ~w30510;
assign w30512 = w17421 & ~w30511;
assign w30513 = ~pi1962 & ~w17421;
assign w30514 = ~w30512 & ~w30513;
assign w30515 = w8240 & w14856;
assign w30516 = ~w15899 & ~w30515;
assign w30517 = ~w17425 & w30516;
assign w30518 = w7965 & w17425;
assign w30519 = ~w30517 & ~w30518;
assign w30520 = w17421 & ~w30519;
assign w30521 = ~pi1963 & ~w17421;
assign w30522 = ~w30520 & ~w30521;
assign w30523 = w1639 & w14856;
assign w30524 = ~w16669 & ~w30523;
assign w30525 = ~w17425 & w30524;
assign w30526 = w1132 & w17425;
assign w30527 = ~w30525 & ~w30526;
assign w30528 = w17421 & ~w30527;
assign w30529 = ~pi1964 & ~w17421;
assign w30530 = ~w30528 & ~w30529;
assign w30531 = w1308 & w14856;
assign w30532 = ~w16860 & ~w30531;
assign w30533 = ~w17425 & w30532;
assign w30534 = w5557 & w17425;
assign w30535 = ~w30533 & ~w30534;
assign w30536 = w17421 & ~w30535;
assign w30537 = ~pi1965 & ~w17421;
assign w30538 = ~w30536 & ~w30537;
assign w30539 = w5635 & w14856;
assign w30540 = ~w16882 & ~w30539;
assign w30541 = ~w17425 & w30540;
assign w30542 = w4949 & w17425;
assign w30543 = ~w30541 & ~w30542;
assign w30544 = w17421 & ~w30543;
assign w30545 = ~pi1966 & ~w17421;
assign w30546 = ~w30544 & ~w30545;
assign w30547 = w5053 & w14856;
assign w30548 = ~w17050 & ~w30547;
assign w30549 = ~w17425 & w30548;
assign w30550 = w4068 & w17425;
assign w30551 = ~w30549 & ~w30550;
assign w30552 = w17421 & ~w30551;
assign w30553 = ~pi1967 & ~w17421;
assign w30554 = ~w30552 & ~w30553;
assign w30555 = pi1968 & ~w29987;
assign w30556 = ~pi0034 & w29987;
assign w30557 = ~w30555 & ~w30556;
assign w30558 = pi1969 & ~w29987;
assign w30559 = ~pi0005 & w29987;
assign w30560 = ~w30558 & ~w30559;
assign w30561 = pi1970 & ~w29987;
assign w30562 = ~pi0003 & w29987;
assign w30563 = ~w30561 & ~w30562;
assign w30564 = w381 & w6971;
assign w30565 = ~w343 & w30564;
assign w30566 = w380 & w7099;
assign w30567 = w23334 & w30566;
assign w30568 = ~w30565 & ~w30567;
assign w30569 = ~pi1971 & w30568;
assign w30570 = ~w30444 & ~w30569;
assign w30571 = ~w30444 & w30568;
assign w30572 = ~pi1972 & w30571;
assign w30573 = pi0405 & ~w30571;
assign w30574 = ~w30572 & ~w30573;
assign w30575 = ~pi1973 & w30571;
assign w30576 = pi0422 & ~w30571;
assign w30577 = ~w30575 & ~w30576;
assign w30578 = ~pi1974 & w30571;
assign w30579 = pi0423 & ~w30571;
assign w30580 = ~w30578 & ~w30579;
assign w30581 = ~pi1975 & w30571;
assign w30582 = pi0424 & ~w30571;
assign w30583 = ~w30581 & ~w30582;
assign w30584 = w849 & ~w23420;
assign w30585 = ~pi1976 & ~w849;
assign w30586 = ~w30584 & ~w30585;
assign w30587 = pi1977 & ~w849;
assign w30588 = w849 & ~w8802;
assign w30589 = ~w30587 & ~w30588;
assign w30590 = w849 & ~w23437;
assign w30591 = ~pi1978 & ~w849;
assign w30592 = ~w30590 & ~w30591;
assign w30593 = w849 & w8745;
assign w30594 = ~w23457 & ~w30593;
assign w30595 = w849 & w8699;
assign w30596 = ~w8704 & ~w30595;
assign w30597 = pi1981 & ~w849;
assign w30598 = w849 & ~w8667;
assign w30599 = ~w30597 & ~w30598;
assign w30600 = pi1982 & ~w849;
assign w30601 = w849 & ~w23496;
assign w30602 = ~w30600 & ~w30601;
assign w30603 = w849 & ~w22214;
assign w30604 = ~pi1983 & ~w849;
assign w30605 = ~w30603 & ~w30604;
assign w30606 = w849 & ~w22222;
assign w30607 = ~w23239 & ~w30606;
assign w30608 = w849 & ~w8560;
assign w30609 = ~pi1985 & ~w849;
assign w30610 = ~w30608 & ~w30609;
assign w30611 = pi1986 & ~w29897;
assign w30612 = pi3398 & w29897;
assign w30613 = ~w30611 & ~w30612;
assign w30614 = pi1987 & ~w29897;
assign w30615 = pi3520 & w29897;
assign w30616 = ~w30614 & ~w30615;
assign w30617 = pi1988 & ~w29897;
assign w30618 = pi3392 & w29897;
assign w30619 = ~w30617 & ~w30618;
assign w30620 = ~pi3394 & w29897;
assign w30621 = pi1989 & ~w29897;
assign w30622 = ~w30620 & ~w30621;
assign w30623 = ~pi2514 & w29897;
assign w30624 = pi1990 & ~w29897;
assign w30625 = ~w30623 & ~w30624;
assign w30626 = pi1991 & ~w29897;
assign w30627 = pi3512 & w29897;
assign w30628 = ~w30626 & ~w30627;
assign w30629 = pi1992 & ~w29897;
assign w30630 = pi3513 & w29897;
assign w30631 = ~w30629 & ~w30630;
assign w30632 = pi1993 & ~w29897;
assign w30633 = pi3514 & w29897;
assign w30634 = ~w30632 & ~w30633;
assign w30635 = pi1994 & ~w29897;
assign w30636 = pi3518 & w29897;
assign w30637 = ~w30635 & ~w30636;
assign w30638 = pi1995 & ~w29897;
assign w30639 = pi3516 & w29897;
assign w30640 = ~w30638 & ~w30639;
assign w30641 = ~pi3330 & w29579;
assign w30642 = pi1996 & ~w29579;
assign w30643 = ~w30641 & ~w30642;
assign w30644 = ~pi3394 & w29579;
assign w30645 = pi1997 & ~w29579;
assign w30646 = ~w30644 & ~w30645;
assign w30647 = pi1998 & ~w29901;
assign w30648 = pi3511 & w29901;
assign w30649 = ~w30647 & ~w30648;
assign w30650 = pi1999 & ~w29901;
assign w30651 = pi3392 & w29901;
assign w30652 = ~w30650 & ~w30651;
assign w30653 = ~pi3394 & w29901;
assign w30654 = pi2000 & ~w29901;
assign w30655 = ~w30653 & ~w30654;
assign w30656 = ~pi2514 & w29901;
assign w30657 = pi2001 & ~w29901;
assign w30658 = ~w30656 & ~w30657;
assign w30659 = pi2002 & ~w29901;
assign w30660 = pi3512 & w29901;
assign w30661 = ~w30659 & ~w30660;
assign w30662 = pi2003 & ~w29901;
assign w30663 = pi3514 & w29901;
assign w30664 = ~w30662 & ~w30663;
assign w30665 = pi2004 & ~w29901;
assign w30666 = pi3516 & w29901;
assign w30667 = ~w30665 & ~w30666;
assign w30668 = pi2005 & ~w29901;
assign w30669 = pi3517 & w29901;
assign w30670 = ~w30668 & ~w30669;
assign w30671 = pi2006 & ~w29901;
assign w30672 = pi3509 & w29901;
assign w30673 = ~w30671 & ~w30672;
assign w30674 = pi2007 & ~w29901;
assign w30675 = pi3521 & w29901;
assign w30676 = ~w30674 & ~w30675;
assign w30677 = pi1797 & pi1798;
assign w30678 = w29891 & w30677;
assign w30679 = ~pi3330 & w30678;
assign w30680 = pi2008 & ~w30678;
assign w30681 = ~w30679 & ~w30680;
assign w30682 = ~pi3394 & w30678;
assign w30683 = pi2009 & ~w30678;
assign w30684 = ~w30682 & ~w30683;
assign w30685 = ~pi2010 & w342;
assign w30686 = w422 & w24445;
assign w30687 = w4423 & ~w30686;
assign w30688 = w382 & ~w30687;
assign w30689 = pi0425 & w29980;
assign w30690 = ~w342 & ~w30689;
assign w30691 = ~w30688 & w30690;
assign w30692 = ~w30685 & ~w30691;
assign w30693 = ~pi2011 & w342;
assign w30694 = w422 & w23437;
assign w30695 = w6446 & ~w30694;
assign w30696 = w382 & ~w30695;
assign w30697 = pi0409 & w29980;
assign w30698 = ~w342 & ~w30697;
assign w30699 = ~w30696 & w30698;
assign w30700 = ~w30693 & ~w30699;
assign w30701 = ~pi2012 & w342;
assign w30702 = w422 & w8745;
assign w30703 = w8752 & ~w30702;
assign w30704 = w382 & ~w30703;
assign w30705 = pi0410 & w29980;
assign w30706 = ~w342 & ~w30705;
assign w30707 = ~w30704 & w30706;
assign w30708 = ~w30701 & ~w30707;
assign w30709 = ~pi2013 & w342;
assign w30710 = pi0411 & w29980;
assign w30711 = ~w342 & ~w30710;
assign w30712 = ~w30709 & ~w30711;
assign w30713 = w422 & w8699;
assign w30714 = w8707 & ~w30713;
assign w30715 = w382 & ~w30709;
assign w30716 = ~w30714 & w30715;
assign w30717 = ~w30712 & ~w30716;
assign w30718 = ~pi2014 & w342;
assign w30719 = w422 & ~w8667;
assign w30720 = w8674 & ~w30719;
assign w30721 = w382 & ~w30720;
assign w30722 = pi0412 & w29980;
assign w30723 = ~w342 & ~w30722;
assign w30724 = ~w30721 & w30723;
assign w30725 = ~w30718 & ~w30724;
assign w30726 = ~pi2015 & w342;
assign w30727 = w422 & ~w23496;
assign w30728 = w8609 & ~w30727;
assign w30729 = w382 & ~w30728;
assign w30730 = pi0413 & w29980;
assign w30731 = ~w342 & ~w30730;
assign w30732 = ~w30729 & w30731;
assign w30733 = ~w30726 & ~w30732;
assign w30734 = ~pi2016 & w342;
assign w30735 = pi0408 & w29980;
assign w30736 = ~w342 & ~w30735;
assign w30737 = ~w30734 & ~w30736;
assign w30738 = w422 & w8560;
assign w30739 = w8567 & ~w30738;
assign w30740 = w382 & ~w30734;
assign w30741 = ~w30739 & w30740;
assign w30742 = ~w30737 & ~w30741;
assign w30743 = pi2017 & ~w23792;
assign w30744 = w23800 & w23801;
assign w30745 = w27127 & w30744;
assign w30746 = ~w30743 & ~w30745;
assign w30747 = pi2018 & ~w23792;
assign w30748 = w23796 & w23804;
assign w30749 = w27127 & w30748;
assign w30750 = ~w30747 & ~w30749;
assign w30751 = pi2019 & ~w23792;
assign w30752 = w23795 & w23805;
assign w30753 = w27127 & w30752;
assign w30754 = ~w30751 & ~w30753;
assign w30755 = ~pi2020 & w6684;
assign w30756 = ~w29429 & w30445;
assign w30757 = ~w30755 & ~w30756;
assign w30758 = pi0405 & w376;
assign w30759 = w379 & w30758;
assign w30760 = ~w2234 & ~w30759;
assign w30761 = w21968 & ~w30760;
assign w30762 = ~pi2021 & w6684;
assign w30763 = ~w30761 & ~w30762;
assign w30764 = pi2022 & ~w29987;
assign w30765 = ~pi0002 & w29987;
assign w30766 = ~w30764 & ~w30765;
assign w30767 = pi2023 & ~w29987;
assign w30768 = ~pi0011 & w29987;
assign w30769 = ~w30767 & ~w30768;
assign w30770 = pi2024 & ~w29987;
assign w30771 = ~pi0010 & w29987;
assign w30772 = ~w30770 & ~w30771;
assign w30773 = pi2025 & ~w29987;
assign w30774 = ~pi0009 & w29987;
assign w30775 = ~w30773 & ~w30774;
assign w30776 = pi2026 & ~w29987;
assign w30777 = ~pi0008 & w29987;
assign w30778 = ~w30776 & ~w30777;
assign w30779 = pi2027 & ~w29987;
assign w30780 = ~pi0006 & w29987;
assign w30781 = ~w30779 & ~w30780;
assign w30782 = pi2028 & ~w29987;
assign w30783 = ~pi0004 & w29987;
assign w30784 = ~w30782 & ~w30783;
assign w30785 = pi2029 & ~w29987;
assign w30786 = pi3353 & ~w6749;
assign w30787 = ~w6750 & ~w30786;
assign w30788 = w29987 & w30787;
assign w30789 = ~w30785 & ~w30788;
assign w30790 = pi2030 & ~w29987;
assign w30791 = pi3355 & ~w6749;
assign w30792 = ~w6751 & ~w30791;
assign w30793 = w29987 & w30792;
assign w30794 = ~w30790 & ~w30793;
assign w30795 = pi2031 & ~w29987;
assign w30796 = ~pi0028 & w29987;
assign w30797 = ~w30795 & ~w30796;
assign w30798 = pi2032 & ~w29987;
assign w30799 = ~pi0037 & w29987;
assign w30800 = ~w30798 & ~w30799;
assign w30801 = pi2033 & ~w29987;
assign w30802 = ~pi0035 & w29987;
assign w30803 = ~w30801 & ~w30802;
assign w30804 = pi2034 & ~w29987;
assign w30805 = ~pi0033 & w29987;
assign w30806 = ~w30804 & ~w30805;
assign w30807 = pi2035 & ~w29987;
assign w30808 = ~pi0031 & w29987;
assign w30809 = ~w30807 & ~w30808;
assign w30810 = pi2036 & ~w29987;
assign w30811 = ~pi0029 & w29987;
assign w30812 = ~w30810 & ~w30811;
assign w30813 = pi2037 & ~w29987;
assign w30814 = ~pi0022 & w29987;
assign w30815 = ~w30813 & ~w30814;
assign w30816 = pi2038 & ~w29987;
assign w30817 = ~pi0021 & w29987;
assign w30818 = ~w30816 & ~w30817;
assign w30819 = pi2039 & ~w29987;
assign w30820 = ~pi0020 & w29987;
assign w30821 = ~w30819 & ~w30820;
assign w30822 = pi2040 & ~w29987;
assign w30823 = ~pi0018 & w29987;
assign w30824 = ~w30822 & ~w30823;
assign w30825 = pi2041 & ~w29987;
assign w30826 = ~pi0017 & w29987;
assign w30827 = ~w30825 & ~w30826;
assign w30828 = pi2042 & ~w29987;
assign w30829 = ~pi0016 & w29987;
assign w30830 = ~w30828 & ~w30829;
assign w30831 = pi2043 & ~w29987;
assign w30832 = ~pi0027 & w29987;
assign w30833 = ~w30831 & ~w30832;
assign w30834 = pi2044 & ~w29987;
assign w30835 = ~pi0026 & w29987;
assign w30836 = ~w30834 & ~w30835;
assign w30837 = pi2045 & ~w29987;
assign w30838 = ~pi0025 & w29987;
assign w30839 = ~w30837 & ~w30838;
assign w30840 = pi2046 & ~w29987;
assign w30841 = ~w7047 & ~w30791;
assign w30842 = w29987 & w30841;
assign w30843 = ~w30840 & ~w30842;
assign w30844 = pi2047 & ~w29987;
assign w30845 = ~w7048 & ~w30786;
assign w30846 = w29987 & w30845;
assign w30847 = ~w30844 & ~w30846;
assign w30848 = w2890 & w22040;
assign w30849 = ~pi2048 & w30848;
assign w30850 = pi2048 & ~w30848;
assign w30851 = ~w30849 & ~w30850;
assign w30852 = w165 & w177;
assign w30853 = w114 & w30852;
assign w30854 = ~pi1860 & w13;
assign w30855 = w97 & w30854;
assign w30856 = w133 & w30855;
assign w30857 = pi3199 & w30856;
assign w30858 = pi2759 & w30857;
assign w30859 = pi2049 & w30858;
assign w30860 = ~pi2049 & ~w30858;
assign w30861 = ~w30859 & ~w30860;
assign w30862 = ~w30853 & w30861;
assign w30863 = pi2050 & ~w29987;
assign w30864 = ~pi0014 & w29987;
assign w30865 = ~w30863 & ~w30864;
assign w30866 = pi2051 & ~w30253;
assign w30867 = w5053 & w30253;
assign w30868 = ~w30866 & ~w30867;
assign w30869 = pi2052 & ~w30253;
assign w30870 = w4749 & w30253;
assign w30871 = ~w30869 & ~w30870;
assign w30872 = pi2053 & ~w30253;
assign w30873 = w1308 & w30253;
assign w30874 = ~w30872 & ~w30873;
assign w30875 = pi2054 & ~w30253;
assign w30876 = w6413 & w30253;
assign w30877 = ~w30875 & ~w30876;
assign w30878 = pi2055 & ~w30253;
assign w30879 = w3195 & w30253;
assign w30880 = ~w30878 & ~w30879;
assign w30881 = ~pi1919 & w29781;
assign w30882 = ~w30374 & ~w30881;
assign w30883 = ~w20671 & ~w30882;
assign w30884 = pi2056 & ~w30372;
assign w30885 = ~w30883 & ~w30884;
assign w30886 = pi2057 & ~w30253;
assign w30887 = w4141 & w30253;
assign w30888 = ~w30886 & ~w30887;
assign w30889 = w5914 & w23862;
assign w30890 = ~pi2058 & ~w23866;
assign w30891 = ~w23867 & ~w30890;
assign w30892 = ~w23862 & w30891;
assign w30893 = ~w30889 & ~w30892;
assign w30894 = w3711 & w23862;
assign w30895 = ~pi2059 & ~w30041;
assign w30896 = pi2059 & w30041;
assign w30897 = ~w30895 & ~w30896;
assign w30898 = ~w23862 & w30897;
assign w30899 = ~w30894 & ~w30898;
assign w30900 = pi2060 & ~w29987;
assign w30901 = ~pi0024 & w29987;
assign w30902 = ~w30900 & ~w30901;
assign w30903 = w4749 & w23862;
assign w30904 = ~pi2061 & ~w23865;
assign w30905 = ~w23866 & ~w30904;
assign w30906 = ~w23862 & w30905;
assign w30907 = ~w30903 & ~w30906;
assign w30908 = pi2062 & ~w29987;
assign w30909 = ~pi0015 & w29987;
assign w30910 = ~w30908 & ~w30909;
assign w30911 = pi2063 & ~w29987;
assign w30912 = ~pi0030 & w29987;
assign w30913 = ~w30911 & ~w30912;
assign w30914 = pi2064 & ~w29987;
assign w30915 = ~pi0019 & w29987;
assign w30916 = ~w30914 & ~w30915;
assign w30917 = pi2065 & ~w29987;
assign w30918 = ~pi0023 & w29987;
assign w30919 = ~w30917 & ~w30918;
assign w30920 = pi2066 & ~w29987;
assign w30921 = ~pi0032 & w29987;
assign w30922 = ~w30920 & ~w30921;
assign w30923 = pi2067 & ~w21638;
assign w30924 = w6177 & w21638;
assign w30925 = ~w30923 & ~w30924;
assign w30926 = pi2068 & ~w21634;
assign w30927 = w4749 & w21634;
assign w30928 = ~w30926 & ~w30927;
assign w30929 = pi2069 & ~w30678;
assign w30930 = pi3516 & w30678;
assign w30931 = ~w30929 & ~w30930;
assign w30932 = pi2070 & ~w29579;
assign w30933 = pi3519 & w29579;
assign w30934 = ~w30932 & ~w30933;
assign w30935 = pi2071 & ~w29579;
assign w30936 = pi3392 & w29579;
assign w30937 = ~w30935 & ~w30936;
assign w30938 = pi2072 & ~w30678;
assign w30939 = pi3504 & w30678;
assign w30940 = ~w30938 & ~w30939;
assign w30941 = pi2073 & ~w29579;
assign w30942 = pi3511 & w29579;
assign w30943 = ~w30941 & ~w30942;
assign w30944 = pi2074 & ~w29897;
assign w30945 = pi3504 & w29897;
assign w30946 = ~w30944 & ~w30945;
assign w30947 = pi2075 & ~w29897;
assign w30948 = pi3511 & w29897;
assign w30949 = ~w30947 & ~w30948;
assign w30950 = pi2076 & ~w30678;
assign w30951 = pi3519 & w30678;
assign w30952 = ~w30950 & ~w30951;
assign w30953 = pi2077 & ~w29897;
assign w30954 = pi3519 & w29897;
assign w30955 = ~w30953 & ~w30954;
assign w30956 = pi2078 & ~w30421;
assign w30957 = pi3688 & w30421;
assign w30958 = ~w30956 & ~w30957;
assign w30959 = ~pi0406 & w29879;
assign w30960 = ~pi0413 & ~w30959;
assign w30961 = pi0408 & ~w30960;
assign w30962 = w21945 & w30959;
assign w30963 = w30961 & ~w30962;
assign w30964 = w29872 & ~w30963;
assign w30965 = pi2079 & ~w29872;
assign w30966 = ~w30964 & ~w30965;
assign w30967 = pi0411 & ~pi0425;
assign w30968 = pi0406 & w30967;
assign w30969 = ~pi0413 & ~w30968;
assign w30970 = pi0408 & ~w30969;
assign w30971 = w21945 & w30968;
assign w30972 = w30970 & ~w30971;
assign w30973 = w29872 & ~w30972;
assign w30974 = pi2080 & ~w29872;
assign w30975 = ~w30973 & ~w30974;
assign w30976 = ~w21945 & w30968;
assign w30977 = w30970 & ~w30976;
assign w30978 = w29872 & ~w30977;
assign w30979 = pi2081 & ~w29872;
assign w30980 = ~w30978 & ~w30979;
assign w30981 = w86 & w113;
assign w30982 = ~w115 & ~w30981;
assign w30983 = w165 & ~w30982;
assign w30984 = w108 & ~w30981;
assign w30985 = ~w165 & w30984;
assign w30986 = w177 & ~w30985;
assign w30987 = ~w30983 & w30986;
assign w30988 = ~w14 & ~w115;
assign w30989 = pi2798 & ~w30988;
assign w30990 = pi2825 & w30989;
assign w30991 = pi2799 & w30990;
assign w30992 = pi2600 & w30991;
assign w30993 = ~pi2082 & ~w30992;
assign w30994 = pi2082 & w30992;
assign w30995 = ~w30993 & ~w30994;
assign w30996 = ~w30987 & w30995;
assign w30997 = ~pi0411 & ~pi0425;
assign w30998 = ~pi0406 & w30997;
assign w30999 = ~pi0413 & ~w30998;
assign w31000 = pi0408 & ~w30999;
assign w31001 = ~w21945 & w30998;
assign w31002 = w31000 & ~w31001;
assign w31003 = w29872 & ~w31002;
assign w31004 = pi2083 & ~w29872;
assign w31005 = ~w31003 & ~w31004;
assign w31006 = pi2084 & ~w21642;
assign w31007 = w6413 & w21642;
assign w31008 = ~w31006 & ~w31007;
assign w31009 = ~pi0598 & w40209;
assign w31010 = ~w30484 & w31009;
assign w31011 = pi2085 & ~w31009;
assign w31012 = ~w31010 & ~w31011;
assign w31013 = pi0406 & w30997;
assign w31014 = ~pi0413 & ~w31013;
assign w31015 = pi0408 & ~w31014;
assign w31016 = w21945 & w31013;
assign w31017 = w31015 & ~w31016;
assign w31018 = w29872 & ~w31017;
assign w31019 = pi2086 & ~w29872;
assign w31020 = ~w31018 & ~w31019;
assign w31021 = pi2087 & ~w21642;
assign w31022 = w4380 & w21642;
assign w31023 = ~w31021 & ~w31022;
assign w31024 = pi2088 & ~w21638;
assign w31025 = w5635 & w21638;
assign w31026 = ~w31024 & ~w31025;
assign w31027 = pi2089 & ~w21642;
assign w31028 = w6177 & w21642;
assign w31029 = ~w31027 & ~w31028;
assign w31030 = ~w4141 & w30202;
assign w31031 = pi2090 & ~w30202;
assign w31032 = ~w31030 & ~w31031;
assign w31033 = ~w6177 & w30202;
assign w31034 = pi2091 & ~w30202;
assign w31035 = ~w31033 & ~w31034;
assign w31036 = ~w40134 & w30202;
assign w31037 = pi2092 & ~w30202;
assign w31038 = ~w31036 & ~w31037;
assign w31039 = ~w4380 & w30202;
assign w31040 = pi2093 & ~w30202;
assign w31041 = ~w31039 & ~w31040;
assign w31042 = ~w5914 & w30202;
assign w31043 = pi2094 & ~w30202;
assign w31044 = ~w31042 & ~w31043;
assign w31045 = ~w8240 & w30202;
assign w31046 = pi2095 & ~w30202;
assign w31047 = ~w31045 & ~w31046;
assign w31048 = ~w1308 & w30202;
assign w31049 = pi2096 & ~w30202;
assign w31050 = ~w31048 & ~w31049;
assign w31051 = ~w1639 & w30202;
assign w31052 = pi2097 & ~w30202;
assign w31053 = ~w31051 & ~w31052;
assign w31054 = ~w3711 & w30202;
assign w31055 = pi2098 & ~w30202;
assign w31056 = ~w31054 & ~w31055;
assign w31057 = w10741 & ~w18313;
assign w31058 = pi2099 & ~pi3136;
assign w31059 = w1639 & w30284;
assign w31060 = w1274 & w23861;
assign w31061 = ~w1639 & w31060;
assign w31062 = ~pi3243 & pi3317;
assign w31063 = pi3243 & ~pi3317;
assign w31064 = ~w31062 & ~w31063;
assign w31065 = pi1749 & ~pi1761;
assign w31066 = ~w31064 & w31065;
assign w31067 = ~pi2101 & ~w31066;
assign w31068 = ~w31060 & w31067;
assign w31069 = ~w31061 & ~w31068;
assign w31070 = ~w1308 & w31060;
assign w31071 = ~pi3219 & pi3318;
assign w31072 = pi3219 & ~pi3318;
assign w31073 = ~w31071 & ~w31072;
assign w31074 = pi1750 & ~pi1762;
assign w31075 = ~w31073 & w31074;
assign w31076 = ~pi2102 & ~w31075;
assign w31077 = ~w31060 & w31076;
assign w31078 = ~w31070 & ~w31077;
assign w31079 = ~w3195 & w31060;
assign w31080 = ~pi3241 & pi3351;
assign w31081 = pi3241 & ~pi3351;
assign w31082 = ~w31080 & ~w31081;
assign w31083 = pi1751 & ~pi1857;
assign w31084 = ~w31082 & w31083;
assign w31085 = ~pi2103 & ~w31084;
assign w31086 = ~w31060 & w31085;
assign w31087 = ~w31079 & ~w31086;
assign w31088 = ~w40134 & w31060;
assign w31089 = ~pi3220 & pi3349;
assign w31090 = pi3220 & ~pi3349;
assign w31091 = ~w31089 & ~w31090;
assign w31092 = pi1752 & ~pi1763;
assign w31093 = ~w31091 & w31092;
assign w31094 = ~pi2104 & ~w31093;
assign w31095 = ~w31060 & w31094;
assign w31096 = ~w31088 & ~w31095;
assign w31097 = ~w6413 & w31060;
assign w31098 = ~pi3242 & pi3346;
assign w31099 = pi3242 & ~pi3346;
assign w31100 = ~w31098 & ~w31099;
assign w31101 = pi1753 & ~pi1764;
assign w31102 = ~w31100 & w31101;
assign w31103 = ~pi2105 & ~w31102;
assign w31104 = ~w31060 & w31103;
assign w31105 = ~w31097 & ~w31104;
assign w31106 = ~w4380 & w31060;
assign w31107 = ~pi3221 & pi3345;
assign w31108 = pi3221 & ~pi3345;
assign w31109 = ~w31107 & ~w31108;
assign w31110 = pi1754 & ~pi1765;
assign w31111 = ~w31109 & w31110;
assign w31112 = ~pi2106 & ~w31111;
assign w31113 = ~w31060 & w31112;
assign w31114 = ~w31106 & ~w31113;
assign w31115 = ~w5320 & w31060;
assign w31116 = ~pi3218 & pi3348;
assign w31117 = pi3218 & ~pi3348;
assign w31118 = ~w31116 & ~w31117;
assign w31119 = pi1755 & ~pi1858;
assign w31120 = ~w31118 & w31119;
assign w31121 = ~pi2107 & ~w31120;
assign w31122 = ~w31060 & w31121;
assign w31123 = ~w31115 & ~w31122;
assign w31124 = ~w4749 & w31060;
assign w31125 = ~pi3223 & pi3320;
assign w31126 = pi3223 & ~pi3320;
assign w31127 = ~w31125 & ~w31126;
assign w31128 = pi1757 & ~pi1767;
assign w31129 = ~w31127 & w31128;
assign w31130 = ~pi2108 & ~w31129;
assign w31131 = ~w31060 & w31130;
assign w31132 = ~w31124 & ~w31131;
assign w31133 = ~w8240 & w31060;
assign w31134 = ~pi3224 & pi3357;
assign w31135 = pi3224 & ~pi3357;
assign w31136 = ~w31134 & ~w31135;
assign w31137 = pi1758 & ~pi1768;
assign w31138 = ~w31136 & w31137;
assign w31139 = ~pi2109 & ~w31138;
assign w31140 = ~w31060 & w31139;
assign w31141 = ~w31133 & ~w31140;
assign w31142 = ~w3711 & w31060;
assign w31143 = ~pi3225 & pi3321;
assign w31144 = pi3225 & ~pi3321;
assign w31145 = ~w31143 & ~w31144;
assign w31146 = pi1760 & ~pi1769;
assign w31147 = ~w31145 & w31146;
assign w31148 = ~pi2110 & ~w31147;
assign w31149 = ~w31060 & w31148;
assign w31150 = ~w31142 & ~w31149;
assign w31151 = pi2111 & ~w30315;
assign w31152 = w1308 & w30315;
assign w31153 = ~w31151 & ~w31152;
assign w31154 = pi2112 & w30364;
assign w31155 = w6598 & ~w30364;
assign w31156 = w4797 & w31155;
assign w31157 = ~w31154 & ~w31156;
assign w31158 = pi2113 & w30994;
assign w31159 = ~pi2113 & ~w30994;
assign w31160 = ~w31158 & ~w31159;
assign w31161 = ~w30987 & w31160;
assign w31162 = pi0565 & w28743;
assign w31163 = w28739 & w31162;
assign w31164 = ~pi3216 & ~pi3256;
assign w31165 = w31163 & ~w31164;
assign w31166 = pi2114 & ~w28750;
assign w31167 = ~w28747 & w31166;
assign w31168 = ~w31165 & ~w31167;
assign w31169 = pi2115 & ~w30421;
assign w31170 = pi3690 & w30421;
assign w31171 = ~w31169 & ~w31170;
assign w31172 = pi2116 & ~w30421;
assign w31173 = pi3689 & w30421;
assign w31174 = ~w31172 & ~w31173;
assign w31175 = pi2117 & ~w30421;
assign w31176 = pi3687 & w30421;
assign w31177 = ~w31175 & ~w31176;
assign w31178 = pi2118 & ~w30421;
assign w31179 = pi3686 & w30421;
assign w31180 = ~w31178 & ~w31179;
assign w31181 = pi2119 & ~w30421;
assign w31182 = pi3685 & w30421;
assign w31183 = ~w31181 & ~w31182;
assign w31184 = pi2120 & ~w30421;
assign w31185 = pi3684 & w30421;
assign w31186 = ~w31184 & ~w31185;
assign w31187 = pi2121 & ~w30421;
assign w31188 = pi3683 & w30421;
assign w31189 = ~w31187 & ~w31188;
assign w31190 = pi2122 & ~w21638;
assign w31191 = w1308 & w21638;
assign w31192 = ~w31190 & ~w31191;
assign w31193 = ~w8081 & w31060;
assign w31194 = ~pi3240 & pi3340;
assign w31195 = pi3240 & ~pi3340;
assign w31196 = ~w31194 & ~w31195;
assign w31197 = pi1759 & ~pi1854;
assign w31198 = ~w31196 & w31197;
assign w31199 = ~pi2123 & ~w31198;
assign w31200 = ~w31060 & w31199;
assign w31201 = ~w31193 & ~w31200;
assign w31202 = ~pi0711 & w40209;
assign w31203 = pi2124 & ~w31202;
assign w31204 = w40189 & w31202;
assign w31205 = ~w31203 & ~w31204;
assign w31206 = pi2125 & ~w31202;
assign w31207 = w40191 & w31202;
assign w31208 = ~w31206 & ~w31207;
assign w31209 = pi2126 & ~w31202;
assign w31210 = w40174 & w31202;
assign w31211 = ~w31209 & ~w31210;
assign w31212 = pi2127 & ~w31202;
assign w31213 = w14325 & w31202;
assign w31214 = ~w31212 & ~w31213;
assign w31215 = pi2128 & ~w31202;
assign w31216 = w14962 & w31202;
assign w31217 = ~w31215 & ~w31216;
assign w31218 = pi2129 & ~w31202;
assign w31219 = w40168 & w31202;
assign w31220 = ~w31218 & ~w31219;
assign w31221 = pi2130 & ~w31202;
assign w31222 = w40176 & w31202;
assign w31223 = ~w31221 & ~w31222;
assign w31224 = pi2131 & ~w31202;
assign w31225 = w13916 & w31202;
assign w31226 = ~w31224 & ~w31225;
assign w31227 = pi2132 & ~w31202;
assign w31228 = w40159 & w31202;
assign w31229 = ~w31227 & ~w31228;
assign w31230 = ~w10746 & w31202;
assign w31231 = pi2133 & ~w31202;
assign w31232 = ~w31230 & ~w31231;
assign w31233 = pi2134 & ~w31202;
assign w31234 = w16629 & w31202;
assign w31235 = ~w31233 & ~w31234;
assign w31236 = pi2135 & ~w31202;
assign w31237 = w16739 & w31202;
assign w31238 = ~w31236 & ~w31237;
assign w31239 = pi2136 & ~w31202;
assign w31240 = ~w16842 & w31202;
assign w31241 = ~w31239 & ~w31240;
assign w31242 = pi2137 & ~w31202;
assign w31243 = w15978 & w31202;
assign w31244 = ~w31242 & ~w31243;
assign w31245 = pi2138 & ~w31202;
assign w31246 = w15171 & w31202;
assign w31247 = ~w31245 & ~w31246;
assign w31248 = pi2139 & ~w31202;
assign w31249 = w40171 & w31202;
assign w31250 = ~w31248 & ~w31249;
assign w31251 = ~pi2140 & w6684;
assign w31252 = ~w28578 & w30761;
assign w31253 = ~w31251 & ~w31252;
assign w31254 = ~w5914 & w31060;
assign w31255 = ~pi3222 & pi3319;
assign w31256 = pi3222 & ~pi3319;
assign w31257 = ~w31255 & ~w31256;
assign w31258 = pi1756 & ~pi1766;
assign w31259 = ~w31257 & w31258;
assign w31260 = ~pi2141 & ~w31259;
assign w31261 = ~w31060 & w31260;
assign w31262 = ~w31254 & ~w31261;
assign w31263 = ~pi2142 & w6684;
assign w31264 = ~w30445 & ~w31263;
assign w31265 = pi2143 & w10;
assign w31266 = w10741 & ~w31265;
assign w31267 = w10689 & ~w13946;
assign w31268 = ~w30452 & w31009;
assign w31269 = pi2144 & ~w31009;
assign w31270 = ~w31268 & ~w31269;
assign w31271 = ~w30460 & w31009;
assign w31272 = pi2145 & ~w31009;
assign w31273 = ~w31271 & ~w31272;
assign w31274 = ~w30468 & w31009;
assign w31275 = pi2146 & ~w31009;
assign w31276 = ~w31274 & ~w31275;
assign w31277 = ~w30476 & w31009;
assign w31278 = pi2147 & ~w31009;
assign w31279 = ~w31277 & ~w31278;
assign w31280 = ~w30492 & w31009;
assign w31281 = pi2148 & ~w31009;
assign w31282 = ~w31280 & ~w31281;
assign w31283 = ~w30500 & w31009;
assign w31284 = pi2149 & ~w31009;
assign w31285 = ~w31283 & ~w31284;
assign w31286 = ~w30508 & w31009;
assign w31287 = pi2150 & ~w31009;
assign w31288 = ~w31286 & ~w31287;
assign w31289 = ~w29844 & w31009;
assign w31290 = pi2151 & ~w31009;
assign w31291 = ~w31289 & ~w31290;
assign w31292 = ~w30516 & w31009;
assign w31293 = pi2152 & ~w31009;
assign w31294 = ~w31292 & ~w31293;
assign w31295 = ~w29852 & w31009;
assign w31296 = pi2153 & ~w31009;
assign w31297 = ~w31295 & ~w31296;
assign w31298 = ~w30524 & w31009;
assign w31299 = pi2154 & ~w31009;
assign w31300 = ~w31298 & ~w31299;
assign w31301 = ~w30532 & w31009;
assign w31302 = pi2155 & ~w31009;
assign w31303 = ~w31301 & ~w31302;
assign w31304 = ~w30540 & w31009;
assign w31305 = pi2156 & ~w31009;
assign w31306 = ~w31304 & ~w31305;
assign w31307 = ~w30548 & w31009;
assign w31308 = pi2157 & ~w31009;
assign w31309 = ~w31307 & ~w31308;
assign w31310 = ~w17426 & w31009;
assign w31311 = pi2158 & ~w31009;
assign w31312 = ~w31310 & ~w31311;
assign w31313 = w17601 & ~w29847;
assign w31314 = ~pi2159 & ~w17601;
assign w31315 = ~w31313 & ~w31314;
assign w31316 = w17601 & ~w29855;
assign w31317 = ~pi2160 & ~w17601;
assign w31318 = ~w31316 & ~w31317;
assign w31319 = ~pi0649 & w40209;
assign w31320 = pi2161 & ~w31319;
assign w31321 = w40189 & w31319;
assign w31322 = ~w31320 & ~w31321;
assign w31323 = pi2162 & ~w31319;
assign w31324 = w40191 & w31319;
assign w31325 = ~w31323 & ~w31324;
assign w31326 = pi2163 & ~w31319;
assign w31327 = w40174 & w31319;
assign w31328 = ~w31326 & ~w31327;
assign w31329 = pi2164 & ~w31319;
assign w31330 = w14325 & w31319;
assign w31331 = ~w31329 & ~w31330;
assign w31332 = pi2165 & ~w31319;
assign w31333 = w14962 & w31319;
assign w31334 = ~w31332 & ~w31333;
assign w31335 = pi2166 & ~w31319;
assign w31336 = w40168 & w31319;
assign w31337 = ~w31335 & ~w31336;
assign w31338 = pi2167 & ~w31319;
assign w31339 = w40176 & w31319;
assign w31340 = ~w31338 & ~w31339;
assign w31341 = pi2168 & ~w31319;
assign w31342 = w13916 & w31319;
assign w31343 = ~w31341 & ~w31342;
assign w31344 = pi2169 & ~w31319;
assign w31345 = w40159 & w31319;
assign w31346 = ~w31344 & ~w31345;
assign w31347 = ~w10746 & w31319;
assign w31348 = pi2170 & ~w31319;
assign w31349 = ~w31347 & ~w31348;
assign w31350 = pi2171 & ~w31319;
assign w31351 = w16629 & w31319;
assign w31352 = ~w31350 & ~w31351;
assign w31353 = pi2172 & ~w31319;
assign w31354 = w16739 & w31319;
assign w31355 = ~w31353 & ~w31354;
assign w31356 = pi2173 & ~w31319;
assign w31357 = ~w16842 & w31319;
assign w31358 = ~w31356 & ~w31357;
assign w31359 = pi2174 & ~w31319;
assign w31360 = w15978 & w31319;
assign w31361 = ~w31359 & ~w31360;
assign w31362 = pi2175 & ~w31319;
assign w31363 = w15171 & w31319;
assign w31364 = ~w31362 & ~w31363;
assign w31365 = pi2176 & ~w31319;
assign w31366 = w40171 & w31319;
assign w31367 = ~w31365 & ~w31366;
assign w31368 = ~pi0575 & w40209;
assign w31369 = pi2177 & ~w31368;
assign w31370 = w40189 & w31368;
assign w31371 = ~w31369 & ~w31370;
assign w31372 = pi2178 & ~w31368;
assign w31373 = w40191 & w31368;
assign w31374 = ~w31372 & ~w31373;
assign w31375 = pi2179 & ~w31368;
assign w31376 = w40174 & w31368;
assign w31377 = ~w31375 & ~w31376;
assign w31378 = pi2180 & ~w31368;
assign w31379 = w14325 & w31368;
assign w31380 = ~w31378 & ~w31379;
assign w31381 = pi2181 & ~w31368;
assign w31382 = w14962 & w31368;
assign w31383 = ~w31381 & ~w31382;
assign w31384 = pi2182 & ~w31368;
assign w31385 = w40168 & w31368;
assign w31386 = ~w31384 & ~w31385;
assign w31387 = pi2183 & ~w31368;
assign w31388 = w40176 & w31368;
assign w31389 = ~w31387 & ~w31388;
assign w31390 = pi2184 & ~w31368;
assign w31391 = w13916 & w31368;
assign w31392 = ~w31390 & ~w31391;
assign w31393 = pi2185 & ~w31368;
assign w31394 = w40159 & w31368;
assign w31395 = ~w31393 & ~w31394;
assign w31396 = ~w10746 & w31368;
assign w31397 = pi2186 & ~w31368;
assign w31398 = ~w31396 & ~w31397;
assign w31399 = pi2187 & ~w31368;
assign w31400 = w16629 & w31368;
assign w31401 = ~w31399 & ~w31400;
assign w31402 = pi2188 & ~w31368;
assign w31403 = w16739 & w31368;
assign w31404 = ~w31402 & ~w31403;
assign w31405 = pi2189 & ~w31368;
assign w31406 = ~w16842 & w31368;
assign w31407 = ~w31405 & ~w31406;
assign w31408 = pi2190 & ~w31368;
assign w31409 = w15978 & w31368;
assign w31410 = ~w31408 & ~w31409;
assign w31411 = pi2191 & ~w31368;
assign w31412 = w15171 & w31368;
assign w31413 = ~w31411 & ~w31412;
assign w31414 = pi2192 & ~w31368;
assign w31415 = w40171 & w31368;
assign w31416 = ~w31414 & ~w31415;
assign w31417 = w7051 & ~w19954;
assign w31418 = ~pi2193 & w19954;
assign w31419 = w6682 & ~w31418;
assign w31420 = ~w31417 & w31419;
assign w31421 = ~w21945 & w31013;
assign w31422 = w31015 & ~w31421;
assign w31423 = w29872 & ~w31422;
assign w31424 = pi2194 & ~w29872;
assign w31425 = ~w31423 & ~w31424;
assign w31426 = ~pi0406 & w29863;
assign w31427 = ~pi0413 & ~w31426;
assign w31428 = pi0408 & ~w31427;
assign w31429 = ~w21945 & w31426;
assign w31430 = w31428 & ~w31429;
assign w31431 = w29872 & ~w31430;
assign w31432 = pi2195 & ~w29872;
assign w31433 = ~w31431 & ~w31432;
assign w31434 = w21945 & w31426;
assign w31435 = w31428 & ~w31434;
assign w31436 = w29872 & ~w31435;
assign w31437 = pi2196 & ~w29872;
assign w31438 = ~w31436 & ~w31437;
assign w31439 = ~w21945 & w30959;
assign w31440 = w30961 & ~w31439;
assign w31441 = w29872 & ~w31440;
assign w31442 = pi2197 & ~w29872;
assign w31443 = ~w31441 & ~w31442;
assign w31444 = ~pi0406 & w30967;
assign w31445 = ~pi0413 & ~w31444;
assign w31446 = pi0408 & ~w31445;
assign w31447 = w21945 & w31444;
assign w31448 = w31446 & ~w31447;
assign w31449 = w29872 & ~w31448;
assign w31450 = pi2198 & ~w29872;
assign w31451 = ~w31449 & ~w31450;
assign w31452 = ~w21945 & w31444;
assign w31453 = w31446 & ~w31452;
assign w31454 = w29872 & ~w31453;
assign w31455 = pi2199 & ~w29872;
assign w31456 = ~w31454 & ~w31455;
assign w31457 = w21945 & w30998;
assign w31458 = w31000 & ~w31457;
assign w31459 = w29872 & ~w31458;
assign w31460 = pi2200 & ~w29872;
assign w31461 = ~w31459 & ~w31460;
assign w31462 = pi2201 & ~w21536;
assign w31463 = w4141 & w21536;
assign w31464 = ~w31462 & ~w31463;
assign w31465 = pi2202 & ~w21536;
assign w31466 = w6177 & w21536;
assign w31467 = ~w31465 & ~w31466;
assign w31468 = pi2203 & ~w21536;
assign w31469 = w3195 & w21536;
assign w31470 = ~w31468 & ~w31469;
assign w31471 = pi2204 & ~w21536;
assign w31472 = w40134 & w21536;
assign w31473 = ~w31471 & ~w31472;
assign w31474 = pi2205 & ~w21536;
assign w31475 = w6413 & w21536;
assign w31476 = ~w31474 & ~w31475;
assign w31477 = pi2206 & ~w21536;
assign w31478 = w4380 & w21536;
assign w31479 = ~w31477 & ~w31478;
assign w31480 = pi2207 & ~w21536;
assign w31481 = w5320 & w21536;
assign w31482 = ~w31480 & ~w31481;
assign w31483 = pi2208 & ~w21536;
assign w31484 = w5914 & w21536;
assign w31485 = ~w31483 & ~w31484;
assign w31486 = pi2209 & ~w21536;
assign w31487 = w4749 & w21536;
assign w31488 = ~w31486 & ~w31487;
assign w31489 = pi2210 & ~w21536;
assign w31490 = w1639 & w21536;
assign w31491 = ~w31489 & ~w31490;
assign w31492 = pi2211 & ~w21536;
assign w31493 = w1308 & w21536;
assign w31494 = ~w31492 & ~w31493;
assign w31495 = pi2212 & ~w21536;
assign w31496 = w5635 & w21536;
assign w31497 = ~w31495 & ~w31496;
assign w31498 = pi2213 & ~w21536;
assign w31499 = w5053 & w21536;
assign w31500 = ~w31498 & ~w31499;
assign w31501 = pi2214 & ~w21536;
assign w31502 = w3711 & w21536;
assign w31503 = ~w31501 & ~w31502;
assign w31504 = w4141 & w21533;
assign w31505 = ~w21895 & ~w31504;
assign w31506 = pi2216 & ~w21533;
assign w31507 = w6177 & w21533;
assign w31508 = ~w31506 & ~w31507;
assign w31509 = pi2217 & ~w21533;
assign w31510 = w3195 & w21533;
assign w31511 = ~w31509 & ~w31510;
assign w31512 = pi2218 & ~w21533;
assign w31513 = w40134 & w21533;
assign w31514 = ~w31512 & ~w31513;
assign w31515 = pi2219 & ~w21533;
assign w31516 = w6413 & w21533;
assign w31517 = ~w31515 & ~w31516;
assign w31518 = pi2220 & ~w21533;
assign w31519 = w4380 & w21533;
assign w31520 = ~w31518 & ~w31519;
assign w31521 = pi2221 & ~w21533;
assign w31522 = w5320 & w21533;
assign w31523 = ~w31521 & ~w31522;
assign w31524 = pi2222 & ~w21533;
assign w31525 = w5914 & w21533;
assign w31526 = ~w31524 & ~w31525;
assign w31527 = pi2223 & ~w21533;
assign w31528 = w4749 & w21533;
assign w31529 = ~w31527 & ~w31528;
assign w31530 = pi2224 & ~w21533;
assign w31531 = w1639 & w21533;
assign w31532 = ~w31530 & ~w31531;
assign w31533 = pi2225 & ~w21533;
assign w31534 = w1308 & w21533;
assign w31535 = ~w31533 & ~w31534;
assign w31536 = pi2226 & ~w21533;
assign w31537 = w5635 & w21533;
assign w31538 = ~w31536 & ~w31537;
assign w31539 = pi2227 & ~w21533;
assign w31540 = w5053 & w21533;
assign w31541 = ~w31539 & ~w31540;
assign w31542 = pi2228 & ~w21533;
assign w31543 = w3711 & w21533;
assign w31544 = ~w31542 & ~w31543;
assign w31545 = pi2229 & ~w21530;
assign w31546 = w4141 & w21530;
assign w31547 = ~w31545 & ~w31546;
assign w31548 = pi2230 & ~w21530;
assign w31549 = w6177 & w21530;
assign w31550 = ~w31548 & ~w31549;
assign w31551 = w3195 & w21530;
assign w31552 = ~w22250 & ~w31551;
assign w31553 = pi2232 & ~w21530;
assign w31554 = w40134 & w21530;
assign w31555 = ~w31553 & ~w31554;
assign w31556 = w6413 & w21530;
assign w31557 = ~w21560 & ~w31556;
assign w31558 = w4380 & w21530;
assign w31559 = ~w21573 & ~w31558;
assign w31560 = pi2235 & ~w21530;
assign w31561 = w5320 & w21530;
assign w31562 = ~w31560 & ~w31561;
assign w31563 = w5914 & w21530;
assign w31564 = ~w21598 & ~w31563;
assign w31565 = pi2237 & ~w21530;
assign w31566 = w4749 & w21530;
assign w31567 = ~w31565 & ~w31566;
assign w31568 = pi2238 & ~w21530;
assign w31569 = w1639 & w21530;
assign w31570 = ~w31568 & ~w31569;
assign w31571 = pi2239 & ~w21530;
assign w31572 = w1308 & w21530;
assign w31573 = ~w31571 & ~w31572;
assign w31574 = w5635 & w21530;
assign w31575 = ~w21920 & ~w31574;
assign w31576 = pi2241 & ~w21530;
assign w31577 = w5053 & w21530;
assign w31578 = ~w31576 & ~w31577;
assign w31579 = w3711 & w21530;
assign w31580 = ~w22275 & ~w31579;
assign w31581 = pi2243 & ~w21539;
assign w31582 = w4141 & w21539;
assign w31583 = ~w31581 & ~w31582;
assign w31584 = pi2244 & ~w21539;
assign w31585 = w6177 & w21539;
assign w31586 = ~w31584 & ~w31585;
assign w31587 = pi2245 & ~w21539;
assign w31588 = w3195 & w21539;
assign w31589 = ~w31587 & ~w31588;
assign w31590 = pi2246 & ~w21539;
assign w31591 = w40134 & w21539;
assign w31592 = ~w31590 & ~w31591;
assign w31593 = pi2247 & ~w21539;
assign w31594 = w6413 & w21539;
assign w31595 = ~w31593 & ~w31594;
assign w31596 = pi2248 & ~w21539;
assign w31597 = w4380 & w21539;
assign w31598 = ~w31596 & ~w31597;
assign w31599 = pi2249 & ~w21539;
assign w31600 = w5320 & w21539;
assign w31601 = ~w31599 & ~w31600;
assign w31602 = pi2250 & ~w21539;
assign w31603 = w5914 & w21539;
assign w31604 = ~w31602 & ~w31603;
assign w31605 = pi2251 & ~w21539;
assign w31606 = w4749 & w21539;
assign w31607 = ~w31605 & ~w31606;
assign w31608 = pi2252 & ~w21539;
assign w31609 = w1639 & w21539;
assign w31610 = ~w31608 & ~w31609;
assign w31611 = pi2253 & ~w21539;
assign w31612 = w1308 & w21539;
assign w31613 = ~w31611 & ~w31612;
assign w31614 = pi2254 & ~w21539;
assign w31615 = w5635 & w21539;
assign w31616 = ~w31614 & ~w31615;
assign w31617 = pi2255 & ~w21539;
assign w31618 = w5053 & w21539;
assign w31619 = ~w31617 & ~w31618;
assign w31620 = pi2256 & ~w21539;
assign w31621 = w3711 & w21539;
assign w31622 = ~w31620 & ~w31621;
assign w31623 = ~w23216 & w23420;
assign w31624 = ~w23422 & ~w31623;
assign w31625 = w8802 & ~w23216;
assign w31626 = ~pi2258 & w23216;
assign w31627 = ~w31625 & ~w31626;
assign w31628 = w8745 & ~w23216;
assign w31629 = pi2259 & w23216;
assign w31630 = ~w31628 & ~w31629;
assign w31631 = w8699 & ~w23216;
assign w31632 = ~w23469 & ~w31631;
assign w31633 = w844 & w23420;
assign w31634 = ~w23424 & ~w31633;
assign w31635 = pi2262 & ~w844;
assign w31636 = w844 & ~w8802;
assign w31637 = ~w31635 & ~w31636;
assign w31638 = w844 & ~w23437;
assign w31639 = ~pi2263 & ~w844;
assign w31640 = ~w31638 & ~w31639;
assign w31641 = w844 & ~w8745;
assign w31642 = ~pi2264 & ~w844;
assign w31643 = ~w31641 & ~w31642;
assign w31644 = w844 & ~w8699;
assign w31645 = ~pi2265 & ~w844;
assign w31646 = ~w31644 & ~w31645;
assign w31647 = w844 & ~w8667;
assign w31648 = ~w23481 & ~w31647;
assign w31649 = w844 & ~w23496;
assign w31650 = ~w23498 & ~w31649;
assign w31651 = w844 & w22214;
assign w31652 = ~w23514 & ~w31651;
assign w31653 = pi2269 & ~w844;
assign w31654 = w844 & ~w22222;
assign w31655 = ~w31653 & ~w31654;
assign w31656 = w844 & ~w8560;
assign w31657 = ~pi2270 & ~w844;
assign w31658 = ~w31656 & ~w31657;
assign w31659 = w856 & ~w23420;
assign w31660 = ~pi2271 & ~w856;
assign w31661 = ~w31659 & ~w31660;
assign w31662 = w856 & ~w8802;
assign w31663 = ~w23225 & ~w31662;
assign w31664 = w856 & w8745;
assign w31665 = ~w23455 & ~w31664;
assign w31666 = pi2274 & ~w856;
assign w31667 = w856 & ~w8667;
assign w31668 = ~w31666 & ~w31667;
assign w31669 = w849 & w8826;
assign w31670 = ~w24431 & ~w31669;
assign w31671 = w849 & ~w24445;
assign w31672 = ~pi2276 & ~w849;
assign w31673 = ~w31671 & ~w31672;
assign w31674 = w849 & ~w24462;
assign w31675 = ~pi2277 & ~w849;
assign w31676 = ~w31674 & ~w31675;
assign w31677 = pi2278 & ~w849;
assign w31678 = w849 & ~w24479;
assign w31679 = ~w31677 & ~w31678;
assign w31680 = pi2279 & ~w21634;
assign w31681 = w4141 & w21634;
assign w31682 = ~w31680 & ~w31681;
assign w31683 = pi2280 & ~w21634;
assign w31684 = w6177 & w21634;
assign w31685 = ~w31683 & ~w31684;
assign w31686 = pi2281 & ~w21634;
assign w31687 = w3195 & w21634;
assign w31688 = ~w31686 & ~w31687;
assign w31689 = pi2282 & ~w21634;
assign w31690 = w40134 & w21634;
assign w31691 = ~w31689 & ~w31690;
assign w31692 = pi2283 & ~w21634;
assign w31693 = w6413 & w21634;
assign w31694 = ~w31692 & ~w31693;
assign w31695 = pi2284 & ~w21634;
assign w31696 = w4380 & w21634;
assign w31697 = ~w31695 & ~w31696;
assign w31698 = pi2285 & ~w21634;
assign w31699 = w5320 & w21634;
assign w31700 = ~w31698 & ~w31699;
assign w31701 = pi2286 & ~w21634;
assign w31702 = w5914 & w21634;
assign w31703 = ~w31701 & ~w31702;
assign w31704 = pi2287 & ~w21634;
assign w31705 = w1639 & w21634;
assign w31706 = ~w31704 & ~w31705;
assign w31707 = pi2288 & ~w21634;
assign w31708 = w1308 & w21634;
assign w31709 = ~w31707 & ~w31708;
assign w31710 = pi2289 & ~w21634;
assign w31711 = w5635 & w21634;
assign w31712 = ~w31710 & ~w31711;
assign w31713 = pi2290 & ~w21634;
assign w31714 = w5053 & w21634;
assign w31715 = ~w31713 & ~w31714;
assign w31716 = pi2291 & ~w21634;
assign w31717 = w3711 & w21634;
assign w31718 = ~w31716 & ~w31717;
assign w31719 = pi2292 & ~w21638;
assign w31720 = w4141 & w21638;
assign w31721 = ~w31719 & ~w31720;
assign w31722 = pi2293 & ~w21638;
assign w31723 = w3195 & w21638;
assign w31724 = ~w31722 & ~w31723;
assign w31725 = pi2294 & ~w21638;
assign w31726 = w40134 & w21638;
assign w31727 = ~w31725 & ~w31726;
assign w31728 = pi2295 & ~w21638;
assign w31729 = w6413 & w21638;
assign w31730 = ~w31728 & ~w31729;
assign w31731 = pi2296 & ~w21638;
assign w31732 = w4380 & w21638;
assign w31733 = ~w31731 & ~w31732;
assign w31734 = pi2297 & ~w21638;
assign w31735 = w5320 & w21638;
assign w31736 = ~w31734 & ~w31735;
assign w31737 = pi2298 & ~w21638;
assign w31738 = w5914 & w21638;
assign w31739 = ~w31737 & ~w31738;
assign w31740 = pi2299 & ~w21638;
assign w31741 = w4749 & w21638;
assign w31742 = ~w31740 & ~w31741;
assign w31743 = pi2300 & ~w21638;
assign w31744 = w1639 & w21638;
assign w31745 = ~w31743 & ~w31744;
assign w31746 = pi2301 & ~w21638;
assign w31747 = w5053 & w21638;
assign w31748 = ~w31746 & ~w31747;
assign w31749 = pi2302 & ~w21638;
assign w31750 = w3711 & w21638;
assign w31751 = ~w31749 & ~w31750;
assign w31752 = w4141 & w21642;
assign w31753 = ~w21650 & ~w31752;
assign w31754 = pi2304 & ~w21642;
assign w31755 = w3195 & w21642;
assign w31756 = ~w31754 & ~w31755;
assign w31757 = pi2305 & ~w21642;
assign w31758 = w40134 & w21642;
assign w31759 = ~w31757 & ~w31758;
assign w31760 = pi2306 & ~w21642;
assign w31761 = w5320 & w21642;
assign w31762 = ~w31760 & ~w31761;
assign w31763 = pi2307 & ~w21642;
assign w31764 = w5914 & w21642;
assign w31765 = ~w31763 & ~w31764;
assign w31766 = w4749 & w21642;
assign w31767 = ~w21724 & ~w31766;
assign w31768 = w1639 & w21642;
assign w31769 = ~w21737 & ~w31768;
assign w31770 = w1308 & w21642;
assign w31771 = ~w22447 & ~w31770;
assign w31772 = pi2311 & ~w21642;
assign w31773 = w5635 & w21642;
assign w31774 = ~w31772 & ~w31773;
assign w31775 = pi2312 & ~w21642;
assign w31776 = w5053 & w21642;
assign w31777 = ~w31775 & ~w31776;
assign w31778 = pi2313 & ~w21642;
assign w31779 = w3711 & w21642;
assign w31780 = ~w31778 & ~w31779;
assign w31781 = pi2314 & ~w21632;
assign w31782 = w4141 & w21632;
assign w31783 = ~w31781 & ~w31782;
assign w31784 = pi2315 & ~w21632;
assign w31785 = w6177 & w21632;
assign w31786 = ~w31784 & ~w31785;
assign w31787 = pi2316 & ~w21632;
assign w31788 = w3195 & w21632;
assign w31789 = ~w31787 & ~w31788;
assign w31790 = pi2317 & ~w21632;
assign w31791 = w40134 & w21632;
assign w31792 = ~w31790 & ~w31791;
assign w31793 = pi2318 & ~w21632;
assign w31794 = w6413 & w21632;
assign w31795 = ~w31793 & ~w31794;
assign w31796 = pi2319 & ~w21632;
assign w31797 = w4380 & w21632;
assign w31798 = ~w31796 & ~w31797;
assign w31799 = pi2320 & ~w21632;
assign w31800 = w5320 & w21632;
assign w31801 = ~w31799 & ~w31800;
assign w31802 = w5914 & w21632;
assign w31803 = ~w21711 & ~w31802;
assign w31804 = pi2322 & ~w21632;
assign w31805 = w4749 & w21632;
assign w31806 = ~w31804 & ~w31805;
assign w31807 = pi2323 & ~w21632;
assign w31808 = w1639 & w21632;
assign w31809 = ~w31807 & ~w31808;
assign w31810 = w1308 & w21632;
assign w31811 = ~w22444 & ~w31810;
assign w31812 = pi2325 & ~w21632;
assign w31813 = w5635 & w21632;
assign w31814 = ~w31812 & ~w31813;
assign w31815 = pi2326 & ~w21632;
assign w31816 = w5053 & w21632;
assign w31817 = ~w31815 & ~w31816;
assign w31818 = w3711 & w21632;
assign w31819 = ~w21774 & ~w31818;
assign w31820 = ~pi2472 & w29897;
assign w31821 = pi2328 & ~w29897;
assign w31822 = ~w31820 & ~w31821;
assign w31823 = ~pi2400 & w29897;
assign w31824 = pi2329 & ~w29897;
assign w31825 = ~w31823 & ~w31824;
assign w31826 = pi2330 & ~w29897;
assign w31827 = pi3517 & w29897;
assign w31828 = ~w31826 & ~w31827;
assign w31829 = pi2331 & ~w29897;
assign w31830 = pi3508 & w29897;
assign w31831 = ~w31829 & ~w31830;
assign w31832 = pi2332 & ~w29897;
assign w31833 = pi3509 & w29897;
assign w31834 = ~w31832 & ~w31833;
assign w31835 = pi2333 & ~w29897;
assign w31836 = pi3521 & w29897;
assign w31837 = ~w31835 & ~w31836;
assign w31838 = pi2334 & ~w29897;
assign w31839 = pi3510 & w29897;
assign w31840 = ~w31838 & ~w31839;
assign w31841 = ~pi2408 & w29897;
assign w31842 = pi2335 & ~w29897;
assign w31843 = ~w31841 & ~w31842;
assign w31844 = pi2336 & ~w29579;
assign w31845 = pi3520 & w29579;
assign w31846 = ~w31844 & ~w31845;
assign w31847 = pi2337 & ~w29579;
assign w31848 = pi3398 & w29579;
assign w31849 = ~w31847 & ~w31848;
assign w31850 = ~pi2514 & w29579;
assign w31851 = pi2338 & ~w29579;
assign w31852 = ~w31850 & ~w31851;
assign w31853 = pi2339 & ~w29579;
assign w31854 = pi3512 & w29579;
assign w31855 = ~w31853 & ~w31854;
assign w31856 = ~pi2400 & w29579;
assign w31857 = pi2340 & ~w29579;
assign w31858 = ~w31856 & ~w31857;
assign w31859 = pi2341 & ~w29579;
assign w31860 = pi3513 & w29579;
assign w31861 = ~w31859 & ~w31860;
assign w31862 = pi2342 & ~w29579;
assign w31863 = pi3504 & w29579;
assign w31864 = ~w31862 & ~w31863;
assign w31865 = pi2343 & ~w29579;
assign w31866 = pi3514 & w29579;
assign w31867 = ~w31865 & ~w31866;
assign w31868 = pi2344 & ~w29579;
assign w31869 = pi3518 & w29579;
assign w31870 = ~w31868 & ~w31869;
assign w31871 = pi2345 & ~w29579;
assign w31872 = pi3516 & w29579;
assign w31873 = ~w31871 & ~w31872;
assign w31874 = pi2346 & ~w29579;
assign w31875 = pi3517 & w29579;
assign w31876 = ~w31874 & ~w31875;
assign w31877 = pi2347 & ~w29579;
assign w31878 = pi3508 & w29579;
assign w31879 = ~w31877 & ~w31878;
assign w31880 = pi2348 & ~w29579;
assign w31881 = pi3509 & w29579;
assign w31882 = ~w31880 & ~w31881;
assign w31883 = pi2349 & ~w29579;
assign w31884 = pi3521 & w29579;
assign w31885 = ~w31883 & ~w31884;
assign w31886 = pi2350 & ~w29579;
assign w31887 = pi3510 & w29579;
assign w31888 = ~w31886 & ~w31887;
assign w31889 = pi2351 & ~w29901;
assign w31890 = pi3520 & w29901;
assign w31891 = ~w31889 & ~w31890;
assign w31892 = pi2352 & ~w29901;
assign w31893 = pi3398 & w29901;
assign w31894 = ~w31892 & ~w31893;
assign w31895 = ~pi2472 & w29901;
assign w31896 = pi2353 & ~w29901;
assign w31897 = ~w31895 & ~w31896;
assign w31898 = ~pi2400 & w29901;
assign w31899 = pi2354 & ~w29901;
assign w31900 = ~w31898 & ~w31899;
assign w31901 = pi2355 & ~w29901;
assign w31902 = pi3504 & w29901;
assign w31903 = ~w31901 & ~w31902;
assign w31904 = pi2356 & ~w29901;
assign w31905 = pi3518 & w29901;
assign w31906 = ~w31904 & ~w31905;
assign w31907 = pi2357 & ~w29901;
assign w31908 = pi3508 & w29901;
assign w31909 = ~w31907 & ~w31908;
assign w31910 = ~pi2408 & w29901;
assign w31911 = pi2358 & ~w29901;
assign w31912 = ~w31910 & ~w31911;
assign w31913 = pi2359 & ~w30678;
assign w31914 = pi3520 & w30678;
assign w31915 = ~w31913 & ~w31914;
assign w31916 = pi2360 & ~w30678;
assign w31917 = pi3398 & w30678;
assign w31918 = ~w31916 & ~w31917;
assign w31919 = pi2361 & ~w30678;
assign w31920 = pi3392 & w30678;
assign w31921 = ~w31919 & ~w31920;
assign w31922 = ~pi2514 & w30678;
assign w31923 = pi2362 & ~w30678;
assign w31924 = ~w31922 & ~w31923;
assign w31925 = pi2363 & ~w30678;
assign w31926 = pi3512 & w30678;
assign w31927 = ~w31925 & ~w31926;
assign w31928 = ~pi2400 & w30678;
assign w31929 = pi2364 & ~w30678;
assign w31930 = ~w31928 & ~w31929;
assign w31931 = pi2365 & ~w30678;
assign w31932 = pi3513 & w30678;
assign w31933 = ~w31931 & ~w31932;
assign w31934 = pi2366 & ~w30678;
assign w31935 = pi3514 & w30678;
assign w31936 = ~w31934 & ~w31935;
assign w31937 = pi2367 & ~w30678;
assign w31938 = pi3518 & w30678;
assign w31939 = ~w31937 & ~w31938;
assign w31940 = pi2368 & ~w30678;
assign w31941 = pi3517 & w30678;
assign w31942 = ~w31940 & ~w31941;
assign w31943 = pi2369 & ~w30678;
assign w31944 = pi3508 & w30678;
assign w31945 = ~w31943 & ~w31944;
assign w31946 = pi2370 & ~w30678;
assign w31947 = pi3509 & w30678;
assign w31948 = ~w31946 & ~w31947;
assign w31949 = pi2371 & ~w30678;
assign w31950 = pi3521 & w30678;
assign w31951 = ~w31949 & ~w31950;
assign w31952 = pi2372 & ~w30678;
assign w31953 = pi3510 & w30678;
assign w31954 = ~w31952 & ~w31953;
assign w31955 = ~pi2373 & w342;
assign w31956 = w422 & w8826;
assign w31957 = w6538 & ~w31956;
assign w31958 = w382 & ~w31957;
assign w31959 = pi0406 & w29980;
assign w31960 = ~w342 & ~w31959;
assign w31961 = ~w31958 & w31960;
assign w31962 = ~w31955 & ~w31961;
assign w31963 = ~pi2374 & w342;
assign w31964 = w422 & ~w8802;
assign w31965 = w2863 & ~w31964;
assign w31966 = w382 & ~w31965;
assign w31967 = pi0426 & w29980;
assign w31968 = ~w342 & ~w31967;
assign w31969 = ~w31966 & w31968;
assign w31970 = ~w31963 & ~w31969;
assign w31971 = ~pi2375 & w342;
assign w31972 = w382 & ~w22216;
assign w31973 = pi0421 & w29980;
assign w31974 = ~w342 & ~w31973;
assign w31975 = ~w31972 & w31974;
assign w31976 = ~w31971 & ~w31975;
assign w31977 = ~pi2376 & w342;
assign w31978 = w422 & ~w22222;
assign w31979 = w883 & ~w31978;
assign w31980 = w382 & ~w31979;
assign w31981 = pi0405 & w29980;
assign w31982 = ~w342 & ~w31981;
assign w31983 = ~w31980 & w31982;
assign w31984 = ~w31977 & ~w31983;
assign w31985 = ~pi2377 & w342;
assign w31986 = w422 & w24462;
assign w31987 = w5650 & ~w31986;
assign w31988 = w382 & ~w31987;
assign w31989 = pi0422 & w29980;
assign w31990 = ~w342 & ~w31989;
assign w31991 = ~w31988 & w31990;
assign w31992 = ~w31985 & ~w31991;
assign w31993 = ~pi2378 & w342;
assign w31994 = w422 & ~w24479;
assign w31995 = w4826 & ~w31994;
assign w31996 = w382 & ~w31995;
assign w31997 = pi0423 & w29980;
assign w31998 = ~w342 & ~w31997;
assign w31999 = ~w31996 & w31998;
assign w32000 = ~w31993 & ~w31999;
assign w32001 = w10564 & w28486;
assign w32002 = ~pi2379 & ~w32001;
assign w32003 = pi2380 & w27073;
assign w32004 = ~w17569 & ~w27342;
assign w32005 = w10687 & w32004;
assign w32006 = ~w32003 & ~w32005;
assign w32007 = ~pi3213 & ~pi3328;
assign w32008 = pi2777 & ~w6682;
assign w32009 = pi2381 & ~pi3375;
assign w32010 = pi3328 & ~w32009;
assign w32011 = ~pi3213 & ~pi3541;
assign w32012 = ~w32010 & ~w32011;
assign w32013 = pi2974 & ~w32012;
assign w32014 = ~w32008 & w32013;
assign w32015 = ~w32007 & ~w32014;
assign w32016 = pi2382 & w6684;
assign w32017 = w6682 & ~w21496;
assign w32018 = ~w32016 & ~w32017;
assign w32019 = ~pi2383 & w6684;
assign w32020 = w2231 & w21969;
assign w32021 = w22006 & w32020;
assign w32022 = pi0414 & w32021;
assign w32023 = ~w32019 & ~w32022;
assign w32024 = pi2384 & w6684;
assign w32025 = ~w22020 & ~w32024;
assign w32026 = ~pi3425 & pi3677;
assign w32027 = w24168 & w32026;
assign w32028 = w24215 & w32027;
assign w32029 = pi2385 & ~w32028;
assign w32030 = pi0853 & w32028;
assign w32031 = ~w32029 & ~w32030;
assign w32032 = ~pi1835 & w10;
assign w32033 = ~pi1836 & pi2507;
assign w32034 = pi1836 & ~pi2507;
assign w32035 = ~w32033 & ~w32034;
assign w32036 = ~pi1828 & pi2771;
assign w32037 = pi1828 & ~pi2771;
assign w32038 = ~w32036 & ~w32037;
assign w32039 = ~pi1792 & pi2770;
assign w32040 = pi1792 & ~pi2770;
assign w32041 = ~w32039 & ~w32040;
assign w32042 = ~w32038 & ~w32041;
assign w32043 = ~w32035 & w32042;
assign w32044 = ~pi1837 & ~pi2772;
assign w32045 = ~pi1705 & ~pi2506;
assign w32046 = pi1705 & pi2506;
assign w32047 = ~w32045 & ~w32046;
assign w32048 = ~w32044 & w32047;
assign w32049 = pi1838 & pi2760;
assign w32050 = pi1829 & pi2523;
assign w32051 = ~w32049 & ~w32050;
assign w32052 = ~pi1838 & ~pi2760;
assign w32053 = pi1837 & pi2772;
assign w32054 = ~w32052 & ~w32053;
assign w32055 = w32051 & w32054;
assign w32056 = w32048 & w32055;
assign w32057 = w32043 & w32056;
assign w32058 = ~pi1829 & ~pi2523;
assign w32059 = w32057 & ~w32058;
assign w32060 = ~pi2386 & w32059;
assign w32061 = pi2386 & ~w32059;
assign w32062 = ~w32060 & ~w32061;
assign w32063 = pi2388 & ~w29901;
assign w32064 = pi3510 & w29901;
assign w32065 = ~w32063 & ~w32064;
assign w32066 = pi2389 & ~w30678;
assign w32067 = pi3511 & w30678;
assign w32068 = ~w32066 & ~w32067;
assign w32069 = pi2390 & ~w29901;
assign w32070 = pi3519 & w29901;
assign w32071 = ~w32069 & ~w32070;
assign w32072 = pi2391 & ~w29901;
assign w32073 = pi3513 & w29901;
assign w32074 = ~w32072 & ~w32073;
assign w32075 = ~pi2392 & w342;
assign w32076 = w422 & w23420;
assign w32077 = w3878 & ~w32076;
assign w32078 = w382 & ~w32077;
assign w32079 = pi0424 & w29980;
assign w32080 = ~w342 & ~w32079;
assign w32081 = ~w32078 & w32080;
assign w32082 = ~w32075 & ~w32081;
assign w32083 = ~w6413 & w30202;
assign w32084 = pi2393 & ~w30202;
assign w32085 = ~w32083 & ~w32084;
assign w32086 = ~w8081 & w30202;
assign w32087 = pi2394 & ~w30202;
assign w32088 = ~w32086 & ~w32087;
assign w32089 = ~w5053 & w30202;
assign w32090 = pi2395 & ~w30202;
assign w32091 = ~w32089 & ~w32090;
assign w32092 = ~w4749 & w30202;
assign w32093 = pi2396 & ~w30202;
assign w32094 = ~w32092 & ~w32093;
assign w32095 = ~w5320 & w30202;
assign w32096 = pi2397 & ~w30202;
assign w32097 = ~w32095 & ~w32096;
assign w32098 = ~w3195 & w30202;
assign w32099 = pi2398 & ~w30202;
assign w32100 = ~w32098 & ~w32099;
assign w32101 = ~pi0944 & w6668;
assign w32102 = ~w4749 & w32101;
assign w32103 = ~w5914 & w32101;
assign w32104 = ~w3711 & w32101;
assign w32105 = ~w32103 & ~w32104;
assign w32106 = ~w5320 & w32101;
assign w32107 = ~pi2400 & ~w32106;
assign w32108 = w32105 & w32107;
assign w32109 = ~w32102 & ~w32108;
assign w32110 = ~pi3212 & ~pi3361;
assign w32111 = ~pi3212 & ~pi3543;
assign w32112 = pi3189 & ~w32111;
assign w32113 = ~pi1931 & ~w32112;
assign w32114 = pi2401 & ~w32113;
assign w32115 = pi3361 & ~w32114;
assign w32116 = w22068 & w32115;
assign w32117 = ~w32110 & ~w32116;
assign w32118 = pi3269 & ~w6682;
assign w32119 = ~pi3442 & ~pi3537;
assign w32120 = ~pi2100 & pi2402;
assign w32121 = ~w32119 & w32120;
assign w32122 = ~w32118 & ~w32121;
assign w32123 = ~pi3232 & ~pi3360;
assign w32124 = ~pi3232 & ~pi3542;
assign w32125 = pi3226 & ~w32124;
assign w32126 = ~pi1931 & ~w32125;
assign w32127 = pi2403 & ~w32126;
assign w32128 = pi3360 & ~w32127;
assign w32129 = w22284 & w32128;
assign w32130 = ~w32123 & ~w32129;
assign w32131 = ~w6413 & w32101;
assign w32132 = ~w3195 & w32101;
assign w32133 = ~w40134 & w32101;
assign w32134 = ~w32132 & ~w32133;
assign w32135 = ~w4380 & w32101;
assign w32136 = ~pi2404 & ~w32135;
assign w32137 = w32134 & w32136;
assign w32138 = ~w32131 & ~w32137;
assign w32139 = ~pi2405 & ~w32131;
assign w32140 = w32134 & w32139;
assign w32141 = ~w32135 & ~w32140;
assign w32142 = ~pi2472 & w29579;
assign w32143 = pi2406 & ~w29579;
assign w32144 = ~w32142 & ~w32143;
assign w32145 = ~pi2472 & w30678;
assign w32146 = pi2407 & ~w30678;
assign w32147 = ~w32145 & ~w32146;
assign w32148 = ~w32102 & ~w32106;
assign w32149 = ~pi2408 & ~w32103;
assign w32150 = w32148 & w32149;
assign w32151 = ~w32104 & ~w32150;
assign w32152 = ~w32131 & ~w32135;
assign w32153 = ~pi2409 & ~w32133;
assign w32154 = w32152 & w32153;
assign w32155 = ~w32132 & ~w32154;
assign w32156 = ~w2875 & w23731;
assign w32157 = ~w23733 & ~w32156;
assign w32158 = ~w2875 & ~w24020;
assign w32159 = ~w5941 & ~w32158;
assign w32160 = ~w2875 & w23682;
assign w32161 = ~w6475 & ~w32160;
assign w32162 = ~w2875 & w23938;
assign w32163 = ~w3853 & ~w32162;
assign w32164 = pi2414 & ~w30421;
assign w32165 = pi3691 & w30421;
assign w32166 = ~w32164 & ~w32165;
assign w32167 = ~w357 & ~w370;
assign w32168 = pi2415 & ~w32167;
assign w32169 = ~pi1029 & ~pi3245;
assign w32170 = ~pi2796 & pi3245;
assign w32171 = ~w32169 & ~w32170;
assign w32172 = w32167 & w32171;
assign w32173 = ~w32168 & ~w32172;
assign w32174 = pi2416 & ~w27275;
assign w32175 = ~w27276 & ~w32174;
assign w32176 = ~pi2417 & w343;
assign w32177 = ~w26817 & ~w32176;
assign w32178 = pi2418 & ~w30421;
assign w32179 = pi3692 & w30421;
assign w32180 = ~w32178 & ~w32179;
assign w32181 = pi3256 & w31163;
assign w32182 = pi2419 & ~w28747;
assign w32183 = ~w29835 & w32182;
assign w32184 = ~w32181 & ~w32183;
assign w32185 = w17601 & ~w30455;
assign w32186 = ~pi2420 & ~w17601;
assign w32187 = ~w32185 & ~w32186;
assign w32188 = w17601 & ~w30463;
assign w32189 = ~pi2421 & ~w17601;
assign w32190 = ~w32188 & ~w32189;
assign w32191 = w17601 & ~w30471;
assign w32192 = ~pi2422 & ~w17601;
assign w32193 = ~w32191 & ~w32192;
assign w32194 = w17601 & ~w30479;
assign w32195 = ~pi2423 & ~w17601;
assign w32196 = ~w32194 & ~w32195;
assign w32197 = w17601 & ~w30487;
assign w32198 = ~pi2424 & ~w17601;
assign w32199 = ~w32197 & ~w32198;
assign w32200 = w17601 & ~w30495;
assign w32201 = ~pi2425 & ~w17601;
assign w32202 = ~w32200 & ~w32201;
assign w32203 = w17601 & ~w30503;
assign w32204 = ~pi2426 & ~w17601;
assign w32205 = ~w32203 & ~w32204;
assign w32206 = w17601 & ~w30511;
assign w32207 = ~pi2427 & ~w17601;
assign w32208 = ~w32206 & ~w32207;
assign w32209 = w17601 & ~w30519;
assign w32210 = ~pi2428 & ~w17601;
assign w32211 = ~w32209 & ~w32210;
assign w32212 = w17601 & ~w30527;
assign w32213 = ~pi2429 & ~w17601;
assign w32214 = ~w32212 & ~w32213;
assign w32215 = w17601 & ~w30535;
assign w32216 = ~pi2430 & ~w17601;
assign w32217 = ~w32215 & ~w32216;
assign w32218 = w17601 & ~w30551;
assign w32219 = ~pi2431 & ~w17601;
assign w32220 = ~w32218 & ~w32219;
assign w32221 = ~w23216 & w23437;
assign w32222 = ~w23443 & ~w32221;
assign w32223 = ~w8667 & ~w23216;
assign w32224 = ~w23486 & ~w32223;
assign w32225 = ~w23216 & ~w23496;
assign w32226 = ~w23503 & ~w32225;
assign w32227 = w22214 & ~w23216;
assign w32228 = ~w23512 & ~w32227;
assign w32229 = ~w22222 & ~w23216;
assign w32230 = pi2436 & w23216;
assign w32231 = ~w32229 & ~w32230;
assign w32232 = w8560 & ~w23216;
assign w32233 = ~w23526 & ~w32232;
assign w32234 = w844 & ~w8826;
assign w32235 = ~pi2438 & ~w844;
assign w32236 = ~w32234 & ~w32235;
assign w32237 = w844 & ~w24445;
assign w32238 = ~pi2439 & ~w844;
assign w32239 = ~w32237 & ~w32238;
assign w32240 = w844 & w24462;
assign w32241 = ~w24466 & ~w32240;
assign w32242 = pi2441 & ~w844;
assign w32243 = w844 & ~w24479;
assign w32244 = ~w32242 & ~w32243;
assign w32245 = w856 & w23437;
assign w32246 = ~w23439 & ~w32245;
assign w32247 = w856 & w8699;
assign w32248 = ~w23467 & ~w32247;
assign w32249 = pi2444 & ~w856;
assign w32250 = w856 & ~w23496;
assign w32251 = ~w32249 & ~w32250;
assign w32252 = w856 & ~w22214;
assign w32253 = ~pi2445 & ~w856;
assign w32254 = ~w32252 & ~w32253;
assign w32255 = pi2446 & ~w856;
assign w32256 = w856 & ~w22222;
assign w32257 = ~w32255 & ~w32256;
assign w32258 = w856 & ~w8560;
assign w32259 = ~pi2447 & ~w856;
assign w32260 = ~w32258 & ~w32259;
assign w32261 = pi2448 & ~w32167;
assign w32262 = ~pi1028 & ~pi3245;
assign w32263 = ~pi2794 & pi3245;
assign w32264 = ~w32262 & ~w32263;
assign w32265 = w32167 & w32264;
assign w32266 = ~w32261 & ~w32265;
assign w32267 = pi2449 & ~w32167;
assign w32268 = ~pi1030 & ~pi3245;
assign w32269 = ~pi2644 & pi3245;
assign w32270 = ~w32268 & ~w32269;
assign w32271 = w32167 & w32270;
assign w32272 = ~w32267 & ~w32271;
assign w32273 = pi2450 & ~w32167;
assign w32274 = ~pi1031 & ~pi3245;
assign w32275 = ~pi2797 & pi3245;
assign w32276 = ~w32274 & ~w32275;
assign w32277 = w32167 & w32276;
assign w32278 = ~w32273 & ~w32277;
assign w32279 = pi2451 & ~w32167;
assign w32280 = ~pi1013 & ~pi3245;
assign w32281 = ~pi2645 & pi3245;
assign w32282 = ~w32280 & ~w32281;
assign w32283 = w32167 & w32282;
assign w32284 = ~w32279 & ~w32283;
assign w32285 = w2294 & w23938;
assign w32286 = ~w3855 & ~w32285;
assign w32287 = w2294 & w23954;
assign w32288 = ~w2930 & ~w32287;
assign w32289 = w2294 & w23971;
assign w32290 = ~w2883 & ~w32289;
assign w32291 = w2294 & w23988;
assign w32292 = ~w3903 & ~w32291;
assign w32293 = w2294 & w24004;
assign w32294 = ~w5353 & ~w32293;
assign w32295 = w2294 & w23714;
assign w32296 = ~w4474 & ~w32295;
assign w32297 = w2294 & w23731;
assign w32298 = ~w3724 & ~w32297;
assign w32299 = w2294 & ~w23763;
assign w32300 = ~w5663 & ~w32299;
assign w32301 = w2294 & ~w23779;
assign w32302 = ~w4839 & ~w32301;
assign w32303 = ~w2875 & w23954;
assign w32304 = ~w23956 & ~w32303;
assign w32305 = ~w2875 & w23971;
assign w32306 = ~w23973 & ~w32305;
assign w32307 = ~w2875 & w23698;
assign w32308 = ~w6423 & ~w32307;
assign w32309 = ~w2875 & w23988;
assign w32310 = ~w3901 & ~w32309;
assign w32311 = ~w2875 & w24004;
assign w32312 = ~w5351 & ~w32311;
assign w32313 = ~w2875 & w23714;
assign w32314 = pi2466 & w2875;
assign w32315 = ~w32313 & ~w32314;
assign w32316 = ~w2875 & ~w23748;
assign w32317 = ~w4759 & ~w32316;
assign w32318 = ~w2875 & ~w23763;
assign w32319 = ~w5661 & ~w32318;
assign w32320 = ~w2875 & ~w23779;
assign w32321 = ~w4837 & ~w32320;
assign w32322 = ~w2875 & w24037;
assign w32323 = ~w3763 & ~w32322;
assign w32324 = pi2471 & ~w30678;
assign w32325 = ~pi2408 & w30678;
assign w32326 = ~w32324 & ~w32325;
assign w32327 = ~pi2472 & ~w32102;
assign w32328 = w32105 & w32327;
assign w32329 = ~w32106 & ~w32328;
assign w32330 = ~pi2473 & ~w32132;
assign w32331 = w32152 & w32330;
assign w32332 = ~w32133 & ~w32331;
assign w32333 = pi2474 & ~w23792;
assign w32334 = w23798 & w23799;
assign w32335 = w27127 & w32334;
assign w32336 = ~w32333 & ~w32335;
assign w32337 = pi3432 & ~w19954;
assign w32338 = pi2475 & w19954;
assign w32339 = ~w32337 & ~w32338;
assign w32340 = pi3453 & ~w19954;
assign w32341 = pi2476 & w19954;
assign w32342 = ~w32340 & ~w32341;
assign w32343 = pi3454 & ~w19954;
assign w32344 = pi2477 & w19954;
assign w32345 = ~w32343 & ~w32344;
assign w32346 = pi3455 & ~w19954;
assign w32347 = pi2478 & w19954;
assign w32348 = ~w32346 & ~w32347;
assign w32349 = pi3434 & ~w19954;
assign w32350 = pi2479 & w19954;
assign w32351 = ~w32349 & ~w32350;
assign w32352 = pi3456 & ~w19954;
assign w32353 = pi2480 & w19954;
assign w32354 = ~w32352 & ~w32353;
assign w32355 = pi3457 & ~w19954;
assign w32356 = pi2481 & w19954;
assign w32357 = ~w32355 & ~w32356;
assign w32358 = pi3433 & ~w19954;
assign w32359 = pi2482 & w19954;
assign w32360 = ~w32358 & ~w32359;
assign w32361 = pi3437 & ~w19954;
assign w32362 = pi2483 & w19954;
assign w32363 = ~w32361 & ~w32362;
assign w32364 = pi3458 & ~w19954;
assign w32365 = pi2484 & w19954;
assign w32366 = ~w32364 & ~w32365;
assign w32367 = pi3450 & ~w19954;
assign w32368 = pi2485 & w19954;
assign w32369 = ~w32367 & ~w32368;
assign w32370 = ~pi2486 & w6684;
assign w32371 = ~pi0405 & w2374;
assign w32372 = w21968 & w32371;
assign w32373 = ~w32370 & ~w32372;
assign w32374 = ~pi2487 & w6684;
assign w32375 = ~w32021 & ~w32374;
assign w32376 = pi2488 & w6684;
assign w32377 = w6682 & w21620;
assign w32378 = ~w32376 & ~w32377;
assign w32379 = w6975 & w21969;
assign w32380 = w21969 & ~w29981;
assign w32381 = pi2489 & w6684;
assign w32382 = ~w32380 & ~w32381;
assign w32383 = ~w32379 & w32382;
assign w32384 = ~pi0408 & w32379;
assign w32385 = pi2490 & w6684;
assign w32386 = ~w32380 & ~w32385;
assign w32387 = ~w32384 & w32386;
assign w32388 = ~pi2491 & w6684;
assign w32389 = ~pi0408 & w381;
assign w32390 = w32380 & ~w32389;
assign w32391 = ~w32388 & ~w32390;
assign w32392 = ~pi3337 & ~pi3389;
assign w32393 = pi3568 & w32392;
assign w32394 = ~pi3417 & ~w25373;
assign w32395 = w10741 & ~w32394;
assign w32396 = w32393 & w32395;
assign w32397 = pi3398 & w6692;
assign w32398 = w6676 & w32397;
assign w32399 = pi2492 & pi3481;
assign w32400 = ~w32398 & ~w32399;
assign w32401 = w1274 & w24374;
assign w32402 = pi2493 & ~w32401;
assign w32403 = w4141 & w32401;
assign w32404 = ~w32402 & ~w32403;
assign w32405 = pi2494 & ~w32401;
assign w32406 = w6177 & w32401;
assign w32407 = ~w32405 & ~w32406;
assign w32408 = pi2495 & ~w32401;
assign w32409 = w3195 & w32401;
assign w32410 = ~w32408 & ~w32409;
assign w32411 = pi2496 & ~w32401;
assign w32412 = w40134 & w32401;
assign w32413 = ~w32411 & ~w32412;
assign w32414 = pi2497 & ~w32401;
assign w32415 = w6413 & w32401;
assign w32416 = ~w32414 & ~w32415;
assign w32417 = pi2498 & ~w32401;
assign w32418 = w5320 & w32401;
assign w32419 = ~w32417 & ~w32418;
assign w32420 = pi2499 & ~w32401;
assign w32421 = w4749 & w32401;
assign w32422 = ~w32420 & ~w32421;
assign w32423 = pi2500 & ~w32401;
assign w32424 = w5635 & w32401;
assign w32425 = ~w32423 & ~w32424;
assign w32426 = pi2501 & ~w32401;
assign w32427 = w5053 & w32401;
assign w32428 = ~w32426 & ~w32427;
assign w32429 = pi2502 & ~w32401;
assign w32430 = w3711 & w32401;
assign w32431 = ~w32429 & ~w32430;
assign w32432 = w1215 & w24374;
assign w32433 = ~pi2503 & ~w32432;
assign w32434 = ~w3195 & ~w40134;
assign w32435 = ~w4380 & w32434;
assign w32436 = ~w6413 & w32435;
assign w32437 = ~w3195 & w32432;
assign w32438 = ~w32436 & w32437;
assign w32439 = ~w32433 & ~w32438;
assign w32440 = ~pi2504 & ~w32432;
assign w32441 = ~w40134 & w32432;
assign w32442 = ~w32436 & w32441;
assign w32443 = ~w32440 & ~w32442;
assign w32444 = ~pi2505 & ~w32432;
assign w32445 = ~w4380 & w32432;
assign w32446 = ~w32436 & w32445;
assign w32447 = ~w32444 & ~w32446;
assign w32448 = ~pi2523 & ~pi2771;
assign w32449 = pi2506 & ~w32448;
assign w32450 = ~pi2506 & w32448;
assign w32451 = ~w32449 & ~w32450;
assign w32452 = ~w32059 & w32451;
assign w32453 = ~pi2760 & w32450;
assign w32454 = ~pi2772 & w32453;
assign w32455 = pi2507 & ~w32454;
assign w32456 = ~pi2507 & w32454;
assign w32457 = ~w32455 & ~w32456;
assign w32458 = ~w32059 & w32457;
assign w32459 = ~pi3247 & w27273;
assign w32460 = ~pi2824 & w32459;
assign w32461 = pi2510 & ~w32460;
assign w32462 = ~w27274 & ~w32461;
assign w32463 = w17601 & ~w30543;
assign w32464 = ~pi2511 & ~w17601;
assign w32465 = ~w32463 & ~w32464;
assign w32466 = pi2512 & ~w32401;
assign w32467 = w5914 & w32401;
assign w32468 = ~w32466 & ~w32467;
assign w32469 = pi2513 & ~w32401;
assign w32470 = w4380 & w32401;
assign w32471 = ~w32469 & ~w32470;
assign w32472 = ~pi2514 & ~w32104;
assign w32473 = w32148 & w32472;
assign w32474 = ~w32103 & ~w32473;
assign w32475 = pi2515 & ~w19038;
assign w32476 = ~w29771 & ~w32475;
assign w32477 = pi3460 & ~w19954;
assign w32478 = pi2516 & w19954;
assign w32479 = ~w32477 & ~w32478;
assign w32480 = pi3459 & ~w19954;
assign w32481 = pi2517 & w19954;
assign w32482 = ~w32480 & ~w32481;
assign w32483 = pi3478 & ~w19954;
assign w32484 = pi2518 & w19954;
assign w32485 = ~w32483 & ~w32484;
assign w32486 = pi2519 & ~w29579;
assign w32487 = ~pi2408 & w29579;
assign w32488 = ~w32486 & ~w32487;
assign w32489 = w2294 & w23682;
assign w32490 = ~w6477 & ~w32489;
assign w32491 = ~pi2522 & ~w32432;
assign w32492 = ~w6413 & w32432;
assign w32493 = ~w32435 & w32492;
assign w32494 = ~w32491 & ~w32493;
assign w32495 = pi2523 & ~w32057;
assign w32496 = w2294 & w24037;
assign w32497 = ~w3770 & ~w32496;
assign w32498 = w2294 & ~w23748;
assign w32499 = ~w4766 & ~w32498;
assign w32500 = w2294 & ~w24020;
assign w32501 = ~w5943 & ~w32500;
assign w32502 = w2294 & w23698;
assign w32503 = ~w6425 & ~w32502;
assign w32504 = w40134 & w23280;
assign w32505 = ~w23570 & ~w32504;
assign w32506 = w21489 & ~w31979;
assign w32507 = pi2529 & ~w21489;
assign w32508 = ~w32506 & ~w32507;
assign w32509 = w2323 & w23731;
assign w32510 = ~w23735 & ~w32509;
assign w32511 = w3195 & w23280;
assign w32512 = ~w23555 & ~w32511;
assign w32513 = w3711 & w23273;
assign w32514 = ~w23373 & ~w32513;
assign w32515 = w2315 & ~w23748;
assign w32516 = ~w4761 & ~w32515;
assign w32517 = w5635 & w23273;
assign w32518 = ~w23650 & ~w32517;
assign w32519 = w2315 & w23682;
assign w32520 = ~w6480 & ~w32519;
assign w32521 = w6413 & w23273;
assign w32522 = ~w23590 & ~w32521;
assign w32523 = ~pi0597 & w40144;
assign w32524 = pi2537 & ~w32523;
assign w32525 = w40171 & w32523;
assign w32526 = ~w32524 & ~w32525;
assign w32527 = pi2538 & ~w32523;
assign w32528 = w15978 & w32523;
assign w32529 = ~w32527 & ~w32528;
assign w32530 = ~w23216 & w24462;
assign w32531 = pi2539 & w23216;
assign w32532 = ~w32530 & ~w32531;
assign w32533 = w21489 & ~w30739;
assign w32534 = pi2540 & ~w21489;
assign w32535 = ~w32533 & ~w32534;
assign w32536 = pi2541 & ~w32523;
assign w32537 = w40176 & w32523;
assign w32538 = ~w32536 & ~w32537;
assign w32539 = pi2542 & ~w23262;
assign w32540 = w3711 & w23262;
assign w32541 = ~w32539 & ~w32540;
assign w32542 = pi2543 & ~w23262;
assign w32543 = w1308 & w23262;
assign w32544 = ~w32542 & ~w32543;
assign w32545 = w2323 & ~w23763;
assign w32546 = ~w23768 & ~w32545;
assign w32547 = pi2545 & ~w23262;
assign w32548 = w5635 & w23262;
assign w32549 = ~w32547 & ~w32548;
assign w32550 = w4380 & w23262;
assign w32551 = ~w23603 & ~w32550;
assign w32552 = pi2547 & ~w23262;
assign w32553 = w5914 & w23262;
assign w32554 = ~w32552 & ~w32553;
assign w32555 = w3195 & w23262;
assign w32556 = ~w23558 & ~w32555;
assign w32557 = w21489 & ~w30728;
assign w32558 = pi2549 & ~w21489;
assign w32559 = ~w32557 & ~w32558;
assign w32560 = w4141 & w22961;
assign w32561 = ~w22962 & ~w32560;
assign w32562 = w21489 & ~w30714;
assign w32563 = pi2551 & ~w21489;
assign w32564 = ~w32562 & ~w32563;
assign w32565 = w3711 & w23259;
assign w32566 = ~w23377 & ~w32565;
assign w32567 = w21489 & ~w30703;
assign w32568 = pi2553 & ~w21489;
assign w32569 = ~w32567 & ~w32568;
assign w32570 = pi2554 & ~w32167;
assign w32571 = ~pi1039 & ~pi3245;
assign w32572 = ~pi2540 & pi3245;
assign w32573 = ~w32571 & ~w32572;
assign w32574 = w32167 & w32573;
assign w32575 = ~w32570 & ~w32574;
assign w32576 = pi0955 & ~pi3250;
assign w32577 = pi2556 & ~w32167;
assign w32578 = ~pi1033 & ~pi3245;
assign w32579 = ~pi2551 & pi3245;
assign w32580 = ~w32578 & ~w32579;
assign w32581 = w32167 & w32580;
assign w32582 = ~w32577 & ~w32581;
assign w32583 = pi2557 & ~w32167;
assign w32584 = ~pi1036 & ~pi3245;
assign w32585 = ~pi2529 & pi3245;
assign w32586 = ~w32584 & ~w32585;
assign w32587 = w32167 & w32586;
assign w32588 = ~w32583 & ~w32587;
assign w32589 = pi2558 & ~w32167;
assign w32590 = ~pi1035 & ~pi3245;
assign w32591 = ~pi2647 & pi3245;
assign w32592 = ~w32590 & ~w32591;
assign w32593 = w32167 & w32592;
assign w32594 = ~w32589 & ~w32593;
assign w32595 = pi2559 & ~w32167;
assign w32596 = ~pi1012 & ~pi3245;
assign w32597 = ~pi2549 & pi3245;
assign w32598 = ~w32596 & ~w32597;
assign w32599 = w32167 & w32598;
assign w32600 = ~w32595 & ~w32599;
assign w32601 = w5914 & w23259;
assign w32602 = ~w23633 & ~w32601;
assign w32603 = w1639 & w23259;
assign w32604 = ~w23294 & ~w32603;
assign w32605 = w3711 & w22954;
assign w32606 = ~w23206 & ~w32605;
assign w32607 = w40134 & w22954;
assign w32608 = ~w23146 & ~w32607;
assign w32609 = w5635 & w23280;
assign w32610 = ~w23644 & ~w32609;
assign w32611 = w6177 & w23259;
assign w32612 = ~w23278 & ~w32611;
assign w32613 = ~pi0758 & w6668;
assign w32614 = ~pi3424 & ~w32613;
assign w32615 = w6177 & ~w32614;
assign w32616 = pi2568 & w32614;
assign w32617 = ~w32615 & ~w32616;
assign w32618 = w3195 & ~w32614;
assign w32619 = pi2569 & w32614;
assign w32620 = ~w32618 & ~w32619;
assign w32621 = w40134 & ~w32614;
assign w32622 = pi2570 & w32614;
assign w32623 = ~w32621 & ~w32622;
assign w32624 = w6413 & ~w32614;
assign w32625 = pi2571 & w32614;
assign w32626 = ~w32624 & ~w32625;
assign w32627 = w4380 & ~w32614;
assign w32628 = pi2572 & w32614;
assign w32629 = ~w32627 & ~w32628;
assign w32630 = w5320 & ~w32614;
assign w32631 = pi2573 & w32614;
assign w32632 = ~w32630 & ~w32631;
assign w32633 = w5914 & ~w32614;
assign w32634 = pi2574 & w32614;
assign w32635 = ~w32633 & ~w32634;
assign w32636 = w4749 & ~w32614;
assign w32637 = pi2575 & w32614;
assign w32638 = ~w32636 & ~w32637;
assign w32639 = w8240 & ~w32614;
assign w32640 = pi2576 & w32614;
assign w32641 = ~w32639 & ~w32640;
assign w32642 = w8081 & ~w32614;
assign w32643 = pi2577 & w32614;
assign w32644 = ~w32642 & ~w32643;
assign w32645 = w1639 & ~w32614;
assign w32646 = pi2578 & w32614;
assign w32647 = ~w32645 & ~w32646;
assign w32648 = w1308 & ~w32614;
assign w32649 = pi2579 & w32614;
assign w32650 = ~w32648 & ~w32649;
assign w32651 = w5635 & ~w32614;
assign w32652 = pi2580 & w32614;
assign w32653 = ~w32651 & ~w32652;
assign w32654 = w5053 & ~w32614;
assign w32655 = pi2581 & w32614;
assign w32656 = ~w32654 & ~w32655;
assign w32657 = w3711 & ~w32614;
assign w32658 = pi2582 & w32614;
assign w32659 = ~w32657 & ~w32658;
assign w32660 = ~pi0581 & pi3535;
assign w32661 = ~pi0982 & w6668;
assign w32662 = ~w32660 & w32661;
assign w32663 = ~w4141 & w32662;
assign w32664 = pi0478 & w32660;
assign w32665 = ~w32660 & ~w32661;
assign w32666 = ~pi2583 & w32665;
assign w32667 = ~w32664 & ~w32666;
assign w32668 = ~w32663 & w32667;
assign w32669 = ~w6177 & w32662;
assign w32670 = pi0477 & w32660;
assign w32671 = ~pi2584 & w32665;
assign w32672 = ~w32670 & ~w32671;
assign w32673 = ~w32669 & w32672;
assign w32674 = ~w3195 & w32662;
assign w32675 = pi0476 & w32660;
assign w32676 = ~pi2585 & w32665;
assign w32677 = ~w32675 & ~w32676;
assign w32678 = ~w32674 & w32677;
assign w32679 = ~w40134 & w32662;
assign w32680 = pi0475 & w32660;
assign w32681 = ~pi2586 & w32665;
assign w32682 = ~w32680 & ~w32681;
assign w32683 = ~w32679 & w32682;
assign w32684 = ~w4380 & w32662;
assign w32685 = pi0474 & w32660;
assign w32686 = ~pi2587 & w32665;
assign w32687 = ~w32685 & ~w32686;
assign w32688 = ~w32684 & w32687;
assign w32689 = ~w5320 & w32662;
assign w32690 = pi0473 & w32660;
assign w32691 = ~pi2588 & w32665;
assign w32692 = ~w32690 & ~w32691;
assign w32693 = ~w32689 & w32692;
assign w32694 = ~w5914 & w32662;
assign w32695 = pi0472 & w32660;
assign w32696 = ~pi2589 & w32665;
assign w32697 = ~w32695 & ~w32696;
assign w32698 = ~w32694 & w32697;
assign w32699 = ~w4749 & w32662;
assign w32700 = pi0697 & w32660;
assign w32701 = ~pi2590 & w32665;
assign w32702 = ~w32700 & ~w32701;
assign w32703 = ~w32699 & w32702;
assign w32704 = ~w8240 & w32662;
assign w32705 = pi0471 & w32660;
assign w32706 = ~pi2591 & w32665;
assign w32707 = ~w32705 & ~w32706;
assign w32708 = ~w32704 & w32707;
assign w32709 = ~w8081 & w32662;
assign w32710 = pi0470 & w32660;
assign w32711 = ~pi2592 & w32665;
assign w32712 = ~w32710 & ~w32711;
assign w32713 = ~w32709 & w32712;
assign w32714 = ~w1639 & w32662;
assign w32715 = pi0469 & w32660;
assign w32716 = ~pi2593 & w32665;
assign w32717 = ~w32715 & ~w32716;
assign w32718 = ~w32714 & w32717;
assign w32719 = ~w1308 & w32662;
assign w32720 = pi0468 & w32660;
assign w32721 = ~pi2594 & w32665;
assign w32722 = ~w32720 & ~w32721;
assign w32723 = ~w32719 & w32722;
assign w32724 = ~w5635 & w32662;
assign w32725 = pi0467 & w32660;
assign w32726 = ~pi2595 & w32665;
assign w32727 = ~w32725 & ~w32726;
assign w32728 = ~w32724 & w32727;
assign w32729 = ~w5053 & w32662;
assign w32730 = pi0466 & w32660;
assign w32731 = ~pi2596 & w32665;
assign w32732 = ~w32730 & ~w32731;
assign w32733 = ~w32729 & w32732;
assign w32734 = ~w3711 & w32662;
assign w32735 = pi0696 & w32660;
assign w32736 = ~pi2597 & w32665;
assign w32737 = ~w32735 & ~w32736;
assign w32738 = ~w32734 & w32737;
assign w32739 = ~pi3429 & ~pi3639;
assign w32740 = pi1738 & pi3647;
assign w32741 = ~w32665 & w32740;
assign w32742 = ~pi2598 & ~w32741;
assign w32743 = ~pi2600 & ~w30991;
assign w32744 = ~w30992 & ~w32743;
assign w32745 = ~w30987 & w32744;
assign w32746 = pi3428 & ~pi3556;
assign w32747 = pi2769 & ~w20669;
assign w32748 = w24805 & w32747;
assign w32749 = ~w19033 & w29771;
assign w32750 = ~pi2601 & ~w32749;
assign w32751 = ~w32748 & w32750;
assign w32752 = w4141 & w22954;
assign w32753 = ~w22955 & ~w32752;
assign w32754 = pi2603 & ~w22957;
assign w32755 = w3711 & w22957;
assign w32756 = ~w32754 & ~w32755;
assign w32757 = w0 & ~w32394;
assign w32758 = pi2492 & pi3441;
assign w32759 = ~pi2604 & ~w32758;
assign w32760 = ~pi0596 & w40209;
assign w32761 = ~w30452 & w32760;
assign w32762 = pi2605 & ~w32760;
assign w32763 = ~w32761 & ~w32762;
assign w32764 = ~w30460 & w32760;
assign w32765 = pi2606 & ~w32760;
assign w32766 = ~w32764 & ~w32765;
assign w32767 = ~w30524 & w32760;
assign w32768 = pi2607 & ~w32760;
assign w32769 = ~w32767 & ~w32768;
assign w32770 = ~w30532 & w32760;
assign w32771 = pi2608 & ~w32760;
assign w32772 = ~w32770 & ~w32771;
assign w32773 = ~w30540 & w32760;
assign w32774 = pi2609 & ~w32760;
assign w32775 = ~w32773 & ~w32774;
assign w32776 = ~w30548 & w32760;
assign w32777 = pi2610 & ~w32760;
assign w32778 = ~w32776 & ~w32777;
assign w32779 = ~pi0596 & w40144;
assign w32780 = ~w30452 & w32779;
assign w32781 = pi2611 & ~w32779;
assign w32782 = ~w32780 & ~w32781;
assign w32783 = ~w30460 & w32779;
assign w32784 = pi2612 & ~w32779;
assign w32785 = ~w32783 & ~w32784;
assign w32786 = ~w30524 & w32779;
assign w32787 = pi2613 & ~w32779;
assign w32788 = ~w32786 & ~w32787;
assign w32789 = ~w30532 & w32779;
assign w32790 = pi2614 & ~w32779;
assign w32791 = ~w32789 & ~w32790;
assign w32792 = pi2615 & ~w22957;
assign w32793 = w5635 & w22957;
assign w32794 = ~w32792 & ~w32793;
assign w32795 = ~w30540 & w32779;
assign w32796 = pi2616 & ~w32779;
assign w32797 = ~w32795 & ~w32796;
assign w32798 = ~w30548 & w32779;
assign w32799 = pi2617 & ~w32779;
assign w32800 = ~w32798 & ~w32799;
assign w32801 = ~pi0580 & w40209;
assign w32802 = ~w30452 & w32801;
assign w32803 = pi2618 & ~w32801;
assign w32804 = ~w32802 & ~w32803;
assign w32805 = ~w30460 & w32801;
assign w32806 = pi2619 & ~w32801;
assign w32807 = ~w32805 & ~w32806;
assign w32808 = ~w30524 & w32801;
assign w32809 = pi2620 & ~w32801;
assign w32810 = ~w32808 & ~w32809;
assign w32811 = ~w30532 & w32801;
assign w32812 = pi2621 & ~w32801;
assign w32813 = ~w32811 & ~w32812;
assign w32814 = ~w30540 & w32801;
assign w32815 = pi2622 & ~w32801;
assign w32816 = ~w32814 & ~w32815;
assign w32817 = ~w30548 & w32801;
assign w32818 = pi2623 & ~w32801;
assign w32819 = ~w32817 & ~w32818;
assign w32820 = ~pi0580 & w40144;
assign w32821 = ~w30452 & w32820;
assign w32822 = pi2624 & ~w32820;
assign w32823 = ~w32821 & ~w32822;
assign w32824 = ~w30460 & w32820;
assign w32825 = pi2625 & ~w32820;
assign w32826 = ~w32824 & ~w32825;
assign w32827 = ~w30524 & w32820;
assign w32828 = pi2626 & ~w32820;
assign w32829 = ~w32827 & ~w32828;
assign w32830 = ~w30532 & w32820;
assign w32831 = pi2627 & ~w32820;
assign w32832 = ~w32830 & ~w32831;
assign w32833 = ~w30540 & w32820;
assign w32834 = pi2628 & ~w32820;
assign w32835 = ~w32833 & ~w32834;
assign w32836 = ~w30548 & w32820;
assign w32837 = pi2629 & ~w32820;
assign w32838 = ~w32836 & ~w32837;
assign w32839 = pi2630 & ~w32523;
assign w32840 = w40189 & w32523;
assign w32841 = ~w32839 & ~w32840;
assign w32842 = pi2631 & ~w32523;
assign w32843 = w40191 & w32523;
assign w32844 = ~w32842 & ~w32843;
assign w32845 = pi2632 & ~w32523;
assign w32846 = w40174 & w32523;
assign w32847 = ~w32845 & ~w32846;
assign w32848 = pi2633 & ~w32523;
assign w32849 = w14325 & w32523;
assign w32850 = ~w32848 & ~w32849;
assign w32851 = pi2634 & ~w32523;
assign w32852 = w14962 & w32523;
assign w32853 = ~w32851 & ~w32852;
assign w32854 = pi2635 & ~w32523;
assign w32855 = w40168 & w32523;
assign w32856 = ~w32854 & ~w32855;
assign w32857 = pi2636 & ~w32523;
assign w32858 = w13916 & w32523;
assign w32859 = ~w32857 & ~w32858;
assign w32860 = pi2637 & ~w32523;
assign w32861 = w40159 & w32523;
assign w32862 = ~w32860 & ~w32861;
assign w32863 = ~w10746 & w32523;
assign w32864 = pi2638 & ~w32523;
assign w32865 = ~w32863 & ~w32864;
assign w32866 = pi2639 & ~w32523;
assign w32867 = w16629 & w32523;
assign w32868 = ~w32866 & ~w32867;
assign w32869 = pi2640 & ~w32523;
assign w32870 = w16739 & w32523;
assign w32871 = ~w32869 & ~w32870;
assign w32872 = pi2641 & ~w32523;
assign w32873 = ~w16842 & w32523;
assign w32874 = ~w32872 & ~w32873;
assign w32875 = pi2642 & ~w32523;
assign w32876 = w15171 & w32523;
assign w32877 = ~w32875 & ~w32876;
assign w32878 = w24250 & w32027;
assign w32879 = pi2643 & ~w32878;
assign w32880 = ~pi0731 & w32878;
assign w32881 = ~w32879 & ~w32880;
assign w32882 = w21489 & ~w30687;
assign w32883 = pi2644 & ~w21489;
assign w32884 = ~w32882 & ~w32883;
assign w32885 = w21489 & ~w30695;
assign w32886 = pi2645 & ~w21489;
assign w32887 = ~w32885 & ~w32886;
assign w32888 = w21489 & ~w30720;
assign w32889 = pi2646 & ~w21489;
assign w32890 = ~w32888 & ~w32889;
assign w32891 = w21489 & ~w22216;
assign w32892 = pi2647 & ~w21489;
assign w32893 = ~w32891 & ~w32892;
assign w32894 = w6177 & w22961;
assign w32895 = ~w23404 & ~w32894;
assign w32896 = w3195 & w22961;
assign w32897 = ~w23126 & ~w32896;
assign w32898 = w40134 & w22961;
assign w32899 = ~w23142 & ~w32898;
assign w32900 = w6413 & w22961;
assign w32901 = ~w24314 & ~w32900;
assign w32902 = w4380 & w22961;
assign w32903 = ~w23161 & ~w32902;
assign w32904 = w5320 & w22961;
assign w32905 = ~w23109 & ~w32904;
assign w32906 = w5914 & w22961;
assign w32907 = ~w23172 & ~w32906;
assign w32908 = w4749 & w22961;
assign w32909 = ~w23191 & ~w32908;
assign w32910 = w1639 & w22961;
assign w32911 = ~w24422 & ~w32910;
assign w32912 = w1308 & w22961;
assign w32913 = ~w22974 & ~w32912;
assign w32914 = w5635 & w22961;
assign w32915 = ~w22993 & ~w32914;
assign w32916 = w5053 & w22961;
assign w32917 = ~w24299 & ~w32916;
assign w32918 = w3711 & w22961;
assign w32919 = ~w23202 & ~w32918;
assign w32920 = w4141 & w22964;
assign w32921 = ~w22965 & ~w32920;
assign w32922 = w6177 & w22964;
assign w32923 = ~w23402 & ~w32922;
assign w32924 = w3195 & w22964;
assign w32925 = ~w23133 & ~w32924;
assign w32926 = w40134 & w22964;
assign w32927 = ~w23148 & ~w32926;
assign w32928 = w6413 & w22964;
assign w32929 = ~w24308 & ~w32928;
assign w32930 = w4380 & w22964;
assign w32931 = ~w23157 & ~w32930;
assign w32932 = w5320 & w22964;
assign w32933 = ~w23116 & ~w32932;
assign w32934 = w5914 & w22964;
assign w32935 = ~w23176 & ~w32934;
assign w32936 = w4749 & w22964;
assign w32937 = ~w23187 & ~w32936;
assign w32938 = w1639 & w22964;
assign w32939 = ~w24416 & ~w32938;
assign w32940 = w1308 & w22964;
assign w32941 = ~w22978 & ~w32940;
assign w32942 = w5635 & w22964;
assign w32943 = ~w22989 & ~w32942;
assign w32944 = w5053 & w22964;
assign w32945 = ~w24297 & ~w32944;
assign w32946 = w3711 & w22964;
assign w32947 = ~w23208 & ~w32946;
assign w32948 = pi2675 & ~w22957;
assign w32949 = w4141 & w22957;
assign w32950 = ~w32948 & ~w32949;
assign w32951 = w6177 & w22957;
assign w32952 = ~w23407 & ~w32951;
assign w32953 = w3195 & w22957;
assign w32954 = ~w23131 & ~w32953;
assign w32955 = pi2678 & ~w22957;
assign w32956 = w40134 & w22957;
assign w32957 = ~w32955 & ~w32956;
assign w32958 = pi2679 & ~w22957;
assign w32959 = w6413 & w22957;
assign w32960 = ~w32958 & ~w32959;
assign w32961 = pi2680 & ~w22957;
assign w32962 = w4380 & w22957;
assign w32963 = ~w32961 & ~w32962;
assign w32964 = w5320 & w22957;
assign w32965 = ~w23114 & ~w32964;
assign w32966 = pi2682 & ~w22957;
assign w32967 = w5914 & w22957;
assign w32968 = ~w32966 & ~w32967;
assign w32969 = pi2683 & ~w22957;
assign w32970 = w4749 & w22957;
assign w32971 = ~w32969 & ~w32970;
assign w32972 = pi2684 & ~w22957;
assign w32973 = w1639 & w22957;
assign w32974 = ~w32972 & ~w32973;
assign w32975 = pi2685 & ~w22957;
assign w32976 = w1308 & w22957;
assign w32977 = ~w32975 & ~w32976;
assign w32978 = pi2686 & ~w22957;
assign w32979 = w5053 & w22957;
assign w32980 = ~w32978 & ~w32979;
assign w32981 = w6177 & w22954;
assign w32982 = ~w23409 & ~w32981;
assign w32983 = w3195 & w22954;
assign w32984 = ~w23128 & ~w32983;
assign w32985 = w6413 & w22954;
assign w32986 = ~w24312 & ~w32985;
assign w32987 = w4380 & w22954;
assign w32988 = ~w23163 & ~w32987;
assign w32989 = w5320 & w22954;
assign w32990 = ~w23111 & ~w32989;
assign w32991 = w5914 & w22954;
assign w32992 = ~w23178 & ~w32991;
assign w32993 = w4749 & w22954;
assign w32994 = ~w23193 & ~w32993;
assign w32995 = w1639 & w22954;
assign w32996 = ~w24420 & ~w32995;
assign w32997 = w1308 & w22954;
assign w32998 = ~w22980 & ~w32997;
assign w32999 = w5635 & w22954;
assign w33000 = ~w22995 & ~w32999;
assign w33001 = w5053 & w22954;
assign w33002 = ~w24293 & ~w33001;
assign w33003 = w8826 & ~w23216;
assign w33004 = pi2698 & w23216;
assign w33005 = ~w33003 & ~w33004;
assign w33006 = ~w23216 & w24445;
assign w33007 = ~w24447 & ~w33006;
assign w33008 = ~w23216 & ~w24479;
assign w33009 = ~w24486 & ~w33008;
assign w33010 = w856 & ~w8826;
assign w33011 = ~pi2701 & ~w856;
assign w33012 = ~w33010 & ~w33011;
assign w33013 = w856 & w24445;
assign w33014 = ~w24449 & ~w33013;
assign w33015 = w856 & w24462;
assign w33016 = ~w24468 & ~w33015;
assign w33017 = pi2704 & ~w32167;
assign w33018 = ~pi1032 & ~pi3245;
assign w33019 = ~pi2553 & pi3245;
assign w33020 = ~w33018 & ~w33019;
assign w33021 = w32167 & w33020;
assign w33022 = ~w33017 & ~w33021;
assign w33023 = pi2705 & ~w32167;
assign w33024 = ~pi1034 & ~pi3245;
assign w33025 = ~pi2646 & pi3245;
assign w33026 = ~w33024 & ~w33025;
assign w33027 = w32167 & w33026;
assign w33028 = ~w33023 & ~w33027;
assign w33029 = pi2706 & ~w32167;
assign w33030 = ~pi1037 & ~pi3245;
assign w33031 = ~pi2953 & pi3245;
assign w33032 = ~w33030 & ~w33031;
assign w33033 = w32167 & w33032;
assign w33034 = ~w33029 & ~w33033;
assign w33035 = pi2707 & ~w32167;
assign w33036 = ~pi1038 & ~pi3245;
assign w33037 = ~pi2788 & pi3245;
assign w33038 = ~w33036 & ~w33037;
assign w33039 = w32167 & w33038;
assign w33040 = ~w33035 & ~w33039;
assign w33041 = w4141 & w23273;
assign w33042 = ~w23545 & ~w33041;
assign w33043 = w6177 & w23273;
assign w33044 = ~w23274 & ~w33043;
assign w33045 = w3195 & w23273;
assign w33046 = ~w23560 & ~w33045;
assign w33047 = w40134 & w23273;
assign w33048 = ~w23575 & ~w33047;
assign w33049 = w4380 & w23273;
assign w33050 = ~w23605 & ~w33049;
assign w33051 = w5320 & w23273;
assign w33052 = ~w23388 & ~w33051;
assign w33053 = w5914 & w23273;
assign w33054 = ~w23635 & ~w33053;
assign w33055 = w4749 & w23273;
assign w33056 = ~w23620 & ~w33055;
assign w33057 = w1639 & w23273;
assign w33058 = ~w23296 & ~w33057;
assign w33059 = w1308 & w23273;
assign w33060 = ~w23311 & ~w33059;
assign w33061 = w5053 & w23273;
assign w33062 = ~w23660 & ~w33061;
assign w33063 = w4141 & w23280;
assign w33064 = ~w23540 & ~w33063;
assign w33065 = w6177 & w23280;
assign w33066 = ~w23281 & ~w33065;
assign w33067 = w6413 & w23280;
assign w33068 = ~w23584 & ~w33067;
assign w33069 = w4380 & w23280;
assign w33070 = ~w23599 & ~w33069;
assign w33071 = w5320 & w23280;
assign w33072 = ~w23393 & ~w33071;
assign w33073 = w5914 & w23280;
assign w33074 = ~w23630 & ~w33073;
assign w33075 = w1308 & w23280;
assign w33076 = ~w23306 & ~w33075;
assign w33077 = w5053 & w23280;
assign w33078 = ~w23665 & ~w33077;
assign w33079 = w3711 & w23280;
assign w33080 = ~w23379 & ~w33079;
assign w33081 = w4141 & w23259;
assign w33082 = ~w23543 & ~w33081;
assign w33083 = pi2729 & ~w23259;
assign w33084 = w3195 & w23259;
assign w33085 = ~w33083 & ~w33084;
assign w33086 = w40134 & w23259;
assign w33087 = ~w23573 & ~w33086;
assign w33088 = w6413 & w23259;
assign w33089 = ~w23588 & ~w33088;
assign w33090 = pi2732 & ~w23259;
assign w33091 = w4380 & w23259;
assign w33092 = ~w33090 & ~w33091;
assign w33093 = pi2733 & ~w23259;
assign w33094 = w5320 & w23259;
assign w33095 = ~w33093 & ~w33094;
assign w33096 = w4749 & w23259;
assign w33097 = ~w23618 & ~w33096;
assign w33098 = w1308 & w23259;
assign w33099 = ~w23309 & ~w33098;
assign w33100 = w5635 & w23259;
assign w33101 = ~w23648 & ~w33100;
assign w33102 = pi2737 & ~w23259;
assign w33103 = w5053 & w23259;
assign w33104 = ~w33102 & ~w33103;
assign w33105 = pi2738 & ~w23262;
assign w33106 = w4141 & w23262;
assign w33107 = ~w33105 & ~w33106;
assign w33108 = pi2739 & ~w23262;
assign w33109 = w6177 & w23262;
assign w33110 = ~w33108 & ~w33109;
assign w33111 = pi2740 & ~w23262;
assign w33112 = w40134 & w23262;
assign w33113 = ~w33111 & ~w33112;
assign w33114 = pi2741 & ~w23262;
assign w33115 = w6413 & w23262;
assign w33116 = ~w33114 & ~w33115;
assign w33117 = pi2742 & ~w23262;
assign w33118 = w5320 & w23262;
assign w33119 = ~w33117 & ~w33118;
assign w33120 = pi2743 & ~w23262;
assign w33121 = w4749 & w23262;
assign w33122 = ~w33120 & ~w33121;
assign w33123 = pi2744 & ~w23262;
assign w33124 = w1639 & w23262;
assign w33125 = ~w33123 & ~w33124;
assign w33126 = w5053 & w23262;
assign w33127 = ~w23663 & ~w33126;
assign w33128 = w2315 & ~w23698;
assign w33129 = ~pi2746 & ~w2315;
assign w33130 = ~w33128 & ~w33129;
assign w33131 = w2315 & w23714;
assign w33132 = ~w23718 & ~w33131;
assign w33133 = w2315 & w23731;
assign w33134 = ~w3727 & ~w33133;
assign w33135 = pi2749 & ~w2315;
assign w33136 = w2315 & ~w23763;
assign w33137 = ~w33135 & ~w33136;
assign w33138 = pi2750 & ~w2315;
assign w33139 = w2315 & ~w23779;
assign w33140 = ~w33138 & ~w33139;
assign w33141 = w856 & ~w24479;
assign w33142 = ~w24481 & ~w33141;
assign w33143 = w2323 & w23682;
assign w33144 = ~w23686 & ~w33143;
assign w33145 = w2323 & w23698;
assign w33146 = ~w23702 & ~w33145;
assign w33147 = w2323 & w23714;
assign w33148 = ~w23720 & ~w33147;
assign w33149 = w2323 & ~w23748;
assign w33150 = ~w4764 & ~w33149;
assign w33151 = w2323 & ~w23779;
assign w33152 = ~w23783 & ~w33151;
assign w33153 = ~pi2757 & w6684;
assign w33154 = ~pi0419 & w21798;
assign w33155 = w21968 & w33154;
assign w33156 = ~w33153 & ~w33155;
assign w33157 = ~pi2758 & w343;
assign w33158 = ~w30567 & ~w33157;
assign w33159 = w6682 & ~w33158;
assign w33160 = ~pi2759 & ~w30857;
assign w33161 = ~w30858 & ~w33160;
assign w33162 = ~w30853 & w33161;
assign w33163 = pi2760 & ~w32450;
assign w33164 = ~w32453 & ~w33163;
assign w33165 = ~w32059 & w33164;
assign w33166 = pi2761 & ~w32878;
assign w33167 = ~pi0730 & w32878;
assign w33168 = ~w33166 & ~w33167;
assign w33169 = pi2762 & ~w32878;
assign w33170 = ~pi0938 & w32878;
assign w33171 = ~w33169 & ~w33170;
assign w33172 = pi2763 & w6684;
assign w33173 = ~w32380 & ~w33172;
assign w33174 = ~w6413 & w32662;
assign w33175 = pi0465 & w32660;
assign w33176 = ~pi2764 & w32665;
assign w33177 = ~w33175 & ~w33176;
assign w33178 = ~w33174 & w33177;
assign w33179 = ~w26523 & w26524;
assign w33180 = ~pi2766 & ~w33179;
assign w33181 = pi2767 & ~w29573;
assign w33182 = ~w29566 & ~w33181;
assign w33183 = ~w6758 & w29567;
assign w33184 = ~w33182 & ~w33183;
assign w33185 = w4141 & ~w32614;
assign w33186 = pi2768 & w32614;
assign w33187 = ~w33185 & ~w33186;
assign w33188 = pi2769 & ~w24808;
assign w33189 = ~w29781 & ~w33188;
assign w33190 = ~pi2770 & w32456;
assign w33191 = pi2770 & ~w32456;
assign w33192 = ~w32059 & ~w33191;
assign w33193 = ~w33190 & w33192;
assign w33194 = pi2523 & pi2771;
assign w33195 = ~w32448 & ~w33194;
assign w33196 = ~w32059 & w33195;
assign w33197 = pi2772 & ~w32453;
assign w33198 = ~w32454 & ~w33197;
assign w33199 = ~w32059 & w33198;
assign w33200 = w4749 & w23280;
assign w33201 = ~w23614 & ~w33200;
assign w33202 = w1639 & w23280;
assign w33203 = ~w23291 & ~w33202;
assign w33204 = w24233 & w32027;
assign w33205 = pi2775 & ~w33204;
assign w33206 = ~pi0824 & w33204;
assign w33207 = ~w33205 & ~w33206;
assign w33208 = w2315 & ~w24020;
assign w33209 = ~w24023 & ~w33208;
assign w33210 = pi2777 & ~w23792;
assign w33211 = pi2402 & w23797;
assign w33212 = w27127 & w33211;
assign w33213 = ~w33210 & ~w33212;
assign w33214 = ~pi0598 & w40144;
assign w33215 = ~w30540 & w33214;
assign w33216 = pi2778 & ~w33214;
assign w33217 = ~w33215 & ~w33216;
assign w33218 = w21821 & w22169;
assign w33219 = pi2779 & w343;
assign w33220 = ~w33218 & ~w33219;
assign w33221 = w2315 & ~w24004;
assign w33222 = ~pi2780 & ~w2315;
assign w33223 = ~w33221 & ~w33222;
assign w33224 = ~w29844 & w32779;
assign w33225 = pi2781 & ~w32779;
assign w33226 = ~w33224 & ~w33225;
assign w33227 = ~w30492 & w32779;
assign w33228 = pi2782 & ~w32779;
assign w33229 = ~w33227 & ~w33228;
assign w33230 = ~pi0575 & w40144;
assign w33231 = pi2783 & ~w33230;
assign w33232 = w40159 & w33230;
assign w33233 = ~w33231 & ~w33232;
assign w33234 = pi2784 & ~w33230;
assign w33235 = w40174 & w33230;
assign w33236 = ~w33234 & ~w33235;
assign w33237 = ~pi3146 & w31162;
assign w33238 = pi2785 & ~w28758;
assign w33239 = ~w28747 & w33238;
assign w33240 = ~w33237 & ~w33239;
assign w33241 = w24210 & w32027;
assign w33242 = pi2786 & ~w33241;
assign w33243 = ~pi0858 & w33241;
assign w33244 = ~w33242 & ~w33243;
assign w33245 = ~w30484 & w33214;
assign w33246 = pi2787 & ~w33214;
assign w33247 = ~w33245 & ~w33246;
assign w33248 = w21489 & ~w31995;
assign w33249 = pi2788 & ~w21489;
assign w33250 = ~w33248 & ~w33249;
assign w33251 = pi2789 & w343;
assign w33252 = w2230 & w22856;
assign w33253 = ~w33251 & ~w33252;
assign w33254 = w24196 & w32027;
assign w33255 = pi2790 & ~w33254;
assign w33256 = ~pi0851 & w33254;
assign w33257 = ~w33255 & ~w33256;
assign w33258 = w24236 & w32027;
assign w33259 = pi2791 & ~w33258;
assign w33260 = ~pi0938 & w33258;
assign w33261 = ~w33259 & ~w33260;
assign w33262 = w24217 & w32027;
assign w33263 = pi2792 & ~w33262;
assign w33264 = ~pi0823 & w33262;
assign w33265 = ~w33263 & ~w33264;
assign w33266 = ~pi0649 & w40144;
assign w33267 = pi2793 & ~w33266;
assign w33268 = w40176 & w33266;
assign w33269 = ~w33267 & ~w33268;
assign w33270 = w21489 & ~w32077;
assign w33271 = pi2794 & ~w21489;
assign w33272 = ~w33270 & ~w33271;
assign w33273 = pi2795 & w343;
assign w33274 = w21489 & ~w31957;
assign w33275 = pi2796 & ~w21489;
assign w33276 = ~w33274 & ~w33275;
assign w33277 = w21489 & ~w31965;
assign w33278 = pi2797 & ~w21489;
assign w33279 = ~w33277 & ~w33278;
assign w33280 = ~pi2798 & w30988;
assign w33281 = ~w30989 & ~w33280;
assign w33282 = ~w30987 & w33281;
assign w33283 = ~pi2799 & ~w30990;
assign w33284 = ~w30991 & ~w33283;
assign w33285 = ~w30987 & w33284;
assign w33286 = ~w25373 & w27117;
assign w33287 = w20527 & w33286;
assign w33288 = pi2801 & ~w33266;
assign w33289 = w15978 & w33266;
assign w33290 = ~w33288 & ~w33289;
assign w33291 = ~pi2802 & w343;
assign w33292 = ~w21489 & ~w33291;
assign w33293 = pi2803 & ~w33266;
assign w33294 = ~w16842 & w33266;
assign w33295 = ~w33293 & ~w33294;
assign w33296 = pi2804 & ~w33266;
assign w33297 = w16629 & w33266;
assign w33298 = ~w33296 & ~w33297;
assign w33299 = ~w10746 & w33266;
assign w33300 = pi2805 & ~w33266;
assign w33301 = ~w33299 & ~w33300;
assign w33302 = pi2806 & ~w33258;
assign w33303 = ~pi0785 & w33258;
assign w33304 = ~w33302 & ~w33303;
assign w33305 = pi2807 & ~w33266;
assign w33306 = w14962 & w33266;
assign w33307 = ~w33305 & ~w33306;
assign w33308 = pi2808 & ~w33266;
assign w33309 = w14325 & w33266;
assign w33310 = ~w33308 & ~w33309;
assign w33311 = pi2809 & ~w33266;
assign w33312 = w40191 & w33266;
assign w33313 = ~w33311 & ~w33312;
assign w33314 = w2323 & w24004;
assign w33315 = ~w24008 & ~w33314;
assign w33316 = pi2811 & ~w33258;
assign w33317 = ~pi0852 & w33258;
assign w33318 = ~w33316 & ~w33317;
assign w33319 = ~w343 & ~w13981;
assign w33320 = ~pi2812 & w343;
assign w33321 = w17481 & ~w33320;
assign w33322 = ~w33319 & w33321;
assign w33323 = pi2813 & ~w6684;
assign w33324 = w88 & w110;
assign w33325 = ~w91 & ~w33324;
assign w33326 = ~w86 & w33325;
assign w33327 = pi3682 & w177;
assign w33328 = ~w113 & w33327;
assign w33329 = ~w33326 & w33328;
assign w33330 = ~w165 & w33329;
assign w33331 = ~pi3682 & w30981;
assign w33332 = w165 & w33331;
assign w33333 = ~pi2813 & ~w33332;
assign w33334 = ~w33330 & w33333;
assign w33335 = ~w33323 & ~w33334;
assign w33336 = w1257 & w24374;
assign w33337 = pi2815 & ~w33254;
assign w33338 = ~pi0824 & w33254;
assign w33339 = ~w33337 & ~w33338;
assign w33340 = ~pi2779 & ~pi3257;
assign w33341 = ~w28745 & ~w33340;
assign w33342 = w86 & w33341;
assign w33343 = ~w183 & w33342;
assign w33344 = pi2816 & ~w33343;
assign w33345 = pi3698 & w33343;
assign w33346 = ~w33344 & ~w33345;
assign w33347 = pi2817 & ~w33343;
assign w33348 = pi3696 & w33343;
assign w33349 = ~w33347 & ~w33348;
assign w33350 = pi2818 & ~w33204;
assign w33351 = ~pi0821 & w33204;
assign w33352 = ~w33350 & ~w33351;
assign w33353 = pi2819 & ~w33343;
assign w33354 = pi3689 & w33343;
assign w33355 = ~w33353 & ~w33354;
assign w33356 = ~pi0955 & w18003;
assign w33357 = ~w18366 & ~w33356;
assign w33358 = pi3635 & ~w33357;
assign w33359 = w24194 & w32027;
assign w33360 = pi2821 & ~w33359;
assign w33361 = ~pi0938 & w33359;
assign w33362 = ~w33360 & ~w33361;
assign w33363 = pi2822 & ~w33359;
assign w33364 = ~pi0851 & w33359;
assign w33365 = ~w33363 & ~w33364;
assign w33366 = pi2823 & ~w33262;
assign w33367 = ~pi0857 & w33262;
assign w33368 = ~w33366 & ~w33367;
assign w33369 = pi2824 & ~w32459;
assign w33370 = ~w32460 & ~w33369;
assign w33371 = ~pi2825 & ~w30989;
assign w33372 = ~w30990 & ~w33371;
assign w33373 = ~w30987 & w33372;
assign w33374 = pi2826 & ~w33343;
assign w33375 = pi3690 & w33343;
assign w33376 = ~w33374 & ~w33375;
assign w33377 = pi2827 & ~w33343;
assign w33378 = pi3688 & w33343;
assign w33379 = ~w33377 & ~w33378;
assign w33380 = pi2828 & ~w33343;
assign w33381 = pi3687 & w33343;
assign w33382 = ~w33380 & ~w33381;
assign w33383 = pi2829 & ~w33343;
assign w33384 = pi3686 & w33343;
assign w33385 = ~w33383 & ~w33384;
assign w33386 = pi2830 & ~w33343;
assign w33387 = pi3685 & w33343;
assign w33388 = ~w33386 & ~w33387;
assign w33389 = pi2831 & ~w33343;
assign w33390 = pi3684 & w33343;
assign w33391 = ~w33389 & ~w33390;
assign w33392 = pi2832 & ~w33343;
assign w33393 = pi3697 & w33343;
assign w33394 = ~w33392 & ~w33393;
assign w33395 = pi2833 & ~w33343;
assign w33396 = pi3695 & w33343;
assign w33397 = ~w33395 & ~w33396;
assign w33398 = pi2834 & ~w33343;
assign w33399 = pi3694 & w33343;
assign w33400 = ~w33398 & ~w33399;
assign w33401 = pi2835 & ~w33343;
assign w33402 = pi3693 & w33343;
assign w33403 = ~w33401 & ~w33402;
assign w33404 = pi2836 & ~w33343;
assign w33405 = pi3683 & w33343;
assign w33406 = ~w33404 & ~w33405;
assign w33407 = pi2837 & ~w33254;
assign w33408 = ~pi0785 & w33254;
assign w33409 = ~w33407 & ~w33408;
assign w33410 = pi2838 & ~w33359;
assign w33411 = ~pi0852 & w33359;
assign w33412 = ~w33410 & ~w33411;
assign w33413 = pi2839 & ~w33359;
assign w33414 = ~pi0860 & w33359;
assign w33415 = ~w33413 & ~w33414;
assign w33416 = ~pi0579 & w40144;
assign w33417 = pi2840 & ~w33416;
assign w33418 = w15171 & w33416;
assign w33419 = ~w33417 & ~w33418;
assign w33420 = ~pi0711 & w40144;
assign w33421 = pi2841 & ~w33420;
assign w33422 = w40189 & w33420;
assign w33423 = ~w33421 & ~w33422;
assign w33424 = pi2842 & ~w33420;
assign w33425 = w40191 & w33420;
assign w33426 = ~w33424 & ~w33425;
assign w33427 = pi2843 & ~w33420;
assign w33428 = w40174 & w33420;
assign w33429 = ~w33427 & ~w33428;
assign w33430 = pi2844 & ~w33420;
assign w33431 = w14325 & w33420;
assign w33432 = ~w33430 & ~w33431;
assign w33433 = pi2845 & ~w33420;
assign w33434 = w14962 & w33420;
assign w33435 = ~w33433 & ~w33434;
assign w33436 = pi2846 & ~w33420;
assign w33437 = w40168 & w33420;
assign w33438 = ~w33436 & ~w33437;
assign w33439 = pi2847 & ~w33420;
assign w33440 = w40176 & w33420;
assign w33441 = ~w33439 & ~w33440;
assign w33442 = pi2848 & ~w33420;
assign w33443 = w13916 & w33420;
assign w33444 = ~w33442 & ~w33443;
assign w33445 = pi2849 & ~w33420;
assign w33446 = w40159 & w33420;
assign w33447 = ~w33445 & ~w33446;
assign w33448 = ~w10746 & w33420;
assign w33449 = pi2850 & ~w33420;
assign w33450 = ~w33448 & ~w33449;
assign w33451 = pi2851 & ~w33420;
assign w33452 = w16629 & w33420;
assign w33453 = ~w33451 & ~w33452;
assign w33454 = pi2852 & ~w33420;
assign w33455 = w16739 & w33420;
assign w33456 = ~w33454 & ~w33455;
assign w33457 = pi2853 & ~w33420;
assign w33458 = ~w16842 & w33420;
assign w33459 = ~w33457 & ~w33458;
assign w33460 = pi2854 & ~w33420;
assign w33461 = w15978 & w33420;
assign w33462 = ~w33460 & ~w33461;
assign w33463 = pi2855 & ~w33420;
assign w33464 = w15171 & w33420;
assign w33465 = ~w33463 & ~w33464;
assign w33466 = pi2856 & ~w33420;
assign w33467 = w40171 & w33420;
assign w33468 = ~w33466 & ~w33467;
assign w33469 = pi2857 & ~w33359;
assign w33470 = ~pi0825 & w33359;
assign w33471 = ~w33469 & ~w33470;
assign w33472 = pi2858 & ~w33359;
assign w33473 = ~pi0854 & w33359;
assign w33474 = ~w33472 & ~w33473;
assign w33475 = w24185 & w32027;
assign w33476 = pi2859 & ~w33475;
assign w33477 = ~pi0860 & w33475;
assign w33478 = ~w33476 & ~w33477;
assign w33479 = w24624 & w32027;
assign w33480 = pi2860 & ~w33479;
assign w33481 = ~pi0855 & w33479;
assign w33482 = ~w33480 & ~w33481;
assign w33483 = ~w29852 & w32760;
assign w33484 = pi2861 & ~w32760;
assign w33485 = ~w33483 & ~w33484;
assign w33486 = ~w30468 & w32779;
assign w33487 = pi2862 & ~w32779;
assign w33488 = ~w33486 & ~w33487;
assign w33489 = ~w30476 & w32779;
assign w33490 = pi2863 & ~w32779;
assign w33491 = ~w33489 & ~w33490;
assign w33492 = ~w30484 & w32779;
assign w33493 = pi2864 & ~w32779;
assign w33494 = ~w33492 & ~w33493;
assign w33495 = ~w30500 & w32779;
assign w33496 = pi2865 & ~w32779;
assign w33497 = ~w33495 & ~w33496;
assign w33498 = ~w30508 & w32779;
assign w33499 = pi2866 & ~w32779;
assign w33500 = ~w33498 & ~w33499;
assign w33501 = ~w30516 & w32779;
assign w33502 = pi2867 & ~w32779;
assign w33503 = ~w33501 & ~w33502;
assign w33504 = ~w29852 & w32779;
assign w33505 = pi2868 & ~w32779;
assign w33506 = ~w33504 & ~w33505;
assign w33507 = ~w29852 & w32801;
assign w33508 = pi2869 & ~w32801;
assign w33509 = ~w33507 & ~w33508;
assign w33510 = ~w30468 & w32820;
assign w33511 = pi2870 & ~w32820;
assign w33512 = ~w33510 & ~w33511;
assign w33513 = ~w30476 & w32820;
assign w33514 = pi2871 & ~w32820;
assign w33515 = ~w33513 & ~w33514;
assign w33516 = ~w30484 & w32820;
assign w33517 = pi2872 & ~w32820;
assign w33518 = ~w33516 & ~w33517;
assign w33519 = ~w30492 & w32820;
assign w33520 = pi2873 & ~w32820;
assign w33521 = ~w33519 & ~w33520;
assign w33522 = ~w30500 & w32820;
assign w33523 = pi2874 & ~w32820;
assign w33524 = ~w33522 & ~w33523;
assign w33525 = ~w30508 & w32820;
assign w33526 = pi2875 & ~w32820;
assign w33527 = ~w33525 & ~w33526;
assign w33528 = ~w29844 & w32820;
assign w33529 = pi2876 & ~w32820;
assign w33530 = ~w33528 & ~w33529;
assign w33531 = ~w30516 & w32820;
assign w33532 = pi2877 & ~w32820;
assign w33533 = ~w33531 & ~w33532;
assign w33534 = ~w29852 & w32820;
assign w33535 = pi2878 & ~w32820;
assign w33536 = ~w33534 & ~w33535;
assign w33537 = ~w17426 & w32820;
assign w33538 = pi2879 & ~w32820;
assign w33539 = ~w33537 & ~w33538;
assign w33540 = pi2880 & ~w33359;
assign w33541 = ~pi0824 & w33359;
assign w33542 = ~w33540 & ~w33541;
assign w33543 = pi2881 & ~w33262;
assign w33544 = ~pi0730 & w33262;
assign w33545 = ~w33543 & ~w33544;
assign w33546 = pi2882 & ~w33204;
assign w33547 = pi0937 & w33204;
assign w33548 = ~w33546 & ~w33547;
assign w33549 = pi2883 & ~w33262;
assign w33550 = ~pi0858 & w33262;
assign w33551 = ~w33549 & ~w33550;
assign w33552 = pi2884 & ~w33359;
assign w33553 = ~pi0731 & w33359;
assign w33554 = ~w33552 & ~w33553;
assign w33555 = pi2885 & ~w33254;
assign w33556 = ~pi0856 & w33254;
assign w33557 = ~w33555 & ~w33556;
assign w33558 = pi2886 & ~w33241;
assign w33559 = ~pi0856 & w33241;
assign w33560 = ~w33558 & ~w33559;
assign w33561 = w24212 & w32027;
assign w33562 = pi2887 & ~w33561;
assign w33563 = ~pi0825 & w33561;
assign w33564 = ~w33562 & ~w33563;
assign w33565 = pi2888 & ~w33416;
assign w33566 = w40189 & w33416;
assign w33567 = ~w33565 & ~w33566;
assign w33568 = pi2889 & ~w33416;
assign w33569 = w40191 & w33416;
assign w33570 = ~w33568 & ~w33569;
assign w33571 = pi2890 & ~w33416;
assign w33572 = w14325 & w33416;
assign w33573 = ~w33571 & ~w33572;
assign w33574 = pi2891 & ~w33416;
assign w33575 = w40176 & w33416;
assign w33576 = ~w33574 & ~w33575;
assign w33577 = pi2892 & ~w33416;
assign w33578 = w13916 & w33416;
assign w33579 = ~w33577 & ~w33578;
assign w33580 = pi2893 & ~w33416;
assign w33581 = w40159 & w33416;
assign w33582 = ~w33580 & ~w33581;
assign w33583 = ~w10746 & w33416;
assign w33584 = pi2894 & ~w33416;
assign w33585 = ~w33583 & ~w33584;
assign w33586 = pi2895 & ~w33416;
assign w33587 = ~w16842 & w33416;
assign w33588 = ~w33586 & ~w33587;
assign w33589 = pi2896 & ~w33416;
assign w33590 = w15978 & w33416;
assign w33591 = ~w33589 & ~w33590;
assign w33592 = pi2897 & ~w33416;
assign w33593 = w40171 & w33416;
assign w33594 = ~w33592 & ~w33593;
assign w33595 = pi2898 & ~w33258;
assign w33596 = ~pi0730 & w33258;
assign w33597 = ~w33595 & ~w33596;
assign w33598 = pi2899 & ~w33204;
assign w33599 = ~pi0823 & w33204;
assign w33600 = ~w33598 & ~w33599;
assign w33601 = pi2900 & ~w33561;
assign w33602 = ~pi0731 & w33561;
assign w33603 = ~w33601 & ~w33602;
assign w33604 = pi2901 & ~w33561;
assign w33605 = ~pi0856 & w33561;
assign w33606 = ~w33604 & ~w33605;
assign w33607 = pi2902 & ~w33258;
assign w33608 = ~pi0853 & w33258;
assign w33609 = ~w33607 & ~w33608;
assign w33610 = pi2903 & ~w33262;
assign w33611 = ~pi0938 & w33262;
assign w33612 = ~w33610 & ~w33611;
assign w33613 = pi2904 & ~w33258;
assign w33614 = ~pi0855 & w33258;
assign w33615 = ~w33613 & ~w33614;
assign w33616 = pi2905 & ~w33262;
assign w33617 = ~pi0860 & w33262;
assign w33618 = ~w33616 & ~w33617;
assign w33619 = pi2906 & ~w33254;
assign w33620 = ~pi0855 & w33254;
assign w33621 = ~w33619 & ~w33620;
assign w33622 = pi2907 & ~w33561;
assign w33623 = ~pi0852 & w33561;
assign w33624 = ~w33622 & ~w33623;
assign w33625 = pi2908 & ~w33561;
assign w33626 = ~pi0854 & w33561;
assign w33627 = ~w33625 & ~w33626;
assign w33628 = pi2909 & ~w33254;
assign w33629 = ~pi0854 & w33254;
assign w33630 = ~w33628 & ~w33629;
assign w33631 = pi2910 & ~w33254;
assign w33632 = ~pi0825 & w33254;
assign w33633 = ~w33631 & ~w33632;
assign w33634 = ~w343 & ~w13989;
assign w33635 = ~pi2911 & w343;
assign w33636 = w17481 & ~w33635;
assign w33637 = ~w33634 & w33636;
assign w33638 = ~w343 & ~w13960;
assign w33639 = ~pi2912 & w343;
assign w33640 = w17481 & ~w33639;
assign w33641 = ~w33638 & w33640;
assign w33642 = ~w343 & ~w13969;
assign w33643 = ~pi2913 & w343;
assign w33644 = w17481 & ~w33643;
assign w33645 = ~w33642 & w33644;
assign w33646 = pi2914 & ~w33416;
assign w33647 = w16629 & w33416;
assign w33648 = ~w33646 & ~w33647;
assign w33649 = pi2915 & ~w33204;
assign w33650 = ~pi0857 & w33204;
assign w33651 = ~w33649 & ~w33650;
assign w33652 = ~w30452 & w33214;
assign w33653 = pi2916 & ~w33214;
assign w33654 = ~w33652 & ~w33653;
assign w33655 = ~w30460 & w33214;
assign w33656 = pi2917 & ~w33214;
assign w33657 = ~w33655 & ~w33656;
assign w33658 = ~w30468 & w33214;
assign w33659 = pi2918 & ~w33214;
assign w33660 = ~w33658 & ~w33659;
assign w33661 = ~w30476 & w33214;
assign w33662 = pi2919 & ~w33214;
assign w33663 = ~w33661 & ~w33662;
assign w33664 = ~w30492 & w33214;
assign w33665 = pi2920 & ~w33214;
assign w33666 = ~w33664 & ~w33665;
assign w33667 = ~w30500 & w33214;
assign w33668 = pi2921 & ~w33214;
assign w33669 = ~w33667 & ~w33668;
assign w33670 = ~w30508 & w33214;
assign w33671 = pi2922 & ~w33214;
assign w33672 = ~w33670 & ~w33671;
assign w33673 = ~w29844 & w33214;
assign w33674 = pi2923 & ~w33214;
assign w33675 = ~w33673 & ~w33674;
assign w33676 = ~w30516 & w33214;
assign w33677 = pi2924 & ~w33214;
assign w33678 = ~w33676 & ~w33677;
assign w33679 = ~w29852 & w33214;
assign w33680 = pi2925 & ~w33214;
assign w33681 = ~w33679 & ~w33680;
assign w33682 = ~w30524 & w33214;
assign w33683 = pi2926 & ~w33214;
assign w33684 = ~w33682 & ~w33683;
assign w33685 = ~w30532 & w33214;
assign w33686 = pi2927 & ~w33214;
assign w33687 = ~w33685 & ~w33686;
assign w33688 = ~w30548 & w33214;
assign w33689 = pi2928 & ~w33214;
assign w33690 = ~w33688 & ~w33689;
assign w33691 = ~w17426 & w33214;
assign w33692 = pi2929 & ~w33214;
assign w33693 = ~w33691 & ~w33692;
assign w33694 = pi2930 & ~w33204;
assign w33695 = ~pi0825 & w33204;
assign w33696 = ~w33694 & ~w33695;
assign w33697 = pi2931 & ~w33266;
assign w33698 = w40189 & w33266;
assign w33699 = ~w33697 & ~w33698;
assign w33700 = pi2932 & ~w33266;
assign w33701 = w40174 & w33266;
assign w33702 = ~w33700 & ~w33701;
assign w33703 = pi2933 & ~w33266;
assign w33704 = w40168 & w33266;
assign w33705 = ~w33703 & ~w33704;
assign w33706 = pi2934 & ~w33266;
assign w33707 = w13916 & w33266;
assign w33708 = ~w33706 & ~w33707;
assign w33709 = pi2935 & ~w33266;
assign w33710 = w40159 & w33266;
assign w33711 = ~w33709 & ~w33710;
assign w33712 = pi2936 & ~w33266;
assign w33713 = w16739 & w33266;
assign w33714 = ~w33712 & ~w33713;
assign w33715 = pi2937 & ~w33266;
assign w33716 = w15171 & w33266;
assign w33717 = ~w33715 & ~w33716;
assign w33718 = pi2938 & ~w33266;
assign w33719 = w40171 & w33266;
assign w33720 = ~w33718 & ~w33719;
assign w33721 = pi2939 & ~w33230;
assign w33722 = w40189 & w33230;
assign w33723 = ~w33721 & ~w33722;
assign w33724 = pi2940 & ~w33230;
assign w33725 = w40191 & w33230;
assign w33726 = ~w33724 & ~w33725;
assign w33727 = pi2941 & ~w33230;
assign w33728 = w14325 & w33230;
assign w33729 = ~w33727 & ~w33728;
assign w33730 = pi2942 & ~w33230;
assign w33731 = w14962 & w33230;
assign w33732 = ~w33730 & ~w33731;
assign w33733 = pi2943 & ~w33230;
assign w33734 = w40168 & w33230;
assign w33735 = ~w33733 & ~w33734;
assign w33736 = pi2944 & ~w33230;
assign w33737 = w40176 & w33230;
assign w33738 = ~w33736 & ~w33737;
assign w33739 = pi2945 & ~w33230;
assign w33740 = w13916 & w33230;
assign w33741 = ~w33739 & ~w33740;
assign w33742 = ~w10746 & w33230;
assign w33743 = pi2946 & ~w33230;
assign w33744 = ~w33742 & ~w33743;
assign w33745 = pi2947 & ~w33230;
assign w33746 = w16629 & w33230;
assign w33747 = ~w33745 & ~w33746;
assign w33748 = pi2948 & ~w33230;
assign w33749 = w16739 & w33230;
assign w33750 = ~w33748 & ~w33749;
assign w33751 = pi2949 & ~w33230;
assign w33752 = ~w16842 & w33230;
assign w33753 = ~w33751 & ~w33752;
assign w33754 = pi2950 & ~w33230;
assign w33755 = w40171 & w33230;
assign w33756 = ~w33754 & ~w33755;
assign w33757 = pi1930 & ~w343;
assign w33758 = pi1826 & w33757;
assign w33759 = ~pi2951 & ~w33757;
assign w33760 = w6682 & ~w33759;
assign w33761 = ~w33758 & w33760;
assign w33762 = pi1825 & w33757;
assign w33763 = ~pi2952 & ~w33757;
assign w33764 = w6682 & ~w33763;
assign w33765 = ~w33762 & w33764;
assign w33766 = w21489 & ~w31987;
assign w33767 = pi2953 & ~w21489;
assign w33768 = ~w33766 & ~w33767;
assign w33769 = pi2954 & ~w33561;
assign w33770 = ~pi0824 & w33561;
assign w33771 = ~w33769 & ~w33770;
assign w33772 = pi2955 & ~w33561;
assign w33773 = ~pi0859 & w33561;
assign w33774 = ~w33772 & ~w33773;
assign w33775 = pi2956 & ~w33254;
assign w33776 = ~pi0731 & w33254;
assign w33777 = ~w33775 & ~w33776;
assign w33778 = pi2957 & ~w33204;
assign w33779 = ~pi0860 & w33204;
assign w33780 = ~w33778 & ~w33779;
assign w33781 = pi2958 & ~w33204;
assign w33782 = ~pi0852 & w33204;
assign w33783 = ~w33781 & ~w33782;
assign w33784 = pi2959 & ~w33241;
assign w33785 = ~pi0857 & w33241;
assign w33786 = ~w33784 & ~w33785;
assign w33787 = w2315 & w23938;
assign w33788 = ~w3858 & ~w33787;
assign w33789 = w2315 & w23954;
assign w33790 = ~w2926 & ~w33789;
assign w33791 = w2315 & w23971;
assign w33792 = ~w2878 & ~w33791;
assign w33793 = w2315 & w23988;
assign w33794 = ~w23992 & ~w33793;
assign w33795 = w2315 & w24037;
assign w33796 = ~w3765 & ~w33795;
assign w33797 = w2323 & w23938;
assign w33798 = ~w23943 & ~w33797;
assign w33799 = w2323 & ~w23988;
assign w33800 = ~pi2966 & ~w2323;
assign w33801 = ~w33799 & ~w33800;
assign w33802 = w2323 & ~w24020;
assign w33803 = ~w24025 & ~w33802;
assign w33804 = w2323 & w24037;
assign w33805 = ~w3768 & ~w33804;
assign w33806 = pi2969 & ~w33416;
assign w33807 = w16739 & w33416;
assign w33808 = ~w33806 & ~w33807;
assign w33809 = pi2970 & ~w33258;
assign w33810 = ~pi0851 & w33258;
assign w33811 = ~w33809 & ~w33810;
assign w33812 = pi2971 & ~w33204;
assign w33813 = ~pi0851 & w33204;
assign w33814 = ~w33812 & ~w33813;
assign w33815 = pi2972 & ~w33241;
assign w33816 = ~pi0825 & w33241;
assign w33817 = ~w33815 & ~w33816;
assign w33818 = pi2973 & ~w33262;
assign w33819 = ~pi0821 & w33262;
assign w33820 = ~w33818 & ~w33819;
assign w33821 = ~pi0833 & ~w370;
assign w33822 = w40134 & w33821;
assign w33823 = ~pi2974 & pi3237;
assign w33824 = ~w33821 & w33823;
assign w33825 = ~w33822 & ~w33824;
assign w33826 = w5914 & w33821;
assign w33827 = ~pi2975 & pi3239;
assign w33828 = ~w33821 & w33827;
assign w33829 = ~w33826 & ~w33828;
assign w33830 = w3711 & w33821;
assign w33831 = ~pi2976 & pi3227;
assign w33832 = ~w33821 & w33831;
assign w33833 = ~w33830 & ~w33832;
assign w33834 = pi2977 & ~w33241;
assign w33835 = ~pi0852 & w33241;
assign w33836 = ~w33834 & ~w33835;
assign w33837 = ~pi1000 & w6668;
assign w33838 = pi2978 & ~w33837;
assign w33839 = w5320 & w33837;
assign w33840 = ~w33838 & ~w33839;
assign w33841 = pi2979 & ~w33837;
assign w33842 = w5914 & w33837;
assign w33843 = ~w33841 & ~w33842;
assign w33844 = pi2980 & ~w33837;
assign w33845 = w4749 & w33837;
assign w33846 = ~w33844 & ~w33845;
assign w33847 = pi2981 & ~w33837;
assign w33848 = w3711 & w33837;
assign w33849 = ~w33847 & ~w33848;
assign w33850 = pi2982 & w343;
assign w33851 = w6682 & ~w29978;
assign w33852 = ~w33850 & w33851;
assign w33853 = ~pi2983 & w6684;
assign w33854 = pi0422 & w21820;
assign w33855 = w21968 & w33854;
assign w33856 = ~w33853 & ~w33855;
assign w33857 = pi2984 & ~w33241;
assign w33858 = ~pi0854 & w33241;
assign w33859 = ~w33857 & ~w33858;
assign w33860 = w156 & w896;
assign w33861 = pi2985 & ~w33860;
assign w33862 = pi3686 & w33860;
assign w33863 = ~w33861 & ~w33862;
assign w33864 = pi2986 & ~w32432;
assign w33865 = w4749 & w32432;
assign w33866 = ~w33864 & ~w33865;
assign w33867 = pi2987 & ~w32432;
assign w33868 = w8081 & w32432;
assign w33869 = ~w33867 & ~w33868;
assign w33870 = pi2988 & ~w32432;
assign w33871 = w1639 & w32432;
assign w33872 = ~w33870 & ~w33871;
assign w33873 = pi2989 & ~w32432;
assign w33874 = w1308 & w32432;
assign w33875 = ~w33873 & ~w33874;
assign w33876 = pi2990 & ~w32432;
assign w33877 = w3711 & w32432;
assign w33878 = ~w33876 & ~w33877;
assign w33879 = pi2991 & ~w33241;
assign w33880 = ~pi0851 & w33241;
assign w33881 = ~w33879 & ~w33880;
assign w33882 = pi2994 & ~w33561;
assign w33883 = ~pi0823 & w33561;
assign w33884 = ~w33882 & ~w33883;
assign w33885 = pi2995 & ~w33561;
assign w33886 = ~pi0730 & w33561;
assign w33887 = ~w33885 & ~w33886;
assign w33888 = pi2996 & ~w33561;
assign w33889 = ~pi0853 & w33561;
assign w33890 = ~w33888 & ~w33889;
assign w33891 = pi2997 & ~w33561;
assign w33892 = ~pi0785 & w33561;
assign w33893 = ~w33891 & ~w33892;
assign w33894 = pi2998 & ~w33561;
assign w33895 = ~pi0855 & w33561;
assign w33896 = ~w33894 & ~w33895;
assign w33897 = pi2999 & ~w33561;
assign w33898 = ~pi0857 & w33561;
assign w33899 = ~w33897 & ~w33898;
assign w33900 = pi3000 & ~w33561;
assign w33901 = ~pi0858 & w33561;
assign w33902 = ~w33900 & ~w33901;
assign w33903 = pi3001 & ~w33561;
assign w33904 = ~pi0821 & w33561;
assign w33905 = ~w33903 & ~w33904;
assign w33906 = pi3002 & ~w33359;
assign w33907 = ~pi0823 & w33359;
assign w33908 = ~w33906 & ~w33907;
assign w33909 = pi3003 & ~w33359;
assign w33910 = ~pi0859 & w33359;
assign w33911 = ~w33909 & ~w33910;
assign w33912 = pi3004 & ~w33359;
assign w33913 = ~pi0730 & w33359;
assign w33914 = ~w33912 & ~w33913;
assign w33915 = pi3005 & ~w33359;
assign w33916 = ~pi0853 & w33359;
assign w33917 = ~w33915 & ~w33916;
assign w33918 = pi3006 & ~w33359;
assign w33919 = ~pi0785 & w33359;
assign w33920 = ~w33918 & ~w33919;
assign w33921 = pi3007 & ~w33359;
assign w33922 = ~pi0855 & w33359;
assign w33923 = ~w33921 & ~w33922;
assign w33924 = pi3008 & ~w33359;
assign w33925 = ~pi0821 & w33359;
assign w33926 = ~w33924 & ~w33925;
assign w33927 = pi3009 & ~w33241;
assign w33928 = ~pi0824 & w33241;
assign w33929 = ~w33927 & ~w33928;
assign w33930 = pi3010 & ~w33241;
assign w33931 = ~pi0823 & w33241;
assign w33932 = ~w33930 & ~w33931;
assign w33933 = pi3011 & ~w33241;
assign w33934 = ~pi0730 & w33241;
assign w33935 = ~w33933 & ~w33934;
assign w33936 = pi3012 & ~w33241;
assign w33937 = ~pi0860 & w33241;
assign w33938 = ~w33936 & ~w33937;
assign w33939 = pi3013 & ~w33241;
assign w33940 = ~pi0853 & w33241;
assign w33941 = ~w33939 & ~w33940;
assign w33942 = pi3014 & ~w33241;
assign w33943 = ~pi0785 & w33241;
assign w33944 = ~w33942 & ~w33943;
assign w33945 = pi3015 & ~w33241;
assign w33946 = ~pi0855 & w33241;
assign w33947 = ~w33945 & ~w33946;
assign w33948 = pi3016 & ~w33241;
assign w33949 = ~pi0821 & w33241;
assign w33950 = ~w33948 & ~w33949;
assign w33951 = pi3017 & ~w33254;
assign w33952 = ~pi0823 & w33254;
assign w33953 = ~w33951 & ~w33952;
assign w33954 = pi3018 & ~w33254;
assign w33955 = ~pi0730 & w33254;
assign w33956 = ~w33954 & ~w33955;
assign w33957 = pi3019 & ~w33254;
assign w33958 = ~pi0938 & w33254;
assign w33959 = ~w33957 & ~w33958;
assign w33960 = pi3020 & ~w33254;
assign w33961 = ~pi0860 & w33254;
assign w33962 = ~w33960 & ~w33961;
assign w33963 = pi3021 & ~w33254;
assign w33964 = ~pi0852 & w33254;
assign w33965 = ~w33963 & ~w33964;
assign w33966 = pi3022 & ~w33254;
assign w33967 = ~pi0853 & w33254;
assign w33968 = ~w33966 & ~w33967;
assign w33969 = pi3023 & ~w33254;
assign w33970 = ~pi0857 & w33254;
assign w33971 = ~w33969 & ~w33970;
assign w33972 = pi3024 & ~w33254;
assign w33973 = ~pi0858 & w33254;
assign w33974 = ~w33972 & ~w33973;
assign w33975 = pi3025 & ~w33254;
assign w33976 = ~pi0821 & w33254;
assign w33977 = ~w33975 & ~w33976;
assign w33978 = pi3026 & ~w33475;
assign w33979 = ~pi0824 & w33475;
assign w33980 = ~w33978 & ~w33979;
assign w33981 = pi3027 & ~w33475;
assign w33982 = ~pi0731 & w33475;
assign w33983 = ~w33981 & ~w33982;
assign w33984 = pi3028 & ~w33475;
assign w33985 = ~pi0852 & w33475;
assign w33986 = ~w33984 & ~w33985;
assign w33987 = pi3029 & ~w33475;
assign w33988 = ~pi0854 & w33475;
assign w33989 = ~w33987 & ~w33988;
assign w33990 = pi3030 & ~w33475;
assign w33991 = ~pi0856 & w33475;
assign w33992 = ~w33990 & ~w33991;
assign w33993 = pi3031 & ~w33475;
assign w33994 = ~pi0858 & w33475;
assign w33995 = ~w33993 & ~w33994;
assign w33996 = pi3032 & ~w33475;
assign w33997 = ~pi0821 & w33475;
assign w33998 = ~w33996 & ~w33997;
assign w33999 = pi3033 & ~w33262;
assign w34000 = ~pi0824 & w33262;
assign w34001 = ~w33999 & ~w34000;
assign w34002 = pi3034 & ~w33262;
assign w34003 = ~pi0859 & w33262;
assign w34004 = ~w34002 & ~w34003;
assign w34005 = pi3035 & ~w33262;
assign w34006 = ~pi0731 & w33262;
assign w34007 = ~w34005 & ~w34006;
assign w34008 = pi3036 & ~w33262;
assign w34009 = ~pi0851 & w33262;
assign w34010 = ~w34008 & ~w34009;
assign w34011 = pi3037 & ~w33262;
assign w34012 = ~pi0852 & w33262;
assign w34013 = ~w34011 & ~w34012;
assign w34014 = pi3038 & ~w33262;
assign w34015 = ~pi0854 & w33262;
assign w34016 = ~w34014 & ~w34015;
assign w34017 = pi3039 & ~w33262;
assign w34018 = ~pi0825 & w33262;
assign w34019 = ~w34017 & ~w34018;
assign w34020 = pi3040 & ~w33258;
assign w34021 = ~pi0823 & w33258;
assign w34022 = ~w34020 & ~w34021;
assign w34023 = pi3041 & ~w33258;
assign w34024 = ~pi0860 & w33258;
assign w34025 = ~w34023 & ~w34024;
assign w34026 = pi3042 & ~w33258;
assign w34027 = ~pi0821 & w33258;
assign w34028 = ~w34026 & ~w34027;
assign w34029 = pi3043 & ~w33258;
assign w34030 = ~pi0854 & w33258;
assign w34031 = ~w34029 & ~w34030;
assign w34032 = pi3044 & ~w33258;
assign w34033 = ~pi0825 & w33258;
assign w34034 = ~w34032 & ~w34033;
assign w34035 = pi3045 & ~w33258;
assign w34036 = ~pi0856 & w33258;
assign w34037 = ~w34035 & ~w34036;
assign w34038 = pi3046 & ~w33258;
assign w34039 = ~pi0858 & w33258;
assign w34040 = ~w34038 & ~w34039;
assign w34041 = pi3047 & ~w33258;
assign w34042 = pi0937 & w33258;
assign w34043 = ~w34041 & ~w34042;
assign w34044 = pi3048 & ~w33204;
assign w34045 = ~pi0859 & w33204;
assign w34046 = ~w34044 & ~w34045;
assign w34047 = pi3049 & ~w33204;
assign w34048 = ~pi0730 & w33204;
assign w34049 = ~w34047 & ~w34048;
assign w34050 = pi3050 & ~w33204;
assign w34051 = ~pi0731 & w33204;
assign w34052 = ~w34050 & ~w34051;
assign w34053 = pi3051 & ~w33204;
assign w34054 = ~pi0853 & w33204;
assign w34055 = ~w34053 & ~w34054;
assign w34056 = pi3052 & ~w33204;
assign w34057 = ~pi0854 & w33204;
assign w34058 = ~w34056 & ~w34057;
assign w34059 = pi3053 & ~w33204;
assign w34060 = ~pi0785 & w33204;
assign w34061 = ~w34059 & ~w34060;
assign w34062 = pi3054 & ~w33204;
assign w34063 = ~pi0855 & w33204;
assign w34064 = ~w34062 & ~w34063;
assign w34065 = pi3055 & ~w33479;
assign w34066 = pi0853 & w33479;
assign w34067 = ~w34065 & ~w34066;
assign w34068 = pi3056 & ~w33241;
assign w34069 = ~pi0731 & w33241;
assign w34070 = ~w34068 & ~w34069;
assign w34071 = pi3057 & ~w33475;
assign w34072 = ~pi0785 & w33475;
assign w34073 = ~w34071 & ~w34072;
assign w34074 = pi3058 & ~w33475;
assign w34075 = ~pi0825 & w33475;
assign w34076 = ~w34074 & ~w34075;
assign w34077 = pi3059 & ~w33416;
assign w34078 = w40168 & w33416;
assign w34079 = ~w34077 & ~w34078;
assign w34080 = pi3060 & ~w33475;
assign w34081 = ~pi0851 & w33475;
assign w34082 = ~w34080 & ~w34081;
assign w34083 = pi3061 & ~w33258;
assign w34084 = ~pi0824 & w33258;
assign w34085 = ~w34083 & ~w34084;
assign w34086 = pi3062 & ~w33475;
assign w34087 = ~pi0938 & w33475;
assign w34088 = ~w34086 & ~w34087;
assign w34089 = pi3063 & ~w32432;
assign w34090 = w5053 & w32432;
assign w34091 = ~w34089 & ~w34090;
assign w34092 = pi3064 & ~w33262;
assign w34093 = ~pi0855 & w33262;
assign w34094 = ~w34092 & ~w34093;
assign w34095 = ~pi3065 & w343;
assign w34096 = ~w30565 & ~w34095;
assign w34097 = w6682 & ~w34096;
assign w34098 = pi3066 & ~w33254;
assign w34099 = ~pi0859 & w33254;
assign w34100 = ~w34098 & ~w34099;
assign w34101 = pi3067 & ~w33561;
assign w34102 = ~pi0851 & w33561;
assign w34103 = ~w34101 & ~w34102;
assign w34104 = w4380 & w33821;
assign w34105 = ~pi3068 & pi3217;
assign w34106 = ~w33821 & w34105;
assign w34107 = ~w34104 & ~w34106;
assign w34108 = pi3069 & ~w33204;
assign w34109 = ~pi0858 & w33204;
assign w34110 = ~w34108 & ~w34109;
assign w34111 = pi3070 & ~w33475;
assign w34112 = ~pi0855 & w33475;
assign w34113 = ~w34111 & ~w34112;
assign w34114 = pi3071 & ~w33262;
assign w34115 = ~pi0856 & w33262;
assign w34116 = ~w34114 & ~w34115;
assign w34117 = pi3072 & ~w33561;
assign w34118 = ~pi0938 & w33561;
assign w34119 = ~w34117 & ~w34118;
assign w34120 = pi3073 & ~w33561;
assign w34121 = ~pi0860 & w33561;
assign w34122 = ~w34120 & ~w34121;
assign w34123 = pi3074 & ~w33416;
assign w34124 = w14962 & w33416;
assign w34125 = ~w34123 & ~w34124;
assign w34126 = pi3075 & ~w33416;
assign w34127 = w40174 & w33416;
assign w34128 = ~w34126 & ~w34127;
assign w34129 = pi1827 & w33757;
assign w34130 = ~pi3076 & ~w33757;
assign w34131 = w6682 & ~w34130;
assign w34132 = ~w34129 & w34131;
assign w34133 = pi3077 & ~w33359;
assign w34134 = ~pi0857 & w33359;
assign w34135 = ~w34133 & ~w34134;
assign w34136 = pi3078 & ~w33475;
assign w34137 = ~pi0857 & w33475;
assign w34138 = ~w34136 & ~w34137;
assign w34139 = pi3079 & ~w33230;
assign w34140 = w15978 & w33230;
assign w34141 = ~w34139 & ~w34140;
assign w34142 = pi3080 & ~w33204;
assign w34143 = ~pi0856 & w33204;
assign w34144 = ~w34142 & ~w34143;
assign w34145 = pi3081 & ~w33475;
assign w34146 = ~pi0823 & w33475;
assign w34147 = ~w34145 & ~w34146;
assign w34148 = pi3082 & ~w33262;
assign w34149 = ~pi0853 & w33262;
assign w34150 = ~w34148 & ~w34149;
assign w34151 = pi3083 & ~w33475;
assign w34152 = ~pi0853 & w33475;
assign w34153 = ~w34151 & ~w34152;
assign w34154 = ~w17426 & w32779;
assign w34155 = pi3084 & ~w32779;
assign w34156 = ~w34154 & ~w34155;
assign w34157 = pi3085 & ~w33359;
assign w34158 = ~pi0858 & w33359;
assign w34159 = ~w34157 & ~w34158;
assign w34160 = pi0853 & pi3086;
assign w34161 = w24189 & w34160;
assign w34162 = w32027 & w34161;
assign w34163 = pi3087 & ~w33475;
assign w34164 = ~pi0859 & w33475;
assign w34165 = ~w34163 & ~w34164;
assign w34166 = pi3088 & ~w33258;
assign w34167 = ~pi0857 & w33258;
assign w34168 = ~w34166 & ~w34167;
assign w34169 = pi3089 & ~w33262;
assign w34170 = ~pi0785 & w33262;
assign w34171 = ~w34169 & ~w34170;
assign w34172 = pi3090 & ~w33475;
assign w34173 = ~pi0730 & w33475;
assign w34174 = ~w34172 & ~w34173;
assign w34175 = pi3091 & ~w32432;
assign w34176 = w5635 & w32432;
assign w34177 = ~w34175 & ~w34176;
assign w34178 = pi3092 & ~w33258;
assign w34179 = ~pi0731 & w33258;
assign w34180 = ~w34178 & ~w34179;
assign w34181 = w2323 & w23971;
assign w34182 = ~w23975 & ~w34181;
assign w34183 = pi3094 & ~w33359;
assign w34184 = ~pi0856 & w33359;
assign w34185 = ~w34183 & ~w34184;
assign w34186 = pi3095 & ~w33241;
assign w34187 = ~pi0859 & w33241;
assign w34188 = ~w34186 & ~w34187;
assign w34189 = w2323 & w23954;
assign w34190 = ~w23958 & ~w34189;
assign w34191 = pi3097 & ~w32432;
assign w34192 = w8240 & w32432;
assign w34193 = ~w34191 & ~w34192;
assign w34194 = pi3098 & ~w33479;
assign w34195 = ~pi0825 & w33479;
assign w34196 = ~w34194 & ~w34195;
assign w34197 = pi3099 & ~w32432;
assign w34198 = w5914 & w32432;
assign w34199 = ~w34197 & ~w34198;
assign w34200 = pi3100 & ~w32432;
assign w34201 = w5320 & w32432;
assign w34202 = ~w34200 & ~w34201;
assign w34203 = pi3101 & ~w32432;
assign w34204 = w6177 & w32432;
assign w34205 = ~w34203 & ~w34204;
assign w34206 = pi3102 & ~w33860;
assign w34207 = pi3687 & w33860;
assign w34208 = ~w34206 & ~w34207;
assign w34209 = pi3103 & ~w33258;
assign w34210 = ~pi0859 & w33258;
assign w34211 = ~w34209 & ~w34210;
assign w34212 = pi3104 & ~w33860;
assign w34213 = pi3685 & w33860;
assign w34214 = ~w34212 & ~w34213;
assign w34215 = pi3105 & ~w33860;
assign w34216 = pi3684 & w33860;
assign w34217 = ~w34215 & ~w34216;
assign w34218 = pi3106 & ~w33860;
assign w34219 = pi3683 & w33860;
assign w34220 = ~w34218 & ~w34219;
assign w34221 = pi3107 & ~w32432;
assign w34222 = w4141 & w32432;
assign w34223 = ~w34221 & ~w34222;
assign w34224 = pi3108 & ~w33241;
assign w34225 = ~pi0938 & w33241;
assign w34226 = ~w34224 & ~w34225;
assign w34227 = pi3109 & ~w33860;
assign w34228 = pi3688 & w33860;
assign w34229 = ~w34227 & ~w34228;
assign w34230 = pi3110 & ~w33204;
assign w34231 = ~pi0938 & w33204;
assign w34232 = ~w34230 & ~w34231;
assign w34233 = pi3111 & ~w33860;
assign w34234 = pi3689 & w33860;
assign w34235 = ~w34233 & ~w34234;
assign w34236 = pi3112 & ~w33860;
assign w34237 = pi3690 & w33860;
assign w34238 = ~w34236 & ~w34237;
assign w34239 = pi3113 & ~w33230;
assign w34240 = w15171 & w33230;
assign w34241 = ~w34239 & ~w34240;
assign w34242 = pi3114 & ~w33757;
assign w34243 = ~pi0408 & w6975;
assign w34244 = pi2047 & ~w34243;
assign w34245 = pi2029 & w34243;
assign w34246 = ~w34244 & ~w34245;
assign w34247 = w33757 & w34246;
assign w34248 = ~w34242 & ~w34247;
assign w34249 = pi3115 & ~w33757;
assign w34250 = ~pi2045 & ~w34243;
assign w34251 = w33757 & w34250;
assign w34252 = ~w34249 & ~w34251;
assign w34253 = pi3116 & ~w33757;
assign w34254 = ~pi2065 & ~w34243;
assign w34255 = w33757 & w34254;
assign w34256 = ~w34253 & ~w34255;
assign w34257 = pi3117 & ~w33757;
assign w34258 = ~pi2037 & ~w34243;
assign w34259 = w33757 & w34258;
assign w34260 = ~w34257 & ~w34259;
assign w34261 = pi3118 & ~w33757;
assign w34262 = pi2046 & ~w34243;
assign w34263 = pi2030 & w34243;
assign w34264 = ~w34262 & ~w34263;
assign w34265 = w33757 & w34264;
assign w34266 = ~w34261 & ~w34265;
assign w34267 = ~pi0579 & w40209;
assign w34268 = pi3119 & ~w34267;
assign w34269 = w16739 & w34267;
assign w34270 = ~w34268 & ~w34269;
assign w34271 = pi3120 & w6684;
assign w34272 = w6971 & w22006;
assign w34273 = w21969 & w34272;
assign w34274 = ~w34271 & ~w34273;
assign w34275 = pi3121 & w6684;
assign w34276 = ~w32384 & ~w34275;
assign w34277 = pi3122 & ~w34267;
assign w34278 = w13916 & w34267;
assign w34279 = ~w34277 & ~w34278;
assign w34280 = pi3123 & ~w34267;
assign w34281 = w40159 & w34267;
assign w34282 = ~w34280 & ~w34281;
assign w34283 = pi3124 & ~w33757;
assign w34284 = ~pi2062 & ~w34243;
assign w34285 = w33757 & w34284;
assign w34286 = ~w34283 & ~w34285;
assign w34287 = pi3125 & ~w34267;
assign w34288 = w40174 & w34267;
assign w34289 = ~w34287 & ~w34288;
assign w34290 = pi3126 & ~w34267;
assign w34291 = w40189 & w34267;
assign w34292 = ~w34290 & ~w34291;
assign w34293 = ~pi0597 & w40209;
assign w34294 = pi3127 & ~w34293;
assign w34295 = w40171 & w34293;
assign w34296 = ~w34294 & ~w34295;
assign w34297 = pi3128 & ~w34293;
assign w34298 = w40159 & w34293;
assign w34299 = ~w34297 & ~w34298;
assign w34300 = ~pi3130 & w343;
assign w34301 = w9066 & w14359;
assign w34302 = ~w34300 & ~w34301;
assign w34303 = pi3131 & ~w34293;
assign w34304 = w40176 & w34293;
assign w34305 = ~w34303 & ~w34304;
assign w34306 = pi3132 & ~w34293;
assign w34307 = w40168 & w34293;
assign w34308 = ~w34306 & ~w34307;
assign w34309 = pi3133 & ~w34293;
assign w34310 = w14325 & w34293;
assign w34311 = ~w34309 & ~w34310;
assign w34312 = pi3134 & ~w34293;
assign w34313 = w14962 & w34293;
assign w34314 = ~w34312 & ~w34313;
assign w34315 = pi3135 & ~w33757;
assign w34316 = ~pi2040 & ~w34243;
assign w34317 = w33757 & w34316;
assign w34318 = ~w34315 & ~w34317;
assign w34319 = w24321 & w29785;
assign w34320 = pi1754 & pi2106;
assign w34321 = pi1755 & pi2107;
assign w34322 = ~w34320 & ~w34321;
assign w34323 = pi1751 & pi2103;
assign w34324 = pi1752 & pi2104;
assign w34325 = ~w34323 & ~w34324;
assign w34326 = w34322 & w34325;
assign w34327 = pi1749 & pi2101;
assign w34328 = pi1758 & pi2109;
assign w34329 = ~w34327 & ~w34328;
assign w34330 = pi1757 & pi2108;
assign w34331 = pi1760 & pi2110;
assign w34332 = ~w34330 & ~w34331;
assign w34333 = w34329 & w34332;
assign w34334 = pi1756 & pi2141;
assign w34335 = pi1759 & pi2123;
assign w34336 = ~w34334 & ~w34335;
assign w34337 = pi1753 & pi2105;
assign w34338 = pi1750 & pi2102;
assign w34339 = ~w34337 & ~w34338;
assign w34340 = w34336 & w34339;
assign w34341 = w34333 & w34340;
assign w34342 = w34326 & w34341;
assign w34343 = pi3138 & w370;
assign w34344 = ~w13946 & ~w34343;
assign w34345 = pi3139 & ~w33757;
assign w34346 = ~pi2041 & ~w34243;
assign w34347 = w33757 & w34346;
assign w34348 = ~w34345 & ~w34347;
assign w34349 = ~w30516 & w32801;
assign w34350 = pi3140 & ~w32801;
assign w34351 = ~w34349 & ~w34350;
assign w34352 = pi3143 & ~w34267;
assign w34353 = ~w16842 & w34267;
assign w34354 = ~w34352 & ~w34353;
assign w34355 = ~pi3145 & w370;
assign w34356 = pi2983 & w13945;
assign w34357 = ~w34355 & ~w34356;
assign w34358 = ~pi3146 & w343;
assign w34359 = ~w33218 & ~w34358;
assign w34360 = ~w30377 & ~w30382;
assign w34361 = ~pi3526 & w342;
assign w34362 = ~pi3663 & ~w34361;
assign w34363 = pi3148 & w7173;
assign w34364 = w6681 & w34363;
assign w34365 = w34361 & w34364;
assign w34366 = ~w34362 & ~w34365;
assign w34367 = pi3149 & ~w33343;
assign w34368 = pi3692 & w33343;
assign w34369 = ~w34367 & ~w34368;
assign w34370 = pi3150 & ~w33343;
assign w34371 = pi3691 & w33343;
assign w34372 = ~w34370 & ~w34371;
assign w34373 = ~w30468 & w32760;
assign w34374 = pi3151 & ~w32760;
assign w34375 = ~w34373 & ~w34374;
assign w34376 = ~w30476 & w32760;
assign w34377 = pi3152 & ~w32760;
assign w34378 = ~w34376 & ~w34377;
assign w34379 = ~w30484 & w32760;
assign w34380 = pi3153 & ~w32760;
assign w34381 = ~w34379 & ~w34380;
assign w34382 = ~w30492 & w32760;
assign w34383 = pi3154 & ~w32760;
assign w34384 = ~w34382 & ~w34383;
assign w34385 = ~w30500 & w32760;
assign w34386 = pi3155 & ~w32760;
assign w34387 = ~w34385 & ~w34386;
assign w34388 = ~w30508 & w32760;
assign w34389 = pi3156 & ~w32760;
assign w34390 = ~w34388 & ~w34389;
assign w34391 = ~w29844 & w32760;
assign w34392 = pi3157 & ~w32760;
assign w34393 = ~w34391 & ~w34392;
assign w34394 = ~w30516 & w32760;
assign w34395 = pi3158 & ~w32760;
assign w34396 = ~w34394 & ~w34395;
assign w34397 = ~w17426 & w32760;
assign w34398 = pi3159 & ~w32760;
assign w34399 = ~w34397 & ~w34398;
assign w34400 = ~w30468 & w32801;
assign w34401 = pi3160 & ~w32801;
assign w34402 = ~w34400 & ~w34401;
assign w34403 = ~w30476 & w32801;
assign w34404 = pi3161 & ~w32801;
assign w34405 = ~w34403 & ~w34404;
assign w34406 = ~w30484 & w32801;
assign w34407 = pi3162 & ~w32801;
assign w34408 = ~w34406 & ~w34407;
assign w34409 = ~w30500 & w32801;
assign w34410 = pi3163 & ~w32801;
assign w34411 = ~w34409 & ~w34410;
assign w34412 = ~w30508 & w32801;
assign w34413 = pi3164 & ~w32801;
assign w34414 = ~w34412 & ~w34413;
assign w34415 = ~w29844 & w32801;
assign w34416 = pi3165 & ~w32801;
assign w34417 = ~w34415 & ~w34416;
assign w34418 = ~w17426 & w32801;
assign w34419 = pi3166 & ~w32801;
assign w34420 = ~w34418 & ~w34419;
assign w34421 = pi3167 & ~w34293;
assign w34422 = w40189 & w34293;
assign w34423 = ~w34421 & ~w34422;
assign w34424 = pi3168 & ~w34293;
assign w34425 = w40191 & w34293;
assign w34426 = ~w34424 & ~w34425;
assign w34427 = pi3169 & ~w34293;
assign w34428 = w40174 & w34293;
assign w34429 = ~w34427 & ~w34428;
assign w34430 = pi3170 & ~w34293;
assign w34431 = w13916 & w34293;
assign w34432 = ~w34430 & ~w34431;
assign w34433 = ~w10746 & w34293;
assign w34434 = pi3171 & ~w34293;
assign w34435 = ~w34433 & ~w34434;
assign w34436 = pi3172 & ~w34293;
assign w34437 = w16629 & w34293;
assign w34438 = ~w34436 & ~w34437;
assign w34439 = pi3173 & ~w34293;
assign w34440 = w16739 & w34293;
assign w34441 = ~w34439 & ~w34440;
assign w34442 = pi3174 & ~w34293;
assign w34443 = ~w16842 & w34293;
assign w34444 = ~w34442 & ~w34443;
assign w34445 = pi3175 & ~w34293;
assign w34446 = w15978 & w34293;
assign w34447 = ~w34445 & ~w34446;
assign w34448 = pi3176 & ~w34293;
assign w34449 = w15171 & w34293;
assign w34450 = ~w34448 & ~w34449;
assign w34451 = pi3177 & ~w34267;
assign w34452 = w40191 & w34267;
assign w34453 = ~w34451 & ~w34452;
assign w34454 = pi3178 & ~w34267;
assign w34455 = w14325 & w34267;
assign w34456 = ~w34454 & ~w34455;
assign w34457 = pi3179 & ~w34267;
assign w34458 = w14962 & w34267;
assign w34459 = ~w34457 & ~w34458;
assign w34460 = pi3180 & ~w34267;
assign w34461 = w40168 & w34267;
assign w34462 = ~w34460 & ~w34461;
assign w34463 = pi3181 & ~w34267;
assign w34464 = w40176 & w34267;
assign w34465 = ~w34463 & ~w34464;
assign w34466 = ~w10746 & w34267;
assign w34467 = pi3182 & ~w34267;
assign w34468 = ~w34466 & ~w34467;
assign w34469 = pi3183 & ~w34267;
assign w34470 = w16629 & w34267;
assign w34471 = ~w34469 & ~w34470;
assign w34472 = pi3184 & ~w34267;
assign w34473 = w15978 & w34267;
assign w34474 = ~w34472 & ~w34473;
assign w34475 = pi3185 & ~w34267;
assign w34476 = w15171 & w34267;
assign w34477 = ~w34475 & ~w34476;
assign w34478 = w5053 & w33821;
assign w34479 = ~pi3186 & pi3226;
assign w34480 = ~w33821 & w34479;
assign w34481 = ~w34478 & ~w34480;
assign w34482 = pi3187 & ~w33757;
assign w34483 = ~pi2064 & ~w34243;
assign w34484 = w33757 & w34483;
assign w34485 = ~w34482 & ~w34484;
assign w34486 = pi0854 & pi3188;
assign w34487 = w33479 & w34486;
assign w34488 = w6177 & w33821;
assign w34489 = ~pi3189 & pi3238;
assign w34490 = ~w33821 & w34489;
assign w34491 = ~w34488 & ~w34490;
assign w34492 = pi3190 & w6684;
assign w34493 = w32020 & w32389;
assign w34494 = ~w34492 & ~w34493;
assign w34495 = ~pi3191 & w6684;
assign w34496 = w21969 & w22005;
assign w34497 = ~w34495 & ~w34496;
assign w34498 = pi3192 & ~w33757;
assign w34499 = ~pi2038 & ~w34243;
assign w34500 = w33757 & w34499;
assign w34501 = ~w34498 & ~w34500;
assign w34502 = pi3193 & ~w33757;
assign w34503 = ~pi2039 & ~w34243;
assign w34504 = w33757 & w34503;
assign w34505 = ~w34502 & ~w34504;
assign w34506 = pi3194 & ~w33757;
assign w34507 = ~pi2042 & ~w34243;
assign w34508 = w33757 & w34507;
assign w34509 = ~w34506 & ~w34508;
assign w34510 = pi3195 & ~w33757;
assign w34511 = ~pi2050 & ~w34243;
assign w34512 = w33757 & w34511;
assign w34513 = ~w34510 & ~w34512;
assign w34514 = pi3196 & ~w33757;
assign w34515 = ~pi2043 & ~w34243;
assign w34516 = w33757 & w34515;
assign w34517 = ~w34514 & ~w34516;
assign w34518 = pi3197 & ~w33757;
assign w34519 = ~pi2044 & ~w34243;
assign w34520 = w33757 & w34519;
assign w34521 = ~w34518 & ~w34520;
assign w34522 = pi3198 & ~w33757;
assign w34523 = ~pi2060 & ~w34243;
assign w34524 = w33757 & w34523;
assign w34525 = ~w34522 & ~w34524;
assign w34526 = ~pi3199 & ~w30856;
assign w34527 = ~w30857 & ~w34526;
assign w34528 = ~w30853 & w34527;
assign w34529 = pi0856 & pi3200;
assign w34530 = w33479 & w34529;
assign w34531 = ~w30492 & w32801;
assign w34532 = pi3201 & ~w32801;
assign w34533 = ~w34531 & ~w34532;
assign w34534 = pi3202 & ~w34267;
assign w34535 = w40171 & w34267;
assign w34536 = ~w34534 & ~w34535;
assign w34537 = pi3510 & w27062;
assign w34538 = ~pi3203 & ~w34537;
assign w34539 = w25108 & w27062;
assign w34540 = ~w34538 & ~w34539;
assign w34541 = pi0615 & w23005;
assign w34542 = ~pi3204 & ~w34541;
assign w34543 = pi0785 & pi3205;
assign w34544 = w33479 & w34543;
assign w34545 = pi3206 & ~w33757;
assign w34546 = pi2034 & ~w34243;
assign w34547 = pi1954 & w34243;
assign w34548 = ~w34546 & ~w34547;
assign w34549 = w33757 & w34548;
assign w34550 = ~w34545 & ~w34549;
assign w34551 = pi3207 & ~w33757;
assign w34552 = pi2066 & ~w34243;
assign w34553 = pi2027 & w34243;
assign w34554 = ~w34552 & ~w34553;
assign w34555 = w33757 & w34554;
assign w34556 = ~w34551 & ~w34555;
assign w34557 = pi3208 & ~w33757;
assign w34558 = pi2036 & ~w34243;
assign w34559 = pi1970 & w34243;
assign w34560 = ~w34558 & ~w34559;
assign w34561 = w33757 & w34560;
assign w34562 = ~w34557 & ~w34561;
assign w34563 = pi3209 & ~w33757;
assign w34564 = pi2031 & ~w34243;
assign w34565 = pi2022 & w34243;
assign w34566 = ~w34564 & ~w34565;
assign w34567 = w33757 & w34566;
assign w34568 = ~w34563 & ~w34567;
assign w34569 = pi3210 & w6684;
assign w34570 = pi0408 & w32379;
assign w34571 = ~w34569 & ~w34570;
assign w34572 = ~pi3211 & w6684;
assign w34573 = ~w32379 & ~w34572;
assign w34574 = pi3212 & pi3488;
assign w34575 = pi3534 & ~w34574;
assign w34576 = ~pi3212 & ~pi3488;
assign w34577 = ~w34575 & ~w34576;
assign w34578 = pi3213 & pi3486;
assign w34579 = pi3532 & ~w34578;
assign w34580 = ~pi3213 & ~pi3486;
assign w34581 = ~w34579 & ~w34580;
assign w34582 = pi3214 & pi3485;
assign w34583 = pi3531 & ~w34582;
assign w34584 = ~pi3214 & ~pi3485;
assign w34585 = ~w34583 & ~w34584;
assign w34586 = w2246 & w22169;
assign w34587 = w361 & w34586;
assign w34588 = ~w6606 & w22169;
assign w34589 = w2361 & w34588;
assign w34590 = pi3215 & w343;
assign w34591 = ~w34589 & ~w34590;
assign w34592 = ~w34587 & w34591;
assign w34593 = pi3216 & w343;
assign w34594 = ~w21809 & w22169;
assign w34595 = ~w34593 & ~w34594;
assign w34596 = w6413 & w33821;
assign w34597 = pi3068 & ~pi3217;
assign w34598 = ~w33821 & w34597;
assign w34599 = ~w34596 & ~w34598;
assign w34600 = pi3998 & ~w26891;
assign w34601 = ~pi3325 & w34600;
assign w34602 = pi3218 & ~w34601;
assign w34603 = pi3325 & ~pi3998;
assign w34604 = ~w26891 & w34603;
assign w34605 = ~w34602 & ~w34604;
assign w34606 = pi4003 & ~w26497;
assign w34607 = ~pi3356 & w34606;
assign w34608 = pi3219 & ~w34607;
assign w34609 = pi3356 & ~pi4003;
assign w34610 = ~w26497 & w34609;
assign w34611 = ~w34608 & ~w34610;
assign w34612 = pi4001 & ~w26873;
assign w34613 = ~pi3341 & w34612;
assign w34614 = pi3220 & ~w34613;
assign w34615 = pi3341 & ~pi4001;
assign w34616 = ~w26873 & w34615;
assign w34617 = ~w34614 & ~w34616;
assign w34618 = pi3999 & ~w26882;
assign w34619 = ~pi3301 & w34618;
assign w34620 = pi3221 & ~w34619;
assign w34621 = pi3301 & ~pi3999;
assign w34622 = ~w26882 & w34621;
assign w34623 = ~w34620 & ~w34622;
assign w34624 = pi3997 & ~w26891;
assign w34625 = ~pi3327 & w34624;
assign w34626 = pi3222 & ~w34625;
assign w34627 = pi3327 & ~pi3997;
assign w34628 = ~w26891 & w34627;
assign w34629 = ~w34626 & ~w34628;
assign w34630 = pi3996 & ~w26900;
assign w34631 = ~pi3334 & w34630;
assign w34632 = pi3223 & ~w34631;
assign w34633 = pi3334 & ~pi3996;
assign w34634 = ~w26900 & w34633;
assign w34635 = ~w34632 & ~w34634;
assign w34636 = pi4006 & ~w26909;
assign w34637 = ~pi3335 & w34636;
assign w34638 = pi3224 & ~w34637;
assign w34639 = pi3335 & ~pi4006;
assign w34640 = ~w26909 & w34639;
assign w34641 = ~w34638 & ~w34640;
assign w34642 = pi3995 & ~w26900;
assign w34643 = ~pi3333 & w34642;
assign w34644 = pi3225 & ~w34643;
assign w34645 = pi3333 & ~pi3995;
assign w34646 = ~w26900 & w34645;
assign w34647 = ~w34644 & ~w34646;
assign w34648 = w5635 & w33821;
assign w34649 = pi3186 & ~pi3226;
assign w34650 = ~w33821 & w34649;
assign w34651 = ~w34648 & ~w34650;
assign w34652 = w4749 & w33821;
assign w34653 = pi2976 & ~pi3227;
assign w34654 = ~w33821 & w34653;
assign w34655 = ~w34652 & ~w34654;
assign w34656 = pi3228 & ~w33757;
assign w34657 = pi2032 & ~w34243;
assign w34658 = pi2023 & w34243;
assign w34659 = ~w34657 & ~w34658;
assign w34660 = w33757 & w34659;
assign w34661 = ~w34656 & ~w34660;
assign w34662 = pi3229 & ~w33757;
assign w34663 = pi1863 & ~w34243;
assign w34664 = pi2024 & w34243;
assign w34665 = ~w34663 & ~w34664;
assign w34666 = w33757 & w34665;
assign w34667 = ~w34662 & ~w34666;
assign w34668 = pi3230 & ~w33757;
assign w34669 = pi2033 & ~w34243;
assign w34670 = pi2025 & w34243;
assign w34671 = ~w34669 & ~w34670;
assign w34672 = w33757 & w34671;
assign w34673 = ~w34668 & ~w34672;
assign w34674 = pi3231 & ~w33757;
assign w34675 = pi1968 & ~w34243;
assign w34676 = pi2026 & w34243;
assign w34677 = ~w34675 & ~w34676;
assign w34678 = w33757 & w34677;
assign w34679 = ~w34674 & ~w34678;
assign w34680 = pi3232 & pi3487;
assign w34681 = pi3533 & ~w34680;
assign w34682 = ~pi3232 & ~pi3487;
assign w34683 = ~w34681 & ~w34682;
assign w34684 = ~pi3233 & w343;
assign w34685 = ~w23341 & ~w34684;
assign w34686 = pi3234 & ~w33757;
assign w34687 = pi2035 & ~w34243;
assign w34688 = pi1969 & w34243;
assign w34689 = ~w34687 & ~w34688;
assign w34690 = w33757 & w34689;
assign w34691 = ~w34686 & ~w34690;
assign w34692 = pi3235 & ~w33757;
assign w34693 = pi2063 & ~w34243;
assign w34694 = pi2028 & w34243;
assign w34695 = ~w34693 & ~w34694;
assign w34696 = w33757 & w34695;
assign w34697 = ~w34692 & ~w34696;
assign w34698 = pi3236 & w6684;
assign w34699 = w6682 & w6972;
assign w34700 = w30566 & w34699;
assign w34701 = ~w34698 & ~w34700;
assign w34702 = w3195 & w33821;
assign w34703 = pi2974 & ~pi3237;
assign w34704 = ~w33821 & w34703;
assign w34705 = ~w34702 & ~w34704;
assign w34706 = w4141 & w33821;
assign w34707 = pi3189 & ~pi3238;
assign w34708 = ~w33821 & w34707;
assign w34709 = ~w34706 & ~w34708;
assign w34710 = w5320 & w33821;
assign w34711 = pi2975 & ~pi3239;
assign w34712 = ~w33821 & w34711;
assign w34713 = ~w34710 & ~w34712;
assign w34714 = pi4005 & ~w26909;
assign w34715 = ~pi3336 & w34714;
assign w34716 = pi3240 & ~w34715;
assign w34717 = pi3336 & ~pi4005;
assign w34718 = ~w26909 & w34717;
assign w34719 = ~w34716 & ~w34718;
assign w34720 = pi4002 & ~w26873;
assign w34721 = ~pi3339 & w34720;
assign w34722 = pi3241 & ~w34721;
assign w34723 = pi3339 & ~pi4002;
assign w34724 = ~w26873 & w34723;
assign w34725 = ~w34722 & ~w34724;
assign w34726 = pi4000 & ~w26882;
assign w34727 = ~pi3338 & w34726;
assign w34728 = pi3242 & ~w34727;
assign w34729 = pi3338 & ~pi4000;
assign w34730 = ~w26882 & w34729;
assign w34731 = ~w34728 & ~w34730;
assign w34732 = pi4004 & ~w26497;
assign w34733 = ~pi3342 & w34732;
assign w34734 = pi3243 & ~w34733;
assign w34735 = pi3342 & ~pi4004;
assign w34736 = ~w26497 & w34735;
assign w34737 = ~w34734 & ~w34736;
assign w34738 = ~w343 & w21509;
assign w34739 = ~pi3244 & w343;
assign w34740 = ~w34738 & ~w34739;
assign w34741 = pi3245 & w6684;
assign w34742 = w6682 & w21792;
assign w34743 = ~w34741 & ~w34742;
assign w34744 = pi3425 & ~pi3502;
assign w34745 = ~pi3677 & w34744;
assign w34746 = pi3246 & ~w34745;
assign w34747 = pi3266 & w34745;
assign w34748 = ~w34746 & ~w34747;
assign w34749 = pi3247 & ~w27273;
assign w34750 = ~w32459 & ~w34749;
assign w34751 = ~pi0427 & ~w343;
assign w34752 = pi3248 & w343;
assign w34753 = ~w34751 & ~w34752;
assign w34754 = w17481 & ~w34753;
assign w34755 = pi3099 & ~pi3199;
assign w34756 = pi3585 & w34755;
assign w34757 = ~pi2049 & ~pi2759;
assign w34758 = w133 & w34757;
assign w34759 = w34756 & w34758;
assign w34760 = ~pi3994 & w33330;
assign w34761 = pi3253 & ~w33330;
assign w34762 = ~w34760 & ~w34761;
assign w34763 = pi3255 & ~w34745;
assign w34764 = pi3678 & w34745;
assign w34765 = ~w34763 & ~w34764;
assign w34766 = ~w2253 & ~w34586;
assign w34767 = ~w6608 & ~w34588;
assign w34768 = ~pi3692 & w33330;
assign w34769 = pi3258 & ~w33330;
assign w34770 = ~w34768 & ~w34769;
assign w34771 = ~pi3691 & w33330;
assign w34772 = pi3259 & ~w33330;
assign w34773 = ~w34771 & ~w34772;
assign w34774 = ~pi3686 & w33330;
assign w34775 = pi3260 & ~w33330;
assign w34776 = ~w34774 & ~w34775;
assign w34777 = ~pi3992 & w33330;
assign w34778 = pi3261 & ~w33330;
assign w34779 = ~w34777 & ~w34778;
assign w34780 = ~pi3684 & w33330;
assign w34781 = pi3262 & ~w33330;
assign w34782 = ~w34780 & ~w34781;
assign w34783 = ~pi3989 & w33330;
assign w34784 = pi3263 & ~w33330;
assign w34785 = ~w34783 & ~w34784;
assign w34786 = ~pi3987 & w33330;
assign w34787 = pi3264 & ~w33330;
assign w34788 = ~w34786 & ~w34787;
assign w34789 = ~pi3693 & w33330;
assign w34790 = pi3265 & ~w33330;
assign w34791 = ~w34789 & ~w34790;
assign w34792 = pi3266 & ~w34745;
assign w34793 = pi3271 & w34745;
assign w34794 = ~w34792 & ~w34793;
assign w34795 = ~pi0407 & ~w343;
assign w34796 = pi3267 & w343;
assign w34797 = ~w34795 & ~w34796;
assign w34798 = w17481 & ~w34797;
assign w34799 = pi3268 & w6684;
assign w34800 = pi2193 & w21968;
assign w34801 = ~w34799 & ~w34800;
assign w34802 = pi3269 & ~w23792;
assign w34803 = ~pi2402 & w27127;
assign w34804 = ~w34802 & ~w34803;
assign w34805 = ~pi3424 & ~pi3639;
assign w34806 = ~pi3588 & pi3647;
assign w34807 = ~w27425 & w34806;
assign w34808 = pi1735 & w34807;
assign w34809 = pi3270 & ~w34808;
assign w34810 = pi3271 & ~w34745;
assign w34811 = pi3255 & w34745;
assign w34812 = ~w34810 & ~w34811;
assign w34813 = ~pi3993 & w33330;
assign w34814 = pi3272 & ~w33330;
assign w34815 = ~w34813 & ~w34814;
assign w34816 = ~pi3990 & w33330;
assign w34817 = pi3273 & ~w33330;
assign w34818 = ~w34816 & ~w34817;
assign w34819 = ~pi3698 & w33330;
assign w34820 = pi3274 & ~w33330;
assign w34821 = ~w34819 & ~w34820;
assign w34822 = ~pi3695 & w33330;
assign w34823 = pi3275 & ~w33330;
assign w34824 = ~w34822 & ~w34823;
assign w34825 = ~pi3694 & w33330;
assign w34826 = pi3276 & ~w33330;
assign w34827 = ~w34825 & ~w34826;
assign w34828 = ~pi3683 & w33330;
assign w34829 = pi3277 & ~w33330;
assign w34830 = ~w34828 & ~w34829;
assign w34831 = ~pi3427 & ~pi3638;
assign w34832 = ~pi3554 & pi3635;
assign w34833 = ~w28384 & w34832;
assign w34834 = pi1444 & w34833;
assign w34835 = pi3278 & ~w34834;
assign w34836 = ~pi3696 & w33330;
assign w34837 = pi3279 & ~w33330;
assign w34838 = ~w34836 & ~w34837;
assign w34839 = ~pi3697 & w33330;
assign w34840 = pi3280 & ~w33330;
assign w34841 = ~w34839 & ~w34840;
assign w34842 = pi3343 & w30855;
assign w34843 = ~pi3281 & ~w34842;
assign w34844 = ~w30856 & ~w34843;
assign w34845 = ~w30853 & w34844;
assign w34846 = ~pi3988 & w33330;
assign w34847 = pi3282 & ~w33330;
assign w34848 = ~w34846 & ~w34847;
assign w34849 = ~pi3991 & w33330;
assign w34850 = pi3283 & ~w33330;
assign w34851 = ~w34849 & ~w34850;
assign w34852 = ~pi3685 & w33330;
assign w34853 = pi3284 & ~w33330;
assign w34854 = ~w34852 & ~w34853;
assign w34855 = pi1798 & w29570;
assign w34856 = w29573 & w34855;
assign w34857 = ~pi3285 & ~w34856;
assign w34858 = ~pi3690 & w33330;
assign w34859 = pi3286 & ~w33330;
assign w34860 = ~w34858 & ~w34859;
assign w34861 = ~pi3689 & w33330;
assign w34862 = pi3287 & ~w33330;
assign w34863 = ~w34861 & ~w34862;
assign w34864 = ~pi3687 & w33330;
assign w34865 = pi3288 & ~w33330;
assign w34866 = ~w34864 & ~w34865;
assign w34867 = ~pi3688 & w33330;
assign w34868 = pi3289 & ~w33330;
assign w34869 = ~w34867 & ~w34868;
assign w34870 = pi3290 & ~w27272;
assign w34871 = ~w27273 & ~w34870;
assign w34872 = pi3291 & w6683;
assign w34873 = ~pi1823 & w6682;
assign w34874 = w19964 & w34873;
assign w34875 = ~w34872 & ~w34874;
assign w34876 = ~w343 & w21524;
assign w34877 = ~pi3292 & w343;
assign w34878 = ~w34876 & ~w34877;
assign w34879 = ~pi0834 & ~w370;
assign w34880 = pi3293 & ~w34879;
assign w34881 = w4380 & w34879;
assign w34882 = ~w34880 & ~w34881;
assign w34883 = w358 & ~w370;
assign w34884 = ~pi3295 & ~w34883;
assign w34885 = ~pi3216 & ~w5630;
assign w34886 = pi3216 & w7824;
assign w34887 = w34883 & ~w34886;
assign w34888 = ~w34885 & w34887;
assign w34889 = ~w34884 & ~w34888;
assign w34890 = ~pi3296 & ~w34883;
assign w34891 = ~pi3216 & ~w1303;
assign w34892 = pi3216 & w7856;
assign w34893 = w34883 & ~w34892;
assign w34894 = ~w34891 & w34893;
assign w34895 = ~w34890 & ~w34894;
assign w34896 = ~pi3297 & ~w34883;
assign w34897 = ~pi3216 & ~w5893;
assign w34898 = pi3216 & w7533;
assign w34899 = w34883 & ~w34898;
assign w34900 = ~w34897 & w34899;
assign w34901 = ~w34896 & ~w34900;
assign w34902 = ~pi3298 & ~w34883;
assign w34903 = ~pi3216 & ~w3411;
assign w34904 = pi3216 & w7664;
assign w34905 = w34883 & ~w34904;
assign w34906 = ~w34903 & w34905;
assign w34907 = ~w34902 & ~w34906;
assign w34908 = ~pi0415 & ~w343;
assign w34909 = ~pi3299 & w343;
assign w34910 = w17481 & ~w34909;
assign w34911 = ~w34908 & w34910;
assign w34912 = ~pi3301 & w26882;
assign w34913 = ~w34618 & ~w34912;
assign w34914 = pi3647 & w32660;
assign w34915 = pi0890 & pi1931;
assign w34916 = pi3569 & w34915;
assign w34917 = pi3270 & ~w34916;
assign w34918 = ~pi0418 & w7238;
assign w34919 = pi3305 & w343;
assign w34920 = ~w34918 & ~w34919;
assign w34921 = ~pi3306 & ~w34883;
assign w34922 = ~pi3216 & ~w4136;
assign w34923 = pi3216 & w7760;
assign w34924 = w34883 & ~w34923;
assign w34925 = ~w34922 & w34924;
assign w34926 = ~w34921 & ~w34925;
assign w34927 = ~pi3307 & ~w34883;
assign w34928 = ~pi3216 & ~w6172;
assign w34929 = pi3216 & w7728;
assign w34930 = w34883 & ~w34929;
assign w34931 = ~w34928 & w34930;
assign w34932 = ~w34927 & ~w34931;
assign w34933 = ~pi3308 & ~w34883;
assign w34934 = ~pi3216 & ~w3190;
assign w34935 = pi3216 & w7696;
assign w34936 = w34883 & ~w34935;
assign w34937 = ~w34934 & w34936;
assign w34938 = ~w34933 & ~w34937;
assign w34939 = pi3309 & ~w34883;
assign w34940 = ~pi3216 & w6351;
assign w34941 = ~w941 & ~w34940;
assign w34942 = ~w6409 & ~w34941;
assign w34943 = pi3216 & ~w7631;
assign w34944 = w34883 & ~w34943;
assign w34945 = ~w34942 & w34944;
assign w34946 = ~w34939 & ~w34945;
assign w34947 = ~pi3310 & ~w34883;
assign w34948 = ~pi3216 & ~w4375;
assign w34949 = pi3216 & w7598;
assign w34950 = w34883 & ~w34949;
assign w34951 = ~w34948 & w34950;
assign w34952 = ~w34947 & ~w34951;
assign w34953 = ~pi3311 & ~w34883;
assign w34954 = ~pi3216 & ~w5315;
assign w34955 = pi3216 & w7566;
assign w34956 = w34883 & ~w34955;
assign w34957 = ~w34954 & w34956;
assign w34958 = ~w34953 & ~w34957;
assign w34959 = ~pi3312 & ~w34883;
assign w34960 = ~pi3216 & ~w4743;
assign w34961 = pi3216 & w7501;
assign w34962 = w34883 & ~w34961;
assign w34963 = ~w34960 & w34962;
assign w34964 = ~w34959 & ~w34963;
assign w34965 = pi3313 & ~w34883;
assign w34966 = ~pi3216 & w8235;
assign w34967 = pi3216 & ~w8262;
assign w34968 = w34883 & ~w34967;
assign w34969 = ~w34966 & w34968;
assign w34970 = ~w34965 & ~w34969;
assign w34971 = pi3314 & ~w34883;
assign w34972 = ~pi3216 & w8077;
assign w34973 = pi3216 & ~w7990;
assign w34974 = w34883 & ~w34973;
assign w34975 = ~w34972 & w34974;
assign w34976 = ~w34971 & ~w34975;
assign w34977 = ~pi3315 & ~w34883;
assign w34978 = ~pi3216 & ~w5048;
assign w34979 = pi3216 & w7792;
assign w34980 = w34883 & ~w34979;
assign w34981 = ~w34978 & w34980;
assign w34982 = ~w34977 & ~w34981;
assign w34983 = ~pi3316 & ~w34883;
assign w34984 = ~pi3216 & ~w3706;
assign w34985 = pi3216 & w7424;
assign w34986 = w34883 & ~w34985;
assign w34987 = ~w34984 & w34986;
assign w34988 = ~w34983 & ~w34987;
assign w34989 = pi3243 & ~w26497;
assign w34990 = pi3317 & w26497;
assign w34991 = ~w34989 & ~w34990;
assign w34992 = pi3219 & ~w26497;
assign w34993 = pi3318 & w26497;
assign w34994 = ~w34992 & ~w34993;
assign w34995 = pi3222 & ~w26891;
assign w34996 = pi3319 & w26891;
assign w34997 = ~w34995 & ~w34996;
assign w34998 = pi3223 & ~w26900;
assign w34999 = pi3320 & w26900;
assign w35000 = ~w34998 & ~w34999;
assign w35001 = pi3225 & ~w26900;
assign w35002 = pi3321 & w26900;
assign w35003 = ~w35001 & ~w35002;
assign w35004 = ~pi3325 & w26891;
assign w35005 = ~w34600 & ~w35004;
assign w35006 = pi0414 & ~w343;
assign w35007 = pi3326 & w343;
assign w35008 = ~w35006 & ~w35007;
assign w35009 = w17481 & ~w35008;
assign w35010 = ~pi3327 & w26891;
assign w35011 = ~w34624 & ~w35010;
assign w35012 = pi3328 & ~w34879;
assign w35013 = w5914 & w34879;
assign w35014 = ~w35012 & ~w35013;
assign w35015 = pi3329 & w343;
assign w35016 = pi0419 & ~w343;
assign w35017 = w14358 & w35016;
assign w35018 = ~w35015 & ~w35017;
assign w35019 = ~pi3330 & w343;
assign w35020 = ~w34795 & ~w35019;
assign w35021 = pi1930 & ~w370;
assign w35022 = pi3331 & ~w35021;
assign w35023 = pi3402 & w35021;
assign w35024 = ~w35022 & ~w35023;
assign w35025 = pi3332 & ~w35021;
assign w35026 = pi3400 & w35021;
assign w35027 = ~w35025 & ~w35026;
assign w35028 = ~pi3333 & w26900;
assign w35029 = ~w34642 & ~w35028;
assign w35030 = ~pi3334 & w26900;
assign w35031 = ~w34630 & ~w35030;
assign w35032 = ~pi3335 & w26909;
assign w35033 = ~w34636 & ~w35032;
assign w35034 = ~pi3336 & w26909;
assign w35035 = ~w34714 & ~w35034;
assign w35036 = pi3337 & pi3389;
assign w35037 = ~pi3338 & w26882;
assign w35038 = ~w34726 & ~w35037;
assign w35039 = ~pi3339 & w26873;
assign w35040 = ~w34720 & ~w35039;
assign w35041 = pi3240 & ~w26909;
assign w35042 = pi3340 & w26909;
assign w35043 = ~w35041 & ~w35042;
assign w35044 = ~pi3341 & w26873;
assign w35045 = ~w34612 & ~w35044;
assign w35046 = ~pi3342 & w26497;
assign w35047 = ~w34732 & ~w35046;
assign w35048 = ~pi3343 & ~w30855;
assign w35049 = ~w34842 & ~w35048;
assign w35050 = ~w30853 & w35049;
assign w35051 = pi3344 & w6684;
assign w35052 = ~w22336 & ~w35051;
assign w35053 = pi3221 & ~w26882;
assign w35054 = pi3345 & w26882;
assign w35055 = ~w35053 & ~w35054;
assign w35056 = pi3242 & ~w26882;
assign w35057 = pi3346 & w26882;
assign w35058 = ~w35056 & ~w35057;
assign w35059 = pi3347 & ~w35021;
assign w35060 = pi3403 & w35021;
assign w35061 = ~w35059 & ~w35060;
assign w35062 = pi3218 & ~w26891;
assign w35063 = pi3348 & w26891;
assign w35064 = ~w35062 & ~w35063;
assign w35065 = pi3220 & ~w26873;
assign w35066 = pi3349 & w26873;
assign w35067 = ~w35065 & ~w35066;
assign w35068 = w165 & w33326;
assign w35069 = w33328 & w35068;
assign w35070 = pi3682 & w105;
assign w35071 = w170 & w35070;
assign w35072 = pi3350 & ~w35071;
assign w35073 = ~w35069 & ~w35072;
assign w35074 = pi3241 & ~w26873;
assign w35075 = pi3351 & w26873;
assign w35076 = ~w35074 & ~w35075;
assign w35077 = pi3352 & ~w35021;
assign w35078 = pi3404 & w35021;
assign w35079 = ~w35077 & ~w35078;
assign w35080 = pi3353 & ~w35021;
assign w35081 = ~w9819 & w35021;
assign w35082 = ~w35080 & ~w35081;
assign w35083 = pi3354 & ~w35021;
assign w35084 = pi3414 & w35021;
assign w35085 = ~w35083 & ~w35084;
assign w35086 = pi3355 & ~w35021;
assign w35087 = ~w9817 & w35021;
assign w35088 = ~w35086 & ~w35087;
assign w35089 = ~pi3356 & w26497;
assign w35090 = ~w34606 & ~w35089;
assign w35091 = pi3224 & ~w26909;
assign w35092 = pi3357 & w26909;
assign w35093 = ~w35091 & ~w35092;
assign w35094 = ~pi3358 & ~w34883;
assign w35095 = ~pi3216 & ~w1617;
assign w35096 = pi3216 & w7888;
assign w35097 = w34883 & ~w35096;
assign w35098 = ~w35095 & w35097;
assign w35099 = ~w35094 & ~w35098;
assign w35100 = w6615 & ~w6652;
assign w35101 = w6655 & w35100;
assign w35102 = pi3360 & ~w34879;
assign w35103 = w4749 & w34879;
assign w35104 = ~w35102 & ~w35103;
assign w35105 = pi3361 & ~w34879;
assign w35106 = w3711 & w34879;
assign w35107 = ~w35105 & ~w35106;
assign w35108 = w6615 & w6652;
assign w35109 = w6661 & w35108;
assign w35110 = w6661 & w35100;
assign w35111 = w6663 & w35100;
assign w35112 = ~w1657 & ~w2256;
assign w35113 = w2267 & w35112;
assign w35114 = w1338 & w35113;
assign w35115 = ~w343 & w416;
assign w35116 = pi3367 & w343;
assign w35117 = ~w35115 & ~w35116;
assign w35118 = w1351 & w35112;
assign w35119 = w2276 & w35118;
assign w35120 = w2273 & w35112;
assign w35121 = w1338 & w35120;
assign w35122 = ~pi3481 & w2260;
assign w35123 = pi3216 & ~w370;
assign w35124 = ~w35122 & ~w35123;
assign w35125 = ~pi0540 & ~w370;
assign w35126 = ~pi3371 & w370;
assign w35127 = w6682 & ~w35126;
assign w35128 = ~w35125 & w35127;
assign w35129 = w8081 & w33821;
assign w35130 = w1639 & w33821;
assign w35131 = w1308 & w33821;
assign w35132 = w8240 & w33821;
assign w35133 = pi0796 & pi2111;
assign w35134 = pi3570 & w35133;
assign w35135 = pi3278 & ~w35134;
assign w35136 = pi0491 & pi3377;
assign w35137 = ~pi1771 & w21341;
assign w35138 = ~w35136 & ~w35137;
assign w35139 = pi2789 & ~w370;
assign w35140 = ~pi3481 & w6622;
assign w35141 = ~w35139 & ~w35140;
assign w35142 = w2276 & w35120;
assign w35143 = w2270 & w35112;
assign w35144 = w2276 & w35143;
assign w35145 = w2276 & w35113;
assign w35146 = w0 & w32393;
assign w35147 = pi3382 & ~pi3410;
assign w35148 = pi3481 & ~w35147;
assign w35149 = w1338 & w35143;
assign w35150 = w1338 & w35118;
assign w35151 = w6663 & w35108;
assign w35152 = w6646 & w35100;
assign w35153 = w6655 & w35108;
assign w35154 = ~w3817 & w6615;
assign w35155 = ~w6599 & w35154;
assign w35156 = pi3337 & ~pi3389;
assign w35157 = pi3390 & w343;
assign w35158 = ~w7238 & ~w35157;
assign w35159 = ~w343 & w408;
assign w35160 = pi3391 & w343;
assign w35161 = ~w35159 & ~w35160;
assign w35162 = ~pi3392 & w343;
assign w35163 = ~w34908 & ~w35162;
assign w35164 = pi3393 & w343;
assign w35165 = ~w35016 & ~w35164;
assign w35166 = ~pi3394 & w343;
assign w35167 = ~w34751 & ~w35166;
assign w35168 = ~pi3395 & w8407;
assign w35169 = pi0420 & ~w343;
assign w35170 = pi3396 & w343;
assign w35171 = ~w35169 & ~w35170;
assign w35172 = ~pi3583 & w27271;
assign w35173 = ~w32398 & ~w35172;
assign w35174 = pi3398 & w343;
assign w35175 = ~w35006 & ~w35174;
assign w35176 = w6646 & w35108;
assign w35177 = pi3400 & w342;
assign w35178 = pi2516 & ~w342;
assign w35179 = ~w35177 & ~w35178;
assign w35180 = pi3401 & w342;
assign w35181 = pi2517 & ~w342;
assign w35182 = ~w35180 & ~w35181;
assign w35183 = pi3402 & w342;
assign w35184 = pi2482 & ~w342;
assign w35185 = ~w35183 & ~w35184;
assign w35186 = pi3403 & w342;
assign w35187 = pi2483 & ~w342;
assign w35188 = ~w35186 & ~w35187;
assign w35189 = pi3404 & w342;
assign w35190 = pi2481 & ~w342;
assign w35191 = ~w35189 & ~w35190;
assign w35192 = pi3405 & w342;
assign w35193 = pi2479 & ~w342;
assign w35194 = ~w35192 & ~w35193;
assign w35195 = pi3406 & w342;
assign w35196 = pi2477 & ~w342;
assign w35197 = ~w35195 & ~w35196;
assign w35198 = pi3407 & ~w34879;
assign w35199 = ~w370 & w2227;
assign w35200 = pi3408 & w370;
assign w35201 = ~w35199 & ~w35200;
assign w35202 = ~pi0783 & ~w6682;
assign w35203 = w10741 & ~w35202;
assign w35204 = pi3411 & w342;
assign w35205 = pi2476 & ~w342;
assign w35206 = ~w35204 & ~w35205;
assign w35207 = ~pi3412 & w370;
assign w35208 = ~w361 & ~w2361;
assign w35209 = ~w370 & w35208;
assign w35210 = ~w35207 & ~w35209;
assign w35211 = pi3413 & w342;
assign w35212 = pi2478 & ~w342;
assign w35213 = ~w35211 & ~w35212;
assign w35214 = pi3414 & w342;
assign w35215 = pi2480 & ~w342;
assign w35216 = ~w35214 & ~w35215;
assign w35217 = pi2492 & ~pi3415;
assign w35218 = ~pi0936 & pi3415;
assign w35219 = ~w35217 & ~w35218;
assign w35220 = ~pi3398 & w6692;
assign w35221 = w6676 & w35220;
assign w35222 = pi3481 & w336;
assign w35223 = ~w35221 & ~w35222;
assign w35224 = ~pi3419 & w889;
assign w35225 = ~w350 & w35224;
assign w35226 = pi3420 & w342;
assign w35227 = pi2475 & ~w342;
assign w35228 = ~w35226 & ~w35227;
assign w35229 = pi3421 & w342;
assign w35230 = pi2485 & ~w342;
assign w35231 = ~w35229 & ~w35230;
assign w35232 = pi3422 & w342;
assign w35233 = pi2518 & ~w342;
assign w35234 = ~w35232 & ~w35233;
assign w35235 = ~pi1930 & ~pi3423;
assign w35236 = pi1930 & ~w9853;
assign w35237 = ~w9929 & w35236;
assign w35238 = ~w35235 & ~w35237;
assign w35239 = ~pi3424 & w828;
assign w35240 = ~w8406 & w35239;
assign w35241 = w0 & w24174;
assign w35242 = ~pi3426 & w343;
assign w35243 = ~w22169 & ~w35242;
assign w35244 = ~pi3427 & w830;
assign w35245 = ~w8406 & w35244;
assign w35246 = pi3641 & w350;
assign w35247 = pi3428 & w938;
assign w35248 = ~w35246 & w35247;
assign w35249 = ~pi3429 & w8409;
assign w35250 = pi3430 & w342;
assign w35251 = pi2484 & ~w342;
assign w35252 = ~w35250 & ~w35251;
assign w35253 = ~w6683 & w9553;
assign w35254 = ~pi3432 & w6683;
assign w35255 = ~w35253 & ~w35254;
assign w35256 = ~w6683 & w9349;
assign w35257 = ~pi3434 & w6683;
assign w35258 = ~w35256 & ~w35257;
assign w35259 = w358 & ~w839;
assign w35260 = pi3435 & ~w358;
assign w35261 = ~w35259 & ~w35260;
assign w35262 = w358 & ~w833;
assign w35263 = pi3436 & ~w358;
assign w35264 = ~w35262 & ~w35263;
assign w35265 = pi1908 & pi2492;
assign w35266 = pi3415 & w35265;
assign w35267 = ~pi3674 & pi3708;
assign w35268 = ~pi3445 & pi3674;
assign w35269 = ~w35267 & ~w35268;
assign w35270 = ~pi3674 & pi3702;
assign w35271 = ~pi3446 & pi3674;
assign w35272 = ~w35270 & ~w35271;
assign w35273 = ~pi3674 & pi3711;
assign w35274 = ~pi3447 & pi3674;
assign w35275 = ~w35273 & ~w35274;
assign w35276 = ~pi3674 & pi3709;
assign w35277 = ~pi3448 & pi3674;
assign w35278 = ~w35276 & ~w35277;
assign w35279 = ~w7107 & w35069;
assign w35280 = pi3449 & ~w35069;
assign w35281 = ~w35279 & ~w35280;
assign w35282 = ~w6683 & w7095;
assign w35283 = ~pi3450 & w6683;
assign w35284 = ~w35282 & ~w35283;
assign w35285 = w358 & ~w864;
assign w35286 = pi3451 & ~w358;
assign w35287 = ~w35285 & ~w35286;
assign w35288 = w28741 & w34363;
assign w35289 = ~w6683 & w9507;
assign w35290 = ~pi3453 & w6683;
assign w35291 = ~w35289 & ~w35290;
assign w35292 = ~w6683 & w9445;
assign w35293 = ~pi3454 & w6683;
assign w35294 = ~w35292 & ~w35293;
assign w35295 = ~w6683 & w9394;
assign w35296 = ~pi3455 & w6683;
assign w35297 = ~w35295 & ~w35296;
assign w35298 = ~w6683 & w7156;
assign w35299 = ~pi3458 & w6683;
assign w35300 = ~w35298 & ~w35299;
assign w35301 = ~w6683 & w9606;
assign w35302 = ~pi3459 & w6683;
assign w35303 = ~w35301 & ~w35302;
assign w35304 = pi2576 & ~w27430;
assign w35305 = pi3473 & w27430;
assign w35306 = ~w35304 & ~w35305;
assign w35307 = ~pi3674 & pi3701;
assign w35308 = ~pi3462 & pi3674;
assign w35309 = ~w35307 & ~w35308;
assign w35310 = ~pi3674 & pi3710;
assign w35311 = ~pi3463 & pi3674;
assign w35312 = ~w35310 & ~w35311;
assign w35313 = ~pi3674 & pi3699;
assign w35314 = ~pi3464 & pi3674;
assign w35315 = ~w35313 & ~w35314;
assign w35316 = ~pi3674 & pi3713;
assign w35317 = ~pi3465 & pi3674;
assign w35318 = ~w35316 & ~w35317;
assign w35319 = ~pi3674 & pi3712;
assign w35320 = ~pi3466 & pi3674;
assign w35321 = ~w35319 & ~w35320;
assign w35322 = ~pi3674 & pi3714;
assign w35323 = ~pi3467 & pi3674;
assign w35324 = ~w35322 & ~w35323;
assign w35325 = ~pi3674 & pi3700;
assign w35326 = ~pi3468 & pi3674;
assign w35327 = ~w35325 & ~w35326;
assign w35328 = ~pi3674 & pi3703;
assign w35329 = ~pi3470 & pi3674;
assign w35330 = ~w35328 & ~w35329;
assign w35331 = ~pi3597 & w27430;
assign w35332 = pi2578 & ~w27430;
assign w35333 = ~w35331 & ~w35332;
assign w35334 = pi2577 & ~w27430;
assign w35335 = pi3471 & w27430;
assign w35336 = ~w35334 & ~w35335;
assign w35337 = ~pi3674 & pi3707;
assign w35338 = ~pi3474 & pi3674;
assign w35339 = ~w35337 & ~w35338;
assign w35340 = ~pi3674 & pi3704;
assign w35341 = ~pi3475 & pi3674;
assign w35342 = ~w35340 & ~w35341;
assign w35343 = ~pi3674 & pi3705;
assign w35344 = ~pi3476 & pi3674;
assign w35345 = ~w35343 & ~w35344;
assign w35346 = ~pi3674 & pi3706;
assign w35347 = ~pi3477 & pi3674;
assign w35348 = ~w35346 & ~w35347;
assign w35349 = ~w6683 & w9666;
assign w35350 = ~pi3478 & w6683;
assign w35351 = ~w35349 & ~w35350;
assign w35352 = w6682 & w10741;
assign w35353 = ~pi3505 & ~pi3524;
assign w35354 = pi3515 & ~w35353;
assign w35355 = ~w9406 & w35069;
assign w35356 = pi3489 & ~w35069;
assign w35357 = ~w35355 & ~w35356;
assign w35358 = ~w9565 & w35069;
assign w35359 = pi3491 & ~w35069;
assign w35360 = ~w35358 & ~w35359;
assign w35361 = ~w9457 & w35069;
assign w35362 = pi3492 & ~w35069;
assign w35363 = ~w35361 & ~w35362;
assign w35364 = ~w9618 & w35069;
assign w35365 = pi3494 & ~w35069;
assign w35366 = ~w35364 & ~w35365;
assign w35367 = ~w9195 & w35069;
assign w35368 = pi3495 & ~w35069;
assign w35369 = ~w35367 & ~w35368;
assign w35370 = ~w9077 & w35069;
assign w35371 = pi3496 & ~w35069;
assign w35372 = ~w35370 & ~w35371;
assign w35373 = ~w9135 & w35069;
assign w35374 = pi3497 & ~w35069;
assign w35375 = ~w35373 & ~w35374;
assign w35376 = ~w9678 & w35069;
assign w35377 = pi3498 & ~w35069;
assign w35378 = ~w35376 & ~w35377;
assign w35379 = ~w9313 & w35069;
assign w35380 = pi3499 & ~w35069;
assign w35381 = ~w35379 & ~w35380;
assign w35382 = ~w9252 & w35069;
assign w35383 = pi3500 & ~w35069;
assign w35384 = ~w35382 & ~w35383;
assign w35385 = ~w9519 & w35069;
assign w35386 = pi3501 & ~w35069;
assign w35387 = ~w35385 & ~w35386;
assign w35388 = w24177 & ~w26311;
assign w35389 = w0 & ~w35388;
assign w35390 = ~w9361 & w35069;
assign w35391 = pi3503 & ~w35069;
assign w35392 = ~w35390 & ~w35391;
assign w35393 = w0 & w26312;
assign w35394 = ~pi3673 & ~pi3674;
assign w35395 = ~w113 & ~w177;
assign w35396 = ~pi3593 & w28389;
assign w35397 = pi1897 & ~w28389;
assign w35398 = ~w35396 & ~w35397;
assign w35399 = pi1866 & ~w28389;
assign w35400 = pi3594 & w28389;
assign w35401 = ~w35399 & ~w35400;
assign w35402 = pi1743 & ~w28389;
assign w35403 = pi3595 & w28389;
assign w35404 = ~w35402 & ~w35403;
assign w35405 = pi1744 & ~w28389;
assign w35406 = pi3596 & w28389;
assign w35407 = ~w35405 & ~w35406;
assign w35408 = pi1714 & ~w28389;
assign w35409 = pi3598 & w28389;
assign w35410 = ~w35408 & ~w35409;
assign w35411 = pi2579 & ~w27430;
assign w35412 = pi3600 & w27430;
assign w35413 = ~w35411 & ~w35412;
assign w35414 = pi1745 & ~w28389;
assign w35415 = pi3599 & w28389;
assign w35416 = ~w35414 & ~w35415;
assign w35417 = pi1742 & ~w28389;
assign w35418 = pi3601 & w28389;
assign w35419 = ~w35417 & ~w35418;
assign w35420 = pi2580 & ~w27430;
assign w35421 = pi3602 & w27430;
assign w35422 = ~w35420 & ~w35421;
assign w35423 = pi1741 & ~w28389;
assign w35424 = pi3603 & w28389;
assign w35425 = ~w35423 & ~w35424;
assign w35426 = pi2581 & ~w27430;
assign w35427 = pi3604 & w27430;
assign w35428 = ~w35426 & ~w35427;
assign w35429 = pi1867 & ~w28389;
assign w35430 = pi3605 & w28389;
assign w35431 = ~w35429 & ~w35430;
assign w35432 = pi2768 & ~w27430;
assign w35433 = pi3606 & w27430;
assign w35434 = ~w35432 & ~w35433;
assign w35435 = pi0368 & ~w28389;
assign w35436 = pi3607 & w28389;
assign w35437 = ~w35435 & ~w35436;
assign w35438 = pi2568 & ~w27430;
assign w35439 = pi3608 & w27430;
assign w35440 = ~w35438 & ~w35439;
assign w35441 = pi0314 & ~w28389;
assign w35442 = pi3609 & w28389;
assign w35443 = ~w35441 & ~w35442;
assign w35444 = pi2569 & ~w27430;
assign w35445 = pi3610 & w27430;
assign w35446 = ~w35444 & ~w35445;
assign w35447 = pi0330 & ~w28389;
assign w35448 = pi3611 & w28389;
assign w35449 = ~w35447 & ~w35448;
assign w35450 = pi2570 & ~w27430;
assign w35451 = pi3612 & w27430;
assign w35452 = ~w35450 & ~w35451;
assign w35453 = pi0072 & ~w28389;
assign w35454 = pi3613 & w28389;
assign w35455 = ~w35453 & ~w35454;
assign w35456 = pi2571 & ~w27430;
assign w35457 = pi3614 & w27430;
assign w35458 = ~w35456 & ~w35457;
assign w35459 = pi0127 & ~w28389;
assign w35460 = pi3615 & w28389;
assign w35461 = ~w35459 & ~w35460;
assign w35462 = pi2572 & ~w27430;
assign w35463 = pi3616 & w27430;
assign w35464 = ~w35462 & ~w35463;
assign w35465 = pi0073 & ~w28389;
assign w35466 = pi3618 & w28389;
assign w35467 = ~w35465 & ~w35466;
assign w35468 = pi2573 & ~w27430;
assign w35469 = pi3617 & w27430;
assign w35470 = ~w35468 & ~w35469;
assign w35471 = pi2574 & ~w27430;
assign w35472 = pi3619 & w27430;
assign w35473 = ~w35471 & ~w35472;
assign w35474 = pi0128 & ~w28389;
assign w35475 = pi2575 & ~w27430;
assign w35476 = pi3623 & w27430;
assign w35477 = ~w35475 & ~w35476;
assign w35478 = ~w113 & ~w33326;
assign w35479 = w30852 & w35478;
assign w35480 = ~w33324 & ~w35479;
assign w35481 = w187 & ~w35480;
assign w35482 = ~w116 & ~w184;
assign w35483 = pi3216 & ~w35482;
assign w35484 = ~pi2789 & ~pi2795;
assign w35485 = w178 & ~w35484;
assign w35486 = w12 & w179;
assign w35487 = ~w35484 & w35486;
assign w35488 = ~w35485 & ~w35487;
assign w35489 = ~w35483 & w35488;
assign w35490 = ~w35481 & w35489;
assign w35491 = w178 & ~w33340;
assign w35492 = ~pi3099 & w35395;
assign w35493 = w35068 & w35492;
assign w35494 = ~w35491 & ~w35493;
assign w35495 = pi3256 & w184;
assign w35496 = ~w187 & w35479;
assign w35497 = ~w35495 & ~w35496;
assign w35498 = w35494 & w35497;
assign w35499 = w187 & w35479;
assign w35500 = pi3216 & w184;
assign w35501 = ~w35485 & ~w35500;
assign w35502 = ~w35499 & w35501;
assign w35503 = pi2582 & ~w27430;
assign w35504 = pi0565 & pi3362;
assign w35505 = ~pi2813 & pi3528;
assign w35506 = ~w35504 & ~w35505;
assign w35507 = ~w918 & w35506;
assign w35508 = w28742 & w35507;
assign w35509 = ~w28744 & ~w35508;
assign w35510 = w6684 & w35509;
assign w35511 = ~pi2143 & w17481;
assign w35512 = ~pi0082 & ~pi0083;
assign w35513 = ~pi0084 & w35512;
assign w35514 = ~pi0043 & ~pi0044;
assign w35515 = ~pi0048 & ~pi0057;
assign w35516 = ~pi0060 & ~pi0061;
assign w35517 = w35515 & w35516;
assign w35518 = w35514 & w35517;
assign w35519 = w35513 & w35518;
assign w35520 = pi0082 & pi0083;
assign w35521 = pi0084 & w35520;
assign w35522 = pi0043 & pi0044;
assign w35523 = pi0048 & pi0057;
assign w35524 = pi0060 & pi0061;
assign w35525 = w35523 & w35524;
assign w35526 = w35522 & w35525;
assign w35527 = w35521 & w35526;
assign w35528 = pi3138 & ~w35527;
assign w35529 = ~w35519 & w35528;
assign w35530 = ~pi1025 & ~w35529;
assign w35531 = w17481 & ~w35530;
assign w35532 = ~pi3672 & ~pi3674;
assign w35533 = pi0939 & pi1609;
assign w35534 = w2 & ~w8;
assign w35535 = w20 & pi2825;
assign w35536 = w26 & ~pi2114;
assign w35537 = pi2799 & ~pi1462;
assign w35538 = ~w20 & ~pi2825;
assign w35539 = w41 & ~pi2114;
assign w35540 = ~pi2114 & ~pi1929;
assign w35541 = w51 & ~pi2114;
assign w35542 = pi1944 & ~w53;
assign w35543 = ~w60 & ~pi2082;
assign w35544 = w66 & pi2113;
assign w35545 = w60 & pi2082;
assign w35546 = ~w66 & ~pi2113;
assign w35547 = ~w40 & w14;
assign w35548 = w96 & w19;
assign w35549 = ~w91 & ~w112;
assign w35550 = ~w40 & ~w120;
assign w35551 = w40 & w14;
assign w35552 = ~w145 & pi3322;
assign w35553 = ~pi3323 & ~w161;
assign w35554 = w114 & ~w177;
assign w35555 = w180 & pi1462;
assign w35556 = w180 & pi2785;
assign w35557 = w114 & w177;
assign w35558 = ~w110 & pi3626;
assign w35559 = pi1781 & pi2785;
assign w35560 = pi1781 & w35556;
assign w35561 = pi1782 & pi1462;
assign w35562 = pi1782 & w35555;
assign w35563 = w185 & pi1783;
assign w35564 = w210 & pi1009;
assign w35565 = w219 & ~pi1009;
assign w35566 = pi1009 & pi0795;
assign w35567 = w225 & ~w205;
assign w35568 = w255 & pi0884;
assign w35569 = w264 & ~pi0884;
assign w35570 = pi0884 & pi0739;
assign w35571 = w270 & ~w250;
assign w35572 = w326 & ~w324;
assign w35573 = pi0541 & w332;
assign w35574 = ~w335 & pi3524;
assign w35575 = w340 & w323;
assign w35576 = w340 & w349;
assign w35577 = ~pi3304 & ~pi2598;
assign w35578 = ~pi3551 & w345;
assign w35579 = ~w35578 & w354;
assign w35580 = w361 & ~w363;
assign w35581 = pi2382 & ~pi3367;
assign w35582 = w35581 & pi3391;
assign w35583 = pi0993 & ~pi3426;
assign w35584 = pi3551 & w369;
assign w35585 = pi3435 & w372;
assign w35586 = ~pi0421 & ~pi0405;
assign w35587 = w35586 & w376;
assign w35588 = w375 & ~pi0412;
assign w35589 = ~w375 & w385;
assign w35590 = w386 & ~w373;
assign w35591 = pi2382 & pi3367;
assign w35592 = pi3391 & ~pi0994;
assign w35593 = pi3551 & w391;
assign w35594 = ~pi3435 & w393;
assign w35595 = w375 & ~pi0411;
assign w35596 = ~w375 & w397;
assign w35597 = w398 & ~w394;
assign w35598 = w35581 & ~pi3391;
assign w35599 = pi0995 & ~pi3426;
assign w35600 = ~pi3435 & w372;
assign w35601 = ~w375 & ~pi0414;
assign w35602 = ~w408 & ~w406;
assign w35603 = w35591 & pi3391;
assign w35604 = pi0992 & ~pi3426;
assign w35605 = ~w375 & ~pi0415;
assign w35606 = pi3435 & w393;
assign w35607 = ~w402 & w362;
assign w35608 = w431 & ~pi0612;
assign w35609 = w435 & ~pi0753;
assign w35610 = ~pi0639 & ~pi0640;
assign w35611 = ~pi0639 & ~pi0641;
assign w35612 = w439 & ~w459;
assign w35613 = ~w442 & ~w462;
assign w35614 = w439 & w426;
assign w35615 = w465 & pi0753;
assign w35616 = ~w437 & ~pi0753;
assign w35617 = ~w437 & ~w35615;
assign w35618 = w465 & ~w438;
assign w35619 = ~w436 & w438;
assign w35620 = ~w436 & ~w35618;
assign w35621 = ~pi0643 & ~pi0534;
assign w35622 = w434 & ~pi0614;
assign w35623 = w465 & ~w439;
assign w35624 = w476 & pi0756;
assign w35625 = ~w442 & w428;
assign w35626 = w430 & ~pi0658;
assign w35627 = w35626 & ~pi0612;
assign w35628 = ~pi0614 & ~pi0735;
assign w35629 = w465 & ~w484;
assign w35630 = ~pi0660 & ~pi0533;
assign w35631 = w465 & ~w483;
assign w35632 = w488 & pi0757;
assign w35633 = w488 & w494;
assign w35634 = w491 & ~w478;
assign w35635 = w473 & ~w472;
assign w35636 = ~w465 & ~w427;
assign w35637 = ~w35636 & pi0665;
assign w35638 = pi0510 & pi0509;
assign w35639 = ~w465 & ~w511;
assign w35640 = ~w464 & pi0664;
assign w35641 = w439 & ~pi0638;
assign w35642 = w465 & pi0634;
assign w35643 = pi0508 & w522;
assign w35644 = ~w465 & ~w428;
assign w35645 = pi0662 & pi0507;
assign w35646 = ~pi0508 & ~w527;
assign w35647 = ~pi0612 & ~pi0658;
assign w35648 = w35647 & ~pi0636;
assign w35649 = w465 & ~w532;
assign w35650 = w465 & pi0637;
assign w35651 = w465 & ~w458;
assign w35652 = pi0661 & pi0506;
assign w35653 = ~pi0661 & ~pi0506;
assign w35654 = ~pi0662 & ~pi0507;
assign w35655 = w35652 & pi0505;
assign w35656 = ~w547 & w549;
assign w35657 = ~pi0755 & ~pi0567;
assign w35658 = w465 & ~w531;
assign w35659 = ~w559 & ~w558;
assign w35660 = pi0535 & ~w473;
assign w35661 = w495 & w562;
assign w35662 = pi0660 & pi0533;
assign w35663 = pi0754 & pi0566;
assign w35664 = pi0755 & pi0567;
assign w35665 = w565 & ~w472;
assign w35666 = ~w573 & ~w500;
assign w35667 = ~pi0663 & ~w580;
assign w35668 = ~pi0641 & ~pi0568;
assign w35669 = ~w35636 & w601;
assign w35670 = pi0667 & ~w606;
assign w35671 = ~w35670 & w609;
assign w35672 = w596 & ~w595;
assign w35673 = ~pi0663 & w614;
assign w35674 = pi0663 & ~w614;
assign w35675 = w623 & ~w622;
assign w35676 = w612 & w626;
assign w35677 = ~w610 & w612;
assign w35678 = w585 & pi0507;
assign w35679 = w585 & ~w35654;
assign w35680 = ~w35663 & ~w650;
assign w35681 = pi0755 & ~pi0636;
assign w35682 = w465 & pi0755;
assign w35683 = pi0636 & ~pi0755;
assign w35684 = pi0636 & ~w35682;
assign w35685 = w35681 & w667;
assign w35686 = w673 & ~w553;
assign w35687 = ~pi0642 & ~pi0637;
assign w35688 = w465 & w690;
assign w35689 = ~pi0642 & ~w691;
assign w35690 = ~pi0505 & w696;
assign w35691 = w673 & ~w699;
assign w35692 = ~w701 & ~w689;
assign w35693 = ~w35652 & ~w696;
assign w35694 = ~w35652 & ~w637;
assign w35695 = w495 & w723;
assign w35696 = ~w35662 & ~w655;
assign w35697 = ~pi0535 & ~w735;
assign w35698 = ~w490 & ~w746;
assign w35699 = w35609 & pi0666;
assign w35700 = ~pi0666 & pi0753;
assign w35701 = w434 & w733;
assign w35702 = w465 & ~pi0568;
assign w35703 = w758 & w757;
assign w35704 = ~w35699 & ~pi0568;
assign w35705 = ~w758 & ~w757;
assign w35706 = ~w495 & w776;
assign w35707 = ~w495 & ~w776;
assign w35708 = w786 & ~w771;
assign w35709 = ~w719 & w755;
assign w35710 = w35699 & ~pi0568;
assign w35711 = ~w799 & w498;
assign w35712 = w575 & w806;
assign w35713 = w729 & ~w754;
assign w35714 = ~w719 & ~w754;
assign w35715 = ~w810 & ~w808;
assign w35716 = ~w807 & w424;
assign w35717 = w821 & pi1732;
assign w35718 = pi3641 & pi1441;
assign w35719 = ~w831 & ~w826;
assign w35720 = w821 & pi1731;
assign w35721 = pi3641 & pi1440;
assign w35722 = ~w837 & ~w835;
assign w35723 = w340 & w842;
assign w35724 = w340 & w847;
assign w35725 = pi3426 & ~w394;
assign w35726 = w340 & w854;
assign w35727 = w821 & pi1730;
assign w35728 = pi3641 & pi1439;
assign w35729 = ~w862 & ~w860;
assign w35730 = w417 & ~w864;
assign w35731 = ~w852 & w363;
assign w35732 = w362 & ~w364;
assign w35733 = w419 & pi2436;
assign w35734 = w410 & pi1984;
assign w35735 = w387 & pi2269;
assign w35736 = w400 & pi2446;
assign w35737 = w35578 & w347;
assign w35738 = ~pi1861 & ~pi1840;
assign w35739 = w35738 & pi3099;
assign w35740 = w344 & w899;
assign w35741 = w344 & w904;
assign w35742 = pi0541 & w906;
assign w35743 = ~pi3589 & pi3644;
assign w35744 = w911 & ~pi3362;
assign w35745 = w910 & pi3148;
assign w35746 = ~w917 & ~w916;
assign w35747 = ~pi3148 & ~w920;
assign w35748 = w922 & pi0541;
assign w35749 = ~pi3522 & ~pi3548;
assign w35750 = ~w923 & w919;
assign w35751 = ~w908 & w932;
assign w35752 = ~w933 & pi2529;
assign w35753 = ~w35737 & ~pi1422;
assign w35754 = ~pi3641 & pi2601;
assign w35755 = pi0819 & pi2601;
assign w35756 = pi0819 & w35754;
assign w35757 = w939 & ~pi1422;
assign w35758 = w939 & w35753;
assign w35759 = ~pi3515 & pi2557;
assign w35760 = ~w942 & ~w35757;
assign w35761 = ~w942 & ~w35758;
assign w35762 = w943 & w905;
assign w35763 = w949 & w950;
assign w35764 = w949 & ~pi3363;
assign w35765 = w979 & pi3983;
assign w35766 = w974 & pi3903;
assign w35767 = w977 & pi3887;
assign w35768 = w966 & pi3967;
assign w35769 = w955 & pi3935;
assign w35770 = w960 & pi3919;
assign w35771 = w971 & pi3855;
assign w35772 = w964 & pi3951;
assign w35773 = ~pi3515 & pi3296;
assign w35774 = pi1014 & pi1312;
assign w35775 = ~pi1043 & ~w1015;
assign w35776 = w1031 & w1030;
assign w35777 = w1017 & pi1331;
assign w35778 = ~w1059 & pi0650;
assign w35779 = ~w1067 & pi0722;
assign w35780 = ~w1090 & pi0539;
assign w35781 = ~w1125 & pi0576;
assign w35782 = ~w1184 & pi0538;
assign w35783 = ~w1199 & ~w1140;
assign w35784 = w1207 & w1215;
assign w35785 = w1205 & pi0688;
assign w35786 = w1207 & w1220;
assign w35787 = w1223 & pi0724;
assign w35788 = w1226 & pi2989;
assign w35789 = w1286 & pi0779;
assign w35790 = pi0796 & pi1844;
assign w35791 = pi0890 & pi1842;
assign w35792 = ~w1293 & ~w1290;
assign w35793 = w1300 & w1230;
assign w35794 = ~w1302 & ~w1003;
assign w35795 = w952 & ~w1305;
assign w35796 = pi1787 & w1306;
assign w35797 = w850 & ~w864;
assign w35798 = ~w417 & ~w864;
assign w35799 = w1311 & pi2436;
assign w35800 = w840 & ~w864;
assign w35801 = w857 & ~w864;
assign w35802 = ~w948 & ~w1320;
assign w35803 = ~w885 & w1322;
assign w35804 = w344 & w938;
assign w35805 = w1328 & ~w938;
assign w35806 = w1328 & ~w35804;
assign w35807 = pi3680 & w1330;
assign w35808 = w1335 & ~w938;
assign w35809 = w1335 & ~w35804;
assign w35810 = w1342 & ~w938;
assign w35811 = w1342 & ~w35804;
assign w35812 = w1348 & ~w938;
assign w35813 = w1348 & ~w35804;
assign w35814 = ~w792 & ~w787;
assign w35815 = w469 & w472;
assign w35816 = w469 & ~w35635;
assign w35817 = ~w572 & w1358;
assign w35818 = w1362 & w472;
assign w35819 = w1362 & ~w35635;
assign w35820 = ~w1360 & ~w1367;
assign w35821 = w1368 & w424;
assign w35822 = w387 & pi2268;
assign w35823 = w419 & pi2435;
assign w35824 = w410 & pi1983;
assign w35825 = w400 & pi2445;
assign w35826 = ~pi3515 & pi3358;
assign w35827 = w1395 & w1036;
assign w35828 = pi1014 & pi1213;
assign w35829 = ~w1394 & pi1331;
assign w35830 = ~w1428 & pi0650;
assign w35831 = ~w1438 & pi0576;
assign w35832 = w1223 & pi0687;
assign w35833 = w1286 & pi0752;
assign w35834 = w1226 & pi2988;
assign w35835 = w1205 & pi0929;
assign w35836 = ~w1561 & pi1934;
assign w35837 = ~w1615 & ~pi1934;
assign w35838 = ~w1615 & ~w35836;
assign w35839 = w1616 & ~w1380;
assign w35840 = w952 & ~w1619;
assign w35841 = pi1787 & w1620;
assign w35842 = w979 & pi3984;
assign w35843 = w974 & pi3904;
assign w35844 = w977 & pi3888;
assign w35845 = w960 & pi3920;
assign w35846 = w964 & pi3952;
assign w35847 = w955 & pi3936;
assign w35848 = w971 & pi3856;
assign w35849 = w966 & pi3968;
assign w35850 = ~w1638 & ~w1620;
assign w35851 = ~w1638 & ~w35841;
assign w35852 = ~w933 & pi2647;
assign w35853 = pi0909 & pi2601;
assign w35854 = pi0909 & w35754;
assign w35855 = w1642 & ~pi1422;
assign w35856 = w1642 & w35753;
assign w35857 = ~pi3515 & pi2558;
assign w35858 = ~w1643 & ~w35855;
assign w35859 = ~w1643 & ~w35856;
assign w35860 = w1644 & w905;
assign w35861 = w1311 & pi2435;
assign w35862 = ~w1379 & w1656;
assign w35863 = pi1014 & pi1212;
assign w35864 = w1669 & ~pi0976;
assign w35865 = w1668 & pi2483;
assign w35866 = pi1014 & pi1304;
assign w35867 = pi1014 & pi1206;
assign w35868 = ~w1704 & ~w1699;
assign w35869 = pi1014 & pi1192;
assign w35870 = w1712 & pi0976;
assign w35871 = ~w1707 & pi2477;
assign w35872 = pi1014 & pi1217;
assign w35873 = w1734 & ~pi0976;
assign w35874 = w1749 & ~w1744;
assign w35875 = w1707 & ~pi2477;
assign w35876 = ~pi1277 & ~pi1014;
assign w35877 = ~w1775 & ~pi0976;
assign w35878 = ~w1793 & ~w1784;
assign w35879 = ~w1668 & ~pi2483;
assign w35880 = w1382 & ~w1899;
assign w35881 = w1897 & pi2480;
assign w35882 = ~w1897 & ~pi2480;
assign w35883 = pi1014 & pi1309;
assign w35884 = pi1014 & pi1211;
assign w35885 = w1928 & ~pi0976;
assign w35886 = w1937 & ~pi2482;
assign w35887 = ~w1937 & pi2482;
assign w35888 = w1017 & ~pi2485;
assign w35889 = ~w1017 & pi2485;
assign w35890 = w1394 & pi2484;
assign w35891 = ~w1394 & ~pi2484;
assign w35892 = ~w1967 & ~pi2763;
assign w35893 = w1965 & w1972;
assign w35894 = w2003 & w1045;
assign w35895 = ~w2002 & ~pi2481;
assign w35896 = pi1014 & pi1302;
assign w35897 = pi1014 & pi1204;
assign w35898 = ~w2036 & ~w2031;
assign w35899 = w1687 & ~w2041;
assign w35900 = ~w2039 & pi2475;
assign w35901 = w2039 & ~pi2475;
assign w35902 = w2002 & pi2481;
assign w35903 = pi2763 & ~w2102;
assign w35904 = ~pi1250 & pi1014;
assign w35905 = ~w2105 & w2104;
assign w35906 = ~pi1320 & ~pi1014;
assign w35907 = ~w2111 & w2110;
assign w35908 = ~w2118 & w1030;
assign w35909 = ~w2133 & pi2479;
assign w35910 = w2133 & ~pi2479;
assign w35911 = w1037 & ~w2151;
assign w35912 = w2149 & pi2476;
assign w35913 = ~w2149 & ~pi2476;
assign w35914 = ~w2136 & ~w2135;
assign w35915 = w1993 & w2173;
assign w35916 = pi2489 & ~pi2490;
assign w35917 = w2178 & pi2912;
assign w35918 = ~w2182 & ~pi2913;
assign w35919 = w2182 & pi2913;
assign w35920 = w2188 & ~pi0045;
assign w35921 = ~w2194 & w2176;
assign w35922 = ~w2178 & pi3267;
assign w35923 = ~pi3248 & ~w2212;
assign w35924 = ~w2213 & ~pi0038;
assign w35925 = pi2490 & ~pi3210;
assign w35926 = w2177 & w2220;
assign w35927 = w2066 & w2171;
assign w35928 = ~w2223 & w2175;
assign w35929 = ~pi0540 & w2229;
assign w35930 = w2231 & pi0421;
assign w35931 = ~w2237 & ~w375;
assign w35932 = ~w2243 & ~w375;
assign w35933 = ~w361 & w2246;
assign w35934 = w35929 & w2247;
assign w35935 = ~pi3551 & pi3256;
assign w35936 = ~w35934 & w2255;
assign w35937 = pi2769 & w938;
assign w35938 = pi2769 & w35804;
assign w35939 = w2257 & w35937;
assign w35940 = w2257 & w35938;
assign w35941 = ~pi3551 & pi3370;
assign w35942 = ~w360 & ~w2260;
assign w35943 = w2263 & w2255;
assign w35944 = w2263 & w35936;
assign w35945 = pi3551 & ~pi3426;
assign w35946 = ~w941 & pi3426;
assign w35947 = ~w941 & ~w35945;
assign w35948 = pi3435 & w2286;
assign w35949 = pi2488 & w2288;
assign w35950 = pi0997 & ~pi3426;
assign w35951 = w340 & w2292;
assign w35952 = ~pi3435 & w2286;
assign w35953 = w864 & ~w2299;
assign w35954 = pi2488 & ~pi3398;
assign w35955 = w35954 & ~pi3392;
assign w35956 = pi0999 & ~pi3426;
assign w35957 = w370 & ~w2300;
assign w35958 = pi2488 & w2307;
assign w35959 = pi0996 & ~pi3426;
assign w35960 = pi3435 & w2310;
assign w35961 = w340 & w2313;
assign w35962 = ~pi3435 & w2310;
assign w35963 = ~pi3392 & ~pi0998;
assign w35964 = pi3426 & ~w2318;
assign w35965 = w340 & w2321;
assign w35966 = ~w2287 & w385;
assign w35967 = ~pi3551 & w385;
assign w35968 = w340 & w2329;
assign w35969 = w2332 & ~pi3551;
assign w35970 = w340 & w2335;
assign w35971 = ~pi3551 & w397;
assign w35972 = w340 & w2340;
assign w35973 = ~w2311 & w2343;
assign w35974 = ~pi3551 & w2343;
assign w35975 = w340 & w2345;
assign w35976 = w2352 & ~w2356;
assign w35977 = pi0418 & ~w375;
assign w35978 = ~w1207 & w2359;
assign w35979 = ~w2362 & ~w874;
assign w35980 = ~w2361 & w2366;
assign w35981 = w402 & ~w354;
assign w35982 = ~w852 & w2358;
assign w35983 = w2231 & ~pi0421;
assign w35984 = ~w874 & w2358;
assign w35985 = ~w2361 & ~w2379;
assign w35986 = pi0830 & w2382;
assign w35987 = ~w2350 & w2384;
assign w35988 = w2385 & ~w363;
assign w35989 = ~w2362 & ~w354;
assign w35990 = w402 & w2389;
assign w35991 = w852 & ~w2363;
assign w35992 = pi0830 & ~w2382;
assign w35993 = w2380 & ~w2395;
assign w35994 = ~w35993 & ~w363;
assign w35995 = w643 & w2400;
assign w35996 = ~w643 & ~w2400;
assign w35997 = ~w537 & pi0642;
assign w35998 = ~w575 & ~w2405;
assign w35999 = ~w546 & w551;
assign w36000 = ~w546 & ~w542;
assign w36001 = w575 & ~w2413;
assign w36002 = ~w2361 & ~w2377;
assign w36003 = w2362 & ~w2384;
assign w36004 = ~w36003 & ~w363;
assign w36005 = ~w2366 & ~w354;
assign w36006 = ~w2366 & ~w35579;
assign w36007 = ~w2350 & w2422;
assign w36008 = ~w2392 & ~w2423;
assign w36009 = ~pi0675 & ~pi0676;
assign w36010 = w2435 & w2453;
assign w36011 = pi0675 & pi0676;
assign w36012 = ~pi0675 & ~pi0668;
assign w36013 = ~w2457 & w2461;
assign w36014 = w2431 & ~pi0671;
assign w36015 = ~w2455 & pi0678;
assign w36016 = ~w2456 & w2428;
assign w36017 = ~w2470 & w2472;
assign w36018 = ~w2466 & pi0513;
assign w36019 = ~pi0672 & ~pi0588;
assign w36020 = w2478 & w2479;
assign w36021 = w2470 & w2483;
assign w36022 = ~w2484 & pi0706;
assign w36023 = w2429 & pi0679;
assign w36024 = ~pi0656 & w2490;
assign w36025 = w2478 & w2470;
assign w36026 = ~w2473 & pi0515;
assign w36027 = ~w2471 & w2502;
assign w36028 = ~w2506 & ~w2476;
assign w36029 = w2508 & w2427;
assign w36030 = w2466 & ~pi0513;
assign w36031 = ~w2456 & ~pi0644;
assign w36032 = ~w2518 & pi0702;
assign w36033 = w2428 & ~pi0668;
assign w36034 = w2521 & ~w2454;
assign w36035 = ~pi0701 & ~pi0511;
assign w36036 = ~w2517 & pi0677;
assign w36037 = pi0512 & pi0520;
assign w36038 = ~w2507 & w2529;
assign w36039 = w2457 & w2452;
assign w36040 = ~w2533 & pi0683;
assign w36041 = pi0701 & pi0511;
assign w36042 = ~w2536 & ~w2534;
assign w36043 = w36042 & ~pi0519;
assign w36044 = ~w2507 & w2547;
assign w36045 = ~w36041 & ~pi0520;
assign w36046 = w2550 & ~pi0519;
assign w36047 = ~pi0676 & w2451;
assign w36048 = ~w36047 & w2450;
assign w36049 = ~w2457 & ~pi0676;
assign w36050 = pi0646 & ~pi0675;
assign w36051 = ~w2560 & ~w2556;
assign w36052 = ~w2558 & w2556;
assign w36053 = ~w2451 & pi0682;
assign w36054 = pi0519 & pi0589;
assign w36055 = pi0519 & ~w4488;
assign w36056 = ~pi0645 & ~w2555;
assign w36057 = ~pi0680 & pi0518;
assign w36058 = w2478 & w2592;
assign w36059 = w2478 & w2599;
assign w36060 = ~w2621 & ~pi0679;
assign w36061 = ~w2621 & ~w36023;
assign w36062 = w2627 & ~pi0679;
assign w36063 = w2627 & ~w36023;
assign w36064 = ~w2635 & ~w2634;
assign w36065 = w2636 & ~w2626;
assign w36066 = ~w2622 & w2638;
assign w36067 = ~w2613 & ~w2612;
assign w36068 = ~w2471 & pi0704;
assign w36069 = ~w2640 & w2656;
assign w36070 = pi0703 & w2673;
assign w36071 = ~pi0703 & ~w2673;
assign w36072 = ~pi0514 & ~w2679;
assign w36073 = ~w36070 & w2687;
assign w36074 = ~w36070 & w2690;
assign w36075 = ~w2428 & w2699;
assign w36076 = w2700 & ~w2699;
assign w36077 = w2700 & ~w36075;
assign w36078 = pi0704 & ~w2701;
assign w36079 = w2703 & ~w2712;
assign w36080 = ~w36070 & ~w2671;
assign w36081 = w2686 & ~w2717;
assign w36082 = ~w2727 & ~w2723;
assign w36083 = pi0677 & ~w2728;
assign w36084 = pi0587 & w2686;
assign w36085 = w2760 & ~w2759;
assign w36086 = w2733 & pi0511;
assign w36087 = w2733 & ~w36035;
assign w36088 = ~w2752 & ~w2750;
assign w36089 = pi0681 & ~w2779;
assign w36090 = ~pi0681 & w2779;
assign w36091 = w2762 & ~w2783;
assign w36092 = ~w2794 & w2784;
assign w36093 = w2776 & pi0589;
assign w36094 = w2776 & ~w4488;
assign w36095 = pi0680 & ~pi0518;
assign w36096 = ~pi0645 & w2801;
assign w36097 = ~w2797 & w2802;
assign w36098 = pi0680 & ~pi0645;
assign w36099 = ~pi0680 & pi0645;
assign w36100 = w2807 & ~pi0518;
assign w36101 = ~w2808 & w2816;
assign w36102 = ~w2773 & w2801;
assign w36103 = w2518 & pi0702;
assign w36104 = ~w2831 & ~w2708;
assign w36105 = w2830 & ~w2712;
assign w36106 = w2682 & w2829;
assign w36107 = ~w2682 & w2836;
assign w36108 = w2507 & w2683;
assign w36109 = ~w2507 & ~w2683;
assign w36110 = w1311 & pi2258;
assign w36111 = w419 & pi2258;
assign w36112 = w400 & pi2272;
assign w36113 = w387 & pi2262;
assign w36114 = w410 & pi1977;
assign w36115 = ~w2856 & w2417;
assign w36116 = w2328 & pi2454;
assign w36117 = w2344 & pi2962;
assign w36118 = w2334 & pi2462;
assign w36119 = w2872 & ~w354;
assign w36120 = pi3551 & w2303;
assign w36121 = ~w2298 & ~w2303;
assign w36122 = ~w2298 & ~w36120;
assign w36123 = w2312 & pi2962;
assign w36124 = w2291 & pi2454;
assign w36125 = w2880 & ~w2877;
assign w36126 = ~w2874 & w2363;
assign w36127 = w344 & ~w2898;
assign w36128 = ~pi3515 & pi2450;
assign w36129 = pi0403 & pi0426;
assign w36130 = ~w2361 & w2902;
assign w36131 = ~w36130 & ~w2900;
assign w36132 = ~w35737 & pi1422;
assign w36133 = pi0904 & pi2601;
assign w36134 = pi0904 & w35754;
assign w36135 = ~w933 & pi1031;
assign w36136 = w2370 & ~w2914;
assign w36137 = w2344 & pi2961;
assign w36138 = w2334 & pi2461;
assign w36139 = w2328 & pi2453;
assign w36140 = w2919 & ~w354;
assign w36141 = w2312 & pi2961;
assign w36142 = w2291 & pi2453;
assign w36143 = w2928 & ~w2925;
assign w36144 = ~w2370 & w2934;
assign w36145 = ~w2849 & w2938;
assign w36146 = ~w2830 & w2944;
assign w36147 = w2830 & w2946;
assign w36148 = w2481 & w2505;
assign w36149 = w979 & pi3978;
assign w36150 = w977 & pi3882;
assign w36151 = w974 & pi3898;
assign w36152 = w960 & pi3914;
assign w36153 = w964 & pi3946;
assign w36154 = w955 & pi3930;
assign w36155 = w971 & pi3850;
assign w36156 = w966 & pi3962;
assign w36157 = ~pi3515 & pi3308;
assign w36158 = w1707 & pi1331;
assign w36159 = ~w2992 & pi0650;
assign w36160 = ~w3000 & pi0722;
assign w36161 = ~w3023 & pi0539;
assign w36162 = ~pi0838 & ~w3084;
assign w36163 = ~w3085 & pi0576;
assign w36164 = w3127 & pi2495;
assign w36165 = w1226 & pi2503;
assign w36166 = w1223 & pi0769;
assign w36167 = w1205 & pi1602;
assign w36168 = w1286 & pi0861;
assign w36169 = ~w3134 & pi1934;
assign w36170 = ~w3189 & ~w2980;
assign w36171 = w952 & ~w3192;
assign w36172 = pi1787 & w3193;
assign w36173 = ~pi3515 & pi3298;
assign w36174 = w3127 & pi2496;
assign w36175 = w1205 & pi1474;
assign w36176 = w1226 & pi2504;
assign w36177 = w1223 & pi0770;
assign w36178 = w1286 & pi0773;
assign w36179 = ~w3204 & pi1934;
assign w36180 = ~pi1331 & w3266;
assign w36181 = ~w3275 & pi0539;
assign w36182 = ~w3298 & pi0722;
assign w36183 = ~pi0768 & ~w3363;
assign w36184 = ~w3364 & pi0576;
assign w36185 = ~w3389 & pi0538;
assign w36186 = ~w3253 & ~w3197;
assign w36187 = w952 & ~w3413;
assign w36188 = pi1787 & w3414;
assign w36189 = w974 & pi3897;
assign w36190 = w979 & pi3977;
assign w36191 = w971 & pi3849;
assign w36192 = w960 & pi3913;
assign w36193 = w955 & pi3929;
assign w36194 = w966 & pi3961;
assign w36195 = w977 & pi3881;
assign w36196 = w964 & pi3945;
assign w36197 = ~w3432 & ~w3414;
assign w36198 = ~w3432 & ~w36188;
assign w36199 = ~w2941 & w3436;
assign w36200 = w2574 & pi0518;
assign w36201 = w2576 & ~pi0518;
assign w36202 = w2576 & ~w36200;
assign w36203 = ~w2794 & ~w2772;
assign w36204 = ~w3445 & w3446;
assign w36205 = pi0645 & ~pi0518;
assign w36206 = ~w36204 & w3449;
assign w36207 = ~w3450 & ~pi0680;
assign w36208 = w2574 & w3454;
assign w36209 = w2797 & ~w3458;
assign w36210 = w3459 & ~w3454;
assign w36211 = w3459 & ~w36208;
assign w36212 = ~w2797 & ~w3462;
assign w36213 = ~w3463 & ~w3460;
assign w36214 = w974 & pi3891;
assign w36215 = w977 & pi3875;
assign w36216 = w979 & pi3971;
assign w36217 = w960 & pi3907;
assign w36218 = w966 & pi3955;
assign w36219 = w955 & pi3923;
assign w36220 = w971 & pi3843;
assign w36221 = w964 & pi3939;
assign w36222 = ~pi3515 & pi3316;
assign w36223 = ~pi1331 & w3502;
assign w36224 = ~w3511 & pi0722;
assign w36225 = ~w3534 & pi0539;
assign w36226 = ~w3569 & pi0538;
assign w36227 = ~pi0838 & ~w3589;
assign w36228 = ~w3590 & pi0576;
assign w36229 = ~w3610 & ~w3585;
assign w36230 = w1286 & pi0749;
assign w36231 = w1226 & pi2990;
assign w36232 = w1223 & pi0787;
assign w36233 = w1205 & pi2059;
assign w36234 = w3127 & pi2502;
assign w36235 = ~w3656 & pi1934;
assign w36236 = ~w3705 & ~w3485;
assign w36237 = w952 & ~w3708;
assign w36238 = pi1787 & w3709;
assign w36239 = w2328 & pi2458;
assign w36240 = w2344 & pi2748;
assign w36241 = w2334 & pi2410;
assign w36242 = w3720 & ~w354;
assign w36243 = w2291 & pi2458;
assign w36244 = w2312 & pi2748;
assign w36245 = w3726 & ~w3723;
assign w36246 = w3712 & w2397;
assign w36247 = ~w3722 & ~w2358;
assign w36248 = ~w933 & pi1035;
assign w36249 = ~w3743 & w3742;
assign w36250 = w2365 & ~w3750;
assign w36251 = w2328 & pi2524;
assign w36252 = w2344 & pi2964;
assign w36253 = w2334 & pi2470;
assign w36254 = w3757 & ~w354;
assign w36255 = w2312 & pi2964;
assign w36256 = w2320 & pi2968;
assign w36257 = w2291 & pi2524;
assign w36258 = ~w2370 & ~w3775;
assign w36259 = ~w1360 & w3780;
assign w36260 = ~w3781 & ~w3784;
assign w36261 = ~w2578 & w3789;
assign w36262 = w2578 & w3791;
assign w36263 = ~w2811 & ~w2814;
assign w36264 = ~w36098 & ~w3794;
assign w36265 = ~pi0707 & ~w3788;
assign w36266 = ~w3796 & w3798;
assign w36267 = pi0521 & ~w3794;
assign w36268 = pi0521 & w36264;
assign w36269 = ~pi0521 & w3794;
assign w36270 = ~pi0521 & ~w36264;
assign w36271 = w2462 & ~w36269;
assign w36272 = w2462 & ~w36270;
assign w36273 = ~pi0656 & ~w3801;
assign w36274 = ~w2811 & w3807;
assign w36275 = ~w2635 & ~w3809;
assign w36276 = w3790 & w3786;
assign w36277 = w569 & ~w565;
assign w36278 = ~w570 & ~w3819;
assign w36279 = w575 & w3821;
assign w36280 = ~w3825 & ~w3824;
assign w36281 = w3823 & ~w3819;
assign w36282 = ~w575 & w3829;
assign w36283 = pi0515 & ~w2472;
assign w36284 = w2471 & pi0704;
assign w36285 = w3835 & ~w3833;
assign w36286 = ~w3837 & w3433;
assign w36287 = ~w2640 & ~w2643;
assign w36288 = ~w2666 & w2643;
assign w36289 = ~w2666 & ~w36287;
assign w36290 = w3840 & w3433;
assign w36291 = w2328 & pi2452;
assign w36292 = w2334 & pi2413;
assign w36293 = w2344 & pi2960;
assign w36294 = w3847 & ~w354;
assign w36295 = w2291 & pi2452;
assign w36296 = w2312 & pi2960;
assign w36297 = w3857 & ~w3854;
assign w36298 = ~w3852 & ~w2358;
assign w36299 = w1311 & pi2257;
assign w36300 = w387 & pi2261;
assign w36301 = w400 & pi2271;
assign w36302 = w419 & pi2257;
assign w36303 = w410 & pi1976;
assign w36304 = ~w3874 & ~w354;
assign w36305 = pi0403 & pi0424;
assign w36306 = w2377 & ~w3881;
assign w36307 = w3864 & w2365;
assign w36308 = pi0902 & pi2601;
assign w36309 = pi0902 & w35754;
assign w36310 = ~w933 & pi1028;
assign w36311 = ~w3887 & w3885;
assign w36312 = ~w3891 & ~w3890;
assign w36313 = w2344 & pi2963;
assign w36314 = w2334 & pi2464;
assign w36315 = w2291 & pi2455;
assign w36316 = w3905 & ~w3902;
assign w36317 = ~w3911 & ~w2397;
assign w36318 = ~w3844 & w3913;
assign w36319 = w3917 & w3918;
assign w36320 = ~w2746 & ~w2789;
assign w36321 = w2790 & ~w3924;
assign w36322 = ~w2507 & ~w2520;
assign w36323 = ~w2539 & ~w2526;
assign w36324 = w2545 & w2526;
assign w36325 = w2545 & ~w36323;
assign w36326 = ~w3924 & ~w36324;
assign w36327 = ~w3924 & ~w36325;
assign w36328 = w3935 & w2397;
assign w36329 = w977 & pi3884;
assign w36330 = w979 & pi3980;
assign w36331 = w974 & pi3900;
assign w36332 = w960 & pi3916;
assign w36333 = w966 & pi3964;
assign w36334 = w955 & pi3932;
assign w36335 = w971 & pi3852;
assign w36336 = w964 & pi3948;
assign w36337 = ~pi3515 & pi3306;
assign w36338 = w2039 & pi1331;
assign w36339 = ~w3963 & pi0650;
assign w36340 = ~w3971 & pi0722;
assign w36341 = ~w3994 & pi0539;
assign w36342 = w4052 & ~pi0979;
assign w36343 = w4057 & pi0979;
assign w36344 = ~w4061 & ~w4056;
assign w36345 = w3127 & pi2493;
assign w36346 = w1205 & pi1066;
assign w36347 = w1223 & pi0723;
assign w36348 = w1226 & pi3107;
assign w36349 = w1286 & pi0845;
assign w36350 = pi0796 & pi1849;
assign w36351 = pi0890 & pi1846;
assign w36352 = w4132 & ~w4123;
assign w36353 = w4133 & w4099;
assign w36354 = ~w4135 & ~w3955;
assign w36355 = w952 & ~w4138;
assign w36356 = pi1787 & w4139;
assign w36357 = w977 & pi3879;
assign w36358 = w979 & pi3975;
assign w36359 = w974 & pi3895;
assign w36360 = w960 & pi3911;
assign w36361 = w964 & pi3943;
assign w36362 = w955 & pi3927;
assign w36363 = w971 & pi3847;
assign w36364 = w966 & pi3959;
assign w36365 = ~pi3515 & pi3310;
assign w36366 = w1286 & pi0775;
assign w36367 = w1223 & pi0782;
assign w36368 = w1226 & pi2505;
assign w36369 = w1205 & pi1467;
assign w36370 = w3127 & pi2513;
assign w36371 = ~w4168 & pi1934;
assign w36372 = ~pi1331 & w4232;
assign w36373 = ~w4241 & pi0539;
assign w36374 = ~w4264 & pi0722;
assign w36375 = ~pi0838 & ~w4294;
assign w36376 = ~w4295 & pi0576;
assign w36377 = ~w4320 & pi0538;
assign w36378 = ~w4336 & ~w4315;
assign w36379 = ~w4373 & ~w941;
assign w36380 = ~w4217 & ~w4161;
assign w36381 = w952 & ~w4377;
assign w36382 = pi1787 & w4378;
assign w36383 = ~w2941 & w4383;
assign w36384 = w643 & ~w715;
assign w36385 = ~w712 & ~w715;
assign w36386 = ~w712 & w36384;
assign w36387 = ~w643 & w4397;
assign w36388 = ~w575 & ~w4399;
assign w36389 = w575 & w4405;
assign w36390 = ~w4406 & ~w4405;
assign w36391 = ~w4406 & ~w36389;
assign w36392 = ~w2924 & ~w2358;
assign w36393 = w1311 & pi2699;
assign w36394 = w387 & pi2439;
assign w36395 = w400 & pi2702;
assign w36396 = w419 & pi2699;
assign w36397 = w410 & pi2276;
assign w36398 = ~w4419 & ~w354;
assign w36399 = pi0403 & pi0425;
assign w36400 = w2377 & ~w4426;
assign w36401 = w4409 & w2365;
assign w36402 = pi0876 & pi2601;
assign w36403 = pi0876 & w35754;
assign w36404 = ~w933 & pi1030;
assign w36405 = ~w4432 & w4430;
assign w36406 = ~w4436 & ~w4435;
assign w36407 = w2397 & w40134;
assign w36408 = ~w2425 & ~w4440;
assign w36409 = ~w2425 & w4443;
assign w36410 = ~w3440 & ~w4449;
assign w36411 = ~pi0656 & w2487;
assign w36412 = w2491 & ~pi0679;
assign w36413 = ~w2429 & pi0679;
assign w36414 = w2328 & pi2457;
assign w36415 = w2344 & pi2747;
assign w36416 = w2334 & pi2466;
assign w36417 = w4470 & ~w354;
assign w36418 = w2291 & pi2457;
assign w36419 = w4476 & ~w4473;
assign w36420 = ~w2425 & w4483;
assign w36421 = ~w4491 & ~w4488;
assign w36422 = ~w4491 & pi0589;
assign w36423 = w3445 & w4496;
assign w36424 = ~w3445 & ~w4496;
assign w36425 = ~w36424 & ~w4498;
assign w36426 = w807 & w3782;
assign w36427 = w979 & pi3972;
assign w36428 = w977 & pi3876;
assign w36429 = w974 & pi3892;
assign w36430 = w960 & pi3908;
assign w36431 = w964 & pi3940;
assign w36432 = w955 & pi3924;
assign w36433 = w971 & pi3844;
assign w36434 = w966 & pi3956;
assign w36435 = w3127 & pi2499;
assign w36436 = w1223 & pi0733;
assign w36437 = w1205 & pi2061;
assign w36438 = w1226 & pi2986;
assign w36439 = w1286 & pi0778;
assign w36440 = ~w4530 & pi1934;
assign w36441 = ~pi1331 & w4596;
assign w36442 = ~w4605 & pi0722;
assign w36443 = ~w4628 & pi0539;
assign w36444 = ~w4663 & pi0538;
assign w36445 = ~pi0768 & ~w4717;
assign w36446 = ~w4718 & pi0576;
assign w36447 = ~w4739 & ~w4678;
assign w36448 = ~w4741 & ~w941;
assign w36449 = ~pi3515 & pi3312;
assign w36450 = ~w4579 & ~w4744;
assign w36451 = w952 & ~w4746;
assign w36452 = pi1787 & w4747;
assign w36453 = w2334 & pi2467;
assign w36454 = w2328 & pi2525;
assign w36455 = w2344 & pi2533;
assign w36456 = w4756 & ~w354;
assign w36457 = w2312 & pi2533;
assign w36458 = w2320 & pi2755;
assign w36459 = w2291 & pi2525;
assign w36460 = ~w882 & ~w354;
assign w36461 = w4505 & w2397;
assign w36462 = ~w4758 & ~w2358;
assign w36463 = w4778 & w2365;
assign w36464 = ~w933 & pi1036;
assign w36465 = ~w4783 & w4782;
assign w36466 = ~w570 & ~w487;
assign w36467 = ~w488 & pi0757;
assign w36468 = ~w570 & w4801;
assign w36469 = w575 & w4803;
assign w36470 = ~w3823 & w4805;
assign w36471 = ~w4807 & ~w4798;
assign w36472 = ~w575 & ~w4810;
assign w36473 = w1311 & pi2700;
assign w36474 = w419 & pi2700;
assign w36475 = w410 & pi2278;
assign w36476 = w387 & pi2441;
assign w36477 = w400 & pi2751;
assign w36478 = ~w4825 & ~w354;
assign w36479 = w2328 & pi2460;
assign w36480 = w2334 & pi2469;
assign w36481 = w2344 & pi2750;
assign w36482 = w4831 & ~w354;
assign w36483 = w2291 & pi2460;
assign w36484 = w4841 & ~w4838;
assign w36485 = w979 & pi3981;
assign w36486 = w974 & pi3901;
assign w36487 = w971 & pi3853;
assign w36488 = w960 & pi3917;
assign w36489 = w964 & pi3949;
assign w36490 = w955 & pi3933;
assign w36491 = w977 & pi3885;
assign w36492 = w966 & pi3965;
assign w36493 = ~pi3515 & pi3315;
assign w36494 = ~pi1331 & w4872;
assign w36495 = ~w4881 & pi0539;
assign w36496 = ~w4904 & pi0722;
assign w36497 = ~w4955 & pi0576;
assign w36498 = ~w4970 & ~w4946;
assign w36499 = w3127 & pi2501;
assign w36500 = w1205 & pi1090;
assign w36501 = w1223 & pi0726;
assign w36502 = w1226 & pi3063;
assign w36503 = w1286 & pi0781;
assign w36504 = pi0890 & pi1702;
assign w36505 = pi0796 & pi1629;
assign w36506 = w5044 & ~w5034;
assign w36507 = w5045 & w5012;
assign w36508 = ~w5047 & ~w4867;
assign w36509 = w952 & ~w5050;
assign w36510 = pi1787 & w5051;
assign w36511 = ~w2397 & w2425;
assign w36512 = ~w4836 & w2363;
assign w36513 = ~pi3515 & pi2707;
assign w36514 = pi0403 & pi0423;
assign w36515 = ~w2361 & w5062;
assign w36516 = ~w36515 & ~w5061;
assign w36517 = pi0910 & pi2601;
assign w36518 = pi0910 & w35754;
assign w36519 = ~w933 & pi1038;
assign w36520 = w974 & pi3894;
assign w36521 = w979 & pi3974;
assign w36522 = w971 & pi3846;
assign w36523 = w960 & pi3910;
assign w36524 = w966 & pi3958;
assign w36525 = w955 & pi3926;
assign w36526 = w977 & pi3878;
assign w36527 = w964 & pi3942;
assign w36528 = ~pi3515 & pi3311;
assign w36529 = ~w2002 & pi1331;
assign w36530 = ~w5111 & pi0650;
assign w36531 = ~w5154 & pi0722;
assign w36532 = ~pi0837 & ~w5172;
assign w36533 = ~w5176 & pi0576;
assign w36534 = ~w5206 & pi0538;
assign w36535 = w1286 & pi0776;
assign w36536 = w1205 & pi1841;
assign w36537 = w1223 & pi0772;
assign w36538 = w1226 & pi3100;
assign w36539 = w3127 & pi2498;
assign w36540 = ~w5232 & pi1934;
assign w36541 = pi3515 & pi0539;
assign w36542 = ~w5296 & w5289;
assign w36543 = w5313 & ~pi1934;
assign w36544 = w5313 & ~w36540;
assign w36545 = w5314 & ~w5093;
assign w36546 = w952 & ~w5317;
assign w36547 = pi1787 & w5318;
assign w36548 = w2397 & w5320;
assign w36549 = ~w5057 & ~w5323;
assign w36550 = ~w2494 & ~pi0588;
assign w36551 = w2494 & pi0588;
assign w36552 = ~pi0705 & ~w5329;
assign w36553 = ~w2817 & ~w5331;
assign w36554 = ~w2578 & w5332;
assign w36555 = w5329 & w2578;
assign w36556 = ~w5333 & w2425;
assign w36557 = w2328 & pi2456;
assign w36558 = w2344 & pi2780;
assign w36559 = w2334 & pi2465;
assign w36560 = w5345 & ~w354;
assign w36561 = w2291 & pi2456;
assign w36562 = w5355 & ~w5352;
assign w36563 = w2533 & pi0683;
assign w36564 = ~w2746 & w5365;
assign w36565 = ~w2746 & w2791;
assign w36566 = w5366 & ~w5364;
assign w36567 = ~w5363 & ~w5324;
assign w36568 = ~w2769 & w2761;
assign w36569 = w2769 & ~w2761;
assign w36570 = ~w2752 & ~w5381;
assign w36571 = w2752 & ~w5385;
assign w36572 = ~w2769 & w5387;
assign w36573 = w2769 & w5389;
assign w36574 = w5391 & ~w5384;
assign w36575 = w2554 & ~w2565;
assign w36576 = ~w2554 & pi0682;
assign w36577 = ~w570 & w5399;
assign w36578 = ~w476 & pi0756;
assign w36579 = ~w799 & w5404;
assign w36580 = w575 & w5406;
assign w36581 = ~w4807 & ~w729;
assign w36582 = ~w729 & ~w5402;
assign w36583 = ~w5407 & w3782;
assign w36584 = ~w5422 & w3786;
assign w36585 = w2484 & pi0706;
assign w36586 = w2638 & ~w5427;
assign w36587 = ~w2397 & ~w5429;
assign w36588 = w979 & pi3982;
assign w36589 = w977 & pi3886;
assign w36590 = w974 & pi3902;
assign w36591 = w960 & pi3918;
assign w36592 = w964 & pi3950;
assign w36593 = w955 & pi3934;
assign w36594 = w971 & pi3854;
assign w36595 = w966 & pi3966;
assign w36596 = w3127 & pi2500;
assign w36597 = w1205 & pi0930;
assign w36598 = w1223 & pi0725;
assign w36599 = w1226 & pi3091;
assign w36600 = w1286 & pi0780;
assign w36601 = pi0796 & pi1687;
assign w36602 = pi0890 & pi1684;
assign w36603 = w5488 & ~w5479;
assign w36604 = w5489 & w5455;
assign w36605 = ~pi1331 & w5496;
assign w36606 = ~w5505 & pi0722;
assign w36607 = ~w5528 & pi0539;
assign w36608 = ~pi0762 & ~w941;
assign w36609 = ~w5563 & pi0576;
assign w36610 = ~w5625 & ~w5579;
assign w36611 = w5631 & ~pi1787;
assign w36612 = w952 & ~w5633;
assign w36613 = ~w5634 & ~w5448;
assign w36614 = w1311 & pi2539;
assign w36615 = w419 & pi2539;
assign w36616 = w410 & pi2277;
assign w36617 = w387 & pi2440;
assign w36618 = w400 & pi2703;
assign w36619 = ~w5649 & ~w354;
assign w36620 = w2344 & pi2749;
assign w36621 = w2334 & pi2468;
assign w36622 = w2328 & pi2459;
assign w36623 = w5655 & ~w354;
assign w36624 = w2291 & pi2459;
assign w36625 = w5665 & ~w5662;
assign w36626 = ~pi3515 & pi3297;
assign w36627 = w1937 & pi1331;
assign w36628 = ~w5691 & pi0650;
assign w36629 = ~w5734 & pi0722;
assign w36630 = ~w5760 & pi0538;
assign w36631 = ~pi0768 & ~w5779;
assign w36632 = ~w5780 & pi0576;
assign w36633 = w1226 & pi3099;
assign w36634 = w1223 & pi0786;
assign w36635 = w3127 & pi2512;
assign w36636 = w3139 & ~w5811;
assign w36637 = w1205 & pi2058;
assign w36638 = w1286 & pi0777;
assign w36639 = w5828 & w5809;
assign w36640 = ~w5866 & w5289;
assign w36641 = ~pi1934 & w5891;
assign w36642 = w5673 & ~pi1787;
assign w36643 = w952 & ~w5894;
assign w36644 = w5895 & pi1787;
assign w36645 = w5895 & ~w36642;
assign w36646 = w974 & pi3893;
assign w36647 = w971 & pi3845;
assign w36648 = w977 & pi3877;
assign w36649 = w966 & pi3957;
assign w36650 = w955 & pi3925;
assign w36651 = w960 & pi3909;
assign w36652 = w979 & pi3973;
assign w36653 = w964 & pi3941;
assign w36654 = ~w5913 & ~w36645;
assign w36655 = ~w5913 & ~w36644;
assign w36656 = w5636 & w2397;
assign w36657 = ~w5660 & w2363;
assign w36658 = pi0820 & pi2601;
assign w36659 = pi0820 & w35754;
assign w36660 = ~w933 & pi1037;
assign w36661 = ~pi3515 & pi2706;
assign w36662 = pi0403 & pi0422;
assign w36663 = ~w2361 & w5924;
assign w36664 = ~w36663 & ~w5923;
assign w36665 = w5925 & ~w5921;
assign w36666 = w2370 & ~w5930;
assign w36667 = w2328 & pi2526;
assign w36668 = w2334 & pi2411;
assign w36669 = w2344 & pi2776;
assign w36670 = w5935 & ~w354;
assign w36671 = w2291 & pi2526;
assign w36672 = w5945 & ~w5942;
assign w36673 = ~w2370 & ~w5950;
assign w36674 = ~w5430 & w5954;
assign w36675 = w545 & ~w544;
assign w36676 = w575 & w5963;
assign w36677 = w589 & ~w645;
assign w36678 = ~w575 & w5967;
assign w36679 = w971 & pi3851;
assign w36680 = w974 & pi3899;
assign w36681 = w977 & pi3883;
assign w36682 = w966 & pi3963;
assign w36683 = w955 & pi3931;
assign w36684 = w964 & pi3947;
assign w36685 = w979 & pi3979;
assign w36686 = w960 & pi3915;
assign w36687 = ~pi3515 & pi3307;
assign w36688 = ~w2149 & pi1331;
assign w36689 = ~w5996 & pi0650;
assign w36690 = ~w6004 & pi0539;
assign w36691 = ~w6027 & pi0722;
assign w36692 = ~w6108 & pi0576;
assign w36693 = w3127 & pi2494;
assign w36694 = w1205 & pi0928;
assign w36695 = w1223 & pi0732;
assign w36696 = w1226 & pi3101;
assign w36697 = w1286 & pi0862;
assign w36698 = pi0890 & pi1847;
assign w36699 = pi0796 & pi1848;
assign w36700 = w6168 & ~w6159;
assign w36701 = w6169 & w6135;
assign w36702 = ~w6171 & ~w5988;
assign w36703 = w952 & ~w6174;
assign w36704 = pi1787 & w6175;
assign w36705 = w977 & pi3880;
assign w36706 = w979 & pi3976;
assign w36707 = w971 & pi3848;
assign w36708 = w960 & pi3912;
assign w36709 = w964 & pi3944;
assign w36710 = w955 & pi3928;
assign w36711 = w974 & pi3896;
assign w36712 = w966 & pi3960;
assign w36713 = w2133 & pi1331;
assign w36714 = ~w6218 & pi0539;
assign w36715 = ~w6241 & pi0722;
assign w36716 = ~pi0838 & ~w6271;
assign w36717 = ~w6272 & pi0576;
assign w36718 = ~w6297 & pi0538;
assign w36719 = ~w6313 & ~w6292;
assign w36720 = ~pi3515 & ~pi3309;
assign w36721 = w1286 & pi0774;
assign w36722 = w1223 & pi0771;
assign w36723 = w3127 & pi2497;
assign w36724 = ~w6360 & pi1934;
assign w36725 = w6409 & ~pi1787;
assign w36726 = w952 & ~w6411;
assign w36727 = ~w6412 & ~w6196;
assign w36728 = w2344 & pi2746;
assign w36729 = w2328 & pi2527;
assign w36730 = w2334 & pi2463;
assign w36731 = w6420 & ~w354;
assign w36732 = w2291 & pi2527;
assign w36733 = w6427 & ~w6424;
assign w36734 = w1311 & pi2432;
assign w36735 = w387 & pi2263;
assign w36736 = w400 & pi2442;
assign w36737 = w419 & pi2432;
assign w36738 = w410 & pi1978;
assign w36739 = ~w6442 & ~w354;
assign w36740 = w6178 & w2397;
assign w36741 = pi0403 & pi0409;
assign w36742 = ~w6422 & ~w2358;
assign w36743 = w6454 & w2365;
assign w36744 = ~pi3515 & pi2451;
assign w36745 = pi0905 & pi2601;
assign w36746 = pi0905 & w35754;
assign w36747 = ~w933 & pi1013;
assign w36748 = ~w6461 & w6459;
assign w36749 = w6456 & ~w6453;
assign w36750 = w2344 & pi2535;
assign w36751 = w2328 & pi2520;
assign w36752 = w2334 & pi2412;
assign w36753 = w6472 & ~w354;
assign w36754 = w2291 & pi2520;
assign w36755 = w2312 & pi2535;
assign w36756 = w6479 & ~w6476;
assign w36757 = ~w2370 & ~w6485;
assign w36758 = ~w3782 & w6489;
assign w36759 = w2667 & w6492;
assign w36760 = w2455 & pi0678;
assign w36761 = w6492 & ~w6494;
assign w36762 = w2481 & ~w2504;
assign w36763 = ~w36762 & ~w2474;
assign w36764 = ~w2537 & ~pi0512;
assign w36765 = w2537 & pi0512;
assign w36766 = ~w3917 & ~w3918;
assign w36767 = ~w6413 & w2397;
assign w36768 = w1311 & pi2698;
assign w36769 = w387 & pi2438;
assign w36770 = w400 & pi2701;
assign w36771 = w419 & pi2698;
assign w36772 = w410 & pi2275;
assign w36773 = ~w6534 & ~w354;
assign w36774 = ~w2941 & w6545;
assign w36775 = w567 & ~w553;
assign w36776 = w575 & ~w6552;
assign w36777 = pi0754 & ~pi0566;
assign w36778 = ~w6555 & w2958;
assign w36779 = ~w6474 & ~w2358;
assign w36780 = pi0403 & pi0406;
assign w36781 = w2377 & ~w6561;
assign w36782 = w6560 & w2365;
assign w36783 = pi0903 & pi2601;
assign w36784 = pi0903 & w35754;
assign w36785 = ~w933 & pi1029;
assign w36786 = ~w6567 & w6565;
assign w36787 = ~w6571 & ~w6570;
assign w36788 = ~w6432 & ~w2397;
assign w36789 = ~w6559 & w6574;
assign w36790 = ~w6496 & w3433;
assign w36791 = ~w702 & ~w715;
assign w36792 = ~w6586 & ~w715;
assign w36793 = ~w6586 & w36791;
assign w36794 = ~w575 & ~w6591;
assign w36795 = ~w344 & ~pi3257;
assign w36796 = pi0405 & ~pi0422;
assign w36797 = pi0403 & ~pi0418;
assign w36798 = ~w2352 & ~pi0419;
assign w36799 = ~w2361 & ~w6606;
assign w36800 = w35929 & w6607;
assign w36801 = ~pi3551 & pi3257;
assign w36802 = w6609 & pi2601;
assign w36803 = w6609 & w35754;
assign w36804 = ~w36801 & ~w6610;
assign w36805 = ~w36800 & w6611;
assign w36806 = w6614 & w6611;
assign w36807 = w6614 & w36805;
assign w36808 = ~w6600 & ~w36806;
assign w36809 = ~w6600 & ~w36807;
assign w36810 = w6616 & pi2601;
assign w36811 = w6616 & w35754;
assign w36812 = ~w2891 & ~w6617;
assign w36813 = w344 & ~w6620;
assign w36814 = ~pi3551 & pi3378;
assign w36815 = ~w2360 & ~w6622;
assign w36816 = w6624 & ~w36808;
assign w36817 = w6624 & ~w36809;
assign w36818 = w6631 & ~w938;
assign w36819 = w6631 & ~w35804;
assign w36820 = w6637 & ~w938;
assign w36821 = w6637 & ~w35804;
assign w36822 = w6633 & w6639;
assign w36823 = w6643 & ~w938;
assign w36824 = w6643 & ~w35804;
assign w36825 = w36822 & w6645;
assign w36826 = w6650 & ~w938;
assign w36827 = w6650 & ~w35804;
assign w36828 = w36822 & ~w6645;
assign w36829 = w6633 & ~w6639;
assign w36830 = w36829 & ~w6645;
assign w36831 = w6669 & ~w6621;
assign w36832 = ~w2352 & ~pi3390;
assign w36833 = pi3548 & pi0404;
assign w36834 = pi3528 & pi0684;
assign w36835 = ~pi3362 & ~w6679;
assign w36836 = w6682 & ~pi3551;
assign w36837 = ~pi3589 & ~pi0684;
assign w36838 = w2175 & w2195;
assign w36839 = pi0540 & w6690;
assign w36840 = ~w6734 & pi1930;
assign w36841 = pi3458 & ~pi1797;
assign w36842 = pi3641 & pi0405;
assign w36843 = w6973 & w6971;
assign w36844 = w6888 & ~w6976;
assign w36845 = w6753 & w6693;
assign w36846 = w6691 & w6687;
assign w36847 = ~pi0540 & w6982;
assign w36848 = w6888 & w6976;
assign w36849 = w36847 & w6983;
assign w36850 = w1031 & w1045;
assign w36851 = ~w6986 & ~w6985;
assign w36852 = w7003 & w7007;
assign w36853 = w2175 & ~w2195;
assign w36854 = w7052 & ~w7010;
assign w36855 = pi3433 & pi3457;
assign w36856 = pi3456 & pi3434;
assign w36857 = w36856 & pi3455;
assign w36858 = pi3454 & pi3453;
assign w36859 = w36858 & pi3432;
assign w36860 = w36859 & pi3459;
assign w36861 = pi3478 & pi3450;
assign w36862 = ~pi3478 & ~pi3450;
assign w36863 = w7053 & w7067;
assign w36864 = pi3236 & pi0815;
assign w36865 = ~w36863 & ~w7069;
assign w36866 = w36847 & w7050;
assign w36867 = ~w2175 & pi0540;
assign w36868 = ~w7077 & w6687;
assign w36869 = pi3402 & pi3404;
assign w36870 = pi3414 & pi3405;
assign w36871 = w36870 & pi3413;
assign w36872 = pi3406 & pi3411;
assign w36873 = w36872 & pi3420;
assign w36874 = w36873 & pi3401;
assign w36875 = pi3422 & pi3421;
assign w36876 = ~pi3422 & ~pi3421;
assign w36877 = w7091 & w6687;
assign w36878 = w7091 & w36868;
assign w36879 = ~w357 & ~w7097;
assign w36880 = pi3551 & pi0405;
assign w36881 = ~pi3551 & pi3512;
assign w36882 = ~w358 & ~w7103;
assign w36883 = ~w6686 & w7106;
assign w36884 = w36866 & pi0027;
assign w36885 = ~w36861 & ~pi3458;
assign w36886 = w36861 & pi3458;
assign w36887 = w7053 & w7113;
assign w36888 = w7003 & w7117;
assign w36889 = pi3236 & pi0814;
assign w36890 = ~w36888 & ~w7118;
assign w36891 = w1395 & w1030;
assign w36892 = w36849 & ~w7148;
assign w36893 = w36875 & pi3430;
assign w36894 = ~w36875 & ~pi3430;
assign w36895 = w7152 & w6687;
assign w36896 = w7152 & w36868;
assign w36897 = ~w357 & ~w7158;
assign w36898 = pi3551 & pi0421;
assign w36899 = ~pi3551 & pi3519;
assign w36900 = ~w358 & ~w7164;
assign w36901 = ~w6686 & w7167;
assign w36902 = ~w908 & w7174;
assign w36903 = w6677 & ~w938;
assign w36904 = ~w6674 & ~pi3682;
assign w36905 = w7182 & w7167;
assign w36906 = w7182 & w36901;
assign w36907 = w7188 & ~w938;
assign w36908 = w7188 & ~w35804;
assign w36909 = w7194 & ~w938;
assign w36910 = w7194 & ~w35804;
assign w36911 = ~w7190 & w7196;
assign w36912 = w7201 & ~w938;
assign w36913 = w7201 & ~w35804;
assign w36914 = w7213 & ~w938;
assign w36915 = w7213 & ~w35804;
assign w36916 = ~w7190 & ~w7196;
assign w36917 = ~pi0909 & ~pi1422;
assign w36918 = w344 & w7234;
assign w36919 = pi3551 & w6673;
assign w36920 = w7172 & pi0418;
assign w36921 = pi3520 & pi2785;
assign w36922 = pi3520 & w35556;
assign w36923 = pi1039 & pi1462;
assign w36924 = pi1039 & w35555;
assign w36925 = w185 & pi2540;
assign w36926 = pi3324 & ~pi0375;
assign w36927 = ~pi3324 & ~pi3496;
assign w36928 = w7242 & pi3626;
assign w36929 = pi1012 & pi1462;
assign w36930 = pi1012 & w35555;
assign w36931 = pi3511 & pi2785;
assign w36932 = pi3511 & w35556;
assign w36933 = w185 & pi2549;
assign w36934 = ~pi3324 & ~pi3497;
assign w36935 = pi3324 & ~pi0374;
assign w36936 = w7253 & pi3626;
assign w36937 = pi3510 & pi2785;
assign w36938 = pi3510 & w35556;
assign w36939 = pi1034 & pi1462;
assign w36940 = pi1034 & w35555;
assign w36941 = w185 & pi2646;
assign w36942 = pi3324 & ~pi0373;
assign w36943 = ~pi3324 & ~pi3495;
assign w36944 = w7264 & pi3626;
assign w36945 = pi1033 & pi1462;
assign w36946 = pi1033 & w35555;
assign w36947 = pi3521 & pi2785;
assign w36948 = pi3521 & w35556;
assign w36949 = w185 & pi2551;
assign w36950 = pi3324 & ~pi0372;
assign w36951 = ~pi3324 & ~pi3500;
assign w36952 = w7275 & pi3626;
assign w36953 = pi3509 & pi2785;
assign w36954 = pi3509 & w35556;
assign w36955 = pi1032 & pi1462;
assign w36956 = pi1032 & w35555;
assign w36957 = w185 & pi2553;
assign w36958 = pi3324 & ~pi0371;
assign w36959 = ~pi3324 & ~pi3499;
assign w36960 = w7286 & pi3626;
assign w36961 = pi1013 & pi1462;
assign w36962 = pi1013 & w35555;
assign w36963 = pi3508 & pi2785;
assign w36964 = pi3508 & w35556;
assign w36965 = w185 & pi2645;
assign w36966 = pi3324 & ~pi0369;
assign w36967 = ~pi3324 & ~pi3503;
assign w36968 = w7297 & pi3626;
assign w36969 = pi3517 & pi2785;
assign w36970 = pi3517 & w35556;
assign w36971 = pi1031 & pi1462;
assign w36972 = pi1031 & w35555;
assign w36973 = w185 & pi2797;
assign w36974 = ~pi3324 & ~pi3489;
assign w36975 = pi3324 & ~pi0380;
assign w36976 = w7308 & pi3626;
assign w36977 = pi3516 & pi2785;
assign w36978 = pi3516 & w35556;
assign w36979 = pi1030 & pi1462;
assign w36980 = pi1030 & w35555;
assign w36981 = w185 & pi2644;
assign w36982 = ~pi3324 & ~pi3492;
assign w36983 = pi3324 & ~pi0379;
assign w36984 = w7319 & pi3626;
assign w36985 = pi1029 & pi1462;
assign w36986 = pi1029 & w35555;
assign w36987 = pi3518 & pi2785;
assign w36988 = pi3518 & w35556;
assign w36989 = w185 & pi2796;
assign w36990 = w7330 & pi3626;
assign w36991 = pi1028 & pi1462;
assign w36992 = pi1028 & w35555;
assign w36993 = pi3514 & pi2785;
assign w36994 = pi3514 & w35556;
assign w36995 = w185 & pi2794;
assign w36996 = w7338 & pi3626;
assign w36997 = pi1038 & pi1462;
assign w36998 = pi1038 & w35555;
assign w36999 = pi3504 & pi2785;
assign w37000 = pi3504 & w35556;
assign w37001 = w185 & pi2788;
assign w37002 = w7346 & pi3626;
assign w37003 = pi1037 & pi1462;
assign w37004 = pi1037 & w35555;
assign w37005 = w185 & pi2953;
assign w37006 = ~w7362 & ~pi3449;
assign w37007 = ~pi3680 & pi3449;
assign w37008 = ~pi3680 & ~w37006;
assign w37009 = ~pi3680 & ~pi3449;
assign w37010 = w7362 & ~pi2408;
assign w37011 = ~w37010 & w7370;
assign w37012 = pi1036 & pi1462;
assign w37013 = pi1036 & w35555;
assign w37014 = w185 & w7377;
assign w37015 = ~pi3626 & ~w7373;
assign w37016 = pi3680 & w7386;
assign w37017 = ~pi3680 & ~pi2400;
assign w37018 = pi2981 & pi1462;
assign w37019 = pi2981 & w35555;
assign w37020 = w185 & w7393;
assign w37021 = ~w7383 & w7395;
assign w37022 = w7362 & ~w7364;
assign w37023 = w185 & w7401;
assign w37024 = w7402 & ~pi3680;
assign w37025 = ~w37022 & w7403;
assign w37026 = w7402 & ~w7410;
assign w37027 = ~w7411 & ~w7412;
assign w37028 = w185 & pi3624;
assign w37029 = ~pi3625 & ~w7417;
assign w37030 = ~w3590 & pi0574;
assign w37031 = w7420 & ~w941;
assign w37032 = pi2419 & w7433;
assign w37033 = w7427 & w7435;
assign w37034 = w7429 & w7437;
assign w37035 = w7427 & w7439;
assign w37036 = w7429 & w7443;
assign w37037 = w7430 & w7449;
assign w37038 = w7430 & w7451;
assign w37039 = ~w7472 & ~w7433;
assign w37040 = ~w7472 & ~w37032;
assign w37041 = ~w3711 & ~w7474;
assign w37042 = ~w4663 & pi0537;
assign w37043 = w7497 & ~w941;
assign w37044 = pi2419 & w7503;
assign w37045 = w7505 & pi3624;
assign w37046 = w7505 & w37028;
assign w37047 = ~w4749 & ~w7506;
assign w37048 = ~w5760 & pi0537;
assign w37049 = ~w5780 & pi0574;
assign w37050 = ~w7531 & ~w7529;
assign w37051 = ~w941 & ~pi2419;
assign w37052 = ~w37051 & w7535;
assign w37053 = w7537 & pi3624;
assign w37054 = w7537 & w37028;
assign w37055 = pi3625 & w5914;
assign w37056 = ~w5206 & pi0537;
assign w37057 = w7562 & ~w941;
assign w37058 = pi2419 & w7568;
assign w37059 = w7570 & pi3624;
assign w37060 = w7570 & w37028;
assign w37061 = ~w5320 & ~w7571;
assign w37062 = ~w4295 & pi0574;
assign w37063 = w7594 & ~w941;
assign w37064 = pi2419 & w7600;
assign w37065 = w7602 & pi3624;
assign w37066 = w7602 & w37028;
assign w37067 = ~w4380 & ~w7603;
assign w37068 = pi3625 & w6413;
assign w37069 = ~w6272 & pi0574;
assign w37070 = w7627 & ~w941;
assign w37071 = pi2419 & w7633;
assign w37072 = w7635 & pi3624;
assign w37073 = w7635 & w37028;
assign w37074 = pi3625 & w40134;
assign w37075 = ~w3364 & pi0574;
assign w37076 = w7660 & ~w941;
assign w37077 = pi2419 & w7666;
assign w37078 = w7668 & pi3624;
assign w37079 = w7668 & w37028;
assign w37080 = ~w3085 & pi0574;
assign w37081 = w7692 & ~w941;
assign w37082 = pi2419 & w7698;
assign w37083 = w7700 & pi3624;
assign w37084 = w7700 & w37028;
assign w37085 = ~w3195 & ~w7701;
assign w37086 = ~w6108 & pi0574;
assign w37087 = ~w1184 & pi0537;
assign w37088 = ~w7726 & ~w7724;
assign w37089 = ~w37051 & w7730;
assign w37090 = w7732 & pi3624;
assign w37091 = w7732 & w37028;
assign w37092 = ~w6177 & ~w7733;
assign w37093 = ~w7757 & ~w7756;
assign w37094 = ~w37051 & w7762;
assign w37095 = w7764 & pi3624;
assign w37096 = w7764 & w37028;
assign w37097 = ~w4141 & ~w7765;
assign w37098 = ~w4955 & pi0574;
assign w37099 = w7788 & ~w941;
assign w37100 = pi2419 & w7794;
assign w37101 = w7796 & pi3624;
assign w37102 = w7796 & w37028;
assign w37103 = ~w5053 & ~w7797;
assign w37104 = w7820 & ~w941;
assign w37105 = pi2419 & w7826;
assign w37106 = w7828 & pi3624;
assign w37107 = w7828 & w37028;
assign w37108 = ~w5635 & ~w7829;
assign w37109 = ~w1125 & pi0574;
assign w37110 = ~w7854 & ~w7852;
assign w37111 = ~w37051 & w7858;
assign w37112 = w7860 & pi3624;
assign w37113 = w7860 & w37028;
assign w37114 = ~w1308 & ~w7861;
assign w37115 = w7884 & ~w941;
assign w37116 = pi2419 & w7890;
assign w37117 = w7892 & pi3624;
assign w37118 = w7892 & w37028;
assign w37119 = pi3625 & w1639;
assign w37120 = ~w7971 & pi0574;
assign w37121 = ~w37051 & w7992;
assign w37122 = w7994 & pi3624;
assign w37123 = w7994 & w37028;
assign w37124 = w977 & pi3889;
assign w37125 = w979 & pi3985;
assign w37126 = w971 & pi3857;
assign w37127 = w964 & pi3953;
assign w37128 = w955 & pi3937;
assign w37129 = w960 & pi3921;
assign w37130 = w974 & pi3905;
assign w37131 = w966 & pi3969;
assign w37132 = ~pi3515 & pi3314;
assign w37133 = w1226 & pi2987;
assign w37134 = w8064 & pi0650;
assign w37135 = w8014 & ~pi1787;
assign w37136 = w952 & ~w8078;
assign w37137 = w8079 & pi1787;
assign w37138 = w8079 & ~w37135;
assign w37139 = pi3625 & w8081;
assign w37140 = w977 & pi3890;
assign w37141 = w979 & pi3986;
assign w37142 = w971 & pi3858;
assign w37143 = w966 & pi3970;
assign w37144 = w955 & pi3938;
assign w37145 = w964 & pi3954;
assign w37146 = w974 & pi3906;
assign w37147 = w960 & pi3922;
assign w37148 = ~pi3515 & pi3313;
assign w37149 = w1226 & pi3097;
assign w37150 = w8186 & pi0650;
assign w37151 = ~w8217 & pi0576;
assign w37152 = ~w8233 & ~w941;
assign w37153 = ~w8234 & ~w8106;
assign w37154 = w952 & ~w8237;
assign w37155 = pi1787 & w8238;
assign w37156 = pi3625 & w8240;
assign w37157 = ~w8217 & pi0574;
assign w37158 = w8258 & ~w941;
assign w37159 = pi2419 & w8264;
assign w37160 = w8266 & pi3624;
assign w37161 = w8266 & w37028;
assign w37162 = pi0434 & pi3641;
assign w37163 = pi0433 & pi3641;
assign w37164 = ~pi0358 & pi3641;
assign w37165 = pi0431 & pi3641;
assign w37166 = pi0430 & pi3641;
assign w37167 = ~pi0355 & pi3641;
assign w37168 = pi0428 & pi3641;
assign w37169 = ~pi0353 & pi3641;
assign w37170 = ~w4744 & w941;
assign w37171 = ~w4744 & ~w37043;
assign w37172 = w941 & ~w5673;
assign w37173 = ~w5093 & w941;
assign w37174 = ~w5093 & ~w37057;
assign w37175 = ~w4161 & w941;
assign w37176 = ~w4161 & ~w37063;
assign w37177 = ~pi3515 & pi3309;
assign w37178 = ~w2980 & w941;
assign w37179 = ~w2980 & ~w37081;
assign w37180 = w941 & ~w5988;
assign w37181 = w941 & ~w3955;
assign w37182 = ~pi3515 & pi3295;
assign w37183 = ~w8374 & w941;
assign w37184 = ~w8374 & ~w37104;
assign w37185 = w941 & ~w1003;
assign w37186 = w941 & ~w8014;
assign w37187 = ~w346 & w825;
assign w37188 = ~w346 & w822;
assign w37189 = w346 & w6618;
assign w37190 = w8414 & ~w8416;
assign w37191 = w8414 & ~w8424;
assign w37192 = w5673 & ~w8414;
assign w37193 = ~w8432 & w8414;
assign w37194 = ~w8432 & ~w37192;
assign w37195 = w8414 & ~w8440;
assign w37196 = w8414 & ~w8448;
assign w37197 = w6409 & ~w8414;
assign w37198 = w8414 & ~w8465;
assign w37199 = w8414 & ~w8473;
assign w37200 = w8414 & ~w8481;
assign w37201 = w8414 & ~w8489;
assign w37202 = w8414 & ~w8497;
assign w37203 = w5631 & ~w8414;
assign w37204 = w8414 & ~w8514;
assign w37205 = w8414 & ~w8522;
assign w37206 = w8014 & ~w8414;
assign w37207 = ~w8530 & w8414;
assign w37208 = ~w8530 & ~w37206;
assign w37209 = w8414 & ~w8538;
assign w37210 = ~w792 & w788;
assign w37211 = ~w607 & ~w8543;
assign w37212 = pi0641 & ~pi0568;
assign w37213 = w756 & w8546;
assign w37214 = w789 & w8545;
assign w37215 = ~w8553 & ~w8551;
assign w37216 = ~w8554 & pi0641;
assign w37217 = ~pi0641 & ~w501;
assign w37218 = w8556 & ~w8543;
assign w37219 = w3484 & w874;
assign w37220 = w874 & ~w8559;
assign w37221 = w387 & pi2270;
assign w37222 = w419 & pi2437;
assign w37223 = w400 & pi2447;
assign w37224 = w410 & pi1985;
assign w37225 = w423 & w8569;
assign w37226 = pi0873 & pi2601;
assign w37227 = pi0873 & w35754;
assign w37228 = w8572 & ~pi1422;
assign w37229 = w8572 & w35753;
assign w37230 = ~pi3515 & pi2554;
assign w37231 = ~w8573 & ~w37228;
assign w37232 = ~w8573 & ~w37229;
assign w37233 = w8574 & w905;
assign w37234 = w364 & ~w8576;
assign w37235 = w1311 & pi2437;
assign w37236 = pi0667 & pi0641;
assign w37237 = ~w37236 & ~w8590;
assign w37238 = ~w597 & ~w8590;
assign w37239 = ~w597 & w37237;
assign w37240 = ~w8593 & ~w505;
assign w37241 = w8593 & pi0665;
assign w37242 = ~w575 & w8596;
assign w37243 = w504 & pi0665;
assign w37244 = w575 & w8600;
assign w37245 = w387 & pi2267;
assign w37246 = w400 & pi2444;
assign w37247 = w419 & pi2434;
assign w37248 = w410 & pi1982;
assign w37249 = ~w424 & w8611;
assign w37250 = w1311 & pi2434;
assign w37251 = ~w933 & pi2549;
assign w37252 = pi0908 & pi2601;
assign w37253 = pi0908 & w35754;
assign w37254 = w8623 & ~pi1422;
assign w37255 = w8623 & w35753;
assign w37256 = ~pi3515 & pi2559;
assign w37257 = ~w8624 & ~w37254;
assign w37258 = ~w8624 & ~w37255;
assign w37259 = w8625 & w905;
assign w37260 = ~w8626 & ~w8621;
assign w37261 = pi0907 & pi2601;
assign w37262 = pi0907 & w35754;
assign w37263 = ~w933 & pi2646;
assign w37264 = ~pi3515 & pi2705;
assign w37265 = ~w8636 & ~w8634;
assign w37266 = w364 & ~w8639;
assign w37267 = w1311 & pi2433;
assign w37268 = w510 & pi0664;
assign w37269 = w575 & w8655;
assign w37270 = w8659 & ~w8661;
assign w37271 = ~w575 & w8663;
assign w37272 = w874 & ~w8666;
assign w37273 = w419 & pi2433;
assign w37274 = w410 & pi1981;
assign w37275 = w387 & pi2266;
assign w37276 = w400 & pi2274;
assign w37277 = w423 & w8676;
assign w37278 = w575 & w8679;
assign w37279 = ~pi0663 & ~w8679;
assign w37280 = ~pi0663 & ~w37278;
assign w37281 = w8679 & w522;
assign w37282 = w623 & ~w595;
assign w37283 = w623 & w35672;
assign w37284 = w610 & ~w8682;
assign w37285 = ~w623 & w595;
assign w37286 = ~w623 & ~w35672;
assign w37287 = ~w622 & ~w37285;
assign w37288 = ~w622 & ~w37286;
assign w37289 = ~w610 & ~w8687;
assign w37290 = ~w514 & ~w8684;
assign w37291 = w628 & ~w8690;
assign w37292 = ~w8689 & ~w8686;
assign w37293 = ~w575 & w8695;
assign w37294 = w8680 & ~w8696;
assign w37295 = w5092 & w874;
assign w37296 = w874 & ~w8698;
assign w37297 = w387 & pi2265;
assign w37298 = w400 & pi2443;
assign w37299 = w419 & pi2260;
assign w37300 = w846 & pi1980;
assign w37301 = w423 & w8709;
assign w37302 = pi0874 & pi2601;
assign w37303 = pi0874 & w35754;
assign w37304 = w8712 & ~pi1422;
assign w37305 = w8712 & w35753;
assign w37306 = ~pi3515 & pi2556;
assign w37307 = ~w8713 & ~w37304;
assign w37308 = ~w8713 & ~w37305;
assign w37309 = w8714 & w905;
assign w37310 = w364 & ~w8716;
assign w37311 = w1311 & pi2260;
assign w37312 = ~w575 & ~w8733;
assign w37313 = w575 & w8741;
assign w37314 = w4160 & w874;
assign w37315 = w874 & ~w8744;
assign w37316 = w387 & pi2264;
assign w37317 = w419 & pi2259;
assign w37318 = w400 & pi2273;
assign w37319 = w410 & pi1979;
assign w37320 = w423 & w8754;
assign w37321 = pi0906 & pi2601;
assign w37322 = pi0906 & w35754;
assign w37323 = w8757 & ~pi1422;
assign w37324 = w8757 & w35753;
assign w37325 = ~pi3515 & pi2704;
assign w37326 = ~w8758 & ~w37323;
assign w37327 = ~w8758 & ~w37324;
assign w37328 = w8759 & w905;
assign w37329 = w364 & ~w8761;
assign w37330 = w1311 & pi2259;
assign w37331 = ~w424 & w8776;
assign w37332 = ~w933 & pi2645;
assign w37333 = ~w6458 & ~w8778;
assign w37334 = w364 & ~w8782;
assign w37335 = ~w933 & pi2797;
assign w37336 = ~w2900 & ~w8791;
assign w37337 = w364 & ~w8795;
assign w37338 = w874 & ~w8801;
assign w37339 = w423 & w8804;
assign w37340 = ~w424 & w8808;
assign w37341 = ~w933 & pi2644;
assign w37342 = ~w4429 & ~w8810;
assign w37343 = w364 & ~w8814;
assign w37344 = w5987 & w874;
assign w37345 = w874 & ~w8825;
assign w37346 = w423 & w8828;
assign w37347 = ~w933 & pi2796;
assign w37348 = w6566 & ~pi1422;
assign w37349 = w6566 & w35753;
assign w37350 = ~w6564 & ~w37348;
assign w37351 = ~w6564 & ~w37349;
assign w37352 = w8832 & w905;
assign w37353 = ~w424 & w8841;
assign w37354 = ~w933 & pi2794;
assign w37355 = ~w3884 & ~w8843;
assign w37356 = w364 & ~w8847;
assign w37357 = ~w424 & w8857;
assign w37358 = ~w933 & pi2788;
assign w37359 = ~w5061 & ~w8859;
assign w37360 = w364 & ~w8863;
assign w37361 = w5407 & w424;
assign w37362 = ~w933 & pi2953;
assign w37363 = ~w5923 & ~w8876;
assign w37364 = w364 & ~w8880;
assign w37365 = ~w8585 & w2417;
assign w37366 = ~w3762 & w2363;
assign w37367 = pi0403 & pi0408;
assign w37368 = ~w2361 & w8896;
assign w37369 = ~w37368 & ~w8573;
assign w37370 = ~w933 & pi1039;
assign w37371 = ~w3433 & w8907;
assign w37372 = ~w3790 & w2941;
assign w37373 = w1639 & w2397;
assign w37374 = ~w4472 & ~w2358;
assign w37375 = ~w8605 & ~w354;
assign w37376 = pi0403 & pi0413;
assign w37377 = w2377 & ~w8924;
assign w37378 = w8921 & w2365;
assign w37379 = w8623 & pi1422;
assign w37380 = w8623 & w36132;
assign w37381 = ~w8624 & ~w37379;
assign w37382 = ~w8624 & ~w37380;
assign w37383 = ~w8929 & ~w2899;
assign w37384 = ~w8931 & ~w8930;
assign w37385 = w4771 & ~w2397;
assign w37386 = ~w3433 & w8934;
assign w37387 = ~w8941 & w2397;
assign w37388 = ~w3440 & ~w8943;
assign w37389 = ~w5940 & ~w2358;
assign w37390 = ~w8673 & ~w354;
assign w37391 = pi0403 & pi0412;
assign w37392 = w2377 & ~w8950;
assign w37393 = w8947 & w2365;
assign w37394 = w8633 & pi1422;
assign w37395 = w8633 & w36132;
assign w37396 = ~w8636 & ~w37394;
assign w37397 = ~w8636 & ~w37395;
assign w37398 = ~w8955 & ~w2899;
assign w37399 = ~w8957 & ~w8956;
assign w37400 = ~w3433 & w8959;
assign w37401 = ~w2941 & w8969;
assign w37402 = ~w2397 & ~w8971;
assign w37403 = pi0403 & pi0411;
assign w37404 = ~w5350 & ~w2358;
assign w37405 = w8975 & w2365;
assign w37406 = ~w8725 & w2417;
assign w37407 = ~w933 & pi1033;
assign w37408 = ~w8982 & w8981;
assign w37409 = ~w8987 & ~w8986;
assign w37410 = ~w3433 & w8989;
assign w37411 = ~w5333 & w2941;
assign w37412 = w5053 & w2397;
assign w37413 = ~w2941 & w9012;
assign w37414 = pi0403 & pi0410;
assign w37415 = ~w8770 & ~w2377;
assign w37416 = w9016 & w2365;
assign w37417 = ~pi1032 & ~w9021;
assign w37418 = ~w9026 & ~w9025;
assign w37419 = ~w3863 & ~w2397;
assign w37420 = ~w2958 & w9029;
assign w37421 = w36866 & pi0014;
assign w37422 = w7053 & ~pi3460;
assign w37423 = w7003 & w9038;
assign w37424 = pi3236 & pi0818;
assign w37425 = ~w37423 & ~w9039;
assign w37426 = ~pi3400 & w6687;
assign w37427 = ~pi3400 & w36868;
assign w37428 = w1734 & pi0976;
assign w37429 = w9051 & ~w9044;
assign w37430 = pi3551 & pi0408;
assign w37431 = ~pi3551 & pi3520;
assign w37432 = ~w358 & ~w9070;
assign w37433 = ~w357 & ~w9074;
assign w37434 = ~w6686 & w9076;
assign w37435 = w1669 & pi0976;
assign w37436 = w36849 & ~w9105;
assign w37437 = w7053 & w9108;
assign w37438 = w7003 & w9112;
assign w37439 = pi3236 & pi0813;
assign w37440 = ~w37438 & ~w9113;
assign w37441 = w9118 & w6687;
assign w37442 = w9118 & w36868;
assign w37443 = w36866 & pi0015;
assign w37444 = pi3551 & pi0413;
assign w37445 = ~pi3551 & pi3511;
assign w37446 = ~w358 & ~w9128;
assign w37447 = ~w357 & ~w9132;
assign w37448 = ~w6686 & w9134;
assign w37449 = w36866 & pi0016;
assign w37450 = w7053 & w9139;
assign w37451 = w7003 & w9143;
assign w37452 = pi3236 & pi0812;
assign w37453 = ~pi3589 & pi0684;
assign w37454 = ~w37451 & w9152;
assign w37455 = w9157 & w6687;
assign w37456 = w9157 & w36868;
assign w37457 = w1928 & pi0976;
assign w37458 = w36849 & ~w9179;
assign w37459 = pi3551 & pi0412;
assign w37460 = ~pi3551 & pi3510;
assign w37461 = ~w358 & ~w9188;
assign w37462 = ~w357 & ~w9192;
assign w37463 = ~w6686 & w9194;
assign w37464 = w36866 & pi0017;
assign w37465 = ~pi3433 & ~pi3457;
assign w37466 = w7053 & w9199;
assign w37467 = w7003 & w9203;
assign w37468 = pi3236 & pi0811;
assign w37469 = ~w37467 & w9209;
assign w37470 = ~pi3402 & ~pi3404;
assign w37471 = w9214 & w6687;
assign w37472 = w9214 & w36868;
assign w37473 = w2003 & w1024;
assign w37474 = w36849 & ~w9236;
assign w37475 = pi3551 & pi0411;
assign w37476 = ~pi3551 & pi3521;
assign w37477 = ~w358 & ~w9245;
assign w37478 = ~w357 & ~w9249;
assign w37479 = ~w6686 & w9251;
assign w37480 = w36849 & ~w9278;
assign w37481 = w7003 & w9282;
assign w37482 = w7053 & w9285;
assign w37483 = pi3236 & pi0810;
assign w37484 = ~w37482 & w9291;
assign w37485 = w9296 & w6687;
assign w37486 = w9296 & w36868;
assign w37487 = w36866 & pi0018;
assign w37488 = pi3551 & pi0410;
assign w37489 = ~pi3551 & pi3509;
assign w37490 = ~w358 & ~w9306;
assign w37491 = ~w357 & ~w9310;
assign w37492 = ~w6686 & w9312;
assign w37493 = w2118 & w1045;
assign w37494 = w9319 & ~w9316;
assign w37495 = w36849 & ~w9326;
assign w37496 = w7003 & w9330;
assign w37497 = ~pi3456 & ~pi3434;
assign w37498 = w7053 & w9333;
assign w37499 = pi3236 & pi0809;
assign w37500 = ~w37498 & w9339;
assign w37501 = ~pi3414 & ~pi3405;
assign w37502 = w9344 & w6687;
assign w37503 = w9344 & w36868;
assign w37504 = w36866 & pi0019;
assign w37505 = pi3551 & pi0409;
assign w37506 = ~pi3551 & pi3508;
assign w37507 = ~w358 & ~w9354;
assign w37508 = ~w357 & ~w9358;
assign w37509 = ~w6686 & w9360;
assign w37510 = ~w1775 & pi0976;
assign w37511 = ~w9364 & ~w9363;
assign w37512 = ~w36856 & ~pi3455;
assign w37513 = w7053 & w9379;
assign w37514 = w7003 & w9383;
assign w37515 = pi3236 & pi0808;
assign w37516 = ~w37514 & ~w9384;
assign w37517 = ~w36870 & ~pi3413;
assign w37518 = w9389 & w6687;
assign w37519 = w9389 & w36868;
assign w37520 = w36866 & pi0020;
assign w37521 = pi3551 & pi0426;
assign w37522 = ~pi3551 & pi3517;
assign w37523 = ~w358 & ~w9399;
assign w37524 = ~w357 & ~w9403;
assign w37525 = ~w6686 & w9405;
assign w37526 = w36849 & ~w9427;
assign w37527 = w7053 & w9430;
assign w37528 = w7003 & w9434;
assign w37529 = pi3236 & pi0807;
assign w37530 = ~w37528 & ~w9435;
assign w37531 = w9440 & w6687;
assign w37532 = w9440 & w36868;
assign w37533 = w36866 & pi0021;
assign w37534 = pi3551 & pi0425;
assign w37535 = ~pi3551 & pi3516;
assign w37536 = ~w358 & ~w9450;
assign w37537 = ~w357 & ~w9454;
assign w37538 = ~w6686 & w9456;
assign w37539 = w36849 & ~w9489;
assign w37540 = ~pi3454 & ~pi3453;
assign w37541 = w7053 & w9492;
assign w37542 = w7003 & w9496;
assign w37543 = pi3236 & pi0806;
assign w37544 = ~w37542 & ~w9497;
assign w37545 = ~pi3406 & ~pi3411;
assign w37546 = w9502 & w6687;
assign w37547 = w9502 & w36868;
assign w37548 = w36866 & pi0022;
assign w37549 = pi3551 & pi0406;
assign w37550 = ~pi3551 & pi3518;
assign w37551 = ~w358 & ~w9512;
assign w37552 = ~w357 & ~w9516;
assign w37553 = ~w6686 & w9518;
assign w37554 = w36849 & ~w9535;
assign w37555 = ~w36858 & ~pi3432;
assign w37556 = w7053 & w9538;
assign w37557 = w7003 & w9542;
assign w37558 = pi3236 & pi0788;
assign w37559 = ~w37557 & ~w9543;
assign w37560 = ~w36872 & ~pi3420;
assign w37561 = w9548 & w6687;
assign w37562 = w9548 & w36868;
assign w37563 = w36866 & pi0023;
assign w37564 = pi3551 & pi0424;
assign w37565 = ~pi3551 & pi3514;
assign w37566 = ~w358 & ~w9558;
assign w37567 = ~w357 & ~w9562;
assign w37568 = ~w6686 & w9564;
assign w37569 = w36849 & ~w9588;
assign w37570 = ~w36859 & ~pi3459;
assign w37571 = w7053 & w9591;
assign w37572 = w7003 & w9595;
assign w37573 = pi3236 & pi0817;
assign w37574 = ~w37572 & ~w9596;
assign w37575 = ~w36873 & ~pi3401;
assign w37576 = w9601 & w6687;
assign w37577 = w9601 & w36868;
assign w37578 = w36866 & pi0024;
assign w37579 = pi3551 & pi0423;
assign w37580 = ~pi3551 & pi3504;
assign w37581 = ~w358 & ~w9611;
assign w37582 = ~w357 & ~w9615;
assign w37583 = ~w6686 & w9617;
assign w37584 = w36866 & pi0025;
assign w37585 = w7053 & w9622;
assign w37586 = w7003 & w9626;
assign w37587 = ~w37586 & ~w9627;
assign w37588 = w9632 & w6687;
assign w37589 = w9632 & w36868;
assign w37590 = w36849 & ~w9662;
assign w37591 = pi3551 & pi0422;
assign w37592 = ~pi3551 & pi3513;
assign w37593 = ~w358 & ~w9671;
assign w37594 = ~w357 & ~w9675;
assign w37595 = ~w6686 & w9677;
assign w37596 = ~pi0844 & ~w938;
assign w37597 = ~pi0433 & pi2601;
assign w37598 = ~pi0433 & w35754;
assign w37599 = ~pi0843 & ~w938;
assign w37600 = ~pi0432 & pi2601;
assign w37601 = ~pi0432 & w35754;
assign w37602 = ~pi0842 & ~w938;
assign w37603 = ~pi0431 & pi2601;
assign w37604 = ~pi0431 & w35754;
assign w37605 = ~pi0864 & ~w938;
assign w37606 = ~pi0430 & pi2601;
assign w37607 = ~pi0430 & w35754;
assign w37608 = ~pi0841 & ~w938;
assign w37609 = ~pi0429 & pi2601;
assign w37610 = ~pi0429 & w35754;
assign w37611 = ~pi0865 & ~w938;
assign w37612 = ~pi0428 & pi2601;
assign w37613 = ~pi0428 & w35754;
assign w37614 = ~pi0840 & ~w938;
assign w37615 = ~pi0435 & pi2601;
assign w37616 = ~pi0435 & w35754;
assign w37617 = ~pi0839 & ~w938;
assign w37618 = ~pi0366 & pi2601;
assign w37619 = ~pi0366 & w35754;
assign w37620 = ~pi1092 & ~w938;
assign w37621 = ~pi0359 & pi2601;
assign w37622 = ~pi0359 & w35754;
assign w37623 = ~pi1060 & ~w938;
assign w37624 = ~pi0358 & pi2601;
assign w37625 = ~pi0358 & w35754;
assign w37626 = ~pi1089 & ~w938;
assign w37627 = ~pi0357 & pi2601;
assign w37628 = ~pi0357 & w35754;
assign w37629 = ~pi1065 & ~w938;
assign w37630 = ~pi0356 & pi2601;
assign w37631 = ~pi0356 & w35754;
assign w37632 = ~pi1064 & ~w938;
assign w37633 = ~pi0355 & pi2601;
assign w37634 = ~pi0355 & w35754;
assign w37635 = ~pi1063 & ~w938;
assign w37636 = ~pi0354 & pi2601;
assign w37637 = ~pi0354 & w35754;
assign w37638 = ~pi1062 & ~w938;
assign w37639 = ~pi0353 & pi2601;
assign w37640 = ~pi0353 & w35754;
assign w37641 = ~pi1061 & ~w938;
assign w37642 = ~pi0352 & pi2601;
assign w37643 = ~pi0352 & w35754;
assign w37644 = ~pi3106 & ~w938;
assign w37645 = ~pi0351 & pi2601;
assign w37646 = ~pi0351 & w35754;
assign w37647 = ~pi3105 & ~w938;
assign w37648 = ~pi0365 & pi2601;
assign w37649 = ~pi0365 & w35754;
assign w37650 = ~pi3104 & ~w938;
assign w37651 = ~pi0364 & pi2601;
assign w37652 = ~pi0364 & w35754;
assign w37653 = ~pi2985 & ~w938;
assign w37654 = ~pi0363 & pi2601;
assign w37655 = ~pi0363 & w35754;
assign w37656 = ~pi3102 & ~w938;
assign w37657 = ~pi0362 & pi2601;
assign w37658 = ~pi0362 & w35754;
assign w37659 = ~pi3109 & ~w938;
assign w37660 = ~pi0361 & pi2601;
assign w37661 = ~pi0361 & w35754;
assign w37662 = ~pi3111 & ~w938;
assign w37663 = ~pi0360 & pi2601;
assign w37664 = ~pi0360 & w35754;
assign w37665 = ~pi3112 & ~w938;
assign w37666 = w6682 & ~pi3460;
assign w37667 = w6682 & ~pi3437;
assign w37668 = w6682 & ~pi3433;
assign w37669 = w6682 & ~pi3457;
assign w37670 = w6682 & ~pi3456;
assign w37671 = ~pi3114 & ~pi0038;
assign w37672 = ~pi3114 & w35924;
assign w37673 = ~pi2952 & ~pi0038;
assign w37674 = ~pi2952 & w35924;
assign w37675 = pi3551 & pi3121;
assign w37676 = ~pi3076 & ~w2214;
assign w37677 = pi2951 & ~pi3195;
assign w37678 = ~pi2951 & ~w9038;
assign w37679 = ~pi2951 & ~w9112;
assign w37680 = pi2951 & ~pi3124;
assign w37681 = ~w37680 & pi2763;
assign w37682 = ~pi2951 & ~w9143;
assign w37683 = pi2951 & ~pi3194;
assign w37684 = ~w37683 & pi2763;
assign w37685 = ~pi2951 & ~w9203;
assign w37686 = pi2951 & ~pi3139;
assign w37687 = ~w37686 & pi2763;
assign w37688 = ~pi2951 & ~w9282;
assign w37689 = pi2951 & ~pi3135;
assign w37690 = ~w37689 & pi2763;
assign w37691 = ~pi2951 & ~w9330;
assign w37692 = pi2951 & ~pi3187;
assign w37693 = ~w37692 & pi2763;
assign w37694 = pi2951 & ~pi3193;
assign w37695 = ~pi2951 & ~w9383;
assign w37696 = pi2951 & ~pi3192;
assign w37697 = ~pi2951 & ~w9434;
assign w37698 = pi2951 & ~pi3117;
assign w37699 = ~pi2951 & ~w9496;
assign w37700 = ~pi2951 & ~w9542;
assign w37701 = pi2951 & ~pi3116;
assign w37702 = ~w37701 & pi2763;
assign w37703 = ~pi2951 & ~w9595;
assign w37704 = pi2951 & ~pi3198;
assign w37705 = ~w37704 & pi2763;
assign w37706 = ~pi2951 & ~w9626;
assign w37707 = pi2951 & ~pi3115;
assign w37708 = ~w37707 & pi2763;
assign w37709 = ~pi2951 & ~w7007;
assign w37710 = pi2951 & ~pi3197;
assign w37711 = ~w37710 & pi2763;
assign w37712 = ~pi2951 & ~w7117;
assign w37713 = pi2951 & ~pi3196;
assign w37714 = pi3509 & w9951;
assign w37715 = w9936 & ~w9953;
assign w37716 = ~w9957 & w9961;
assign w37717 = ~w9965 & w9961;
assign w37718 = ~w9965 & w37716;
assign w37719 = pi1975 & pi3065;
assign w37720 = pi1972 & pi1974;
assign w37721 = w9971 & ~w9981;
assign w37722 = ~w9996 & ~w9988;
assign w37723 = w9996 & w9988;
assign w37724 = w10015 & ~w10025;
assign w37725 = w10031 & w9987;
assign w37726 = ~w10031 & w9988;
assign w37727 = ~pi2982 & pi1793;
assign w37728 = ~w10049 & w9990;
assign w37729 = ~w37728 & w9988;
assign w37730 = w37728 & w9987;
assign w37731 = w10064 & ~w10074;
assign w37732 = ~w10080 & ~w9988;
assign w37733 = w10080 & w9988;
assign w37734 = w10044 & ~w10013;
assign w37735 = ~w10061 & ~w10099;
assign w37736 = w37735 & pi0828;
assign w37737 = w10097 & w10101;
assign w37738 = ~w10013 & w10100;
assign w37739 = w10111 & ~w10121;
assign w37740 = ~w10127 & ~w9988;
assign w37741 = w10127 & w9988;
assign w37742 = ~w9937 & ~pi3508;
assign w37743 = ~pi3509 & w9951;
assign w37744 = w10161 & w9987;
assign w37745 = ~w10161 & w9988;
assign w37746 = w10178 & w9990;
assign w37747 = w9988 & ~w9995;
assign w37748 = w10194 & ~w10204;
assign w37749 = ~w9933 & ~pi3508;
assign w37750 = w10218 & ~w10219;
assign w37751 = w10230 & w9987;
assign w37752 = ~w10230 & w9988;
assign w37753 = w10246 & ~w10256;
assign w37754 = ~pi2982 & pi2198;
assign w37755 = w10262 & w9988;
assign w37756 = ~w10262 & w10274;
assign w37757 = pi3518 & pi3516;
assign w37758 = ~w10282 & ~w10278;
assign w37759 = w10296 & ~w10306;
assign w37760 = ~pi3509 & ~pi3508;
assign w37761 = ~w9930 & ~w9951;
assign w37762 = ~w10317 & w10316;
assign w37763 = ~pi2982 & pi2200;
assign w37764 = w10331 & w9988;
assign w37765 = ~w10331 & w10274;
assign w37766 = ~w10350 & w9961;
assign w37767 = ~w10350 & w37716;
assign w37768 = w10344 & ~w10353;
assign w37769 = w10312 & ~w10277;
assign w37770 = ~w10243 & ~w10277;
assign w37771 = ~w10243 & w37769;
assign w37772 = ~w10359 & ~w10210;
assign w37773 = ~pi2982 & pi2196;
assign w37774 = w10380 & w9988;
assign w37775 = ~w10380 & w10274;
assign w37776 = ~w10394 & ~w10393;
assign w37777 = w10174 & w10398;
assign w37778 = w10401 & ~w10398;
assign w37779 = w10401 & ~w37777;
assign w37780 = ~pi2982 & pi2194;
assign w37781 = w10408 & ~w10404;
assign w37782 = w10439 & w9969;
assign w37783 = w10446 & ~w10456;
assign w37784 = ~w10462 & ~w9988;
assign w37785 = w10462 & w9988;
assign w37786 = w10478 & ~w10488;
assign w37787 = ~pi2982 & pi2081;
assign w37788 = w10494 & w9988;
assign w37789 = ~w10494 & w10274;
assign w37790 = w10509 & ~w10519;
assign w37791 = ~w10525 & ~w9988;
assign w37792 = w10525 & w9988;
assign w37793 = w10543 & w10476;
assign w37794 = ~w10544 & w10551;
assign w37795 = ~w4523 & ~pi0835;
assign w37796 = pi1620 & ~pi1041;
assign w37797 = ~w37795 & ~w10577;
assign w37798 = w10061 & ~w10099;
assign w37799 = ~w10540 & w10106;
assign w37800 = w10098 & w10583;
assign w37801 = ~pi0828 & w10578;
assign w37802 = w10140 & w10589;
assign w37803 = ~w10098 & w10100;
assign w37804 = w10061 & ~w10594;
assign w37805 = w10061 & w10593;
assign w37806 = w10597 & w10099;
assign w37807 = w10098 & w10596;
assign w37808 = w10061 & ~w10605;
assign w37809 = w10106 & w10606;
assign w37810 = w10140 & w10607;
assign w37811 = ~w10098 & w10606;
assign w37812 = ~pi1824 & ~pi0038;
assign w37813 = ~pi1824 & w35924;
assign w37814 = ~pi3426 & ~pi2142;
assign w37815 = ~w10615 & ~w10577;
assign w37816 = ~w10615 & w37797;
assign w37817 = ~w10588 & w10618;
assign w37818 = w10106 & ~w10620;
assign w37819 = w10140 & w10622;
assign w37820 = ~pi0835 & w36655;
assign w37821 = ~pi0835 & w36654;
assign w37822 = w10628 & ~pi1041;
assign w37823 = ~pi1570 & pi1041;
assign w37824 = ~w10634 & w10633;
assign w37825 = ~w10626 & ~w10639;
assign w37826 = ~w10640 & ~w37821;
assign w37827 = ~w10640 & ~w37820;
assign w37828 = w10642 & w10643;
assign w37829 = ~w10642 & w10648;
assign w37830 = ~w10588 & ~w10616;
assign w37831 = w10642 & w10653;
assign w37832 = ~w10642 & w10655;
assign w37833 = ~w10544 & w10550;
assign w37834 = ~w10106 & w10663;
assign w37835 = w37814 & ~w10099;
assign w37836 = ~w10062 & w10665;
assign w37837 = ~w5092 & ~pi0835;
assign w37838 = pi1516 & ~pi1041;
assign w37839 = pi1569 & pi1041;
assign w37840 = ~w10674 & w10673;
assign w37841 = ~w10626 & w10679;
assign w37842 = ~w37837 & ~w10680;
assign w37843 = ~w370 & ~w10626;
assign w37844 = ~w37843 & ~w10686;
assign w37845 = ~w370 & w10691;
assign w37846 = ~w4160 & ~pi0835;
assign w37847 = pi1480 & ~pi1041;
assign w37848 = pi1552 & pi1041;
assign w37849 = ~w10700 & w10699;
assign w37850 = ~w10626 & w10705;
assign w37851 = ~w37846 & ~w10706;
assign w37852 = ~w10692 & pi0659;
assign w37853 = w10693 & w10710;
assign w37854 = w10724 & w397;
assign w37855 = ~w10690 & ~w10731;
assign w37856 = w10733 & ~w10684;
assign w37857 = w10733 & ~w10720;
assign w37858 = w10733 & w10719;
assign w37859 = ~pi3551 & ~pi0038;
assign w37860 = ~w37859 & w10741;
assign w37861 = ~w8105 & ~pi3245;
assign w37862 = ~w8257 & pi3245;
assign w37863 = ~w37861 & ~w10745;
assign w37864 = pi0979 & ~pi3426;
assign w37865 = pi0979 & w35945;
assign w37866 = pi3551 & pi0979;
assign w37867 = ~pi3426 & ~pi1666;
assign w37868 = ~w10750 & ~w10754;
assign w37869 = ~w10749 & w10755;
assign w37870 = w7561 & pi3245;
assign w37871 = w5092 & ~pi3245;
assign w37872 = ~w10758 & pi3245;
assign w37873 = ~w10758 & ~w37871;
assign w37874 = pi0713 & ~pi0039;
assign w37875 = ~w10757 & w10761;
assign w37876 = ~w10824 & ~w10814;
assign w37877 = w10918 & ~w10908;
assign w37878 = (w10934 & ~w10903) | (w10934 & w40063) | (~w10903 & w40063);
assign w37879 = w10829 & ~w10940;
assign w37880 = ~w10941 & w10773;
assign w37881 = w10779 & ~w10804;
assign w37882 = ~w10955 & ~w10951;
assign w37883 = w10955 & w10951;
assign w37884 = w10847 & ~w10969;
assign w37885 = w10946 & w10773;
assign w37886 = w10970 & w10965;
assign w37887 = w10976 & ~w11010;
assign w37888 = w10950 & ~w10960;
assign w37889 = ~w10970 & ~w10965;
assign w37890 = w11100 & ~w11090;
assign w37891 = ~w10934 & ~w11117;
assign w37892 = ~w10934 & w10921;
assign w37893 = w11120 & w11115;
assign w37894 = ~w11126 & ~w11122;
assign w37895 = ~w11134 & w11119;
assign w37896 = w11161 & ~w11151;
assign w37897 = ~pi0056 & ~pi0104;
assign w37898 = w11208 & w11187;
assign w37899 = ~w10774 & w11216;
assign w37900 = pi0067 & ~pi0104;
assign w37901 = w11232 & ~w11238;
assign w37902 = ~w11251 & ~w11210;
assign w37903 = w11208 & ~w11187;
assign w37904 = w10934 & w11117;
assign w37905 = ~w11291 & ~w11083;
assign w37906 = w11139 & ~w11295;
assign w37907 = w11063 & ~w11073;
assign w37908 = (~w11041 & ~w11053) | (~w11041 & w40064) | (~w11053 & w40064);
assign w37909 = w11331 & w11327;
assign w37910 = ~w11331 & ~w11327;
assign w37911 = w11017 & ~w11344;
assign w37912 = w11072 & ~w11009;
assign w37913 = w11345 & w11341;
assign w37914 = ~w11343 & ~w11423;
assign w37915 = w11322 & w11424;
assign w37916 = ~w11345 & ~w11341;
assign w37917 = ~w11299 & w11321;
assign w37918 = w11495 & ~w11378;
assign w37919 = ~w11494 & ~w11501;
assign w37920 = w11321 & ~w11302;
assign w37921 = w11422 & w11493;
assign w37922 = ~w11319 & ~w11417;
assign w37923 = ~w11519 & ~w11520;
assign w37924 = w11451 & w11478;
assign w37925 = w11431 & ~w11527;
assign w37926 = ~w11451 & ~w11478;
assign w37927 = w11299 & ~w11321;
assign w37928 = w11493 & ~w11499;
assign w37929 = w11534 & ~w11637;
assign w37930 = ~w11576 & ~w11566;
assign w37931 = ~w11528 & w11582;
assign w37932 = w11704 & w11693;
assign w37933 = w11599 & ~w11748;
assign w37934 = w11715 & w40065;
assign w37935 = (~w11755 & ~w11715) | (~w11755 & w40066) | (~w11715 & w40066);
assign w37936 = w11760 & ~w11594;
assign w37937 = w11526 & ~w11764;
assign w37938 = w11526 & w11755;
assign w37939 = w11721 & w11768;
assign w37940 = w11422 & w11763;
assign w37941 = ~w37940 & ~w11770;
assign w37942 = w11644 & ~w11778;
assign w37943 = w11818 & w11814;
assign w37944 = ~w11818 & ~w11814;
assign w37945 = w11669 & ~w11683;
assign w37946 = ~w11779 & ~w11829;
assign w37947 = w11807 & ~w11822;
assign w37948 = ~pi0081 & ~pi0104;
assign w37949 = w11785 & ~w11851;
assign w37950 = w11779 & w11829;
assign w37951 = ~w11890 & ~w11894;
assign w37952 = ~w11729 & ~w11924;
assign w37953 = w11810 & w11930;
assign w37954 = ~w11810 & ~w11930;
assign w37955 = w11925 & w11933;
assign w37956 = ~w11905 & ~w11937;
assign w37957 = ~w37953 & ~w11966;
assign w37958 = ~w11528 & ~w11582;
assign w37959 = w11690 & ~w11995;
assign w37960 = w11999 & ~w11994;
assign w37961 = ~w11999 & w11994;
assign w37962 = ~w11720 & ~w11753;
assign w37963 = w11528 & w11582;
assign w37964 = ~w12016 & ~w12020;
assign w37965 = w11721 & w12027;
assign w37966 = ~w11765 & ~w12028;
assign w37967 = w11994 & ~w12011;
assign w37968 = ~w12038 & w40067;
assign w37969 = ~w12045 & ~w12040;
assign w37970 = ~w12055 & ~w12025;
assign w37971 = ~w11526 & ~w11420;
assign w37972 = ~w12074 & ~w11771;
assign w37973 = ~w11526 & ~w11763;
assign w37974 = ~w11420 & ~w11770;
assign w37975 = ~w11759 & w12084;
assign w37976 = ~w11832 & ~w11842;
assign w37977 = w12100 & w11201;
assign w37978 = ~w12104 & ~pi0081;
assign w37979 = w12104 & ~w12100;
assign w37980 = ~w12107 & ~pi0104;
assign w37981 = ~w37980 & w12106;
assign w37982 = w11858 & ~w12119;
assign w37983 = ~w11944 & ~w12157;
assign w37984 = ~w11935 & ~w12214;
assign w37985 = ~w12212 & w12156;
assign w37986 = w12212 & ~w12156;
assign w37987 = ~w12158 & w12207;
assign w37988 = ~w12209 & ~w12229;
assign w37989 = w12158 & ~w12207;
assign w37990 = w12164 & ~w12233;
assign w37991 = w12202 & ~w12201;
assign w37992 = w12120 & w12115;
assign w37993 = ~w12120 & ~w12115;
assign w37994 = ~w12107 & ~w12099;
assign w37995 = ~w37994 & ~w12322;
assign w37996 = ~w12139 & ~w12323;
assign w37997 = w12321 & w12344;
assign w37998 = ~w12321 & ~w12323;
assign w37999 = w12301 & ~w12351;
assign w38000 = ~pi0097 & pi1424;
assign w38001 = pi1424 & pi0081;
assign w38002 = ~w12320 & w40068;
assign w38003 = (w12391 & w12320) | (w12391 & w40069) | (w12320 & w40069);
assign w38004 = w12278 & ~w12277;
assign w38005 = ~w12254 & ~w12429;
assign w38006 = ~w12234 & ~w12284;
assign w38007 = w12232 & ~w12259;
assign w38008 = w12285 & w12259;
assign w38009 = w12470 & ~w12471;
assign w38010 = w11986 & ~w12005;
assign w38011 = ~w12092 & w12504;
assign w38012 = w12518 & ~w12515;
assign w38013 = w12527 & ~w11813;
assign w38014 = w12529 & ~w12525;
assign w38015 = ~w12529 & w12525;
assign w38016 = w12408 & ~w12547;
assign w38017 = w12605 & ~w11561;
assign w38018 = w11558 & w11561;
assign w38019 = w12554 & ~w12576;
assign w38020 = ~w12428 & ~w12450;
assign w38021 = w12663 & w12110;
assign w38022 = w12352 & w12110;
assign w38023 = pi1640 & ~w10830;
assign w38024 = pi1468 & pi0081;
assign w38025 = w12392 & ~w12390;
assign w38026 = w12386 & w40070;
assign w38027 = w12710 & ~w12712;
assign w38028 = ~w12719 & w12713;
assign w38029 = ~w12742 & ~w12755;
assign w38030 = ~w12742 & w12757;
assign w38031 = w12546 & ~w12619;
assign w38032 = w12783 & ~w11561;
assign w38033 = w12611 & ~w12601;
assign w38034 = w12798 & w11813;
assign w38035 = ~w11813 & ~pi0078;
assign w38036 = w12845 & ~w12843;
assign w38037 = w12850 & w12857;
assign w38038 = ~w12828 & w12110;
assign w38039 = w12664 & ~w12860;
assign w38040 = ~pi0081 & ~w12101;
assign w38041 = w12842 & w12882;
assign w38042 = ~w12842 & ~w12882;
assign w38043 = w12902 & ~w11813;
assign w38044 = w12811 & ~w12810;
assign w38045 = ~w12787 & ~w12779;
assign w38046 = ~w12963 & w12856;
assign w38047 = w12963 & ~w12856;
assign w38048 = w12842 & ~w12882;
assign w38049 = w12838 & ~w12882;
assign w38050 = ~w12690 & w12110;
assign w38051 = ~w12851 & w12989;
assign w38052 = ~w12885 & w12990;
assign w38053 = w12984 & w12998;
assign w38054 = ~w12984 & ~w12998;
assign w38055 = ~w12943 & w12909;
assign w38056 = w13026 & ~w11561;
assign w38057 = ~w12920 & ~w12937;
assign w38058 = w13051 & ~w11813;
assign w38059 = ~w12900 & ~w12898;
assign w38060 = ~w12911 & w13059;
assign w38061 = ~w13034 & ~w13058;
assign w38062 = w13079 & ~w13078;
assign w38063 = ~w13030 & ~w13022;
assign w38064 = ~w13049 & ~w13047;
assign w38065 = w13007 & ~w12999;
assign w38066 = ~w13007 & w12999;
assign w38067 = ~w13007 & ~w12999;
assign w38068 = w12838 & w12110;
assign w38069 = w12875 & w12997;
assign w38070 = ~w13166 & w13178;
assign w38071 = w12982 & ~w12761;
assign w38072 = w13202 & ~w11813;
assign w38073 = w13204 & ~w13200;
assign w38074 = w13219 & ~w11813;
assign w38075 = ~w13272 & ~w13227;
assign w38076 = w13221 & ~w13215;
assign w38077 = pi1418 & pi0081;
assign w38078 = w13316 & ~w13315;
assign w38079 = w13272 & ~w13226;
assign w38080 = ~w13334 & w13349;
assign w38081 = w13326 & ~w13169;
assign w38082 = w13290 & ~w13289;
assign w38083 = ~w13300 & w13411;
assign w38084 = w13419 & w13408;
assign w38085 = ~w13419 & ~w13408;
assign w38086 = ~w13119 & ~w13108;
assign w38087 = w13145 & ~w13434;
assign w38088 = ~w13454 & ~w13169;
assign w38089 = w13511 & ~w13510;
assign w38090 = ~w13498 & w13169;
assign w38091 = pi1640 & ~w11808;
assign w38092 = ~w13545 & ~w13544;
assign w38093 = w13401 & ~w13400;
assign w38094 = w13563 & w13565;
assign w38095 = w13557 & ~w13558;
assign w38096 = ~w13585 & w13567;
assign w38097 = ~w13589 & ~w13587;
assign w38098 = ~w13585 & w13588;
assign w38099 = w13585 & w13565;
assign w38100 = ~w13571 & ~w13580;
assign w38101 = ~w13568 & ~w12101;
assign w38102 = w13597 & ~w13567;
assign w38103 = w13618 & ~w13594;
assign w38104 = ~w13575 & w40071;
assign w38105 = (~w13623 & w13575) | (~w13623 & w40072) | (w13575 & w40072);
assign w38106 = ~w13387 & w13316;
assign w38107 = w13387 & w13565;
assign w38108 = w13644 & ~w13650;
assign w38109 = ~w13563 & w13567;
assign w38110 = ~w13387 & ~w13316;
assign w38111 = ~w13604 & w13623;
assign w38112 = ~w13604 & w13600;
assign w38113 = ~w13411 & w13696;
assign w38114 = w13411 & ~w13696;
assign w38115 = ~w13597 & ~w13567;
assign w38116 = ~w13709 & ~w13702;
assign w38117 = w13709 & w13702;
assign w38118 = ~w13741 & w13744;
assign w38119 = ~w13620 & ~w13169;
assign w38120 = ~w13720 & ~w13749;
assign w38121 = w13491 & w13750;
assign w38122 = ~w13525 & ~w13759;
assign w38123 = w13757 & w13772;
assign w38124 = ~w13773 & w13750;
assign w38125 = w12729 & w13787;
assign w38126 = w12397 & w13789;
assign w38127 = w12718 & ~w12712;
assign w38128 = ~w12397 & w13792;
assign w38129 = ~w12746 & w13794;
assign w38130 = ~w13604 & w13696;
assign w38131 = w13811 & ~w13605;
assign w38132 = w13814 & ~w13565;
assign w38133 = ~w13411 & w13820;
assign w38134 = w13411 & ~w13820;
assign w38135 = ~w13786 & ~w13836;
assign w38136 = w13786 & ~w13839;
assign w38137 = w13183 & ~w13839;
assign w38138 = ~w13720 & w13849;
assign w38139 = w13183 & w13850;
assign w38140 = w13737 & ~w13686;
assign w38141 = w13757 & w13858;
assign w38142 = ~w13859 & ~w13863;
assign w38143 = w13491 & ~w13863;
assign w38144 = w13864 & ~w13718;
assign w38145 = w13183 & ~w13718;
assign w38146 = ~w13741 & ~w13743;
assign w38147 = w13183 & w13877;
assign w38148 = w13539 & w40073;
assign w38149 = w13757 & w13882;
assign w38150 = ~w13883 & w13877;
assign w38151 = w13686 & ~w13687;
assign w38152 = w13846 & ~w13893;
assign w38153 = ~w13864 & w13901;
assign w38154 = w13859 & ~w13905;
assign w38155 = ~w13686 & ~w13687;
assign w38156 = ~w38155 & w13904;
assign w38157 = w13183 & w13908;
assign w38158 = w13913 & w10752;
assign w38159 = ~pi3245 & ~w36655;
assign w38160 = ~pi3245 & ~w36654;
assign w38161 = pi0713 & ~pi0040;
assign w38162 = ~w10757 & w13918;
assign w38163 = pi3551 & ~pi0979;
assign w38164 = ~pi0979 & ~pi3426;
assign w38165 = ~pi0979 & w35945;
assign w38166 = ~w13922 & ~w13926;
assign w38167 = ~w13929 & w13927;
assign w38168 = w13931 & ~w37873;
assign w38169 = w13931 & ~w37872;
assign w38170 = pi0713 & ~pi0041;
assign w38171 = w13913 & w13923;
assign w38172 = pi0713 & ~pi0042;
assign w38173 = ~w13931 & w13941;
assign w38174 = ~w370 & pi2384;
assign w38175 = ~w13913 & w13946;
assign w38176 = ~w13961 & w13990;
assign w38177 = ~w10690 & ~w13999;
assign w38178 = w14002 & w10710;
assign w38179 = w14002 & w37853;
assign w38180 = w10690 & ~w13960;
assign w38181 = w14008 & w13995;
assign w38182 = w14012 & w13995;
assign w38183 = ~pi3551 & ~pi0045;
assign w38184 = ~w38183 & w10741;
assign w38185 = w10690 & w13990;
assign w38186 = w10642 & ~w13969;
assign w38187 = ~w10642 & w14024;
assign w38188 = ~w14020 & ~w14026;
assign w38189 = w10642 & ~w14028;
assign w38190 = ~w10642 & ~w14030;
assign w38191 = ~w14032 & w14016;
assign w38192 = w7496 & pi3245;
assign w38193 = w4523 & ~pi3245;
assign w38194 = ~w14036 & pi3245;
assign w38195 = ~w14036 & ~w38193;
assign w38196 = pi0713 & ~pi0046;
assign w38197 = ~w10757 & w14038;
assign w38198 = ~w10756 & ~w10752;
assign w38199 = w13491 & ~w13742;
assign w38200 = ~w13883 & ~w13742;
assign w38201 = ~w14046 & ~w14049;
assign w38202 = w14046 & ~w14052;
assign w38203 = w13183 & ~w14052;
assign w38204 = ~pi0868 & ~w14040;
assign w38205 = w13931 & ~w38195;
assign w38206 = w13931 & ~w38194;
assign w38207 = pi0713 & ~pi0047;
assign w38208 = ~w13930 & ~w13923;
assign w38209 = ~pi0868 & ~w14070;
assign w38210 = ~pi0868 & w13946;
assign w38211 = ~w14046 & ~w14079;
assign w38212 = w14046 & ~w14082;
assign w38213 = w13491 & w13730;
assign w38214 = w13782 & w14093;
assign w38215 = w13757 & w14093;
assign w38216 = ~w14098 & w14100;
assign w38217 = w14098 & w14103;
assign w38218 = w13183 & w14103;
assign w38219 = w14108 & w10752;
assign w38220 = w3484 & ~pi3245;
assign w38221 = ~w14110 & pi3245;
assign w38222 = ~w14110 & ~w38220;
assign w38223 = pi0713 & ~pi0049;
assign w38224 = ~w10757 & w14112;
assign w38225 = w14108 & w13923;
assign w38226 = w13931 & ~w38222;
assign w38227 = w13931 & ~w38221;
assign w38228 = pi0713 & ~pi0050;
assign w38229 = w13604 & ~w13820;
assign w38230 = w14129 & w13565;
assign w38231 = ~w14129 & ~w13565;
assign w38232 = w14125 & w14133;
assign w38233 = ~w14133 & ~w14125;
assign w38234 = w13826 & ~w13169;
assign w38235 = w13757 & w14151;
assign w38236 = ~w14136 & ~w13169;
assign w38237 = ~w13604 & w14125;
assign w38238 = w14161 & w14159;
assign w38239 = ~w14161 & ~w14159;
assign w38240 = w14136 & ~w14161;
assign w38241 = w13604 & ~w14159;
assign w38242 = ~w14198 & ~w14195;
assign w38243 = w14206 & w14210;
assign w38244 = ~w14206 & ~w14210;
assign w38245 = ~w14175 & ~w14173;
assign w38246 = w14152 & ~w14218;
assign w38247 = ~w13808 & ~w14222;
assign w38248 = w13834 & w14147;
assign w38249 = w14223 & ~w14213;
assign w38250 = ~w14227 & w14215;
assign w38251 = w13183 & w14230;
assign w38252 = ~w13169 & ~w14199;
assign w38253 = w13604 & ~w14180;
assign w38254 = ~w13411 & w14180;
assign w38255 = w14126 & ~w14237;
assign w38256 = w13169 & w14199;
assign w38257 = w14185 & w13565;
assign w38258 = ~w14238 & ~w13565;
assign w38259 = ~w14238 & ~w38257;
assign w38260 = ~w14258 & ~w14256;
assign w38261 = w14258 & w14256;
assign w38262 = ~w14255 & w14261;
assign w38263 = w14255 & ~w14261;
assign w38264 = ~w14152 & w14228;
assign w38265 = ~w14274 & w14276;
assign w38266 = w14227 & w14280;
assign w38267 = w13183 & w14281;
assign w38268 = ~w14214 & w10752;
assign w38269 = w7691 & pi3245;
assign w38270 = w2979 & ~pi3245;
assign w38271 = ~w14290 & pi3245;
assign w38272 = ~w14290 & ~w38270;
assign w38273 = pi0713 & ~pi0051;
assign w38274 = ~w10757 & w14292;
assign w38275 = w13183 & w14296;
assign w38276 = ~w14152 & w14296;
assign w38277 = w13540 & w14296;
assign w38278 = ~w14274 & ~pi0868;
assign w38279 = ~w14274 & w14308;
assign w38280 = w14152 & ~w14312;
assign w38281 = ~w14227 & ~w14214;
assign w38282 = w13183 & w14316;
assign w38283 = w7659 & pi3245;
assign w38284 = ~pi3245 & ~w36198;
assign w38285 = ~pi3245 & ~w36197;
assign w38286 = pi0713 & ~pi0052;
assign w38287 = ~w10757 & w14327;
assign w38288 = ~w10747 & ~w38272;
assign w38289 = ~w10747 & ~w38271;
assign w38290 = pi0713 & pi0053;
assign w38291 = ~w13931 & w14333;
assign w38292 = ~w13922 & ~w14335;
assign w38293 = ~w13929 & w14336;
assign w38294 = ~w14214 & ~w14338;
assign w38295 = ~w14337 & ~w13923;
assign w38296 = pi0713 & ~pi0054;
assign w38297 = ~w13931 & w14346;
assign w38298 = pi3516 & pi0541;
assign w38299 = pi3516 & w35748;
assign w38300 = pi3518 & pi0541;
assign w38301 = pi3518 & w35748;
assign w38302 = ~pi0416 & ~pi0418;
assign w38303 = ~pi0419 & pi0408;
assign w38304 = ~pi3130 & pi0541;
assign w38305 = ~pi3130 & w35748;
assign w38306 = w14371 & w14369;
assign w38307 = ~w14385 & w14381;
assign w38308 = ~pi0426 & ~pi0695;
assign w38309 = w14387 & w10747;
assign w38310 = ~pi0409 & w14398;
assign w38311 = w14375 & w14400;
assign w38312 = w38311 & ~pi0410;
assign w38313 = w38312 & w14365;
assign w38314 = w37798 & pi0828;
assign w38315 = ~w10097 & w14402;
assign w38316 = ~w10106 & w14403;
assign w38317 = ~w14406 & w14401;
assign w38318 = w10109 & w14401;
assign w38319 = ~w10276 & ~w10099;
assign w38320 = w10312 & w14411;
assign w38321 = w10312 & ~w10605;
assign w38322 = w10357 & ~w10605;
assign w38323 = w10357 & w38321;
assign w38324 = ~w10276 & w10594;
assign w38325 = ~w14419 & ~w14412;
assign w38326 = w38311 & w14376;
assign w38327 = w9936 & ~w14423;
assign w38328 = w4327 & w6295;
assign w38329 = w38328 & w3392;
assign w38330 = w14427 & ~w1182;
assign w38331 = ~w14427 & w14433;
assign w38332 = ~w38328 & w14427;
assign w38333 = ~pi2486 & pi3510;
assign w38334 = ~w3392 & ~w14440;
assign w38335 = ~w4327 & w14427;
assign w38336 = w14443 & ~w14427;
assign w38337 = w14443 & ~w38335;
assign w38338 = w14444 & w14450;
assign w38339 = w14436 & pi3518;
assign w38340 = ~w5763 & w14427;
assign w38341 = ~pi2486 & pi3398;
assign w38342 = ~w14458 & ~w14459;
assign w38343 = ~pi2486 & pi3330;
assign w38344 = ~w14427 & w14470;
assign w38345 = w14427 & w4327;
assign w38346 = ~w38345 & ~w14472;
assign w38347 = ~pi2486 & pi3392;
assign w38348 = w14480 & w14450;
assign w38349 = ~pi2486 & pi3394;
assign w38350 = ~w14463 & w14450;
assign w38351 = w14436 & ~pi3518;
assign w38352 = ~w14425 & ~w14498;
assign w38353 = ~w14499 & w14487;
assign w38354 = ~w14480 & w14450;
assign w38355 = w38353 & w14505;
assign w38356 = ~w14499 & ~w14487;
assign w38357 = w38356 & w14508;
assign w38358 = w14425 & w14510;
assign w38359 = w14444 & w14487;
assign w38360 = ~w14514 & ~w14442;
assign w38361 = w14486 & w14450;
assign w38362 = w14519 & w14522;
assign w38363 = ~w14436 & w14524;
assign w38364 = w14507 & w14511;
assign w38365 = w14518 & ~w14494;
assign w38366 = w38353 & w14508;
assign w38367 = w38356 & w14548;
assign w38368 = w14450 & ~pi3518;
assign w38369 = w14436 & ~w14487;
assign w38370 = w14511 & w14484;
assign w38371 = ~w14486 & w14450;
assign w38372 = ~w14559 & w14560;
assign w38373 = ~w14559 & w14505;
assign w38374 = w14436 & w14559;
assign w38375 = pi2021 & ~pi3518;
assign w38376 = w14584 & ~w14585;
assign w38377 = w14511 & w14530;
assign w38378 = w14511 & w14592;
assign w38379 = w14595 & w14556;
assign w38380 = ~w14559 & w14513;
assign w38381 = w14600 & w14426;
assign w38382 = w14604 & w14539;
assign w38383 = w10421 & ~w14607;
assign w38384 = ~w14436 & pi3518;
assign w38385 = ~w14559 & w14484;
assign w38386 = w14487 & ~w14612;
assign w38387 = w14611 & w14609;
assign w38388 = w10111 & ~w14618;
assign w38389 = w10446 & ~w14621;
assign w38390 = w10478 & ~w14632;
assign w38391 = w10064 & ~w14635;
assign w38392 = w10015 & ~w14647;
assign w38393 = w9971 & ~w14650;
assign w38394 = w14450 & w14548;
assign w38395 = ~w14660 & w14559;
assign w38396 = w10194 & ~w14663;
assign w38397 = w14450 & w14531;
assign w38398 = ~w14671 & w14559;
assign w38399 = w10363 & ~w14674;
assign w38400 = w10296 & ~w14683;
assign w38401 = w10246 & ~w14686;
assign w38402 = w14526 & ~w14689;
assign w38403 = ~w14670 & ~w14659;
assign w38404 = w10509 & ~w14696;
assign w38405 = w14513 & w14550;
assign w38406 = w10315 & ~w14701;
assign w38407 = w14526 & w14703;
assign w38408 = w14502 & w14524;
assign w38409 = w14436 & w14490;
assign w38410 = ~w14559 & w14592;
assign w38411 = ~w14559 & w14530;
assign w38412 = w14508 & w14522;
assign w38413 = w14600 & w14709;
assign w38414 = ~w14606 & ~pi0709;
assign w38415 = ~w14731 & ~w36655;
assign w38416 = ~w14731 & ~w36654;
assign w38417 = w9941 & pi0541;
assign w38418 = w9941 & w35748;
assign w38419 = ~w14375 & pi0410;
assign w38420 = w14737 & pi0410;
assign w38421 = w14737 & w38419;
assign w38422 = ~pi3426 & ~w923;
assign w38423 = ~w14744 & ~pi0343;
assign w38424 = w9934 & pi0541;
assign w38425 = w9934 & w35748;
assign w38426 = w14748 & pi0410;
assign w38427 = w14748 & w38419;
assign w38428 = w9938 & pi0541;
assign w38429 = w9938 & w35748;
assign w38430 = ~w14375 & ~pi0410;
assign w38431 = w14748 & ~pi0410;
assign w38432 = w14748 & w38430;
assign w38433 = ~w14735 & ~w14734;
assign w38434 = w38312 & w14378;
assign w38435 = w14453 & ~w14763;
assign w38436 = ~w14442 & ~w14766;
assign w38437 = ~w14759 & ~w14509;
assign w38438 = w14490 & ~w14624;
assign w38439 = w14775 & w14710;
assign w38440 = w14774 & w14453;
assign w38441 = ~w14773 & ~w14771;
assign w38442 = w14507 & pi3518;
assign w38443 = w14450 & ~w14689;
assign w38444 = w38311 & ~w14381;
assign w38445 = pi0343 & w14800;
assign w38446 = ~pi3551 & ~w923;
assign w38447 = w9951 & pi0541;
assign w38448 = w9951 & w35748;
assign w38449 = pi3551 & w14811;
assign w38450 = ~w14809 & ~w14811;
assign w38451 = ~w14809 & ~w38449;
assign w38452 = w14805 & w14813;
assign w38453 = w9931 & pi0541;
assign w38454 = w9931 & w35748;
assign w38455 = w14737 & ~pi0410;
assign w38456 = w14737 & w38430;
assign w38457 = w9944 & pi0541;
assign w38458 = w9944 & w35748;
assign w38459 = w14819 & ~pi0410;
assign w38460 = w14819 & w38430;
assign w38461 = w14818 & ~w5758;
assign w38462 = w9946 & pi0541;
assign w38463 = w9946 & w35748;
assign w38464 = w14819 & pi0410;
assign w38465 = w14819 & w38419;
assign w38466 = w14823 & ~w5767;
assign w38467 = w14814 & w14828;
assign w38468 = w14830 & ~w14757;
assign w38469 = ~w14408 & w14364;
assign w38470 = w14841 & pi3245;
assign w38471 = ~w14807 & w14355;
assign w38472 = pi3509 & pi0541;
assign w38473 = pi3509 & w35748;
assign w38474 = ~w14869 & ~w14868;
assign w38475 = ~w14807 & w14872;
assign w38476 = w14812 & w14364;
assign w38477 = w14806 & ~pi0055;
assign w38478 = w14806 & w14884;
assign w38479 = pi3551 & w14374;
assign w38480 = pi2384 & pi0541;
assign w38481 = pi2384 & w35748;
assign w38482 = ~w14841 & ~w14870;
assign w38483 = ~w14888 & pi0056;
assign w38484 = w14889 & w14892;
assign w38485 = ~w14108 & w13946;
assign w38486 = ~w14898 & w10755;
assign w38487 = ~w14898 & w37869;
assign w38488 = w13766 & ~pi0868;
assign w38489 = ~w13758 & w14909;
assign w38490 = ~w14904 & ~w14899;
assign w38491 = ~w14917 & w13927;
assign w38492 = ~w14917 & w38167;
assign w38493 = ~w14904 & ~w14918;
assign w38494 = ~w14214 & w13946;
assign w38495 = w13773 & ~w14933;
assign w38496 = ~w13720 & w14224;
assign w38497 = w13183 & w14937;
assign w38498 = w13833 & ~pi0868;
assign w38499 = w13773 & ~w14943;
assign w38500 = ~w14942 & ~pi0868;
assign w38501 = w13183 & w14946;
assign w38502 = w14274 & pi0868;
assign w38503 = w14951 & w10752;
assign w38504 = w7626 & pi3245;
assign w38505 = ~pi3245 & w6196;
assign w38506 = ~pi3245 & ~w36727;
assign w38507 = ~w14961 & ~w38505;
assign w38508 = ~w14961 & ~w38506;
assign w38509 = pi0713 & ~pi0062;
assign w38510 = ~w10757 & w14964;
assign w38511 = w13746 & pi0868;
assign w38512 = ~w13786 & ~w14970;
assign w38513 = ~w13786 & w14975;
assign w38514 = w13183 & w14978;
assign w38515 = ~pi0868 & w10752;
assign w38516 = w7593 & pi3245;
assign w38517 = w4160 & ~pi3245;
assign w38518 = ~w14987 & pi3245;
assign w38519 = ~w14987 & ~w38517;
assign w38520 = pi0713 & ~pi0063;
assign w38521 = ~w10757 & w14989;
assign w38522 = w14951 & w13923;
assign w38523 = pi0713 & ~pi0064;
assign w38524 = ~w13931 & w14995;
assign w38525 = ~pi0868 & w13923;
assign w38526 = w13931 & ~w38519;
assign w38527 = w13931 & ~w38518;
assign w38528 = pi0713 & ~pi0065;
assign w38529 = w10344 & ~w10099;
assign w38530 = ~w10293 & ~w10594;
assign w38531 = w14611 & ~w15020;
assign w38532 = ~w14660 & w14521;
assign w38533 = w14450 & w14487;
assign w38534 = w14601 & w14709;
assign w38535 = ~w14671 & w14521;
assign w38536 = w14526 & ~w15056;
assign w38537 = w15034 & ~w15021;
assign w38538 = ~pi0709 & w14422;
assign w38539 = w4523 & ~w14731;
assign w38540 = w4685 & w14745;
assign w38541 = ~w15066 & w14735;
assign w38542 = w15075 & ~w15074;
assign w38543 = w14584 & ~w15037;
assign w38544 = w14534 & ~w15020;
assign w38545 = w14502 & w14469;
assign w38546 = w14504 & ~w15051;
assign w38547 = w14502 & w14504;
assign w38548 = w15083 & w14453;
assign w38549 = ~w15079 & w14758;
assign w38550 = ~w38445 & w14813;
assign w38551 = ~w7496 & ~w14805;
assign w38552 = w14823 & ~w4661;
assign w38553 = w14818 & ~w4657;
assign w38554 = ~w7496 & ~w14856;
assign w38555 = ~w15123 & ~w15122;
assign w38556 = ~w4523 & w14852;
assign w38557 = w14806 & pi0066;
assign w38558 = ~w38556 & w15135;
assign w38559 = w15124 & ~w14889;
assign w38560 = (~w13179 & w13779) | (~w13179 & w40074) | (w13779 & w40074);
assign w38561 = w15144 & ~w15145;
assign w38562 = ~w13782 & ~w13757;
assign w38563 = w15152 & w15153;
assign w38564 = w15145 & ~w15144;
assign w38565 = w7787 & pi3245;
assign w38566 = w4866 & ~pi3245;
assign w38567 = ~w15170 & pi3245;
assign w38568 = ~w15170 & ~w38566;
assign w38569 = ~w10750 & ~w15172;
assign w38570 = ~w10749 & w15175;
assign w38571 = w13929 & ~w38568;
assign w38572 = w13929 & ~w38567;
assign w38573 = ~pi3426 & ~pi1667;
assign w38574 = ~w10750 & pi0070;
assign w38575 = ~w13922 & pi0071;
assign w38576 = ~pi0127 & ~pi0072;
assign w38577 = w15196 & ~pi0368;
assign w38578 = w15195 & ~pi1742;
assign w38579 = w38578 & ~pi1745;
assign w38580 = pi1714 & pi1897;
assign w38581 = ~pi1744 & ~pi1897;
assign w38582 = ~pi1744 & ~w38580;
assign w38583 = w15206 & ~w38581;
assign w38584 = w15206 & ~w38582;
assign w38585 = ~w15194 & ~w38584;
assign w38586 = ~w15194 & ~w38583;
assign w38587 = ~w15196 & pi1897;
assign w38588 = w15208 & pi0072;
assign w38589 = w15227 & pi0127;
assign w38590 = pi0314 & pi0330;
assign w38591 = ~pi0128 & w15234;
assign w38592 = ~w15235 & ~pi0330;
assign w38593 = ~w15235 & ~w38590;
assign w38594 = ~pi0330 & w15239;
assign w38595 = ~w15200 & ~w15239;
assign w38596 = ~w15200 & ~w38594;
assign w38597 = w15240 & w15217;
assign w38598 = ~pi1897 & w15243;
assign w38599 = ~w15244 & ~w15248;
assign w38600 = w38599 & ~w15249;
assign w38601 = ~w38578 & pi1897;
assign w38602 = w38600 & ~w15254;
assign w38603 = ~w38602 & ~pi1017;
assign w38604 = w15212 & pi1017;
assign w38605 = w15212 & ~w38603;
assign w38606 = ~w15257 & ~w15258;
assign w38607 = pi1744 & pi1897;
assign w38608 = pi1744 & w38580;
assign w38609 = ~w15259 & ~w15261;
assign w38610 = w38578 & pi1897;
assign w38611 = ~w38600 & w15265;
assign w38612 = ~w15267 & ~pi1017;
assign w38613 = ~w38599 & w15273;
assign w38614 = ~w15278 & ~w38607;
assign w38615 = ~w15278 & ~w38608;
assign w38616 = ~w15279 & ~w15207;
assign w38617 = ~pi1745 & ~w15281;
assign w38618 = ~w15195 & ~pi1017;
assign w38619 = w15283 & pi1017;
assign w38620 = w15283 & ~w38618;
assign w38621 = ~w38600 & ~w15286;
assign w38622 = ~w15195 & w15287;
assign w38623 = ~w15288 & w15286;
assign w38624 = ~w15288 & ~w38621;
assign w38625 = ~w15248 & ~w15249;
assign w38626 = w15244 & ~w15295;
assign w38627 = w15280 & ~w15301;
assign w38628 = ~pi1897 & ~w15306;
assign w38629 = ~w15310 & w15314;
assign w38630 = pi0368 & ~w15239;
assign w38631 = pi0368 & ~w38594;
assign w38632 = ~w15319 & pi1867;
assign w38633 = w15319 & ~pi1867;
assign w38634 = w15320 & ~w15318;
assign w38635 = ~w15240 & ~w15217;
assign w38636 = ~pi0330 & ~pi1017;
assign w38637 = ~w15234 & ~w15336;
assign w38638 = w15330 & w15342;
assign w38639 = w15196 & ~pi1017;
assign w38640 = w15196 & w15210;
assign w38641 = pi1897 & pi0330;
assign w38642 = w15346 & pi1017;
assign w38643 = w15346 & ~w38636;
assign w38644 = ~w15330 & w15353;
assign w38645 = w38600 & ~w15270;
assign w38646 = pi1714 & ~w15273;
assign w38647 = w15360 & ~w15265;
assign w38648 = w15360 & ~w38611;
assign w38649 = w15297 & ~w15362;
assign w38650 = ~w15363 & ~w15330;
assign w38651 = ~w15376 & w15263;
assign w38652 = w15376 & ~w15353;
assign w38653 = ~w15382 & w15386;
assign w38654 = pi0734 & ~pi3427;
assign w38655 = pi0072 & ~pi3427;
assign w38656 = pi0072 & w38654;
assign w38657 = ~pi2555 & ~w38655;
assign w38658 = ~pi2555 & ~w38656;
assign w38659 = ~w15390 & ~w15391;
assign w38660 = ~w15390 & ~w15394;
assign w38661 = w15218 & pi1017;
assign w38662 = w15317 & ~w15407;
assign w38663 = ~w38662 & ~w15398;
assign w38664 = w15221 & ~pi1017;
assign w38665 = w15324 & ~w15424;
assign w38666 = ~w15318 & w15430;
assign w38667 = w15373 & ~w15323;
assign w38668 = w15408 & w15435;
assign w38669 = ~w15436 & ~w15409;
assign w38670 = pi0073 & ~pi3427;
assign w38671 = pi0073 & w38654;
assign w38672 = ~pi2555 & ~w38670;
assign w38673 = ~pi2555 & ~w38671;
assign w38674 = ~w15439 & ~w15391;
assign w38675 = ~w15439 & ~w15394;
assign w38676 = ~w10392 & ~w10593;
assign w38677 = w10174 & w10397;
assign w38678 = w10605 & ~w10593;
assign w38679 = w10393 & ~w10593;
assign w38680 = w14508 & w14709;
assign w38681 = ~w15454 & ~w14700;
assign w38682 = w14654 & w14550;
assign w38683 = w14723 & ~w15458;
assign w38684 = w15460 & w15456;
assign w38685 = w14600 & w14550;
assign w38686 = ~w14716 & ~w15464;
assign w38687 = w14611 & ~w14653;
assign w38688 = ~w14772 & ~w15470;
assign w38689 = w14526 & ~w14666;
assign w38690 = w14600 & ~w14559;
assign w38691 = w14526 & ~w15484;
assign w38692 = w14505 & ~w15486;
assign w38693 = w14600 & w14640;
assign w38694 = w15481 & w15491;
assign w38695 = ~w15493 & ~pi0709;
assign w38696 = ~w14731 & ~w36198;
assign w38697 = ~w14731 & ~w36197;
assign w38698 = w3335 & w14745;
assign w38699 = ~w15497 & w14735;
assign w38700 = ~w14587 & w14517;
assign w38701 = ~w15508 & ~w15507;
assign w38702 = w14511 & w14654;
assign w38703 = w14453 & ~w14653;
assign w38704 = w14763 & ~w15525;
assign w38705 = ~w15506 & w14758;
assign w38706 = ~w7659 & ~w14805;
assign w38707 = w14818 & ~w3387;
assign w38708 = w14823 & ~w3396;
assign w38709 = w15542 & ~w15503;
assign w38710 = ~w7659 & ~w14856;
assign w38711 = ~w15556 & ~w15555;
assign w38712 = w14806 & ~pi0074;
assign w38713 = w14806 & w15568;
assign w38714 = w10395 & ~w10099;
assign w38715 = ~w10173 & w10594;
assign w38716 = ~w15574 & ~w10099;
assign w38717 = ~w15574 & w38714;
assign w38718 = w14611 & ~w15029;
assign w38719 = ~w14487 & ~w15479;
assign w38720 = ~w14486 & ~w14450;
assign w38721 = w14526 & ~w15588;
assign w38722 = w14526 & ~w15024;
assign w38723 = w15056 & ~w15592;
assign w38724 = ~w15581 & ~w15579;
assign w38725 = ~w15462 & ~pi0709;
assign w38726 = w6330 & w14745;
assign w38727 = ~w15603 & w14735;
assign w38728 = w14450 & ~w15045;
assign w38729 = w14490 & ~w15041;
assign w38730 = ~w15619 & w14453;
assign w38731 = ~w14709 & ~w15627;
assign w38732 = w15631 & ~w15610;
assign w38733 = ~w15505 & w14758;
assign w38734 = ~w7626 & ~w14805;
assign w38735 = w14823 & ~w6304;
assign w38736 = w14818 & ~w6308;
assign w38737 = w15643 & ~w15609;
assign w38738 = ~w7626 & ~w14856;
assign w38739 = ~w15656 & ~w15655;
assign w38740 = w14852 & ~w6196;
assign w38741 = w14852 & w36727;
assign w38742 = w14806 & ~pi0075;
assign w38743 = ~w10359 & ~w10099;
assign w38744 = w10594 & w15674;
assign w38745 = w14611 & ~w14638;
assign w38746 = ~w15683 & ~w14700;
assign w38747 = w14584 & w14662;
assign w38748 = w14526 & w14665;
assign w38749 = ~w15692 & ~w15691;
assign w38750 = w14725 & ~w15681;
assign w38751 = w4160 & ~w14731;
assign w38752 = w4357 & w14745;
assign w38753 = ~w15706 & w14735;
assign w38754 = ~w14559 & w14567;
assign w38755 = ~w15717 & ~w15713;
assign w38756 = ~w14620 & ~w15729;
assign w38757 = ~w15732 & w15730;
assign w38758 = ~w15728 & ~w15727;
assign w38759 = ~w7593 & ~w14805;
assign w38760 = w14823 & ~w4323;
assign w38761 = w14818 & ~w4331;
assign w38762 = w15747 & ~w15712;
assign w38763 = ~w4160 & w14852;
assign w38764 = ~w7593 & ~w14856;
assign w38765 = ~w15761 & ~w15760;
assign w38766 = ~w15770 & ~w14806;
assign w38767 = w10592 & w10610;
assign w38768 = w14491 & w14487;
assign w38769 = w14560 & w14521;
assign w38770 = ~w14487 & ~w15715;
assign w38771 = w14563 & w15519;
assign w38772 = w14567 & w14522;
assign w38773 = ~w15809 & w15800;
assign w38774 = w14490 & ~w15045;
assign w38775 = w15822 & w14710;
assign w38776 = w14534 & ~w15037;
assign w38777 = ~w15827 & ~w15821;
assign w38778 = ~w15828 & w14526;
assign w38779 = ~w14709 & ~w15833;
assign w38780 = w15798 & w15835;
assign w38781 = w14611 & ~w15037;
assign w38782 = ~w14577 & ~w15850;
assign w38783 = w14563 & ~w14587;
assign w38784 = w15865 & ~w15839;
assign w38785 = ~w15838 & w14758;
assign w38786 = w2979 & pi0343;
assign w38787 = w14375 & ~w923;
assign w38788 = w38787 & w15873;
assign w38789 = ~w38788 & ~pi0343;
assign w38790 = ~w7691 & w14804;
assign w38791 = ~w38445 & ~w15881;
assign w38792 = ~w8105 & w14734;
assign w38793 = ~w8257 & w14803;
assign w38794 = w14823 & ~w8195;
assign w38795 = w14818 & ~w8203;
assign w38796 = ~w15883 & w15892;
assign w38797 = w15882 & ~w15880;
assign w38798 = ~w8257 & ~w14856;
assign w38799 = ~w15906 & ~w15905;
assign w38800 = w37861 & ~w14851;
assign w38801 = ~w38800 & w15918;
assign w38802 = ~w14888 & ~pi0078;
assign w38803 = ~w14841 & w15923;
assign w38804 = w15922 & ~w14813;
assign w38805 = ~w14888 & ~pi0079;
assign w38806 = ~w14841 & w15928;
assign w38807 = w15927 & ~w14813;
assign w38808 = w15762 & ~w14889;
assign w38809 = ~w14401 & w15896;
assign w38810 = ~w14841 & ~w15907;
assign w38811 = ~w14888 & pi0081;
assign w38812 = w14889 & w15940;
assign w38813 = ~w14951 & w13946;
assign w38814 = ~w14904 & w13946;
assign w38815 = w15152 & w15954;
assign w38816 = w15152 & w15960;
assign w38817 = w15152 & w13539;
assign w38818 = w13183 & pi0868;
assign w38819 = w7819 & pi3245;
assign w38820 = ~pi3245 & w5448;
assign w38821 = ~pi3245 & ~w36613;
assign w38822 = ~w15977 & ~w38820;
assign w38823 = ~w15977 & ~w38821;
assign w38824 = ~w10749 & w15980;
assign w38825 = ~w11635 & ~w11624;
assign w38826 = ~w11635 & w11777;
assign w38827 = w12088 & w15991;
assign w38828 = ~w12088 & ~w15991;
assign w38829 = w11401 & w11634;
assign w38830 = ~pi0868 & ~w16013;
assign w38831 = w11295 & ~w11290;
assign w38832 = w11139 & w11290;
assign w38833 = ~w16020 & w11082;
assign w38834 = w16020 & ~w11082;
assign w38835 = ~pi0868 & ~w16030;
assign w38836 = ~pi0868 & ~w16042;
assign w38837 = ~pi0868 & ~w16046;
assign w38838 = ~pi0868 & ~w16054;
assign w38839 = ~pi0868 & ~w16058;
assign w38840 = ~pi0868 & ~w16063;
assign w38841 = ~w16051 & w16073;
assign w38842 = w16027 & w16078;
assign w38843 = ~w16087 & ~w10752;
assign w38844 = ~w12055 & ~w12089;
assign w38845 = w12055 & ~w12034;
assign w38846 = ~w12090 & w16092;
assign w38847 = ~w12055 & ~w12034;
assign w38848 = ~w16095 & ~pi0868;
assign w38849 = w12092 & w16103;
assign w38850 = ~w12092 & ~w16103;
assign w38851 = ~w16102 & w10752;
assign w38852 = ~w16119 & ~w13923;
assign w38853 = ~w16102 & w13923;
assign w38854 = ~w10750 & ~pi0089;
assign w38855 = ~w14904 & w15185;
assign w38856 = ~w10750 & pi0090;
assign w38857 = ~w10750 & ~pi0091;
assign w38858 = w16102 & w15185;
assign w38859 = ~w13922 & ~pi0092;
assign w38860 = ~w14904 & w15189;
assign w38861 = ~w13922 & pi0093;
assign w38862 = ~w13922 & ~pi0094;
assign w38863 = w16102 & w15189;
assign w38864 = w10140 & ~w10099;
assign w38865 = ~w10474 & ~w10593;
assign w38866 = ~w10474 & ~w10594;
assign w38867 = ~w16156 & ~w10099;
assign w38868 = ~w16156 & w38864;
assign w38869 = w14611 & w14640;
assign w38870 = w14505 & w14550;
assign w38871 = ~w16184 & ~w16185;
assign w38872 = w16187 & ~w16177;
assign w38873 = ~w16168 & w16166;
assign w38874 = w15461 & w15465;
assign w38875 = ~w15517 & ~w14506;
assign w38876 = w16194 & ~w14602;
assign w38877 = ~w14487 & w14703;
assign w38878 = w14453 & w14640;
assign w38879 = w14638 & ~w16213;
assign w38880 = ~w16210 & ~w16209;
assign w38881 = ~w16196 & w14758;
assign w38882 = w1143 & w14745;
assign w38883 = w5987 & ~pi3245;
assign w38884 = ~w16226 & pi3245;
assign w38885 = ~w16226 & ~w38883;
assign w38886 = ~w5987 & w14734;
assign w38887 = w14823 & ~w6087;
assign w38888 = ~w38886 & w16230;
assign w38889 = ~w16227 & ~w16225;
assign w38890 = w14408 & w14882;
assign w38891 = ~w5987 & w14852;
assign w38892 = ~w16250 & ~w16249;
assign w38893 = ~w16259 & ~w14806;
assign w38894 = ~w10139 & w10593;
assign w38895 = w10139 & ~w10594;
assign w38896 = w10392 & ~w10099;
assign w38897 = w16268 & ~w10398;
assign w38898 = w16268 & ~w37777;
assign w38899 = w14518 & ~w15463;
assign w38900 = w14526 & ~w15045;
assign w38901 = w15056 & ~w16278;
assign w38902 = ~w16276 & ~w16275;
assign w38903 = w14450 & ~w15037;
assign w38904 = w15041 & ~w16300;
assign w38905 = w16301 & ~w16299;
assign w38906 = ~w16298 & ~w16297;
assign w38907 = ~w2979 & w14734;
assign w38908 = w14818 & ~w3112;
assign w38909 = ~w38907 & w16317;
assign w38910 = ~w7691 & ~w14805;
assign w38911 = w16318 & ~w16314;
assign w38912 = ~w2979 & w14852;
assign w38913 = ~w7691 & ~w14856;
assign w38914 = ~w16338 & ~w16337;
assign w38915 = ~w16347 & ~w14806;
assign w38916 = w10242 & ~w10594;
assign w38917 = w10242 & w10593;
assign w38918 = w10099 & w16357;
assign w38919 = ~w10099 & w16355;
assign w38920 = w14611 & ~w15041;
assign w38921 = ~w16364 & ~w16363;
assign w38922 = w14724 & w15456;
assign w38923 = w16369 & ~w16362;
assign w38924 = ~w5092 & ~pi0341;
assign w38925 = ~pi0343 & ~pi0342;
assign w38926 = ~w7561 & ~w14805;
assign w38927 = w14818 & ~w5200;
assign w38928 = w14823 & ~w5204;
assign w38929 = w5129 & w14745;
assign w38930 = w5092 & pi0343;
assign w38931 = ~w14499 & w16403;
assign w38932 = ~w14512 & ~w16407;
assign w38933 = w14453 & ~w15041;
assign w38934 = w14450 & ~w15024;
assign w38935 = w16424 & w16426;
assign w38936 = ~w14758 & ~w16402;
assign w38937 = ~w7561 & ~w14856;
assign w38938 = ~w16441 & ~w16440;
assign w38939 = ~w5092 & w14852;
assign w38940 = w14806 & ~pi0097;
assign w38941 = ~w38939 & w16453;
assign w38942 = ~w10140 & ~w10546;
assign w38943 = ~w10474 & ~w10099;
assign w38944 = ~w38942 & w16457;
assign w38945 = ~w10419 & ~w10594;
assign w38946 = ~w16461 & w16457;
assign w38947 = ~w16461 & w38944;
assign w38948 = w14534 & ~w15056;
assign w38949 = w14504 & ~w15037;
assign w38950 = w38532 & pi3518;
assign w38951 = w16470 & w14526;
assign w38952 = w14600 & w14652;
assign w38953 = ~w16495 & ~pi0709;
assign w38954 = w15029 & ~w16501;
assign w38955 = w14426 & w14484;
assign w38956 = ~w16507 & ~w16506;
assign w38957 = w3954 & ~pi3245;
assign w38958 = ~w16524 & pi3245;
assign w38959 = ~w16524 & ~w38957;
assign w38960 = w14818 & ~w4075;
assign w38961 = w14823 & ~w4083;
assign w38962 = ~w3954 & w14734;
assign w38963 = ~w38962 & ~w16527;
assign w38964 = w16532 & ~w15881;
assign w38965 = w16532 & w38791;
assign w38966 = ~w16525 & ~w16523;
assign w38967 = ~w16547 & ~w16546;
assign w38968 = w14806 & ~pi0098;
assign w38969 = ~w3954 & w14852;
assign w38970 = ~w38969 & ~w16558;
assign w38971 = w10044 & ~w10099;
assign w38972 = ~w10012 & ~w10594;
assign w38973 = ~w10012 & w10593;
assign w38974 = w16563 & w16571;
assign w38975 = ~w16563 & ~w16571;
assign w38976 = w16578 & w14583;
assign w38977 = ~w16582 & ~w16587;
assign w38978 = ~w16581 & ~w16577;
assign w38979 = ~w14526 & ~w16591;
assign w38980 = w15798 & w16593;
assign w38981 = w14611 & w14673;
assign w38982 = ~w14523 & ~w14602;
assign w38983 = w15486 & ~w16614;
assign w38984 = w16606 & w16604;
assign w38985 = ~w16598 & w14758;
assign w38986 = w14823 & ~w7950;
assign w38987 = w8013 & ~pi3245;
assign w38988 = ~w8013 & w14734;
assign w38989 = ~w14803 & w14813;
assign w38990 = w14818 & ~w7958;
assign w38991 = ~w16627 & w16637;
assign w38992 = w14364 & ~w15881;
assign w38993 = w14364 & w38791;
assign w38994 = ~w8013 & w14852;
assign w38995 = ~w16654 & ~w16653;
assign w38996 = w14806 & ~pi0099;
assign w38997 = w14806 & w16666;
assign w38998 = ~w7883 & ~w14856;
assign w38999 = ~w16676 & ~w16675;
assign w39000 = w16670 & ~w14806;
assign w39001 = w14852 & ~w35851;
assign w39002 = w14852 & ~w35850;
assign w39003 = w16687 & ~w16688;
assign w39004 = w14519 & w14426;
assign w39005 = w15813 & w16695;
assign w39006 = w14504 & ~w15041;
assign w39007 = w14490 & ~w15024;
assign w39008 = w14534 & ~w15045;
assign w39009 = ~w16702 & w14526;
assign w39010 = ~w14709 & ~w16710;
assign w39011 = ~w16697 & ~pi0709;
assign w39012 = w14611 & ~w15045;
assign w39013 = w15051 & ~w16721;
assign w39014 = ~w16719 & ~w16718;
assign w39015 = w16724 & ~w16717;
assign w39016 = w7883 & pi3245;
assign w39017 = ~pi3245 & ~w35851;
assign w39018 = ~pi3245 & ~w35850;
assign w39019 = ~w7883 & w14803;
assign w39020 = w14823 & ~w1540;
assign w39021 = w14734 & w35851;
assign w39022 = w14734 & w35850;
assign w39023 = w14818 & ~w1548;
assign w39024 = ~w16745 & ~w39022;
assign w39025 = ~w16745 & ~w39021;
assign w39026 = ~w16744 & w16743;
assign w39027 = ~w14758 & w16749;
assign w39028 = w10043 & w10593;
assign w39029 = ~w10043 & ~w10594;
assign w39030 = ~w10093 & w10550;
assign w39031 = ~w10093 & w37833;
assign w39032 = ~w10092 & ~w10099;
assign w39033 = ~w16758 & ~w16756;
assign w39034 = w16750 & ~w16761;
assign w39035 = ~w16689 & w16691;
assign w39036 = w10092 & ~w10594;
assign w39037 = ~w10092 & w10593;
assign w39038 = w16596 & w15519;
assign w39039 = w14611 & w14662;
assign w39040 = ~w14640 & ~w16779;
assign w39041 = w14450 & ~w14638;
assign w39042 = w16606 & ~w16788;
assign w39043 = ~w16776 & w16775;
assign w39044 = w14534 & w14665;
assign w39045 = w14504 & ~w14763;
assign w39046 = w14490 & ~w14689;
assign w39047 = w14524 & ~w14636;
assign w39048 = w14622 & ~pi3518;
assign w39049 = ~w14770 & pi3518;
assign w39050 = ~w15782 & ~w14630;
assign w39051 = ~w1002 & ~pi3245;
assign w39052 = ~w39051 & ~w16841;
assign w39053 = w14823 & ~w1187;
assign w39054 = ~w1002 & w14734;
assign w39055 = w14818 & ~w1191;
assign w39056 = ~w39054 & ~w16845;
assign w39057 = w16850 & ~w15881;
assign w39058 = w16850 & w38791;
assign w39059 = w16851 & ~w16843;
assign w39060 = ~w14422 & w16853;
assign w39061 = w39051 & ~w14851;
assign w39062 = ~w16867 & ~w16866;
assign w39063 = ~w16876 & ~w14806;
assign w39064 = ~w7819 & ~w14856;
assign w39065 = w14852 & ~w5448;
assign w39066 = w14852 & w36613;
assign w39067 = ~w16889 & ~w16888;
assign w39068 = w16883 & ~w14806;
assign w39069 = ~w16899 & w14806;
assign w39070 = ~w16899 & ~w39068;
assign w39071 = w14611 & w15022;
assign w39072 = w15051 & ~w16905;
assign w39073 = ~w16902 & w16775;
assign w39074 = w15037 & ~w16925;
assign w39075 = ~w15822 & ~w16927;
assign w39076 = ~w16930 & w16926;
assign w39077 = ~w16692 & ~w16924;
assign w39078 = ~w14512 & w14559;
assign w39079 = w14542 & ~w16939;
assign w39080 = ~w16941 & ~w16940;
assign w39081 = ~w16945 & ~pi0709;
assign w39082 = w14798 & w38823;
assign w39083 = w14798 & w38822;
assign w39084 = w14818 & ~w5617;
assign w39085 = ~w7819 & w14803;
assign w39086 = w14734 & ~w5448;
assign w39087 = w14734 & w36613;
assign w39088 = w14823 & ~w5613;
assign w39089 = ~w16953 & w16958;
assign w39090 = ~w14422 & w16961;
assign w39091 = w10506 & w10593;
assign w39092 = ~w10506 & ~w10594;
assign w39093 = w10140 & w10476;
assign w39094 = w10548 & ~w10476;
assign w39095 = w10548 & ~w39093;
assign w39096 = ~w10537 & ~w10099;
assign w39097 = w10538 & w16970;
assign w39098 = ~w16968 & ~w16970;
assign w39099 = ~w16968 & ~w39097;
assign w39100 = w10538 & w16972;
assign w39101 = w16900 & w16691;
assign w39102 = ~w10099 & ~w39095;
assign w39103 = ~w10099 & ~w39094;
assign w39104 = ~w10537 & w10593;
assign w39105 = w10537 & ~w10594;
assign w39106 = ~w16981 & w39103;
assign w39107 = ~w16981 & w39102;
assign w39108 = w14666 & ~w16990;
assign w39109 = ~w16993 & w16991;
assign w39110 = w14519 & ~w15486;
assign w39111 = w14763 & ~w16995;
assign w39112 = w15790 & w17001;
assign w39113 = w16989 & w16166;
assign w39114 = ~w15461 & ~pi0709;
assign w39115 = w14653 & ~w17019;
assign w39116 = ~w16195 & w14758;
assign w39117 = w14818 & ~w4933;
assign w39118 = ~w7787 & w14803;
assign w39119 = ~w4866 & w14734;
assign w39120 = ~w39119 & ~w17036;
assign w39121 = w14823 & ~w4941;
assign w39122 = ~w17035 & w17040;
assign w39123 = w17041 & ~w17034;
assign w39124 = ~w4866 & w14852;
assign w39125 = ~w7787 & ~w14856;
assign w39126 = ~w17057 & ~w17056;
assign w39127 = ~w17066 & ~w14806;
assign w39128 = ~w10343 & w17072;
assign w39129 = ~pi1975 & pi1974;
assign w39130 = w17073 & ~w10353;
assign w39131 = ~w10343 & ~w10099;
assign w39132 = w17078 & ~w10351;
assign w39133 = ~w14487 & w15714;
assign w39134 = w14518 & ~w17082;
assign w39135 = w14511 & ~w14559;
assign w39136 = w14450 & ~w14619;
assign w39137 = w17098 & w14495;
assign w39138 = ~w14577 & ~w17105;
assign w39139 = w17111 & w14487;
assign w39140 = ~w17116 & w14610;
assign w39141 = w17087 & w17083;
assign w39142 = ~w3484 & w14734;
assign w39143 = w14823 & ~w3576;
assign w39144 = ~w39142 & ~w17126;
assign w39145 = w14818 & ~w3580;
assign w39146 = w17131 & w14813;
assign w39147 = w17131 & w38550;
assign w39148 = w17132 & ~w17124;
assign w39149 = w3627 & w14745;
assign w39150 = w3484 & pi0343;
assign w39151 = w14544 & w15621;
assign w39152 = w14534 & ~w14622;
assign w39153 = w14504 & w15726;
assign w39154 = w14637 & ~pi3518;
assign w39155 = w17146 & w14557;
assign w39156 = ~w17145 & ~w17144;
assign w39157 = ~w17098 & ~w17156;
assign w39158 = w14666 & ~w17162;
assign w39159 = w17165 & w17151;
assign w39160 = ~w17143 & w14758;
assign w39161 = ~w17181 & ~w17180;
assign w39162 = ~w3484 & w14852;
assign w39163 = w14806 & ~pi0104;
assign w39164 = ~w39162 & w17193;
assign w39165 = w14408 & w14813;
assign w39166 = ~w14841 & w17198;
assign w39167 = w17200 & ~w17198;
assign w39168 = w17200 & ~w39166;
assign w39169 = w16442 & ~w14889;
assign w39170 = ~w14841 & w17209;
assign w39171 = w17211 & ~w17209;
assign w39172 = w17211 & ~w39170;
assign w39173 = ~w14888 & ~pi0108;
assign w39174 = ~w17216 & ~w17214;
assign w39175 = ~w14888 & ~pi0109;
assign w39176 = ~w14841 & w17221;
assign w39177 = w17220 & ~w14813;
assign w39178 = ~w14888 & ~pi0110;
assign w39179 = ~w14841 & w17227;
assign w39180 = w17226 & ~w14813;
assign w39181 = w14813 & w16691;
assign w39182 = w16868 & ~w14889;
assign w39183 = ~w14888 & ~pi0112;
assign w39184 = w14841 & w38823;
assign w39185 = w14841 & w38822;
assign w39186 = ~w17239 & ~w17237;
assign w39187 = ~w14841 & w17245;
assign w39188 = w17247 & ~w17245;
assign w39189 = w17247 & ~w39187;
assign w39190 = ~w14888 & ~pi0114;
assign w39191 = ~w17252 & ~w17250;
assign w39192 = ~w13782 & w17257;
assign w39193 = (~w17261 & w17258) | (~w17261 & w40075) | (w17258 & w40075);
assign w39194 = w13766 & pi0868;
assign w39195 = ~w17266 & ~w17262;
assign w39196 = ~w13758 & w17271;
assign w39197 = ~w17273 & w17275;
assign w39198 = ~w13490 & ~pi0868;
assign w39199 = ~w17281 & w10752;
assign w39200 = ~w10749 & w17285;
assign w39201 = w13490 & pi0868;
assign w39202 = w13183 & ~w17290;
assign w39203 = ~w17258 & w40076;
assign w39204 = (~w17301 & w17258) | (~w17301 & w40077) | (w17258 & w40077);
assign w39205 = w13183 & ~w17301;
assign w39206 = w17306 & w10752;
assign w39207 = ~w10749 & w17309;
assign w39208 = w17296 & ~w17317;
assign w39209 = ~w17296 & ~w17320;
assign w39210 = ~w17316 & w10752;
assign w39211 = w17306 & w13923;
assign w39212 = ~w13929 & w17334;
assign w39213 = ~w17281 & w13923;
assign w39214 = ~w13929 & w17340;
assign w39215 = ~w17316 & w13923;
assign w39216 = w17306 & w15185;
assign w39217 = ~w10750 & pi0121;
assign w39218 = ~w10750 & pi0122;
assign w39219 = ~w17316 & w15185;
assign w39220 = ~w10750 & pi0123;
assign w39221 = ~w17281 & w15185;
assign w39222 = ~w13922 & pi0124;
assign w39223 = ~w17281 & w15189;
assign w39224 = w17306 & w15189;
assign w39225 = ~w13922 & pi0126;
assign w39226 = ~w17316 & w15189;
assign w39227 = w15330 & w17373;
assign w39228 = ~w15330 & w15342;
assign w39229 = ~w15303 & w15317;
assign w39230 = ~w17387 & w15380;
assign w39231 = w15301 & pi2555;
assign w39232 = pi0127 & ~pi3427;
assign w39233 = pi0127 & w38654;
assign w39234 = ~pi2555 & ~w39232;
assign w39235 = ~pi2555 & ~w39233;
assign w39236 = ~w3484 & ~w15388;
assign w39237 = pi0128 & ~pi3427;
assign w39238 = pi0128 & w38654;
assign w39239 = ~pi2555 & ~w39237;
assign w39240 = ~pi2555 & ~w39238;
assign w39241 = w15376 & ~w15424;
assign w39242 = w15316 & pi2555;
assign w39243 = ~w17401 & ~w17399;
assign w39244 = w15330 & w17406;
assign w39245 = ~w15330 & w15424;
assign w39246 = ~w17408 & ~w17407;
assign w39247 = w17409 & w17378;
assign w39248 = ~w15303 & ~w15410;
assign w39249 = ~w17416 & w17417;
assign w39250 = ~w17420 & w37864;
assign w39251 = ~w17420 & w37865;
assign w39252 = pi0129 & ~w39251;
assign w39253 = pi0129 & ~w39250;
assign w39254 = w10049 & ~pi2758;
assign w39255 = ~pi2758 & ~w17423;
assign w39256 = ~w3484 & w14856;
assign w39257 = ~w39256 & ~w17174;
assign w39258 = w17425 & ~w17427;
assign w39259 = ~w17428 & ~w17423;
assign w39260 = ~w17428 & w39255;
assign w39261 = w17425 & ~w17430;
assign w39262 = ~w17429 & w17421;
assign w39263 = ~w12479 & ~w13799;
assign w39264 = ~w12092 & w17435;
assign w39265 = w17438 & w39400;
assign w39266 = ~pi0868 & w12981;
assign w39267 = ~pi0868 & w13775;
assign w39268 = w17440 & w17454;
assign w39269 = w17453 & w12749;
assign w39270 = ~w10749 & w17463;
assign w39271 = ~w13929 & w17468;
assign w39272 = ~w10750 & pi0132;
assign w39273 = ~w13922 & pi0133;
assign w39274 = ~w10690 & ~pi0134;
assign w39275 = ~w17486 & ~w10752;
assign w39276 = ~w17495 & w17499;
assign w39277 = w17495 & w17501;
assign w39278 = w13774 & ~pi0868;
assign w39279 = w17448 & ~pi0868;
assign w39280 = ~w17522 & ~w17524;
assign w39281 = ~w17525 & w17529;
assign w39282 = w17525 & w17531;
assign w39283 = ~w17542 & ~w13923;
assign w39284 = ~w10750 & ~pi0139;
assign w39285 = ~w10750 & pi0140;
assign w39286 = ~w13922 & ~pi0141;
assign w39287 = ~w13922 & pi0142;
assign w39288 = w17570 & ~pi1093;
assign w39289 = ~w10626 & ~w17585;
assign w39290 = pi0835 & ~w17586;
assign w39291 = w370 & w9954;
assign w39292 = w17588 & w17423;
assign w39293 = w17588 & ~w39255;
assign w39294 = w370 & ~w9954;
assign w39295 = ~pi3551 & ~pi0143;
assign w39296 = ~w39295 & w17592;
assign w39297 = w17593 & ~w17589;
assign w39298 = pi0143 & w17481;
assign w39299 = ~w17420 & w38164;
assign w39300 = ~w17420 & w38165;
assign w39301 = pi0144 & ~w39300;
assign w39302 = pi0144 & ~w39299;
assign w39303 = ~w17429 & w17601;
assign w39304 = ~w17607 & ~w10752;
assign w39305 = ~w17495 & w17610;
assign w39306 = w17495 & w17612;
assign w39307 = ~w17525 & w17615;
assign w39308 = w17525 & w17617;
assign w39309 = ~w17625 & ~w13923;
assign w39310 = ~w10750 & ~pi0147;
assign w39311 = ~w13922 & ~pi0148;
assign w39312 = ~w10690 & ~pi0149;
assign w39313 = ~w3484 & ~pi0835;
assign w39314 = w17641 & ~pi1041;
assign w39315 = ~pi1564 & pi1041;
assign w39316 = ~w17647 & w17646;
assign w39317 = ~w10626 & ~w17652;
assign w39318 = ~w39313 & w17654;
assign w39319 = w14420 & ~w15679;
assign w39320 = w15577 & ~w16272;
assign w39321 = w15452 & w16159;
assign w39322 = ~pi3426 & ~w17674;
assign w39323 = ~w10750 & pi0150;
assign w39324 = ~pi0715 & w17676;
assign w39325 = pi0715 & w17679;
assign w39326 = ~w13922 & pi0151;
assign w39327 = ~pi0715 & w17682;
assign w39328 = ~w10615 & w17687;
assign w39329 = pi0152 & w17481;
assign w39330 = ~w10750 & ~pi0153;
assign w39331 = ~w14406 & ~pi0715;
assign w39332 = ~pi0715 & ~w16464;
assign w39333 = ~w39332 & ~w17694;
assign w39334 = ~w10750 & ~pi0154;
assign w39335 = ~pi0715 & ~w16159;
assign w39336 = ~w39335 & ~w17700;
assign w39337 = ~w10750 & ~pi0155;
assign w39338 = ~pi0715 & w16272;
assign w39339 = ~w39338 & ~w17705;
assign w39340 = ~w10750 & pi0156;
assign w39341 = ~pi0715 & w14406;
assign w39342 = ~pi0715 & w15452;
assign w39343 = ~w10750 & ~pi0157;
assign w39344 = ~pi0715 & ~w15577;
assign w39345 = ~w39344 & ~w17718;
assign w39346 = ~w10750 & ~pi0158;
assign w39347 = ~pi0715 & w15679;
assign w39348 = ~w39347 & ~w17723;
assign w39349 = ~w10750 & pi0159;
assign w39350 = pi0715 & ~w37873;
assign w39351 = pi0715 & ~w37872;
assign w39352 = ~pi0715 & ~w16360;
assign w39353 = ~w39352 & ~w17728;
assign w39354 = ~w10750 & pi0160;
assign w39355 = ~pi0715 & w14420;
assign w39356 = ~w39355 & ~w17733;
assign w39357 = ~w10750 & pi0161;
assign w39358 = pi0715 & ~w38195;
assign w39359 = pi0715 & ~w38194;
assign w39360 = ~pi0715 & ~w15014;
assign w39361 = ~w39360 & ~w17738;
assign w39362 = ~w10750 & ~pi0162;
assign w39363 = ~w16574 & ~w17743;
assign w39364 = ~w10750 & ~pi0163;
assign w39365 = w17668 & ~w17748;
assign w39366 = ~w10750 & ~pi0164;
assign w39367 = w16773 & ~w17753;
assign w39368 = ~w10750 & ~pi0165;
assign w39369 = pi0715 & w38823;
assign w39370 = pi0715 & w38822;
assign w39371 = ~pi0715 & ~w17669;
assign w39372 = ~w10750 & ~pi0166;
assign w39373 = ~pi0715 & w16984;
assign w39374 = ~w39373 & ~w17764;
assign w39375 = ~w13922 & ~pi0167;
assign w39376 = ~w13922 & ~pi0168;
assign w39377 = ~w13922 & ~pi0169;
assign w39378 = ~w13922 & pi0170;
assign w39379 = ~w13922 & ~pi0171;
assign w39380 = ~w13922 & ~pi0172;
assign w39381 = ~w13922 & pi0173;
assign w39382 = ~w10750 & pi0174;
assign w39383 = pi0715 & ~w38222;
assign w39384 = pi0715 & ~w38221;
assign w39385 = ~pi0715 & w17080;
assign w39386 = ~w39385 & ~w17792;
assign w39387 = ~w13922 & pi0175;
assign w39388 = ~w13922 & pi0176;
assign w39389 = ~w13922 & ~pi0177;
assign w39390 = ~w13922 & ~pi0178;
assign w39391 = ~w13922 & ~pi0179;
assign w39392 = ~w13922 & ~pi0180;
assign w39393 = ~w13922 & ~pi0181;
assign w39394 = ~w13922 & pi0182;
assign w39395 = ~pi3426 & ~w17820;
assign w39396 = w17823 & w17822;
assign w39397 = ~w10750 & pi0183;
assign w39398 = w17823 & w17827;
assign w39399 = ~w17833 & ~w10752;
assign w39400 = w13799 & w12760;
assign w39401 = ~w17837 & ~w17836;
assign w39402 = ~w13192 & w17836;
assign w39403 = ~w39402 & ~w13799;
assign w39404 = w13192 & w17842;
assign w39405 = w13797 & pi0868;
assign w39406 = ~w17852 & ~w13923;
assign w39407 = ~w10750 & ~pi0187;
assign w39408 = ~w13922 & ~pi0188;
assign w39409 = ~pi0329 & ~w17874;
assign w39410 = ~pi0248 & ~w17873;
assign w39411 = ~w17881 & ~pi0248;
assign w39412 = ~w17889 & ~w17869;
assign w39413 = w17876 & ~pi0329;
assign w39414 = ~w17897 & pi0248;
assign w39415 = pi0278 & ~pi0248;
assign w39416 = w17900 & ~pi1017;
assign w39417 = ~w17872 & ~w17873;
assign w39418 = ~w17872 & w39410;
assign w39419 = w17881 & ~w17885;
assign w39420 = pi0248 & w17872;
assign w39421 = w17909 & ~pi1017;
assign w39422 = ~w17872 & pi0248;
assign w39423 = w17899 & ~pi0248;
assign w39424 = ~w17913 & ~w17869;
assign w39425 = ~w17889 & w17869;
assign w39426 = w17930 & ~w17890;
assign w39427 = ~pi1017 & ~w17933;
assign w39428 = ~pi0248 & w17941;
assign w39429 = w17936 & w17943;
assign w39430 = ~pi0278 & ~pi1017;
assign w39431 = ~w17947 & w17956;
assign w39432 = w17944 & ~pi0247;
assign w39433 = w17961 & pi0248;
assign w39434 = ~w17931 & ~pi0247;
assign w39435 = ~w17929 & ~pi0247;
assign w39436 = ~w17897 & ~pi0248;
assign w39437 = w17913 & w17869;
assign w39438 = ~w17872 & ~w17941;
assign w39439 = ~pi0248 & ~w17875;
assign w39440 = ~w39439 & ~w17873;
assign w39441 = w17930 & w17868;
assign w39442 = ~w17991 & ~w17990;
assign w39443 = w17994 & w17926;
assign w39444 = w17910 & ~w17972;
assign w39445 = w17996 & ~pi1017;
assign w39446 = ~w18001 & w18005;
assign w39447 = ~pi0831 & w18008;
assign w39448 = ~w1002 & w18009;
assign w39449 = pi0831 & w18008;
assign w39450 = pi0189 & w18008;
assign w39451 = pi0189 & w39449;
assign w39452 = ~w18011 & ~w39450;
assign w39453 = ~w18011 & ~w39451;
assign w39454 = ~w17440 & ~w18017;
assign w39455 = ~w17837 & w18022;
assign w39456 = ~w10749 & w18029;
assign w39457 = ~w13929 & w18034;
assign w39458 = w16090 & w10752;
assign w39459 = ~pi0695 & w37864;
assign w39460 = ~pi0695 & w37865;
assign w39461 = ~pi0192 & ~w39459;
assign w39462 = ~pi0192 & ~w39460;
assign w39463 = ~w18039 & w18041;
assign w39464 = w16090 & w13923;
assign w39465 = pi0695 & ~pi0193;
assign w39466 = ~w18046 & w18048;
assign w39467 = ~w10750 & pi0194;
assign w39468 = ~w13922 & pi0195;
assign w39469 = w10681 & ~w10719;
assign w39470 = ~w10690 & ~pi0196;
assign w39471 = w18062 & w17822;
assign w39472 = ~w10750 & pi0197;
assign w39473 = w18062 & w17827;
assign w39474 = ~w9999 & w18074;
assign w39475 = w14661 & w14664;
assign w39476 = w14672 & ~w14675;
assign w39477 = ~w14619 & w14622;
assign w39478 = ~w14661 & ~w14664;
assign w39479 = ~w14672 & w14675;
assign w39480 = w14619 & ~w14622;
assign w39481 = w18088 & w18081;
assign w39482 = ~w18078 & w18075;
assign w39483 = w18124 & w18120;
assign w39484 = w18115 & w18112;
assign w39485 = ~w18111 & w18110;
assign w39486 = w4674 & w3563;
assign w39487 = w4674 & w18110;
assign w39488 = w4674 & w39485;
assign w39489 = ~w18141 & w18110;
assign w39490 = ~w18110 & ~w5217;
assign w39491 = ~w18148 & w18153;
assign w39492 = w18073 & ~w9999;
assign w39493 = w18156 & w18072;
assign w39494 = w18110 & w5217;
assign w39495 = ~w18156 & w1178;
assign w39496 = ~w9999 & pi3518;
assign w39497 = ~pi3426 & w18165;
assign w39498 = ~w18162 & w18167;
assign w39499 = ~w18168 & ~w18167;
assign w39500 = ~w18168 & ~w39498;
assign w39501 = w4160 & pi0867;
assign w39502 = ~w10750 & ~pi0199;
assign w39503 = ~w10750 & pi0200;
assign w39504 = w5092 & pi0867;
assign w39505 = ~w18110 & ~pi0867;
assign w39506 = ~w10750 & pi0201;
assign w39507 = pi0867 & ~w36655;
assign w39508 = pi0867 & ~w36654;
assign w39509 = w10750 & w18184;
assign w39510 = ~w10750 & pi0202;
assign w39511 = w4523 & pi0867;
assign w39512 = w10750 & w18190;
assign w39513 = w13922 & ~w39499;
assign w39514 = w13922 & ~w39500;
assign w39515 = w3484 & pi0867;
assign w39516 = ~pi0867 & w18075;
assign w39517 = ~pi0867 & w39482;
assign w39518 = w10750 & ~w18202;
assign w39519 = ~w10750 & ~pi0205;
assign w39520 = ~w12092 & ~w12502;
assign w39521 = ~w18215 & w10752;
assign w39522 = ~w18215 & w13923;
assign w39523 = ~pi0211 & ~w39459;
assign w39524 = ~pi0211 & ~w39460;
assign w39525 = ~w18039 & w18237;
assign w39526 = pi0695 & ~pi0212;
assign w39527 = ~w18046 & w18243;
assign w39528 = w18215 & w15185;
assign w39529 = ~w10750 & ~pi0213;
assign w39530 = w18215 & w15189;
assign w39531 = ~w13192 & w18253;
assign w39532 = w13187 & ~w12495;
assign w39533 = ~w12092 & w12503;
assign w39534 = w18255 & w18258;
assign w39535 = w13192 & w18260;
assign w39536 = ~w18255 & w18264;
assign w39537 = ~w39536 & w10752;
assign w39538 = ~w18254 & w18265;
assign w39539 = ~w18255 & w18273;
assign w39540 = w18255 & w18275;
assign w39541 = w18277 & w10752;
assign w39542 = ~w10749 & w18280;
assign w39543 = w18277 & w13923;
assign w39544 = ~w13929 & w18285;
assign w39545 = ~w39536 & w13923;
assign w39546 = ~w18254 & w18288;
assign w39547 = ~w10750 & pi0219;
assign w39548 = ~w39536 & w15185;
assign w39549 = ~w18254 & w18296;
assign w39550 = ~w10750 & pi0220;
assign w39551 = w18277 & w15185;
assign w39552 = ~w13922 & pi0221;
assign w39553 = ~w39536 & w15189;
assign w39554 = ~w13922 & pi0222;
assign w39555 = w18277 & w15189;
assign w39556 = w1 & ~pi1426;
assign w39557 = ~pi3681 & pi2095;
assign w39558 = ~pi3641 & ~w18315;
assign w39559 = w18323 & pi0827;
assign w39560 = w18315 & ~pi0849;
assign w39561 = ~pi0699 & ~pi0849;
assign w39562 = ~pi0699 & w39560;
assign w39563 = ~pi0728 & w39561;
assign w39564 = ~pi0728 & w39562;
assign w39565 = pi0822 & ~w18315;
assign w39566 = ~pi0863 & w18315;
assign w39567 = ~pi0863 & ~w39565;
assign w39568 = ~pi0653 & w39566;
assign w39569 = ~pi0653 & w39567;
assign w39570 = ~pi0577 & w39568;
assign w39571 = ~pi0577 & w39569;
assign w39572 = pi0496 & ~w18315;
assign w39573 = ~pi0458 & w18315;
assign w39574 = ~pi0458 & ~w39572;
assign w39575 = ~pi0398 & w39573;
assign w39576 = ~pi0398 & w39574;
assign w39577 = ~pi0367 & w39575;
assign w39578 = ~pi0367 & w39576;
assign w39579 = ~pi0336 & w39577;
assign w39580 = ~pi0336 & w39578;
assign w39581 = w18315 & ~pi0303;
assign w39582 = ~pi0277 & w39581;
assign w39583 = ~pi0246 & w18347;
assign w39584 = ~pi0246 & w39582;
assign w39585 = pi0223 & w39583;
assign w39586 = pi0223 & w39584;
assign w39587 = ~pi0223 & ~w39583;
assign w39588 = ~pi0223 & ~w39584;
assign w39589 = ~w18359 & ~w39587;
assign w39590 = ~w18359 & ~w39588;
assign w39591 = w18358 & pi1722;
assign w39592 = ~w39591 & ~w18313;
assign w39593 = ~pi0248 & ~w17951;
assign w39594 = w18367 & ~w18365;
assign w39595 = w39593 & w18367;
assign w39596 = w18009 & ~w5448;
assign w39597 = w18009 & w36613;
assign w39598 = ~pi2599 & ~pi0955;
assign w39599 = ~w18374 & ~w18008;
assign w39600 = ~w18374 & ~w39449;
assign w39601 = pi0224 & ~w39599;
assign w39602 = pi0224 & ~w39600;
assign w39603 = ~w18373 & ~w39601;
assign w39604 = ~w18373 & ~w39602;
assign w39605 = w18376 & ~w18371;
assign w39606 = w17926 & ~w17983;
assign w39607 = ~w17976 & ~w17978;
assign w39608 = ~w39607 & w17990;
assign w39609 = w18382 & w18367;
assign w39610 = ~w4866 & w18009;
assign w39611 = pi0225 & ~w39599;
assign w39612 = pi0225 & ~w39600;
assign w39613 = ~w18387 & ~w39611;
assign w39614 = ~w18387 & ~w39612;
assign w39615 = w18391 & w17822;
assign w39616 = ~w10750 & pi0226;
assign w39617 = w18391 & w17827;
assign w39618 = ~w16001 & w10752;
assign w39619 = ~pi0228 & ~w39459;
assign w39620 = ~pi0228 & ~w39460;
assign w39621 = ~w18039 & w18400;
assign w39622 = ~w16001 & w13923;
assign w39623 = pi0695 & ~pi0229;
assign w39624 = ~w18046 & w18406;
assign w39625 = ~pi3426 & ~w18410;
assign w39626 = ~w10750 & pi0230;
assign w39627 = ~w13922 & pi0231;
assign w39628 = w18425 & w18366;
assign w39629 = ~w5987 & pi2599;
assign w39630 = ~w39629 & ~w18003;
assign w39631 = ~w18431 & ~w18008;
assign w39632 = ~w18431 & ~w39449;
assign w39633 = pi0709 & w38823;
assign w39634 = pi0709 & w38822;
assign w39635 = ~w18435 & pi0709;
assign w39636 = ~w18435 & ~w39081;
assign w39637 = ~w10750 & pi0233;
assign w39638 = ~w13922 & pi0234;
assign w39639 = ~pi3426 & ~w18443;
assign w39640 = pi0710 & ~w38885;
assign w39641 = pi0710 & ~w38884;
assign w39642 = w16196 & ~pi0710;
assign w39643 = w18446 & w18445;
assign w39644 = ~w10750 & ~pi0235;
assign w39645 = w18446 & w18451;
assign w39646 = w17976 & ~w17993;
assign w39647 = ~w18457 & w18366;
assign w39648 = w3954 & pi2599;
assign w39649 = ~w18463 & ~w18008;
assign w39650 = ~w18463 & ~w39449;
assign w39651 = pi0709 & ~w18467;
assign w39652 = ~w10750 & pi0238;
assign w39653 = ~w13922 & pi0239;
assign w39654 = w16008 & w10752;
assign w39655 = w18039 & ~w16841;
assign w39656 = w18039 & w39052;
assign w39657 = ~pi0240 & ~w39459;
assign w39658 = ~pi0240 & ~w39460;
assign w39659 = ~w18478 & w15173;
assign w39660 = w16008 & w13923;
assign w39661 = w18046 & ~w16841;
assign w39662 = w18046 & w39052;
assign w39663 = pi0695 & ~pi0241;
assign w39664 = ~w18484 & w14336;
assign w39665 = ~w10750 & pi0242;
assign w39666 = ~w10750 & pi0243;
assign w39667 = ~w13922 & pi0244;
assign w39668 = ~w13922 & pi0245;
assign w39669 = ~pi3681 & ~pi2394;
assign w39670 = w18358 & ~pi1723;
assign w39671 = ~w39670 & ~w18313;
assign w39672 = ~w17926 & w17983;
assign w39673 = ~w18514 & pi0955;
assign w39674 = ~w2979 & w18008;
assign w39675 = ~w18521 & ~w18008;
assign w39676 = ~w18521 & ~w39449;
assign w39677 = ~w39674 & w18522;
assign w39678 = w18008 & ~w36198;
assign w39679 = w18008 & ~w36197;
assign w39680 = ~w18530 & ~w18012;
assign w39681 = pi0710 & ~w38959;
assign w39682 = pi0710 & ~w38958;
assign w39683 = w18534 & w18445;
assign w39684 = ~w10750 & ~pi0249;
assign w39685 = pi0710 & ~w38272;
assign w39686 = pi0710 & ~w38271;
assign w39687 = w18539 & w18445;
assign w39688 = ~w10750 & ~pi0250;
assign w39689 = ~w10750 & pi0251;
assign w39690 = ~w15838 & ~pi0710;
assign w39691 = w18545 & w18445;
assign w39692 = w18534 & w18451;
assign w39693 = w18539 & w18451;
assign w39694 = ~w13922 & pi0254;
assign w39695 = w18545 & w18451;
assign w39696 = ~pi0255 & ~w39459;
assign w39697 = ~pi0255 & ~w39460;
assign w39698 = ~w18561 & w15173;
assign w39699 = w16027 & w10752;
assign w39700 = w18039 & ~w38568;
assign w39701 = w18039 & ~w38567;
assign w39702 = ~pi0256 & ~w39459;
assign w39703 = ~pi0256 & ~w39460;
assign w39704 = ~w18567 & w15173;
assign w39705 = pi0695 & ~pi0257;
assign w39706 = ~w18573 & w14336;
assign w39707 = w16027 & w13923;
assign w39708 = pi0695 & ~pi0258;
assign w39709 = ~w18046 & w18578;
assign w39710 = w18582 & w17822;
assign w39711 = ~w10750 & pi0259;
assign w39712 = w18586 & w17822;
assign w39713 = ~w10750 & pi0260;
assign w39714 = w18590 & w17822;
assign w39715 = ~w10750 & pi0261;
assign w39716 = pi0709 & ~w18594;
assign w39717 = ~w10750 & pi0262;
assign w39718 = w18582 & w17827;
assign w39719 = w18586 & w17827;
assign w39720 = w18590 & w17827;
assign w39721 = ~w13922 & pi0266;
assign w39722 = w16019 & w10752;
assign w39723 = w18039 & ~w38959;
assign w39724 = w18039 & ~w38958;
assign w39725 = ~pi0267 & ~w39459;
assign w39726 = ~pi0267 & ~w39460;
assign w39727 = ~w18614 & w15173;
assign w39728 = w16019 & w13923;
assign w39729 = w18046 & ~w38959;
assign w39730 = w18046 & ~w38958;
assign w39731 = pi0695 & ~pi0268;
assign w39732 = ~w18620 & w14336;
assign w39733 = pi0709 & ~w18623;
assign w39734 = ~w10750 & pi0269;
assign w39735 = ~w13922 & pi0270;
assign w39736 = pi0710 & ~w18631;
assign w39737 = ~w10750 & pi0271;
assign w39738 = ~w13922 & pi0272;
assign w39739 = ~w10750 & pi0273;
assign w39740 = w18641 & w18412;
assign w39741 = ~w10750 & pi0274;
assign w39742 = w18645 & w18412;
assign w39743 = ~w13922 & pi0275;
assign w39744 = w18641 & w18419;
assign w39745 = ~w13922 & pi0276;
assign w39746 = w18645 & w18419;
assign w39747 = ~pi3681 & ~pi2097;
assign w39748 = w18358 & ~pi1879;
assign w39749 = ~w39748 & ~w18313;
assign w39750 = w17967 & ~pi0247;
assign w39751 = w17931 & w18367;
assign w39752 = ~pi0278 & ~w39599;
assign w39753 = ~pi0278 & ~w39600;
assign w39754 = ~w18667 & ~w39752;
assign w39755 = ~w18667 & ~w39753;
assign w39756 = w18671 & w17822;
assign w39757 = ~w10750 & pi0279;
assign w39758 = w18671 & w17827;
assign w39759 = pi0710 & ~w18678;
assign w39760 = ~w10750 & ~pi0281;
assign w39761 = pi0710 & ~w38568;
assign w39762 = pi0710 & ~w38567;
assign w39763 = w16195 & ~pi0710;
assign w39764 = w18683 & w18445;
assign w39765 = ~w10750 & ~pi0282;
assign w39766 = w18451 & w18678;
assign w39767 = w18451 & ~w39759;
assign w39768 = ~w13922 & ~pi0283;
assign w39769 = w18683 & w18451;
assign w39770 = pi0709 & ~w18694;
assign w39771 = ~w10750 & pi0285;
assign w39772 = ~w13922 & pi0286;
assign w39773 = w15506 & ~pi0710;
assign w39774 = w18702 & w18445;
assign w39775 = ~w10750 & ~pi0287;
assign w39776 = w15505 & ~pi0710;
assign w39777 = w18707 & w18445;
assign w39778 = ~w10750 & ~pi0288;
assign w39779 = pi0710 & ~w38195;
assign w39780 = pi0710 & ~w38194;
assign w39781 = w15079 & ~pi0710;
assign w39782 = w18712 & w18445;
assign w39783 = ~w10750 & ~pi0289;
assign w39784 = w18702 & w18451;
assign w39785 = w18707 & w18451;
assign w39786 = w18712 & w18451;
assign w39787 = w18039 & ~w38885;
assign w39788 = w18039 & ~w38884;
assign w39789 = ~pi0293 & ~w39459;
assign w39790 = ~pi0293 & ~w39460;
assign w39791 = ~w18729 & w15173;
assign w39792 = w18046 & ~w38885;
assign w39793 = w18046 & ~w38884;
assign w39794 = pi0695 & ~pi0294;
assign w39795 = ~w18735 & w14336;
assign w39796 = ~w10750 & pi0295;
assign w39797 = ~w13922 & pi0296;
assign w39798 = pi0709 & ~w18747;
assign w39799 = ~w10750 & pi0297;
assign w39800 = ~w13922 & pi0298;
assign w39801 = pi0710 & ~w18755;
assign w39802 = ~w10750 & ~pi0299;
assign w39803 = w18451 & w18755;
assign w39804 = w18451 & ~w39801;
assign w39805 = ~w13922 & ~pi0300;
assign w39806 = ~w10750 & pi0301;
assign w39807 = ~w13922 & pi0302;
assign w39808 = ~pi3681 & ~pi2096;
assign w39809 = ~w18315 & pi0303;
assign w39810 = w18358 & ~pi1880;
assign w39811 = ~w39810 & ~w18313;
assign w39812 = pi0709 & ~w18779;
assign w39813 = ~w10750 & pi0304;
assign w39814 = pi0709 & ~w18784;
assign w39815 = ~w10750 & pi0305;
assign w39816 = ~w13922 & pi0306;
assign w39817 = ~w13922 & pi0307;
assign w39818 = pi0710 & ~w18795;
assign w39819 = ~w10750 & ~pi0308;
assign w39820 = pi0710 & ~w38222;
assign w39821 = pi0710 & ~w38221;
assign w39822 = w17143 & ~pi0710;
assign w39823 = w18800 & w18445;
assign w39824 = ~w10750 & ~pi0309;
assign w39825 = w18451 & w18795;
assign w39826 = w18451 & ~w39818;
assign w39827 = ~w13922 & ~pi0310;
assign w39828 = w18800 & w18451;
assign w39829 = w16038 & w10752;
assign w39830 = w18039 & ~w38272;
assign w39831 = w18039 & ~w38271;
assign w39832 = ~pi0312 & ~w39459;
assign w39833 = ~pi0312 & ~w39460;
assign w39834 = ~w18814 & w15173;
assign w39835 = w16038 & w13923;
assign w39836 = w18046 & ~w38272;
assign w39837 = w18046 & ~w38271;
assign w39838 = pi0695 & ~pi0313;
assign w39839 = ~w18820 & w14336;
assign w39840 = w15324 & w15277;
assign w39841 = ~w15388 & ~w6196;
assign w39842 = ~w15388 & w36727;
assign w39843 = pi0314 & ~pi3427;
assign w39844 = pi0314 & w38654;
assign w39845 = ~pi2555 & ~w39843;
assign w39846 = ~pi2555 & ~w39844;
assign w39847 = ~w15391 & ~w18827;
assign w39848 = w18830 & w17822;
assign w39849 = ~w10750 & pi0315;
assign w39850 = w18830 & w17827;
assign w39851 = pi0710 & ~w38519;
assign w39852 = pi0710 & ~w38518;
assign w39853 = w18837 & w18445;
assign w39854 = ~w10750 & ~pi0317;
assign w39855 = w16598 & ~pi0710;
assign w39856 = w18842 & w18445;
assign w39857 = ~w10750 & ~pi0318;
assign w39858 = w18837 & w18451;
assign w39859 = w18842 & w18451;
assign w39860 = ~w10750 & pi0321;
assign w39861 = ~w13922 & pi0322;
assign w39862 = pi0710 & ~w37873;
assign w39863 = pi0710 & ~w37872;
assign w39864 = pi0710 & ~w18862;
assign w39865 = ~w10750 & ~pi0323;
assign w39866 = w18451 & w18862;
assign w39867 = w18451 & ~w39864;
assign w39868 = ~w13922 & ~pi0324;
assign w39869 = w15449 & w17425;
assign w39870 = ~w10750 & ~pi0325;
assign w39871 = ~w13922 & ~pi0326;
assign w39872 = ~pi0327 & ~w39459;
assign w39873 = ~pi0327 & ~w39460;
assign w39874 = ~w18039 & w18881;
assign w39875 = pi0695 & ~pi0328;
assign w39876 = ~w18046 & w18887;
assign w39877 = w4160 & w18008;
assign w39878 = w17967 & pi0955;
assign w39879 = ~w18898 & ~w18008;
assign w39880 = ~w18898 & ~w39449;
assign w39881 = ~w18897 & w18899;
assign w39882 = w15377 & pi2555;
assign w39883 = pi0330 & ~pi3427;
assign w39884 = pi0330 & w38654;
assign w39885 = ~pi2555 & ~w39883;
assign w39886 = ~pi2555 & ~w39884;
assign w39887 = ~w5092 & w18008;
assign w39888 = w17944 & w18367;
assign w39889 = ~w39887 & w18912;
assign w39890 = ~pi2021 & ~pi3518;
assign w39891 = ~w18919 & w18926;
assign w39892 = ~w18927 & w10750;
assign w39893 = ~w18927 & w13922;
assign w39894 = ~pi0334 & ~w39459;
assign w39895 = ~pi0334 & ~w39460;
assign w39896 = ~w18039 & w18941;
assign w39897 = pi0695 & ~pi0335;
assign w39898 = ~w18046 & w18947;
assign w39899 = ~pi3681 & ~pi1881;
assign w39900 = w18358 & ~pi1724;
assign w39901 = ~w39900 & ~w18313;
assign w39902 = ~w10750 & pi0337;
assign w39903 = ~w15449 & ~w17425;
assign w39904 = w18960 & w18412;
assign w39905 = ~w10750 & pi0338;
assign w39906 = ~w13922 & pi0339;
assign w39907 = w18960 & w18419;
assign w39908 = ~w13922 & pi0340;
assign w39909 = ~pi0714 & pi0410;
assign w39910 = w18975 & ~w18978;
assign w39911 = w18984 & ~w18985;
assign w39912 = ~w16051 & w10752;
assign w39913 = w18039 & ~w38519;
assign w39914 = w18039 & ~w38518;
assign w39915 = ~pi0344 & ~w39459;
assign w39916 = ~pi0344 & ~w39460;
assign w39917 = ~w18991 & w15173;
assign w39918 = ~w16051 & w13923;
assign w39919 = pi0695 & ~pi0345;
assign w39920 = ~w18046 & w18996;
assign w39921 = w19001 & w18412;
assign w39922 = ~w10750 & ~pi0346;
assign w39923 = ~w10750 & pi0347;
assign w39924 = w17425 & ~w14412;
assign w39925 = w17425 & w38325;
assign w39926 = w19001 & w18419;
assign w39927 = ~w13922 & pi0349;
assign w39928 = w18008 & w36655;
assign w39929 = w18008 & w36654;
assign w39930 = w19019 & ~w19022;
assign w39931 = ~w17947 & ~w19023;
assign w39932 = w19028 & ~w39929;
assign w39933 = w19028 & ~w39928;
assign w39934 = ~w19037 & pi2515;
assign w39935 = w19041 & ~w19033;
assign w39936 = w3954 & w6609;
assign w39937 = w19047 & pi3563;
assign w39938 = w19049 & pi3560;
assign w39939 = w19047 & pi3565;
assign w39940 = pi3566 & w19067;
assign w39941 = pi3566 & w19069;
assign w39942 = pi3566 & ~pi3560;
assign w39943 = ~w19070 & ~w19068;
assign w39944 = w19050 & pi4072;
assign w39945 = w19053 & pi4048;
assign w39946 = w19060 & pi4144;
assign w39947 = w19063 & pi4096;
assign w39948 = w39940 & pi4168;
assign w39949 = w39941 & pi4192;
assign w39950 = w19071 & pi4216;
assign w39951 = w19073 & pi4120;
assign w39952 = ~w19087 & ~w19086;
assign w39953 = w19092 & w19094;
assign w39954 = ~w19096 & ~w19033;
assign w39955 = ~w19096 & w39935;
assign w39956 = w5987 & w6609;
assign w39957 = w19071 & pi4215;
assign w39958 = w19053 & pi4047;
assign w39959 = w19063 & pi4095;
assign w39960 = w19050 & pi4071;
assign w39961 = w39940 & pi4167;
assign w39962 = w39941 & pi4191;
assign w39963 = w19060 & pi4143;
assign w39964 = w19073 & pi4119;
assign w39965 = ~w19113 & ~w19112;
assign w39966 = w19118 & w19094;
assign w39967 = ~w19121 & ~w19033;
assign w39968 = ~w19121 & w39935;
assign w39969 = w2979 & w6609;
assign w39970 = w7691 & w2251;
assign w39971 = w19060 & pi4142;
assign w39972 = w19053 & pi4046;
assign w39973 = w19063 & pi4094;
assign w39974 = w19050 & pi4070;
assign w39975 = w39941 & pi4190;
assign w39976 = w39940 & pi4166;
assign w39977 = w19071 & pi4214;
assign w39978 = w19073 & pi4118;
assign w39979 = ~w19138 & ~w19137;
assign w39980 = w19143 & w19094;
assign w39981 = ~w19146 & ~w19033;
assign w39982 = ~w19146 & w39935;
assign w39983 = pi1422 & ~w36198;
assign w39984 = pi1422 & ~w36197;
assign w39985 = w7659 & w2257;
assign w39986 = w19050 & pi4069;
assign w39987 = w19071 & pi4213;
assign w39988 = w19060 & pi4141;
assign w39989 = w19063 & pi4093;
assign w39990 = w39941 & pi4189;
assign w39991 = w39940 & pi4165;
assign w39992 = w19053 & pi4045;
assign w39993 = w19073 & pi4117;
assign w39994 = ~w19164 & ~w19163;
assign w39995 = w19169 & w7230;
assign w39996 = ~w19174 & ~w19033;
assign w39997 = ~w19174 & w39935;
assign w39998 = ~w19173 & w19175;
assign w39999 = w7626 & w2251;
assign w40000 = w19050 & pi4068;
assign w40001 = w19053 & pi4044;
assign w40002 = w19060 & pi4140;
assign w40003 = w19063 & pi4092;
assign w40004 = w39941 & pi4188;
assign w40005 = w39940 & pi4164;
assign w40006 = w19071 & pi4212;
assign w40007 = w19073 & pi4116;
assign w40008 = ~w19190 & ~w19189;
assign w40009 = w19195 & w19094;
assign w40010 = ~w19198 & ~w19033;
assign w40011 = ~w19198 & w39935;
assign w40012 = w4160 & w6609;
assign w40013 = w7593 & w2251;
assign w40014 = w19071 & pi4211;
assign w40015 = w19060 & pi4139;
assign w40016 = w19063 & pi4091;
assign w40017 = w19050 & pi4067;
assign w40018 = w39941 & pi4187;
assign w40019 = w39940 & pi4163;
assign w40020 = w19053 & pi4043;
assign w40021 = w19073 & pi4115;
assign w40022 = ~w19215 & ~w19214;
assign w40023 = w19220 & w19094;
assign w40024 = ~w19223 & ~w19033;
assign w40025 = ~w19223 & w39935;
assign w40026 = w5092 & w6609;
assign w40027 = w7561 & w2251;
assign w40028 = w19053 & pi4042;
assign w40029 = w19063 & pi4090;
assign w40030 = w19071 & pi4210;
assign w40031 = w19060 & pi4138;
assign w40032 = w39940 & pi4162;
assign w40033 = w39941 & pi4186;
assign w40034 = w19050 & pi4066;
assign w40035 = w19073 & pi4114;
assign w40036 = ~w19240 & ~w19239;
assign w40037 = w19245 & w19094;
assign w40038 = ~w19248 & ~w19033;
assign w40039 = ~w19248 & w39935;
assign w40040 = pi1422 & ~w36655;
assign w40041 = pi1422 & ~w36654;
assign w40042 = w19050 & pi4065;
assign w40043 = w19071 & pi4209;
assign w40044 = w19060 & pi4137;
assign w40045 = w19063 & pi4089;
assign w40046 = w39940 & pi4161;
assign w40047 = w39941 & pi4185;
assign w40048 = w19053 & pi4041;
assign w40049 = w12139 & w12323;
assign w40050 = ~w12294 & w12332;
assign w40051 = w12294 & ~w12332;
assign w40052 = w12333 & w12399;
assign w40053 = ~w12333 & ~w12399;
assign w40054 = ~w12254 & w12429;
assign w40055 = w12430 & w12449;
assign w40056 = w12742 & w13798;
assign w40057 = w13183 & ~w13893;
assign w40058 = w13183 & ~w14082;
assign w40059 = w13183 & ~w17261;
assign w40060 = ~w17289 & ~w17290;
assign w40061 = w13183 & ~w17320;
assign w40062 = w26725 & w26740;
assign w40063 = ~w10920 & w10934;
assign w40064 = w11045 & ~w11041;
assign w40065 = w11720 & w11755;
assign w40066 = ~w11720 & ~w11755;
assign w40067 = ~w11999 & w12012;
assign w40068 = ~w12139 & w12110;
assign w40069 = w12139 & w12391;
assign w40070 = w12352 & ~w12110;
assign w40071 = w13604 & w13623;
assign w40072 = ~w13604 & ~w13623;
assign w40073 = w13491 & w13877;
assign w40074 = w13780 & ~w13179;
assign w40075 = ~w17260 & ~w17261;
assign w40076 = ~w13760 & ~w17298;
assign w40077 = w13760 & ~w17301;
assign w40078 = w37935 & w12072;
assign w40079 = ~w17514 & ~w17513;
assign w40080 = ~w17518 & w17519;
assign w40081 = ~w17521 & w10752;
assign w40082 = ~w17521 & w13923;
assign w40083 = ~w17521 & w15185;
assign w40084 = ~w17521 & w15189;
assign w40085 = ~w38561 & w15146;
assign w40086 = ~w38561 & ~pi0868;
assign w40087 = ~w38561 & pi0868;
assign w40088 = (~w332 & ~w35573) | (~w332 & ~w331) | (~w35573 & ~w331);
assign w40089 = (~w472 & w35635) | (~w472 & ~w498) | (w35635 & ~w498);
assign w40090 = (w580 & ~w35667) | (w580 & ~w521) | (~w35667 & ~w521);
assign w40091 = (pi0637 & ~w35687) | (pi0637 & ~w536) | (~w35687 & ~w536);
assign w40092 = (~pi0753 & ~w35700) | (~pi0753 & ~w468) | (~w35700 & ~w468);
assign w40093 = (~w498 & ~w35711) | (~w498 & ~w561) | (~w35711 & ~w561);
assign w40094 = (w904 & w35741) | (w904 & ~w886) | (w35741 & ~w886);
assign w40095 = (~w1620 & ~w35841) | (~w1620 & ~w1618) | (~w35841 & ~w1618);
assign w40096 = (~pi2913 & ~w35919) | (~pi2913 & ~w2181) | (~w35919 & ~w2181);
assign w40097 = pi2769 & w1324;
assign w40098 = ~w2264 & ~w1657;
assign w40099 = (w542 & ~w36000) | (w542 & ~w530) | (~w36000 & ~w530);
assign w40100 = (pi0679 & w36023) | (pi0679 & ~w2462) | (w36023 & ~w2462);
assign w40101 = (~w36061 & ~w36060) | (~w36061 & ~w2462) | (~w36060 & ~w2462);
assign w40102 = (pi1422 & w36132) | (pi1422 & ~w342) | (w36132 & ~w342);
assign w40103 = (~w3414 & ~w36188) | (~w3414 & ~w3412) | (~w36188 & ~w3412);
assign w40104 = (~w2643 & w36287) | (~w2643 & ~w2607) | (w36287 & ~w2607);
assign w40105 = (~w36385 & ~w36386) | (~w36385 & ~w647) | (~w36386 & ~w647);
assign w40106 = (w715 & ~w36384) | (w715 & ~w647) | (~w36384 & ~w647);
assign w40107 = (w487 & ~w36466) | (w487 & ~w561) | (~w36466 & ~w561);
assign w40108 = (w2761 & ~w36569) | (w2761 & ~w5366) | (~w36569 & ~w5366);
assign w40109 = (~w36645 & ~w36644) | (~w36645 & ~w5893) | (~w36644 & ~w5893);
assign w40110 = (~pi1331 & ~w36713) | (~pi1331 & ~w2132) | (~w36713 & ~w2132);
assign w40111 = (~w6552 & w36776) | (~w6552 & ~w797) | (w36776 & ~w797);
assign w40112 = (w715 & ~w36791) | (w715 & ~w647) | (~w36791 & ~w647);
assign w40113 = (~w36806 & ~w36807) | (~w36806 & ~w2227) | (~w36807 & ~w2227);
assign w40114 = (~pi0540 & ~w36867) | (~pi0540 & ~w6688) | (~w36867 & ~w6688);
assign w40115 = (~pi2540 & ~w36925) | (~pi2540 & ~w184) | (~w36925 & ~w184);
assign w40116 = (~pi2549 & ~w36933) | (~pi2549 & ~w184) | (~w36933 & ~w184);
assign w40117 = (~pi2646 & ~w36941) | (~pi2646 & ~w184) | (~w36941 & ~w184);
assign w40118 = (~pi2551 & ~w36949) | (~pi2551 & ~w184) | (~w36949 & ~w184);
assign w40119 = (~pi2553 & ~w36957) | (~pi2553 & ~w184) | (~w36957 & ~w184);
assign w40120 = (~pi2645 & ~w36965) | (~pi2645 & ~w184) | (~w36965 & ~w184);
assign w40121 = (~pi2797 & ~w36973) | (~pi2797 & ~w184) | (~w36973 & ~w184);
assign w40122 = (~pi2644 & ~w36981) | (~pi2644 & ~w184) | (~w36981 & ~w184);
assign w40123 = (~pi2796 & ~w36989) | (~pi2796 & ~w184) | (~w36989 & ~w184);
assign w40124 = (~pi2794 & ~w36995) | (~pi2794 & ~w184) | (~w36995 & ~w184);
assign w40125 = (~pi2788 & ~w37001) | (~pi2788 & ~w184) | (~w37001 & ~w184);
assign w40126 = (~pi2953 & ~w37005) | (~pi2953 & ~w184) | (~w37005 & ~w184);
assign w40127 = (~w7393 & ~w37020) | (~w7393 & ~w184) | (~w37020 & ~w184);
assign w40128 = (~w7401 & ~w37023) | (~w7401 & ~w184) | (~w37023 & ~w184);
assign w40129 = w903 & w40094;
assign w40130 = (w35939 & w35940) | (w35939 & ~w886) | (w35940 & ~w886);
assign w40131 = w6616 & w1324;
assign w40132 = w2891 & w40094;
assign w40133 = (w36655 & w36654) | (w36655 & ~w5893) | (w36654 & ~w5893);
assign w40134 = ~w3432 & w40103;
assign w40135 = (w9038 & ~w37678) | (w9038 & ~w9857) | (~w37678 & ~w9857);
assign w40136 = (w9383 & ~w37695) | (w9383 & ~w9857) | (~w37695 & ~w9857);
assign w40137 = (w9434 & ~w37697) | (w9434 & ~w9857) | (~w37697 & ~w9857);
assign w40138 = (w9496 & ~w37699) | (w9496 & ~w9857) | (~w37699 & ~w9857);
assign w40139 = (~w10663 & ~w37834) | (~w10663 & ~w10660) | (~w37834 & ~w10660);
assign w40140 = w10747 & w40209;
assign w40141 = (pi3245 & ~w37871) | (pi3245 & ~w5319) | (~w37871 & ~w5319);
assign w40142 = (w13687 & ~w38151) | (w13687 & ~w13745) | (~w38151 & ~w13745);
assign w40143 = (~w38160 & ~w38159) | (~w38160 & ~w5893) | (~w38159 & ~w5893);
assign w40144 = ~pi0979 & w6668;
assign w40145 = w10747 & w40210;
assign w40146 = ~pi0714 & w40211;
assign w40147 = (~w14024 & ~w38187) | (~w14024 & ~w10625) | (~w38187 & ~w10625);
assign w40148 = (pi3245 & ~w38193) | (pi3245 & ~w4748) | (~w38193 & ~w4748);
assign w40149 = (pi3245 & ~w38220) | (pi3245 & ~w3710) | (~w38220 & ~w3710);
assign w40150 = (pi3245 & ~w38270) | (pi3245 & ~w3194) | (~w38270 & ~w3194);
assign w40151 = (~w38285 & ~w38284) | (~w38285 & ~w3412) | (~w38284 & ~w3412);
assign w40152 = (~w14433 & ~w38331) | (~w14433 & ~w14430) | (~w38331 & ~w14430);
assign w40153 = (w14427 & w38335) | (w14427 & ~w14429) | (w38335 & ~w14429);
assign w40154 = (~w38420 & ~w38421) | (~w38420 & ~w14399) | (~w38421 & ~w14399);
assign w40155 = (~w38426 & ~w38427) | (~w38426 & ~w14399) | (~w38427 & ~w14399);
assign w40156 = (~w38431 & ~w38432) | (~w38431 & ~w14399) | (~w38432 & ~w14399);
assign w40157 = (~w38455 & ~w38456) | (~w38455 & ~w14399) | (~w38456 & ~w14399);
assign w40158 = (pi3245 & ~w38517) | (pi3245 & ~w4379) | (~w38517 & ~w4379);
assign w40159 = ~w14036 & w40148;
assign w40160 = (w14889 & ~w38559) | (w14889 & ~w15139) | (~w38559 & ~w15139);
assign w40161 = (pi3245 & ~w38566) | (pi3245 & ~w5052) | (~w38566 & ~w5052);
assign w40162 = (~w15243 & ~w38598) | (~w15243 & ~w15201) | (~w38598 & ~w15201);
assign w40163 = (pi1897 & w38580) | (pi1897 & ~w15203) | (w38580 & ~w15203);
assign w40164 = (~w38643 & ~w38642) | (~w38643 & ~w15233) | (~w38642 & ~w15233);
assign w40165 = (w10593 & ~w38678) | (w10593 & ~w15447) | (~w38678 & ~w15447);
assign w40166 = (w10593 & ~w38679) | (w10593 & ~w15448) | (~w38679 & ~w15448);
assign w40167 = (w10099 & ~w38714) | (w10099 & ~w10360) | (~w38714 & ~w10360);
assign w40168 = ~w14987 & w40158;
assign w40169 = (~pi0343 & ~w38786) | (~pi0343 & ~w3194) | (~w38786 & ~w3194);
assign w40170 = (w14889 & ~w38808) | (w14889 & ~w15932) | (~w38808 & ~w15932);
assign w40171 = ~w14110 & w40149;
assign w40172 = (w10099 & ~w38864) | (w10099 & ~w10402) | (~w38864 & ~w10402);
assign w40173 = (pi3245 & ~w38883) | (pi3245 & ~w6176) | (~w38883 & ~w6176);
assign w40174 = ~w14290 & w40150;
assign w40175 = (w10277 & ~w37769) | (w10277 & ~w10354) | (~w37769 & ~w10354);
assign w40176 = ~w10758 & w40141;
assign w40177 = (~pi0343 & ~w38930) | (~pi0343 & ~w5319) | (~w38930 & ~w5319);
assign w40178 = (~w16457 & ~w38944) | (~w16457 & ~w10402) | (~w38944 & ~w10402);
assign w40179 = (pi3245 & ~w38957) | (pi3245 & ~w4140) | (~w38957 & ~w4140);
assign w40180 = (pi3245 & ~w38987) | (pi3245 & ~w8080) | (~w38987 & ~w8080);
assign w40181 = (~w39018 & ~w39017) | (~w39018 & ~w1618) | (~w39017 & ~w1618);
assign w40182 = (~w39066 & ~w39065) | (~w39066 & ~w5632) | (~w39065 & ~w5632);
assign w40183 = (~w39086 & ~w39087) | (~w39086 & ~w5632) | (~w39087 & ~w5632);
assign w40184 = (~w10476 & ~w39093) | (~w10476 & ~w10402) | (~w39093 & ~w10402);
assign w40185 = (~w39103 & ~w39102) | (~w39103 & ~w10402) | (~w39102 & ~w10402);
assign w40186 = (~pi0343 & ~w39150) | (~pi0343 & ~w3710) | (~w39150 & ~w3710);
assign w40187 = (w14889 & ~w39169) | (w14889 & ~w17203) | (~w39169 & ~w17203);
assign w40188 = (w14889 & ~w39182) | (w14889 & ~w17232) | (~w39182 & ~w17232);
assign w40189 = ~w16524 & w40179;
assign w40190 = (w39265 & w17439) | (w39265 & ~w13192) | (w17439 & ~w13192);
assign w40191 = ~w16226 & w40173;
assign w40192 = ~w15170 & w40161;
assign w40193 = (~w17842 & ~w39404) | (~w17842 & ~w12505) | (~w39404 & ~w12505);
assign w40194 = (w17873 & ~w39440) | (w17873 & ~w17985) | (~w39440 & ~w17985);
assign w40195 = (~w14622 & ~w39477) | (~w14622 & ~w18085) | (~w39477 & ~w18085);
assign w40196 = (w14622 & ~w39480) | (w14622 & ~w18092) | (~w39480 & ~w18092);
assign w40197 = (~w18167 & ~w39498) | (~w18167 & ~w18154) | (~w39498 & ~w18154);
assign w40198 = (~pi0867 & ~w39501) | (~pi0867 & ~w4379) | (~w39501 & ~w4379);
assign w40199 = (~pi0867 & ~w39504) | (~pi0867 & ~w5319) | (~w39504 & ~w5319);
assign w40200 = (~pi2599 & ~w39648) | (~pi2599 & ~w4140) | (~w39648 & ~w4140);
assign w40201 = (~w18347 & ~w39582) | (~w18347 & ~w18340) | (~w39582 & ~w18340);
assign w40202 = (~w39583 & ~w39584) | (~w39583 & ~w18340) | (~w39584 & ~w18340);
assign w40203 = (~w39679 & ~w39678) | (~w39679 & ~w3412) | (~w39678 & ~w3412);
assign w40204 = (~w6609 & ~w39936) | (~w6609 & ~w4140) | (~w39936 & ~w4140);
assign w40205 = (~w6609 & ~w39956) | (~w6609 & ~w6176) | (~w39956 & ~w6176);
assign w40206 = (~w6609 & ~w39969) | (~w6609 & ~w3194) | (~w39969 & ~w3194);
assign w40207 = (~w6609 & ~w40012) | (~w6609 & ~w4379) | (~w40012 & ~w4379);
assign w40208 = (~w6609 & ~w40026) | (~w6609 & ~w5319) | (~w40026 & ~w5319);
assign w40209 = pi0979 & w6668;
assign w40210 = ~pi0979 & w6668;
assign w40211 = ~pi0979 & w6668;
assign one = 1;
assign po0000 = ~w10;// level 5
assign po0001 = ~w10;// level 5
assign po0002 = ~w10;// level 5
assign po0003 = ~w10;// level 5
assign po0004 = ~w10;// level 5
assign po0005 = ~w10;// level 5
assign po0006 = ~w10;// level 5
assign po0007 = ~w10;// level 5
assign po0008 = ~w10;// level 5
assign po0009 = w11;// level 1
assign po0010 = pi3397;// level 0
assign po0011 = ~w3;// level 2
assign po0012 = ~pi3452;// level 0
assign po0013 = w192;// level 16
assign po0014 = w186;// level 13
assign po0015 = ~w181;// level 13
assign po0016 = pi3626;// level 0
assign po0017 = ~w182;// level 13
assign po0018 = w197;// level 15
assign po0019 = pi3621;// level 0
assign po0020 = ~w200;// level 2
assign po0021 = w201;// level 1
assign po0022 = ~w202;// level 2
assign po0023 = ~w204;// level 2
assign po0024 = ~pi3350;// level 0
assign po0025 = pi3627;// level 0
assign po0026 = w249;// level 9
assign po0027 = w294;// level 9
assign po0028 = ~w297;// level 2
assign po0029 = pi0959;// level 0
assign po0030 = ~w300;// level 2
assign po0031 = pi0887;// level 0
assign po0032 = ~w305;// level 3
assign po0033 = pi0941;// level 0
assign po0034 = ~w309;// level 3
assign po0035 = pi0792;// level 0
assign po0036 = ~w314;// level 3
assign po0037 = pi0790;// level 0
assign po0038 = ~w318;// level 3
assign po0039 = pi0738;// level 0
assign po0040 = pi1771;// level 0
assign po0041 = ~w319;// level 1
assign po0042 = pi3648;// level 0
assign po0043 = w320;// level 1
assign po0044 = w2266;// level 28
assign po0045 = w2269;// level 28
assign po0046 = w2272;// level 28
assign po0047 = w2275;// level 28
assign po0048 = w2277;// level 28
assign po0049 = w2278;// level 28
assign po0050 = w2279;// level 28
assign po0051 = w2280;// level 28
assign po0052 = ~w2285;// level 27
assign po0053 = one;// level 0
assign po0054 = one;// level 0
assign po0055 = one;// level 0
assign po0056 = one;// level 0
assign po0057 = one;// level 0
assign po0058 = one;// level 0
assign po0059 = one;// level 0
assign po0060 = one;// level 0
assign po0061 = w6627;// level 32
assign po0062 = w6654;// level 29
assign po0063 = w6656;// level 29
assign po0064 = w6658;// level 29
assign po0065 = w6659;// level 29
assign po0066 = w6662;// level 30
assign po0067 = w6664;// level 29
assign po0068 = w6665;// level 30
assign po0069 = w6666;// level 29
assign po0070 = ~w6672;// level 32
assign po0071 = one;// level 0
assign po0072 = one;// level 0
assign po0073 = one;// level 0
assign po0074 = one;// level 0
assign po0075 = one;// level 0
assign po0076 = one;// level 0
assign po0077 = one;// level 0
assign po0078 = one;// level 0
assign po0079 = one;// level 0
assign po0080 = w7184;// level 24
assign po0081 = w7217;// level 27
assign po0082 = w7219;// level 27
assign po0083 = w7222;// level 27
assign po0084 = w7224;// level 27
assign po0085 = w7226;// level 27
assign po0086 = w7227;// level 27
assign po0087 = w7228;// level 27
assign po0088 = w7229;// level 27
assign po0089 = w7241;// level 14
assign po0090 = one;// level 0
assign po0091 = one;// level 0
assign po0092 = one;// level 0
assign po0093 = one;// level 0
assign po0094 = one;// level 0
assign po0095 = one;// level 0
assign po0096 = one;// level 0
assign po0097 = one;// level 0
assign po0098 = one;// level 0
assign po0099 = ~w7252;// level 17
assign po0100 = ~w7263;// level 17
assign po0101 = ~w7274;// level 17
assign po0102 = ~w7285;// level 17
assign po0103 = ~w7296;// level 17
assign po0104 = ~w7307;// level 17
assign po0105 = ~w7318;// level 17
assign po0106 = ~w7329;// level 17
assign po0107 = ~w7337;// level 17
assign po0108 = ~w7345;// level 17
assign po0109 = ~w7353;// level 17
assign po0110 = ~w7360;// level 17
assign po0111 = ~w7381;// level 27
assign po0112 = w7397;// level 27
assign po0113 = w7414;// level 26
assign po0114 = ~w7478;// level 19
assign po0115 = ~w7510;// level 19
assign po0116 = ~w7543;// level 20
assign po0117 = ~w7575;// level 19
assign po0118 = ~w7607;// level 19
assign po0119 = ~w7640;// level 20
assign po0120 = ~w7673;// level 20
assign po0121 = ~w7705;// level 19
assign po0122 = ~w7737;// level 19
assign po0123 = ~w7769;// level 19
assign po0124 = ~w7801;// level 19
assign po0125 = ~w7833;// level 19
assign po0126 = ~w7865;// level 19
assign po0127 = ~w7898;// level 20
assign po0128 = ~w8086;// level 19
assign po0129 = ~w8269;// level 17
assign po0130 = w8273;// level 3
assign po0131 = w8276;// level 3
assign po0132 = ~w8279;// level 3
assign po0133 = w8282;// level 3
assign po0134 = w8285;// level 3
assign po0135 = ~w8288;// level 3
assign po0136 = w8291;// level 3
assign po0137 = ~w8294;// level 3
assign po0138 = w8296;// level 3
assign po0139 = w8297;// level 3
assign po0140 = ~w8299;// level 3
assign po0141 = w8300;// level 3
assign po0142 = w8301;// level 3
assign po0143 = ~w8303;// level 3
assign po0144 = w8304;// level 3
assign po0145 = ~w8306;// level 3
assign po0146 = w8312;// level 14
assign po0147 = w8318;// level 14
assign po0148 = w8324;// level 14
assign po0149 = w8330;// level 14
assign po0150 = w8336;// level 14
assign po0151 = w8343;// level 14
assign po0152 = w8349;// level 14
assign po0153 = w8355;// level 14
assign po0154 = w8361;// level 14
assign po0155 = w8367;// level 14
assign po0156 = w8373;// level 14
assign po0157 = w8380;// level 14
assign po0158 = w8386;// level 14
assign po0159 = w8392;// level 14
assign po0160 = w8398;// level 14
assign po0161 = w8404;// level 14
assign po0162 = ~w8418;// level 14
assign po0163 = ~w8426;// level 14
assign po0164 = ~w8434;// level 14
assign po0165 = ~w8442;// level 14
assign po0166 = ~w8450;// level 14
assign po0167 = ~w8459;// level 15
assign po0168 = ~w8467;// level 14
assign po0169 = ~w8475;// level 14
assign po0170 = ~w8483;// level 14
assign po0171 = ~w8491;// level 14
assign po0172 = ~w8499;// level 14
assign po0173 = ~w8508;// level 15
assign po0174 = ~w8516;// level 14
assign po0175 = ~w8524;// level 14
assign po0176 = ~w8532;// level 14
assign po0177 = ~w8540;// level 14
assign po0178 = pi1769;// level 0
assign po0179 = pi1767;// level 0
assign po0180 = pi1766;// level 0
assign po0181 = pi1858;// level 0
assign po0182 = pi1765;// level 0
assign po0183 = pi1764;// level 0
assign po0184 = pi1763;// level 0
assign po0185 = pi1857;// level 0
assign po0186 = pi1762;// level 0
assign po0187 = pi1761;// level 0
assign po0188 = pi1854;// level 0
assign po0189 = pi1768;// level 0
assign po0190 = pi1103;// level 0
assign po0191 = pi1023;// level 0
assign po0192 = pi1101;// level 0
assign po0193 = pi1022;// level 0
assign po0194 = pi1100;// level 0
assign po0195 = pi1021;// level 0
assign po0196 = pi1099;// level 0
assign po0197 = pi1020;// level 0
assign po0198 = pi1019;// level 0
assign po0199 = pi0974;// level 0
assign po0200 = pi1102;// level 0
assign po0201 = pi1024;// level 0
assign po0202 = w8589;// level 28
assign po0203 = ~w8632;// level 25
assign po0204 = w8678;// level 26
assign po0205 = w8729;// level 27
assign po0206 = w8774;// level 26
assign po0207 = ~w8790;// level 25
assign po0208 = w8806;// level 26
assign po0209 = w8822;// level 26
assign po0210 = ~w8839;// level 27
assign po0211 = ~w8855;// level 26
assign po0212 = ~w8871;// level 26
assign po0213 = ~w8888;// level 26
assign po0214 = ~w1323;// level 25
assign po0215 = ~w1657;// level 25
assign po0216 = ~w8919;// level 29
assign po0217 = ~w8945;// level 27
assign po0218 = w8973;// level 27
assign po0219 = ~w9002;// level 27
assign po0220 = w9032;// level 27
assign po0221 = ~w6523;// level 27
assign po0222 = ~w3439;// level 28
assign po0223 = ~w4452;// level 27
assign po0224 = w6596;// level 27
assign po0225 = w4385;// level 27
assign po0226 = ~w5379;// level 27
assign po0227 = ~w5958;// level 26
assign po0228 = ~w4795;// level 27
assign po0229 = ~w3817;// level 27
assign po0230 = ~w9077;// level 22
assign po0231 = ~w9135;// level 22
assign po0232 = ~w9195;// level 22
assign po0233 = ~w9252;// level 22
assign po0234 = ~w9313;// level 22
assign po0235 = ~w9361;// level 22
assign po0236 = ~w9406;// level 22
assign po0237 = ~w9457;// level 22
assign po0238 = ~w9519;// level 22
assign po0239 = ~w9565;// level 22
assign po0240 = ~w9618;// level 22
assign po0241 = ~w9678;// level 22
assign po0242 = ~w7107;// level 22
assign po0243 = ~w7168;// level 22
assign po0244 = w9683;// level 8
assign po0245 = w9688;// level 8
assign po0246 = w9693;// level 8
assign po0247 = w9698;// level 8
assign po0248 = w9703;// level 8
assign po0249 = w9708;// level 8
assign po0250 = w9713;// level 8
assign po0251 = w9718;// level 8
assign po0252 = w9723;// level 8
assign po0253 = w9728;// level 8
assign po0254 = w9733;// level 8
assign po0255 = w9738;// level 8
assign po0256 = w9743;// level 8
assign po0257 = w9748;// level 8
assign po0258 = w9753;// level 8
assign po0259 = w9758;// level 8
assign po0260 = w9763;// level 8
assign po0261 = w9768;// level 8
assign po0262 = w9773;// level 8
assign po0263 = w9778;// level 8
assign po0264 = w9783;// level 8
assign po0265 = w9788;// level 8
assign po0266 = w9793;// level 8
assign po0267 = w9798;// level 8
assign po0268 = w9801;// level 23
assign po0269 = w9804;// level 23
assign po0270 = w9807;// level 23
assign po0271 = w9810;// level 23
assign po0272 = w9813;// level 23
assign po0273 = pi3400;// level 0
assign po0274 = pi3403;// level 0
assign po0275 = pi3402;// level 0
assign po0276 = pi3404;// level 0
assign po0277 = pi3414;// level 0
assign po0278 = ~w9817;// level 9
assign po0279 = ~w9819;// level 9
assign po0280 = ~w9823;// level 3
assign po0281 = ~w9826;// level 4
assign po0282 = ~w9829;// level 4
assign po0283 = ~w9832;// level 4
assign po0284 = ~w9835;// level 4
assign po0285 = ~w9838;// level 4
assign po0286 = ~w9841;// level 4
assign po0287 = ~w9844;// level 4
assign po0288 = ~w9847;// level 4
assign po0289 = ~w9850;// level 4
assign po0290 = ~w9853;// level 9
assign po0291 = w9855;// level 2
assign po0292 = one;// level 0
assign po0293 = ~w9861;// level 19
assign po0294 = ~w9866;// level 18
assign po0295 = ~w9871;// level 18
assign po0296 = ~w9876;// level 18
assign po0297 = ~w9881;// level 18
assign po0298 = ~w9886;// level 18
assign po0299 = ~w9891;// level 19
assign po0300 = ~w9896;// level 19
assign po0301 = ~w9901;// level 19
assign po0302 = ~w9906;// level 18
assign po0303 = ~w9911;// level 18
assign po0304 = ~w9916;// level 18
assign po0305 = ~w9921;// level 18
assign po0306 = ~w9927;// level 19
assign po0307 = ~w9929;// level 10
assign po0308 = w10744;// level 25
assign po0309 = w13876;// level 34
assign po0310 = w13921;// level 34
assign po0311 = w13938;// level 34
assign po0312 = w13944;// level 34
assign po0313 = ~w13949;// level 34
assign po0314 = ~w13952;// level 34
assign po0315 = ~w14035;// level 25
assign po0316 = ~w14065;// level 34
assign po0317 = ~w14074;// level 34
assign po0318 = ~w14078;// level 34
assign po0319 = w14115;// level 34
assign po0320 = w14122;// level 34
assign po0321 = w14295;// level 34
assign po0322 = w14330;// level 34
assign po0323 = w14343;// level 34
assign po0324 = w14349;// level 34
assign po0325 = w14886;// level 24
assign po0326 = w14894;// level 24
assign po0327 = ~w14897;// level 34
assign po0328 = ~w14916;// level 34
assign po0329 = ~w14922;// level 34
assign po0330 = w14927;// level 34
assign po0331 = ~w14930;// level 34
assign po0332 = w14967;// level 34
assign po0333 = w14992;// level 34
assign po0334 = w14998;// level 34
assign po0335 = w15006;// level 34
assign po0336 = w15138;// level 24
assign po0337 = w15143;// level 23
assign po0338 = w15177;// level 34
assign po0339 = ~w15183;// level 34
assign po0340 = w15188;// level 34
assign po0341 = w15192;// level 34
assign po0342 = ~w15397;// level 23
assign po0343 = w15444;// level 23
assign po0344 = w15570;// level 24
assign po0345 = w15672;// level 24
assign po0346 = w15775;// level 24
assign po0347 = w15921;// level 24
assign po0348 = w15926;// level 24
assign po0349 = w15931;// level 24
assign po0350 = w15936;// level 23
assign po0351 = w15942;// level 24
assign po0352 = w15946;// level 34
assign po0353 = ~w15949;// level 34
assign po0354 = ~w15953;// level 34
assign po0355 = w15982;// level 34
assign po0356 = w16110;// level 34
assign po0357 = ~w16116;// level 34
assign po0358 = w16126;// level 34
assign po0359 = ~w16130;// level 34
assign po0360 = w16133;// level 34
assign po0361 = w16139;// level 34
assign po0362 = ~w16143;// level 34
assign po0363 = w16146;// level 34
assign po0364 = w16152;// level 34
assign po0365 = ~w16263;// level 24
assign po0366 = w16352;// level 24
assign po0367 = w16456;// level 24
assign po0368 = ~w16561;// level 24
assign po0369 = w16668;// level 24
assign po0370 = w16766;// level 25
assign po0371 = w16881;// level 24
assign po0372 = w16977;// level 25
assign po0373 = ~w17070;// level 24
assign po0374 = w17196;// level 24
assign po0375 = ~w17202;// level 24
assign po0376 = w17207;// level 23
assign po0377 = ~w17213;// level 24
assign po0378 = w17219;// level 24
assign po0379 = w17225;// level 24
assign po0380 = w17231;// level 25
assign po0381 = w17236;// level 24
assign po0382 = w17243;// level 25
assign po0383 = ~w17249;// level 24
assign po0384 = w17255;// level 23
assign po0385 = w17287;// level 34
assign po0386 = w17311;// level 34
assign po0387 = w17331;// level 34
assign po0388 = w17336;// level 34
assign po0389 = w17342;// level 34
assign po0390 = w17348;// level 34
assign po0391 = w17351;// level 34
assign po0392 = w17354;// level 34
assign po0393 = w17358;// level 34
assign po0394 = w17362;// level 34
assign po0395 = w17365;// level 34
assign po0396 = w17368;// level 34
assign po0397 = w17396;// level 23
assign po0398 = ~w17419;// level 22
assign po0399 = ~w17434;// level 23
assign po0400 = w17465;// level 34
assign po0401 = w17470;// level 34
assign po0402 = w17473;// level 34
assign po0403 = w17476;// level 34
assign po0404 = w17483;// level 23
assign po0405 = ~w17511;// level 34
assign po0406 = w17539;// level 34
assign po0407 = ~w17547;// level 34
assign po0408 = w17553;// level 34
assign po0409 = ~w17557;// level 34
assign po0410 = w17560;// level 34
assign po0411 = ~w17564;// level 34
assign po0412 = w17567;// level 34
assign po0413 = ~w17600;// level 23
assign po0414 = ~w17604;// level 23
assign po0415 = ~w17622;// level 34
assign po0416 = ~w17630;// level 34
assign po0417 = ~w17634;// level 34
assign po0418 = ~w17638;// level 34
assign po0419 = ~w17673;// level 25
assign po0420 = ~w17681;// level 23
assign po0421 = ~w17686;// level 24
assign po0422 = w17690;// level 20
assign po0423 = w17698;// level 24
assign po0424 = w17703;// level 24
assign po0425 = w17708;// level 24
assign po0426 = ~w17716;// level 24
assign po0427 = w17721;// level 24
assign po0428 = w17726;// level 24
assign po0429 = ~w17731;// level 24
assign po0430 = ~w17736;// level 24
assign po0431 = ~w17741;// level 24
assign po0432 = w17746;// level 24
assign po0433 = w17751;// level 24
assign po0434 = w17756;// level 24
assign po0435 = w17762;// level 24
assign po0436 = w17767;// level 24
assign po0437 = w17771;// level 24
assign po0438 = w17774;// level 24
assign po0439 = w17777;// level 24
assign po0440 = ~w17781;// level 24
assign po0441 = w17784;// level 24
assign po0442 = w17787;// level 24
assign po0443 = ~w17790;// level 24
assign po0444 = ~w17795;// level 24
assign po0445 = ~w17798;// level 24
assign po0446 = ~w17801;// level 24
assign po0447 = w17804;// level 24
assign po0448 = w17807;// level 24
assign po0449 = w17810;// level 24
assign po0450 = w17813;// level 24
assign po0451 = w17816;// level 24
assign po0452 = ~w17819;// level 24
assign po0453 = ~w17826;// level 21
assign po0454 = ~w17830;// level 21
assign po0455 = ~w17849;// level 33
assign po0456 = ~w17857;// level 33
assign po0457 = ~w17861;// level 33
assign po0458 = ~w17865;// level 33
assign po0459 = ~w18015;// level 16
assign po0460 = w18031;// level 34
assign po0461 = w18036;// level 34
assign po0462 = w18044;// level 32
assign po0463 = w18051;// level 32
assign po0464 = w18054;// level 34
assign po0465 = w18057;// level 34
assign po0466 = w18061;// level 21
assign po0467 = ~w18065;// level 21
assign po0468 = ~w18068;// level 21
assign po0469 = w18175;// level 22
assign po0470 = ~w18180;// level 22
assign po0471 = ~w18186;// level 21
assign po0472 = ~w18192;// level 21
assign po0473 = w18196;// level 20
assign po0474 = ~w18199;// level 20
assign po0475 = w18205;// level 21
assign po0476 = ~w18208;// level 20
assign po0477 = ~w18211;// level 20
assign po0478 = w18214;// level 20
assign po0479 = w18228;// level 33
assign po0480 = w18234;// level 33
assign po0481 = w18240;// level 32
assign po0482 = w18246;// level 32
assign po0483 = ~w18249;// level 33
assign po0484 = ~w18252;// level 33
assign po0485 = w18271;// level 32
assign po0486 = w18282;// level 33
assign po0487 = w18287;// level 33
assign po0488 = w18294;// level 32
assign po0489 = w18298;// level 32
assign po0490 = w18301;// level 33
assign po0491 = w18305;// level 33
assign po0492 = w18308;// level 33
assign po0493 = w10741;// level 1
assign po0494 = ~w18311;// level 6
assign po0495 = w18364;// level 11
assign po0496 = ~w18378;// level 16
assign po0497 = ~w18390;// level 16
assign po0498 = ~w18394;// level 21
assign po0499 = ~w18397;// level 21
assign po0500 = w18403;// level 31
assign po0501 = w18409;// level 31
assign po0502 = w18418;// level 24
assign po0503 = w18422;// level 24
assign po0504 = ~w18434;// level 17
assign po0505 = ~w18439;// level 21
assign po0506 = ~w18442;// level 21
assign po0507 = w18450;// level 20
assign po0508 = w18454;// level 20
assign po0509 = w18466;// level 18
assign po0510 = ~w18471;// level 22
assign po0511 = ~w18474;// level 22
assign po0512 = w18480;// level 30
assign po0513 = w18486;// level 30
assign po0514 = w18492;// level 24
assign po0515 = w18498;// level 24
assign po0516 = w18501;// level 24
assign po0517 = w18504;// level 24
assign po0518 = ~w18511;// level 12
assign po0519 = w18525;// level 17
assign po0520 = w18533;// level 17
assign po0521 = w18538;// level 20
assign po0522 = w18543;// level 20
assign po0523 = ~w18548;// level 21
assign po0524 = w18551;// level 20
assign po0525 = w18554;// level 20
assign po0526 = ~w18557;// level 21
assign po0527 = w18563;// level 29
assign po0528 = w18569;// level 27
assign po0529 = w18575;// level 29
assign po0530 = w18581;// level 27
assign po0531 = ~w18585;// level 21
assign po0532 = ~w18589;// level 21
assign po0533 = ~w18593;// level 21
assign po0534 = ~w18598;// level 21
assign po0535 = ~w18601;// level 21
assign po0536 = ~w18604;// level 21
assign po0537 = ~w18607;// level 21
assign po0538 = ~w18610;// level 21
assign po0539 = w18616;// level 26
assign po0540 = w18622;// level 26
assign po0541 = ~w18627;// level 21
assign po0542 = ~w18630;// level 21
assign po0543 = ~w18635;// level 21
assign po0544 = ~w18638;// level 21
assign po0545 = w18643;// level 23
assign po0546 = w18648;// level 22
assign po0547 = w18651;// level 23
assign po0548 = w18654;// level 22
assign po0549 = ~w18661;// level 12
assign po0550 = w18670;// level 17
assign po0551 = ~w18674;// level 21
assign po0552 = ~w18677;// level 21
assign po0553 = w18682;// level 21
assign po0554 = w18687;// level 20
assign po0555 = w18690;// level 20
assign po0556 = w18693;// level 20
assign po0557 = ~w18698;// level 22
assign po0558 = ~w18701;// level 22
assign po0559 = w18706;// level 20
assign po0560 = w18711;// level 20
assign po0561 = w18716;// level 19
assign po0562 = w18719;// level 20
assign po0563 = w18722;// level 20
assign po0564 = w18725;// level 19
assign po0565 = w18731;// level 25
assign po0566 = w18737;// level 25
assign po0567 = w18743;// level 22
assign po0568 = w18746;// level 22
assign po0569 = ~w18751;// level 22
assign po0570 = ~w18754;// level 22
assign po0571 = w18759;// level 20
assign po0572 = w18762;// level 19
assign po0573 = w18768;// level 22
assign po0574 = w18771;// level 22
assign po0575 = ~w18778;// level 12
assign po0576 = ~w18783;// level 21
assign po0577 = ~w18788;// level 21
assign po0578 = ~w18791;// level 21
assign po0579 = ~w18794;// level 21
assign po0580 = w18799;// level 21
assign po0581 = w18804;// level 19
assign po0582 = w18807;// level 20
assign po0583 = w18810;// level 19
assign po0584 = w18816;// level 23
assign po0585 = w18822;// level 23
assign po0586 = w18829;// level 18
assign po0587 = ~w18833;// level 21
assign po0588 = ~w18836;// level 21
assign po0589 = w18841;// level 20
assign po0590 = w18846;// level 21
assign po0591 = w18849;// level 20
assign po0592 = w18852;// level 21
assign po0593 = w18858;// level 22
assign po0594 = w18861;// level 22
assign po0595 = w18866;// level 20
assign po0596 = w18869;// level 19
assign po0597 = ~w18875;// level 22
assign po0598 = ~w18878;// level 22
assign po0599 = w18884;// level 22
assign po0600 = w18890;// level 22
assign po0601 = ~w18902;// level 16
assign po0602 = w18907;// level 19
assign po0603 = ~w18916;// level 16
assign po0604 = ~w18934;// level 19
assign po0605 = ~w18938;// level 19
assign po0606 = w18944;// level 20
assign po0607 = w18950;// level 20
assign po0608 = ~w18957;// level 11
assign po0609 = w18962;// level 21
assign po0610 = w18968;// level 21
assign po0611 = w18971;// level 21
assign po0612 = w18974;// level 21
assign po0613 = ~w18977;// level 11
assign po0614 = w18981;// level 11
assign po0615 = ~w18983;// level 11
assign po0616 = ~w18987;// level 11
assign po0617 = w18993;// level 18
assign po0618 = w18999;// level 18
assign po0619 = ~w19004;// level 20
assign po0620 = w19010;// level 20
assign po0621 = ~w19013;// level 20
assign po0622 = w19016;// level 20
assign po0623 = ~w19032;// level 15
assign po0624 = ~w19101;// level 16
assign po0625 = ~w19126;// level 16
assign po0626 = ~w19151;// level 16
assign po0627 = w19177;// level 15
assign po0628 = ~w19203;// level 17
assign po0629 = ~w19228;// level 16
assign po0630 = ~w19253;// level 16
assign po0631 = w19281;// level 16
assign po0632 = w19309;// level 18
assign po0633 = ~w19336;// level 16
assign po0634 = w19363;// level 16
assign po0635 = ~w19390;// level 17
assign po0636 = ~w19418;// level 19
assign po0637 = ~w19445;// level 17
assign po0638 = ~w19472;// level 17
assign po0639 = ~w19499;// level 17
assign po0640 = ~w19507;// level 11
assign po0641 = w19513;// level 17
assign po0642 = ~w19531;// level 14
assign po0643 = w19547;// level 16
assign po0644 = ~w19555;// level 14
assign po0645 = ~w19563;// level 14
assign po0646 = ~w19571;// level 14
assign po0647 = ~w19579;// level 13
assign po0648 = ~w19587;// level 13
assign po0649 = ~w19598;// level 15
assign po0650 = ~w19608;// level 15
assign po0651 = ~w19618;// level 16
assign po0652 = ~w19626;// level 14
assign po0653 = ~w19634;// level 14
assign po0654 = ~w19644;// level 16
assign po0655 = ~w19654;// level 16
assign po0656 = ~w19664;// level 16
assign po0657 = ~w19691;// level 16
assign po0658 = ~w19718;// level 16
assign po0659 = ~w19745;// level 16
assign po0660 = ~w19772;// level 16
assign po0661 = ~w19799;// level 16
assign po0662 = ~w19826;// level 16
assign po0663 = ~w19853;// level 16
assign po0664 = ~w19863;// level 16
assign po0665 = ~w19873;// level 16
assign po0666 = ~w19900;// level 16
assign po0667 = ~w19906;// level 19
assign po0668 = ~w19909;// level 19
assign po0669 = w19916;// level 19
assign po0670 = w19923;// level 19
assign po0671 = ~w19931;// level 11
assign po0672 = ~w19937;// level 18
assign po0673 = ~w19940;// level 18
assign po0674 = w19946;// level 20
assign po0675 = w19949;// level 20
assign po0676 = pi3561;// level 0
assign po0677 = ~w19963;// level 14
assign po0678 = w20529;// level 21
assign po0679 = ~w20535;// level 13
assign po0680 = ~w20541;// level 13
assign po0681 = ~w20547;// level 14
assign po0682 = ~w20553;// level 14
assign po0683 = ~w20559;// level 14
assign po0684 = ~w20565;// level 14
assign po0685 = ~w20571;// level 14
assign po0686 = ~w20577;// level 14
assign po0687 = ~w20583;// level 14
assign po0688 = ~w20589;// level 14
assign po0689 = ~w20595;// level 14
assign po0690 = ~w20601;// level 14
assign po0691 = ~w20607;// level 14
assign po0692 = ~w20613;// level 14
assign po0693 = ~w20619;// level 14
assign po0694 = ~w20625;// level 14
assign po0695 = ~w20631;// level 13
assign po0696 = ~w20637;// level 13
assign po0697 = ~w20643;// level 13
assign po0698 = ~w20649;// level 13
assign po0699 = ~w20655;// level 13
assign po0700 = ~w20661;// level 14
assign po0701 = ~w20667;// level 14
assign po0702 = w20679;// level 13
assign po0703 = w20685;// level 13
assign po0704 = w20691;// level 13
assign po0705 = w20697;// level 13
assign po0706 = w20702;// level 13
assign po0707 = w20707;// level 13
assign po0708 = w20713;// level 13
assign po0709 = w20719;// level 13
assign po0710 = w20725;// level 18
assign po0711 = w20728;// level 18
assign po0712 = w20737;// level 17
assign po0713 = w20745;// level 17
assign po0714 = w20751;// level 17
assign po0715 = w20757;// level 17
assign po0716 = w20763;// level 17
assign po0717 = w20769;// level 17
assign po0718 = w20775;// level 17
assign po0719 = w20781;// level 14
assign po0720 = w20787;// level 14
assign po0721 = w20793;// level 14
assign po0722 = w20799;// level 14
assign po0723 = w20805;// level 17
assign po0724 = w20811;// level 14
assign po0725 = w20817;// level 14
assign po0726 = w20823;// level 13
assign po0727 = w20831;// level 16
assign po0728 = w20839;// level 16
assign po0729 = w20847;// level 17
assign po0730 = w20855;// level 17
assign po0731 = w20863;// level 17
assign po0732 = ~w20871;// level 11
assign po0733 = w20877;// level 17
assign po0734 = w20883;// level 17
assign po0735 = w20891;// level 17
assign po0736 = w20897;// level 13
assign po0737 = w20903;// level 18
assign po0738 = w20906;// level 18
assign po0739 = w20912;// level 4
assign po0740 = ~w20944;// level 15
assign po0741 = ~w20949;// level 15
assign po0742 = ~w20954;// level 15
assign po0743 = ~w20959;// level 15
assign po0744 = ~w20964;// level 15
assign po0745 = ~w20969;// level 15
assign po0746 = ~w20974;// level 15
assign po0747 = ~w20979;// level 15
assign po0748 = ~w20984;// level 15
assign po0749 = ~w20989;// level 15
assign po0750 = ~w20994;// level 15
assign po0751 = ~w20999;// level 15
assign po0752 = ~w21004;// level 15
assign po0753 = ~w21009;// level 15
assign po0754 = ~w21019;// level 18
assign po0755 = ~w21025;// level 19
assign po0756 = ~w21028;// level 19
assign po0757 = ~pi3589;// level 0
assign po0758 = ~w21298;// level 23
assign po0759 = ~w21305;// level 19
assign po0760 = ~w21310;// level 18
assign po0761 = ~w21315;// level 18
assign po0762 = ~w21318;// level 19
assign po0763 = ~w21321;// level 18
assign po0764 = ~w21324;// level 18
assign po0765 = w21331;// level 18
assign po0766 = w21338;// level 18
assign po0767 = w0;// level 1
assign po0768 = ~w21343;// level 3
assign po0769 = pi3647;// level 0
assign po0770 = ~w20912;// level 4
assign po0771 = w21372;// level 16
assign po0772 = ~w21378;// level 17
assign po0773 = ~w21384;// level 19
assign po0774 = ~w21387;// level 19
assign po0775 = ~w21395;// level 11
assign po0776 = ~w21401;// level 17
assign po0777 = ~w21405;// level 17
assign po0778 = pi3635;// level 0
assign po0779 = ~w21411;// level 4
assign po0780 = w21459;// level 16
assign po0781 = ~w21465;// level 17
assign po0782 = ~w21471;// level 17
assign po0783 = ~w21477;// level 17
assign po0784 = ~w21481;// level 17
assign po0785 = ~w21487;// level 17
assign po0786 = pi3584;// level 0
assign po0787 = w21554;// level 17
assign po0788 = w21567;// level 17
assign po0789 = w21580;// level 17
assign po0790 = w21592;// level 17
assign po0791 = w21605;// level 17
assign po0792 = w21617;// level 17
assign po0793 = pi3558;// level 0
assign po0794 = w21657;// level 17
assign po0795 = w21669;// level 17
assign po0796 = w21681;// level 17
assign po0797 = w21693;// level 17
assign po0798 = w21705;// level 17
assign po0799 = w21718;// level 17
assign po0800 = w21731;// level 17
assign po0801 = w21744;// level 17
assign po0802 = w21756;// level 17
assign po0803 = w21768;// level 17
assign po0804 = w21781;// level 17
assign po0805 = w21790;// level 7
assign po0806 = pi3483;// level 0
assign po0807 = ~w21849;// level 16
assign po0808 = ~w21853;// level 16
assign po0809 = w21858;// level 15
assign po0810 = w21863;// level 15
assign po0811 = w21868;// level 15
assign po0812 = w21875;// level 15
assign po0813 = w21877;// level 15
assign po0814 = w21884;// level 15
assign po0815 = w21886;// level 15
assign po0816 = w21889;// level 15
assign po0817 = w21902;// level 17
assign po0818 = w21914;// level 17
assign po0819 = w21927;// level 17
assign po0820 = w21939;// level 17
assign po0821 = ~w21957;// level 15
assign po0822 = ~w21960;// level 15
assign po0823 = ~w21967;// level 11
assign po0824 = ~w22018;// level 21
assign po0825 = ~w22028;// level 12
assign po0826 = ~w22030;// level 15
assign po0827 = w21362;// level 12
assign po0828 = w22038;// level 7
assign po0829 = w22066;// level 14
assign po0830 = w22075;// level 8
assign po0831 = ~w22086;// level 16
assign po0832 = w22090;// level 16
assign po0833 = w22095;// level 15
assign po0834 = w22100;// level 15
assign po0835 = w22105;// level 15
assign po0836 = w22110;// level 15
assign po0837 = w22115;// level 15
assign po0838 = ~w22117;// level 15
assign po0839 = ~w22128;// level 16
assign po0840 = w22132;// level 16
assign po0841 = w22137;// level 15
assign po0842 = w22142;// level 15
assign po0843 = w22147;// level 15
assign po0844 = w22152;// level 15
assign po0845 = ~w22156;// level 16
assign po0846 = w21434;// level 12
assign po0847 = w22161;// level 15
assign po0848 = w22166;// level 15
assign po0849 = ~w22167;// level 1
assign po0850 = ~w22168;// level 1
assign po0851 = ~w22232;// level 32
assign po0852 = w22244;// level 17
assign po0853 = w22257;// level 17
assign po0854 = w22269;// level 17
assign po0855 = w22282;// level 17
assign po0856 = w22292;// level 8
assign po0857 = ~w22295;// level 19
assign po0858 = ~w22298;// level 19
assign po0859 = ~w22301;// level 19
assign po0860 = ~w22311;// level 16
assign po0861 = ~w22339;// level 14
assign po0862 = ~w22342;// level 16
assign po0863 = ~w22350;// level 10
assign po0864 = ~w22353;// level 19
assign po0865 = ~w22361;// level 14
assign po0866 = ~w22370;// level 14
assign po0867 = pi0635;// level 0
assign po0868 = pi0633;// level 0
assign po0869 = w22377;// level 19
assign po0870 = w22384;// level 19
assign po0871 = ~w22386;// level 19
assign po0872 = w22416;// level 17
assign po0873 = w22428;// level 17
assign po0874 = w22440;// level 17
assign po0875 = w22454;// level 17
assign po0876 = ~w22457;// level 19
assign po0877 = ~w22460;// level 19
assign po0878 = ~w22463;// level 19
assign po0879 = ~w22466;// level 19
assign po0880 = ~w22469;// level 19
assign po0881 = ~w22472;// level 19
assign po0882 = ~w22479;// level 14
assign po0883 = ~w22484;// level 14
assign po0884 = ~w22491;// level 14
assign po0885 = ~w22494;// level 14
assign po0886 = ~pi3639;// level 0
assign po0887 = ~w22584;// level 18
assign po0888 = ~pi3638;// level 0
assign po0889 = ~w22674;// level 19
assign po0890 = ~w22677;// level 19
assign po0891 = ~w22680;// level 19
assign po0892 = ~w22683;// level 13
assign po0893 = ~w22690;// level 18
assign po0894 = ~w22697;// level 19
assign po0895 = ~w22704;// level 18
assign po0896 = w21411;// level 4
assign po0897 = w22714;// level 14
assign po0898 = pi3479;// level 0
assign po0899 = w22919;// level 32
assign po0900 = w22924;// level 14
assign po0901 = w22929;// level 14
assign po0902 = w22971;// level 17
assign po0903 = w22986;// level 17
assign po0904 = w23001;// level 17
assign po0905 = ~w23010;// level 15
assign po0906 = w23019;// level 17
assign po0907 = ~w23024;// level 17
assign po0908 = ~w23029;// level 18
assign po0909 = w23042;// level 9
assign po0910 = w23047;// level 9
assign po0911 = w23052;// level 14
assign po0912 = w23057;// level 14
assign po0913 = w23062;// level 14
assign po0914 = w23067;// level 14
assign po0915 = w23072;// level 14
assign po0916 = w23077;// level 14
assign po0917 = w23082;// level 14
assign po0918 = w23087;// level 14
assign po0919 = w23092;// level 14
assign po0920 = w23097;// level 14
assign po0921 = w23102;// level 14
assign po0922 = ~w23105;// level 19
assign po0923 = w23106;// level 15
assign po0924 = w23122;// level 17
assign po0925 = w23123;// level 15
assign po0926 = w23139;// level 17
assign po0927 = w23154;// level 17
assign po0928 = w23169;// level 17
assign po0929 = w23184;// level 17
assign po0930 = w23199;// level 17
assign po0931 = w23214;// level 17
assign po0932 = w23235;// level 27
assign po0933 = w23248;// level 29
assign po0934 = w23287;// level 17
assign po0935 = w23302;// level 17
assign po0936 = w23317;// level 17
assign po0937 = w23324;// level 18
assign po0938 = w23331;// level 7
assign po0939 = ~w23337;// level 14
assign po0940 = w23352;// level 14
assign po0941 = ~w23357;// level 14
assign po0942 = ~w23362;// level 15
assign po0943 = ~w23370;// level 10
assign po0944 = w21363;// level 13
assign po0945 = w21449;// level 13
assign po0946 = w23385;// level 17
assign po0947 = w23399;// level 17
assign po0948 = w23415;// level 17
assign po0949 = w23416;// level 16
assign po0950 = w23433;// level 29
assign po0951 = w23450;// level 28
assign po0952 = w23464;// level 27
assign po0953 = w23478;// level 28
assign po0954 = w23492;// level 27
assign po0955 = w23509;// level 28
assign po0956 = w23523;// level 29
assign po0957 = w23536;// level 29
assign po0958 = w23551;// level 17
assign po0959 = w23566;// level 17
assign po0960 = w23581;// level 17
assign po0961 = w23596;// level 17
assign po0962 = w23611;// level 17
assign po0963 = w23626;// level 17
assign po0964 = w23641;// level 17
assign po0965 = w23656;// level 17
assign po0966 = w23671;// level 17
assign po0967 = w23694;// level 29
assign po0968 = w23710;// level 29
assign po0969 = w23727;// level 29
assign po0970 = w23744;// level 29
assign po0971 = w23759;// level 29
assign po0972 = w23775;// level 29
assign po0973 = w23791;// level 29
assign po0974 = pi3482;// level 0
assign po0975 = ~w23828;// level 19
assign po0976 = w23832;// level 16
assign po0977 = w23837;// level 15
assign po0978 = pi3525;// level 0
assign po0979 = ~w23860;// level 25
assign po0980 = pi3562;// level 0
assign po0981 = ~w23881;// level 23
assign po0982 = ~w23886;// level 13
assign po0983 = ~w23891;// level 14
assign po0984 = w23896;// level 8
assign po0985 = w23899;// level 32
assign po0986 = w23905;// level 14
assign po0987 = w23908;// level 14
assign po0988 = ~w23913;// level 14
assign po0989 = w23919;// level 14
assign po0990 = ~w23921;// level 14
assign po0991 = ~w23926;// level 16
assign po0992 = ~w23934;// level 9
assign po0993 = w21452;// level 14
assign po0994 = w23950;// level 29
assign po0995 = w23967;// level 29
assign po0996 = w23984;// level 29
assign po0997 = w24000;// level 29
assign po0998 = w24016;// level 28
assign po0999 = w24033;// level 29
assign po1000 = w24048;// level 28
assign po1001 = ~w24083;// level 17
assign po1002 = ~w24086;// level 14
assign po1003 = ~w24090;// level 14
assign po1004 = ~w24093;// level 14
assign po1005 = ~w24096;// level 14
assign po1006 = ~w24099;// level 14
assign po1007 = ~w24102;// level 14
assign po1008 = ~w24105;// level 14
assign po1009 = ~w24112;// level 14
assign po1010 = ~w24117;// level 14
assign po1011 = ~w24120;// level 14
assign po1012 = ~w24124;// level 14
assign po1013 = ~w24127;// level 14
assign po1014 = ~w24130;// level 15
assign po1015 = ~w24134;// level 11
assign po1016 = w24139;// level 21
assign po1017 = w24144;// level 24
assign po1018 = w24149;// level 23
assign po1019 = w24154;// level 22
assign po1020 = ~w24159;// level 15
assign po1021 = ~w24167;// level 9
assign po1022 = w21366;// level 14
assign po1023 = pi3676;// level 0
assign po1024 = ~w24230;// level 10
assign po1025 = ~w24270;// level 10
assign po1026 = w24275;// level 20
assign po1027 = w24280;// level 16
assign po1028 = ~w24290;// level 13
assign po1029 = w24305;// level 17
assign po1030 = w24320;// level 17
assign po1031 = w24329;// level 17
assign po1032 = w24339;// level 18
assign po1033 = w24345;// level 18
assign po1034 = w24348;// level 18
assign po1035 = w24352;// level 18
assign po1036 = w24355;// level 17
assign po1037 = w24358;// level 17
assign po1038 = w24361;// level 17
assign po1039 = w24364;// level 17
assign po1040 = w24367;// level 17
assign po1041 = ~w24370;// level 17
assign po1042 = ~w24373;// level 17
assign po1043 = ~w24381;// level 16
assign po1044 = w24388;// level 19
assign po1045 = w24395;// level 19
assign po1046 = ~w24413;// level 25
assign po1047 = w24428;// level 17
assign po1048 = w24441;// level 28
assign po1049 = w24458;// level 29
assign po1050 = w24475;// level 29
assign po1051 = w24492;// level 29
assign po1052 = ~w24496;// level 13
assign po1053 = ~w24500;// level 19
assign po1054 = ~w24508;// level 13
assign po1055 = ~w24511;// level 14
assign po1056 = ~w24515;// level 11
assign po1057 = ~w24519;// level 14
assign po1058 = ~w24523;// level 14
assign po1059 = ~w24527;// level 14
assign po1060 = ~w24530;// level 14
assign po1061 = ~w24533;// level 14
assign po1062 = ~w24536;// level 14
assign po1063 = w24541;// level 19
assign po1064 = w24546;// level 18
assign po1065 = ~w24548;// level 2
assign po1066 = ~w24549;// level 2
assign po1067 = w24554;// level 17
assign po1068 = w24559;// level 16
assign po1069 = ~w24564;// level 18
assign po1070 = ~w24569;// level 17
assign po1071 = ~w24574;// level 16
assign po1072 = ~w24579;// level 16
assign po1073 = ~w24584;// level 16
assign po1074 = ~w24589;// level 16
assign po1075 = ~w24594;// level 24
assign po1076 = ~w24599;// level 23
assign po1077 = ~w24604;// level 22
assign po1078 = w24609;// level 16
assign po1079 = ~w22057;// level 10
assign po1080 = w24610;// level 12
assign po1081 = ~w24647;// level 10
assign po1082 = w24652;// level 16
assign po1083 = w24656;// level 16
assign po1084 = ~w24663;// level 9
assign po1085 = w22681;// level 12
assign po1086 = w24666;// level 18
assign po1087 = w24669;// level 18
assign po1088 = w24679;// level 17
assign po1089 = w24686;// level 17
assign po1090 = w24689;// level 17
assign po1091 = w24693;// level 17
assign po1092 = w24696;// level 15
assign po1093 = w24699;// level 16
assign po1094 = w24702;// level 16
assign po1095 = w24705;// level 16
assign po1096 = w24710;// level 17
assign po1097 = w24713;// level 17
assign po1098 = w24716;// level 17
assign po1099 = w24719;// level 17
assign po1100 = w24722;// level 17
assign po1101 = w24725;// level 17
assign po1102 = ~w24731;// level 9
assign po1103 = ~w24737;// level 9
assign po1104 = ~w24743;// level 9
assign po1105 = ~w24749;// level 9
assign po1106 = ~w24755;// level 9
assign po1107 = ~w24761;// level 9
assign po1108 = ~w24767;// level 9
assign po1109 = ~w24773;// level 9
assign po1110 = ~w24779;// level 9
assign po1111 = ~w24785;// level 9
assign po1112 = ~w24791;// level 9
assign po1113 = ~w24797;// level 9
assign po1114 = ~w24803;// level 9
assign po1115 = ~pi3556;// level 0
assign po1116 = ~w24844;// level 23
assign po1117 = ~w24852;// level 22
assign po1118 = w24884;// level 9
assign po1119 = ~w24892;// level 10
assign po1120 = ~w24927;// level 10
assign po1121 = w24960;// level 9
assign po1122 = ~w24997;// level 10
assign po1123 = ~pi3587;// level 0
assign po1124 = w25027;// level 17
assign po1125 = w25053;// level 17
assign po1126 = w25079;// level 17
assign po1127 = w25105;// level 17
assign po1128 = w25131;// level 17
assign po1129 = ~w25136;// level 13
assign po1130 = ~w25140;// level 20
assign po1131 = ~w25143;// level 20
assign po1132 = ~w25148;// level 20
assign po1133 = ~w25151;// level 13
assign po1134 = ~w25154;// level 14
assign po1135 = ~w25157;// level 14
assign po1136 = ~w25160;// level 15
assign po1137 = ~w25172;// level 10
assign po1138 = ~w25175;// level 10
assign po1139 = ~w25178;// level 10
assign po1140 = ~w25181;// level 10
assign po1141 = ~w25184;// level 10
assign po1142 = ~w25187;// level 10
assign po1143 = ~w25192;// level 21
assign po1144 = w25195;// level 17
assign po1145 = ~w25200;// level 11
assign po1146 = ~w25205;// level 12
assign po1147 = ~w25213;// level 9
assign po1148 = w25216;// level 17
assign po1149 = w25248;// level 9
assign po1150 = w25279;// level 9
assign po1151 = w25319;// level 9
assign po1152 = w25356;// level 9
assign po1153 = ~w25394;// level 10
assign po1154 = ~w25431;// level 10
assign po1155 = ~w25464;// level 10
assign po1156 = w25498;// level 9
assign po1157 = w25531;// level 9
assign po1158 = ~w25562;// level 10
assign po1159 = ~w25567;// level 19
assign po1160 = ~w25572;// level 20
assign po1161 = ~w25580;// level 10
assign po1162 = ~w25583;// level 10
assign po1163 = ~w25586;// level 10
assign po1164 = ~w25591;// level 20
assign po1165 = ~w25594;// level 13
assign po1166 = ~w25620;// level 17
assign po1167 = ~w25623;// level 17
assign po1168 = ~w25627;// level 17
assign po1169 = ~w25630;// level 17
assign po1170 = ~w25633;// level 17
assign po1171 = ~w25641;// level 18
assign po1172 = ~w25649;// level 18
assign po1173 = w25655;// level 25
assign po1174 = ~w25663;// level 18
assign po1175 = w25664;// level 25
assign po1176 = w25665;// level 25
assign po1177 = w25666;// level 25
assign po1178 = ~w25669;// level 18
assign po1179 = ~w25672;// level 18
assign po1180 = ~w25675;// level 18
assign po1181 = ~w25678;// level 18
assign po1182 = ~w25681;// level 18
assign po1183 = ~w25684;// level 18
assign po1184 = ~w25688;// level 18
assign po1185 = ~w25691;// level 18
assign po1186 = ~w25694;// level 18
assign po1187 = ~w25698;// level 18
assign po1188 = w25701;// level 16
assign po1189 = w25704;// level 17
assign po1190 = w25707;// level 17
assign po1191 = w25710;// level 17
assign po1192 = ~w25713;// level 17
assign po1193 = ~w25716;// level 17
assign po1194 = ~w25719;// level 17
assign po1195 = ~w25722;// level 17
assign po1196 = w25804;// level 17
assign po1197 = w25807;// level 17
assign po1198 = ~w25810;// level 16
assign po1199 = w25892;// level 17
assign po1200 = ~w25900;// level 20
assign po1201 = ~w25908;// level 19
assign po1202 = ~w25916;// level 18
assign po1203 = ~w25924;// level 18
assign po1204 = ~w25932;// level 18
assign po1205 = ~w25940;// level 18
assign po1206 = ~w25948;// level 18
assign po1207 = ~w25957;// level 24
assign po1208 = ~w25965;// level 21
assign po1209 = ~w25978;// level 8
assign po1210 = w26010;// level 17
assign po1211 = ~w26033;// level 17
assign po1212 = ~w26055;// level 17
assign po1213 = ~w26077;// level 17
assign po1214 = ~w26104;// level 17
assign po1215 = w26126;// level 17
assign po1216 = ~w26149;// level 17
assign po1217 = ~w26175;// level 18
assign po1218 = ~w26180;// level 12
assign po1219 = ~w26183;// level 20
assign po1220 = w26195;// level 11
assign po1221 = ~w26204;// level 11
assign po1222 = ~w26213;// level 11
assign po1223 = ~w26222;// level 11
assign po1224 = w26231;// level 11
assign po1225 = ~w26240;// level 11
assign po1226 = ~w26245;// level 19
assign po1227 = ~w26251;// level 24
assign po1228 = ~w26256;// level 22
assign po1229 = ~w26261;// level 11
assign po1230 = ~w26266;// level 11
assign po1231 = ~w26271;// level 11
assign po1232 = ~w26276;// level 11
assign po1233 = ~w26281;// level 11
assign po1234 = w26282;// level 2
assign po1235 = w7;// level 3
assign po1236 = w26308;// level 8
assign po1237 = ~w26329;// level 10
assign po1238 = w26364;// level 9
assign po1239 = w26366;// level 4
assign po1240 = w26375;// level 14
assign po1241 = ~w26380;// level 11
assign po1242 = w26383;// level 17
assign po1243 = ~w26392;// level 11
assign po1244 = ~w26401;// level 11
assign po1245 = ~w26406;// level 13
assign po1246 = ~w26410;// level 13
assign po1247 = w26413;// level 16
assign po1248 = ~w26416;// level 16
assign po1249 = ~w26419;// level 17
assign po1250 = ~w26422;// level 17
assign po1251 = ~w26425;// level 17
assign po1252 = ~w26428;// level 17
assign po1253 = ~w26431;// level 17
assign po1254 = ~w26434;// level 17
assign po1255 = ~w26437;// level 17
assign po1256 = ~w26440;// level 17
assign po1257 = ~w26443;// level 17
assign po1258 = ~w26446;// level 17
assign po1259 = ~w26449;// level 17
assign po1260 = ~w26452;// level 17
assign po1261 = ~w26455;// level 17
assign po1262 = ~w26458;// level 17
assign po1263 = ~w26461;// level 16
assign po1264 = ~w26464;// level 16
assign po1265 = ~w26467;// level 16
assign po1266 = ~w26470;// level 16
assign po1267 = ~w26473;// level 16
assign po1268 = ~w26476;// level 16
assign po1269 = ~w26479;// level 17
assign po1270 = ~w26482;// level 17
assign po1271 = ~w26485;// level 17
assign po1272 = ~w26488;// level 17
assign po1273 = ~w26491;// level 17
assign po1274 = w26494;// level 16
assign po1275 = w26504;// level 17
assign po1276 = ~w26510;// level 13
assign po1277 = ~w26531;// level 15
assign po1278 = ~w26534;// level 17
assign po1279 = ~w26537;// level 17
assign po1280 = pi0979;// level 0
assign po1281 = ~w25000;// level 12
assign po1282 = w26560;// level 16
assign po1283 = w26584;// level 17
assign po1284 = ~w26587;// level 17
assign po1285 = ~w26590;// level 13
assign po1286 = ~w26601;// level 13
assign po1287 = ~w26604;// level 13
assign po1288 = ~w26607;// level 13
assign po1289 = ~w26610;// level 13
assign po1290 = ~w26615;// level 12
assign po1291 = ~w26618;// level 12
assign po1292 = ~w26622;// level 12
assign po1293 = ~w26625;// level 13
assign po1294 = ~w26628;// level 13
assign po1295 = ~w26632;// level 13
assign po1296 = ~w26635;// level 13
assign po1297 = ~w26638;// level 13
assign po1298 = ~w26641;// level 13
assign po1299 = ~w26644;// level 13
assign po1300 = ~w26647;// level 13
assign po1301 = ~w26650;// level 12
assign po1302 = ~w26653;// level 13
assign po1303 = ~w26657;// level 13
assign po1304 = ~w26686;// level 10
assign po1305 = ~w26716;// level 10
assign po1306 = w26717;// level 2
assign po1307 = ~w26718;// level 6
assign po1308 = w26760;// level 23
assign po1309 = w26781;// level 26
assign po1310 = w26787;// level 30
assign po1311 = w26801;// level 9
assign po1312 = ~w26804;// level 20
assign po1313 = ~w26807;// level 13
assign po1314 = ~w26810;// level 17
assign po1315 = ~w26813;// level 12
assign po1316 = ~w26816;// level 13
assign po1317 = ~w26838;// level 29
assign po1318 = ~w26841;// level 29
assign po1319 = w26849;// level 16
assign po1320 = w26855;// level 15
assign po1321 = w26858;// level 12
assign po1322 = ~w26861;// level 17
assign po1323 = w26864;// level 12
assign po1324 = w26870;// level 17
assign po1325 = w26879;// level 17
assign po1326 = w26888;// level 17
assign po1327 = w26897;// level 17
assign po1328 = w26906;// level 17
assign po1329 = w26915;// level 17
assign po1330 = w26937;// level 17
assign po1331 = ~w26942;// level 11
assign po1332 = ~w26947;// level 11
assign po1333 = ~w26950;// level 31
assign po1334 = ~w26953;// level 30
assign po1335 = ~w26957;// level 28
assign po1336 = ~w26960;// level 28
assign po1337 = ~w26981;// level 29
assign po1338 = ~w27001;// level 29
assign po1339 = ~w27023;// level 29
assign po1340 = ~w27026;// level 29
assign po1341 = ~w27029;// level 30
assign po1342 = ~w27032;// level 29
assign po1343 = ~w27035;// level 30
assign po1344 = w27056;// level 30
assign po1345 = ~w27061;// level 11
assign po1346 = w27071;// level 16
assign po1347 = ~w27080;// level 15
assign po1348 = ~w27093;// level 17
assign po1349 = ~w27099;// level 17
assign po1350 = ~w27115;// level 10
assign po1351 = w27118;// level 14
assign po1352 = ~w27121;// level 14
assign po1353 = ~w27125;// level 12
assign po1354 = ~w27130;// level 13
assign po1355 = ~w27133;// level 13
assign po1356 = ~w27137;// level 12
assign po1357 = ~w27152;// level 9
assign po1358 = ~w27157;// level 13
assign po1359 = ~w27161;// level 12
assign po1360 = ~w27165;// level 13
assign po1361 = ~w27168;// level 13
assign po1362 = ~w27171;// level 13
assign po1363 = ~w27175;// level 11
assign po1364 = ~w27178;// level 13
assign po1365 = ~w27184;// level 9
assign po1366 = ~w27187;// level 9
assign po1367 = ~w27190;// level 9
assign po1368 = ~w27193;// level 9
assign po1369 = ~w27196;// level 9
assign po1370 = ~w27199;// level 9
assign po1371 = ~w27204;// level 20
assign po1372 = ~w27209;// level 11
assign po1373 = ~w27214;// level 11
assign po1374 = ~w27220;// level 11
assign po1375 = ~w27225;// level 17
assign po1376 = ~w27230;// level 11
assign po1377 = ~w27235;// level 11
assign po1378 = ~w27240;// level 9
assign po1379 = ~w27243;// level 10
assign po1380 = w27245;// level 10
assign po1381 = w27247;// level 28
assign po1382 = w27249;// level 29
assign po1383 = w27253;// level 32
assign po1384 = w27255;// level 15
assign po1385 = ~w27269;// level 9
assign po1386 = w27270;// level 3
assign po1387 = w27284;// level 13
assign po1388 = ~w27298;// level 10
assign po1389 = ~w27303;// level 11
assign po1390 = w27306;// level 33
assign po1391 = ~w27311;// level 12
assign po1392 = w27313;// level 31
assign po1393 = ~w27318;// level 16
assign po1394 = ~w27323;// level 11
assign po1395 = ~w27326;// level 9
assign po1396 = ~w27331;// level 21
assign po1397 = ~w27336;// level 13
assign po1398 = ~w27339;// level 9
assign po1399 = ~w27346;// level 15
assign po1400 = w27349;// level 13
assign po1401 = w27352;// level 13
assign po1402 = pi1641;// level 0
assign po1403 = w27355;// level 14
assign po1404 = w27358;// level 14
assign po1405 = w27364;// level 17
assign po1406 = w27370;// level 17
assign po1407 = w27376;// level 17
assign po1408 = w27382;// level 17
assign po1409 = w27388;// level 17
assign po1410 = ~w27436;// level 16
assign po1411 = w27438;// level 17
assign po1412 = ~w27450;// level 19
assign po1413 = ~w27459;// level 19
assign po1414 = ~w27468;// level 19
assign po1415 = ~w27477;// level 19
assign po1416 = ~w27486;// level 19
assign po1417 = ~w27495;// level 19
assign po1418 = ~w27504;// level 19
assign po1419 = ~w27513;// level 19
assign po1420 = ~w27522;// level 19
assign po1421 = ~w27533;// level 19
assign po1422 = ~w27542;// level 19
assign po1423 = ~w27551;// level 19
assign po1424 = ~w27558;// level 19
assign po1425 = ~w27565;// level 19
assign po1426 = ~w27569;// level 19
assign po1427 = ~w27572;// level 19
assign po1428 = ~w27575;// level 19
assign po1429 = ~w27578;// level 19
assign po1430 = ~w27581;// level 19
assign po1431 = ~w27584;// level 19
assign po1432 = ~w27587;// level 19
assign po1433 = ~w27590;// level 19
assign po1434 = ~w27593;// level 19
assign po1435 = ~w27596;// level 19
assign po1436 = ~w27599;// level 19
assign po1437 = ~w27602;// level 19
assign po1438 = ~w27605;// level 19
assign po1439 = ~w27608;// level 19
assign po1440 = ~w27612;// level 19
assign po1441 = ~w27615;// level 19
assign po1442 = ~w27618;// level 19
assign po1443 = ~w27621;// level 19
assign po1444 = ~w27624;// level 19
assign po1445 = ~w27627;// level 19
assign po1446 = ~w27630;// level 19
assign po1447 = ~w27633;// level 19
assign po1448 = ~w27636;// level 19
assign po1449 = ~w27639;// level 19
assign po1450 = ~w27642;// level 19
assign po1451 = ~w27645;// level 19
assign po1452 = ~w27648;// level 19
assign po1453 = ~w27651;// level 19
assign po1454 = ~w27655;// level 19
assign po1455 = ~w27658;// level 19
assign po1456 = ~w27661;// level 19
assign po1457 = ~w27664;// level 19
assign po1458 = ~w27667;// level 19
assign po1459 = ~w27670;// level 19
assign po1460 = ~w27673;// level 19
assign po1461 = ~w27676;// level 19
assign po1462 = ~w27679;// level 19
assign po1463 = ~w27682;// level 19
assign po1464 = ~w27685;// level 19
assign po1465 = ~w27688;// level 19
assign po1466 = ~w27691;// level 19
assign po1467 = ~w27694;// level 19
assign po1468 = ~w27698;// level 19
assign po1469 = ~w27701;// level 19
assign po1470 = ~w27704;// level 19
assign po1471 = ~w27707;// level 19
assign po1472 = ~w27710;// level 19
assign po1473 = ~w27713;// level 19
assign po1474 = ~w27716;// level 19
assign po1475 = ~w27719;// level 19
assign po1476 = ~w27722;// level 19
assign po1477 = ~w27725;// level 19
assign po1478 = ~w27728;// level 19
assign po1479 = ~w27731;// level 19
assign po1480 = ~w27734;// level 19
assign po1481 = ~w27737;// level 19
assign po1482 = ~w27741;// level 19
assign po1483 = ~w27744;// level 19
assign po1484 = ~w27747;// level 19
assign po1485 = ~w27750;// level 19
assign po1486 = ~w27753;// level 19
assign po1487 = ~w27756;// level 19
assign po1488 = ~w27759;// level 19
assign po1489 = ~w27762;// level 19
assign po1490 = ~w27765;// level 19
assign po1491 = ~w27768;// level 19
assign po1492 = ~w27771;// level 19
assign po1493 = ~w27774;// level 19
assign po1494 = ~w27777;// level 19
assign po1495 = ~w27780;// level 19
assign po1496 = ~w27784;// level 19
assign po1497 = ~w27787;// level 19
assign po1498 = ~w27790;// level 19
assign po1499 = ~w27793;// level 19
assign po1500 = ~w27796;// level 19
assign po1501 = ~w27799;// level 19
assign po1502 = ~w27802;// level 19
assign po1503 = ~w27805;// level 19
assign po1504 = ~w27808;// level 19
assign po1505 = ~w27811;// level 19
assign po1506 = ~w27814;// level 19
assign po1507 = ~w27817;// level 19
assign po1508 = ~w27820;// level 19
assign po1509 = ~w27823;// level 19
assign po1510 = ~w27827;// level 19
assign po1511 = ~w27830;// level 19
assign po1512 = ~w27833;// level 19
assign po1513 = ~w27836;// level 19
assign po1514 = ~w27839;// level 19
assign po1515 = ~w27842;// level 19
assign po1516 = ~w27845;// level 19
assign po1517 = ~w27848;// level 19
assign po1518 = ~w27851;// level 19
assign po1519 = ~w27854;// level 19
assign po1520 = ~w27857;// level 19
assign po1521 = ~w27860;// level 19
assign po1522 = ~w27863;// level 19
assign po1523 = ~w27866;// level 19
assign po1524 = ~w27870;// level 19
assign po1525 = ~w27873;// level 19
assign po1526 = ~w27876;// level 19
assign po1527 = ~w27879;// level 19
assign po1528 = ~w27882;// level 19
assign po1529 = ~w27885;// level 19
assign po1530 = ~w27888;// level 19
assign po1531 = ~w27891;// level 19
assign po1532 = ~w27894;// level 19
assign po1533 = ~w27897;// level 19
assign po1534 = ~w27900;// level 19
assign po1535 = ~w27903;// level 19
assign po1536 = ~w27906;// level 19
assign po1537 = ~w27909;// level 19
assign po1538 = ~w27913;// level 19
assign po1539 = ~w27916;// level 19
assign po1540 = ~w27919;// level 19
assign po1541 = ~w27922;// level 19
assign po1542 = ~w27925;// level 19
assign po1543 = ~w27928;// level 19
assign po1544 = ~w27931;// level 19
assign po1545 = ~w27934;// level 19
assign po1546 = ~w27937;// level 19
assign po1547 = ~w27940;// level 19
assign po1548 = ~w27943;// level 19
assign po1549 = ~w27946;// level 19
assign po1550 = ~w27949;// level 19
assign po1551 = ~w27952;// level 19
assign po1552 = ~w27956;// level 19
assign po1553 = ~w27959;// level 19
assign po1554 = ~w27962;// level 19
assign po1555 = ~w27965;// level 19
assign po1556 = ~w27968;// level 19
assign po1557 = ~w27971;// level 19
assign po1558 = ~w27974;// level 19
assign po1559 = ~w27977;// level 19
assign po1560 = ~w27980;// level 19
assign po1561 = ~w27983;// level 19
assign po1562 = ~w27986;// level 19
assign po1563 = ~w27989;// level 19
assign po1564 = ~w27992;// level 19
assign po1565 = ~w27995;// level 19
assign po1566 = ~w27999;// level 19
assign po1567 = ~w28002;// level 19
assign po1568 = ~w28005;// level 19
assign po1569 = ~w28008;// level 19
assign po1570 = ~w28011;// level 19
assign po1571 = ~w28014;// level 19
assign po1572 = ~w28017;// level 19
assign po1573 = ~w28020;// level 19
assign po1574 = ~w28023;// level 19
assign po1575 = ~w28026;// level 19
assign po1576 = ~w28029;// level 19
assign po1577 = ~w28032;// level 19
assign po1578 = ~w28035;// level 19
assign po1579 = ~w28038;// level 19
assign po1580 = ~w28042;// level 19
assign po1581 = ~w28045;// level 19
assign po1582 = ~w28048;// level 19
assign po1583 = ~w28051;// level 19
assign po1584 = ~w28054;// level 19
assign po1585 = ~w28057;// level 19
assign po1586 = ~w28060;// level 19
assign po1587 = ~w28063;// level 19
assign po1588 = ~w28066;// level 19
assign po1589 = ~w28069;// level 19
assign po1590 = ~w28072;// level 19
assign po1591 = ~w28075;// level 19
assign po1592 = ~w28078;// level 19
assign po1593 = ~w28081;// level 19
assign po1594 = ~w28085;// level 19
assign po1595 = ~w28088;// level 19
assign po1596 = ~w28091;// level 19
assign po1597 = ~w28094;// level 19
assign po1598 = ~w28097;// level 19
assign po1599 = ~w28100;// level 19
assign po1600 = ~w28103;// level 19
assign po1601 = ~w28106;// level 19
assign po1602 = ~w28109;// level 19
assign po1603 = ~w28112;// level 19
assign po1604 = ~w28115;// level 19
assign po1605 = ~w28118;// level 19
assign po1606 = ~w28121;// level 19
assign po1607 = ~w28124;// level 19
assign po1608 = ~w28128;// level 19
assign po1609 = ~w28131;// level 19
assign po1610 = ~w28134;// level 19
assign po1611 = ~w28137;// level 19
assign po1612 = ~w28140;// level 19
assign po1613 = ~w28143;// level 19
assign po1614 = ~w28146;// level 19
assign po1615 = ~w28149;// level 19
assign po1616 = ~w28152;// level 19
assign po1617 = ~w28155;// level 19
assign po1618 = ~w28158;// level 19
assign po1619 = ~w28161;// level 19
assign po1620 = ~w28164;// level 19
assign po1621 = ~w28167;// level 19
assign po1622 = ~w28170;// level 19
assign po1623 = ~w28173;// level 19
assign po1624 = ~w28176;// level 19
assign po1625 = ~w28179;// level 19
assign po1626 = ~w28182;// level 19
assign po1627 = ~w28185;// level 19
assign po1628 = ~w28188;// level 19
assign po1629 = ~w28191;// level 19
assign po1630 = ~w28194;// level 19
assign po1631 = ~w28197;// level 19
assign po1632 = ~w28200;// level 19
assign po1633 = ~w28203;// level 19
assign po1634 = ~w28206;// level 19
assign po1635 = ~w28209;// level 19
assign po1636 = ~w28213;// level 14
assign po1637 = ~w28215;// level 20
assign po1638 = ~w28218;// level 11
assign po1639 = ~w28221;// level 11
assign po1640 = ~w28225;// level 11
assign po1641 = ~w28229;// level 11
assign po1642 = ~w28232;// level 11
assign po1643 = ~w28235;// level 11
assign po1644 = ~w28239;// level 11
assign po1645 = ~w28242;// level 11
assign po1646 = ~w28245;// level 12
assign po1647 = ~w28248;// level 12
assign po1648 = ~w28251;// level 12
assign po1649 = ~w28254;// level 12
assign po1650 = ~w28258;// level 11
assign po1651 = ~w28261;// level 11
assign po1652 = ~w28264;// level 11
assign po1653 = ~w28267;// level 11
assign po1654 = ~w28270;// level 11
assign po1655 = ~w28273;// level 12
assign po1656 = ~w28277;// level 11
assign po1657 = ~w28280;// level 11
assign po1658 = ~w28283;// level 11
assign po1659 = ~w28286;// level 11
assign po1660 = ~w28289;// level 12
assign po1661 = ~w28293;// level 13
assign po1662 = ~w28296;// level 13
assign po1663 = ~w28299;// level 13
assign po1664 = ~w28302;// level 11
assign po1665 = ~w28305;// level 11
assign po1666 = ~w28308;// level 11
assign po1667 = w28310;// level 19
assign po1668 = w28312;// level 20
assign po1669 = w28314;// level 21
assign po1670 = w28316;// level 24
assign po1671 = w28318;// level 23
assign po1672 = w28320;// level 27
assign po1673 = w28322;// level 12
assign po1674 = w28324;// level 16
assign po1675 = w28326;// level 18
assign po1676 = w28331;// level 8
assign po1677 = w28337;// level 15
assign po1678 = ~w28343;// level 16
assign po1679 = ~w28347;// level 16
assign po1680 = w28395;// level 15
assign po1681 = ~w28401;// level 16
assign po1682 = ~w28407;// level 16
assign po1683 = ~w28411;// level 16
assign po1684 = w28455;// level 12
assign po1685 = w28457;// level 12
assign po1686 = w28459;// level 10
assign po1687 = w28461;// level 19
assign po1688 = w28463;// level 11
assign po1689 = w28465;// level 14
assign po1690 = w28467;// level 13
assign po1691 = w28469;// level 25
assign po1692 = w28471;// level 22
assign po1693 = w28473;// level 22
assign po1694 = ~w28479;// level 16
assign po1695 = ~w28485;// level 16
assign po1696 = w28490;// level 15
assign po1697 = w28495;// level 15
assign po1698 = w28499;// level 15
assign po1699 = w28503;// level 15
assign po1700 = w28506;// level 15
assign po1701 = w28510;// level 15
assign po1702 = w28513;// level 15
assign po1703 = w28516;// level 15
assign po1704 = w28519;// level 15
assign po1705 = w28522;// level 15
assign po1706 = w28525;// level 15
assign po1707 = w28528;// level 15
assign po1708 = w28531;// level 15
assign po1709 = w28534;// level 15
assign po1710 = w28537;// level 15
assign po1711 = w28540;// level 15
assign po1712 = w28543;// level 15
assign po1713 = w28547;// level 15
assign po1714 = w28550;// level 15
assign po1715 = w28553;// level 15
assign po1716 = w28556;// level 15
assign po1717 = w28559;// level 15
assign po1718 = w28562;// level 15
assign po1719 = w28565;// level 15
assign po1720 = w28568;// level 15
assign po1721 = w28571;// level 15
assign po1722 = w28574;// level 15
assign po1723 = w28577;// level 15
assign po1724 = ~w28583;// level 10
assign po1725 = w28586;// level 15
assign po1726 = w28589;// level 15
assign po1727 = w28592;// level 15
assign po1728 = w28598;// level 16
assign po1729 = w28601;// level 15
assign po1730 = ~w28603;// level 10
assign po1731 = ~w28605;// level 10
assign po1732 = ~w28610;// level 15
assign po1733 = ~w28613;// level 16
assign po1734 = ~w28616;// level 16
assign po1735 = ~w28619;// level 16
assign po1736 = ~w28622;// level 16
assign po1737 = ~w28625;// level 16
assign po1738 = ~w28628;// level 16
assign po1739 = ~w28631;// level 16
assign po1740 = ~w28634;// level 16
assign po1741 = w28637;// level 10
assign po1742 = ~w28641;// level 16
assign po1743 = ~w28644;// level 16
assign po1744 = ~w28647;// level 16
assign po1745 = ~w28650;// level 16
assign po1746 = ~w28653;// level 16
assign po1747 = ~w28656;// level 16
assign po1748 = ~w28659;// level 16
assign po1749 = ~w28662;// level 16
assign po1750 = ~w28665;// level 16
assign po1751 = ~w28668;// level 16
assign po1752 = ~w28671;// level 16
assign po1753 = ~w28674;// level 16
assign po1754 = w28677;// level 10
assign po1755 = ~w28679;// level 2
assign po1756 = ~w28680;// level 2
assign po1757 = w28696;// level 7
assign po1758 = w28703;// level 18
assign po1759 = w28706;// level 18
assign po1760 = w28709;// level 18
assign po1761 = w28712;// level 18
assign po1762 = w28715;// level 18
assign po1763 = w28718;// level 18
assign po1764 = w28721;// level 18
assign po1765 = w28724;// level 18
assign po1766 = w28727;// level 18
assign po1767 = w28730;// level 18
assign po1768 = w28733;// level 18
assign po1769 = w28736;// level 18
assign po1770 = pi3409;// level 0
assign po1771 = ~w28761;// level 14
assign po1772 = w28764;// level 15
assign po1773 = w28767;// level 15
assign po1774 = w28771;// level 15
assign po1775 = w28774;// level 15
assign po1776 = ~w28779;// level 16
assign po1777 = ~w28781;// level 10
assign po1778 = ~w28783;// level 10
assign po1779 = ~w28785;// level 10
assign po1780 = ~w28787;// level 10
assign po1781 = ~w28793;// level 10
assign po1782 = ~w28795;// level 10
assign po1783 = ~w28800;// level 17
assign po1784 = w28803;// level 15
assign po1785 = w28806;// level 15
assign po1786 = w28809;// level 15
assign po1787 = w28812;// level 15
assign po1788 = w28815;// level 15
assign po1789 = w28818;// level 15
assign po1790 = w28821;// level 15
assign po1791 = w28824;// level 15
assign po1792 = w28827;// level 15
assign po1793 = w28830;// level 15
assign po1794 = w28833;// level 15
assign po1795 = w28836;// level 15
assign po1796 = w28839;// level 15
assign po1797 = w28842;// level 15
assign po1798 = w28845;// level 15
assign po1799 = w28848;// level 15
assign po1800 = w28851;// level 15
assign po1801 = w28854;// level 15
assign po1802 = w28857;// level 15
assign po1803 = w28860;// level 15
assign po1804 = w28863;// level 15
assign po1805 = w28866;// level 15
assign po1806 = w28869;// level 15
assign po1807 = w28872;// level 15
assign po1808 = w28875;// level 15
assign po1809 = w28878;// level 15
assign po1810 = w28881;// level 15
assign po1811 = w28884;// level 15
assign po1812 = w28887;// level 15
assign po1813 = w28890;// level 15
assign po1814 = w28893;// level 15
assign po1815 = w28896;// level 15
assign po1816 = w28899;// level 15
assign po1817 = w28902;// level 15
assign po1818 = w28905;// level 15
assign po1819 = w28908;// level 15
assign po1820 = w28911;// level 15
assign po1821 = w28914;// level 15
assign po1822 = w28917;// level 15
assign po1823 = w28920;// level 15
assign po1824 = w28923;// level 15
assign po1825 = w28926;// level 15
assign po1826 = w28929;// level 15
assign po1827 = w28932;// level 15
assign po1828 = w28935;// level 15
assign po1829 = w28938;// level 15
assign po1830 = w28941;// level 15
assign po1831 = w28944;// level 15
assign po1832 = w28947;// level 15
assign po1833 = w28950;// level 15
assign po1834 = w28953;// level 15
assign po1835 = w28956;// level 15
assign po1836 = w28959;// level 15
assign po1837 = w28962;// level 15
assign po1838 = w28965;// level 15
assign po1839 = w28968;// level 15
assign po1840 = w28971;// level 15
assign po1841 = w28974;// level 15
assign po1842 = w28977;// level 15
assign po1843 = w28980;// level 15
assign po1844 = w28983;// level 15
assign po1845 = w28986;// level 15
assign po1846 = w28989;// level 15
assign po1847 = w28992;// level 15
assign po1848 = w28995;// level 15
assign po1849 = w28998;// level 15
assign po1850 = w29001;// level 15
assign po1851 = w29004;// level 15
assign po1852 = w29007;// level 15
assign po1853 = w29010;// level 15
assign po1854 = w29013;// level 15
assign po1855 = w29016;// level 15
assign po1856 = w29019;// level 15
assign po1857 = w29022;// level 15
assign po1858 = w29025;// level 15
assign po1859 = w29028;// level 15
assign po1860 = w29031;// level 15
assign po1861 = w29034;// level 15
assign po1862 = w29037;// level 15
assign po1863 = w29040;// level 15
assign po1864 = w29043;// level 15
assign po1865 = w29046;// level 15
assign po1866 = w29049;// level 15
assign po1867 = w29052;// level 15
assign po1868 = w29055;// level 15
assign po1869 = w29058;// level 15
assign po1870 = w29061;// level 15
assign po1871 = w29064;// level 15
assign po1872 = w29067;// level 15
assign po1873 = w29070;// level 15
assign po1874 = w29073;// level 15
assign po1875 = w29076;// level 15
assign po1876 = w29079;// level 15
assign po1877 = w29082;// level 15
assign po1878 = w29085;// level 15
assign po1879 = w29088;// level 15
assign po1880 = w29091;// level 15
assign po1881 = w29094;// level 15
assign po1882 = w29097;// level 15
assign po1883 = w29100;// level 15
assign po1884 = w29103;// level 15
assign po1885 = w29106;// level 15
assign po1886 = w29109;// level 15
assign po1887 = w29112;// level 15
assign po1888 = w29115;// level 15
assign po1889 = w29118;// level 15
assign po1890 = w29121;// level 15
assign po1891 = w29124;// level 15
assign po1892 = w29127;// level 15
assign po1893 = w29130;// level 15
assign po1894 = w29133;// level 15
assign po1895 = w29136;// level 15
assign po1896 = w29139;// level 15
assign po1897 = w29142;// level 15
assign po1898 = w29145;// level 15
assign po1899 = w29148;// level 15
assign po1900 = w29151;// level 15
assign po1901 = w29154;// level 15
assign po1902 = w29157;// level 15
assign po1903 = w29160;// level 15
assign po1904 = w29163;// level 15
assign po1905 = ~w29167;// level 3
assign po1906 = ~w29171;// level 11
assign po1907 = ~w29175;// level 11
assign po1908 = ~w29178;// level 11
assign po1909 = ~w29181;// level 11
assign po1910 = ~w29196;// level 7
assign po1911 = ~w29201;// level 18
assign po1912 = ~w29206;// level 16
assign po1913 = w29211;// level 26
assign po1914 = w29217;// level 7
assign po1915 = w29224;// level 7
assign po1916 = w29234;// level 14
assign po1917 = ~w29242;// level 14
assign po1918 = ~w29245;// level 7
assign po1919 = w29248;// level 11
assign po1920 = w29251;// level 15
assign po1921 = w29254;// level 15
assign po1922 = w29257;// level 15
assign po1923 = w29260;// level 15
assign po1924 = w29263;// level 15
assign po1925 = w29266;// level 15
assign po1926 = w29269;// level 15
assign po1927 = w29272;// level 15
assign po1928 = w29275;// level 15
assign po1929 = w29278;// level 15
assign po1930 = w29281;// level 15
assign po1931 = w29284;// level 15
assign po1932 = w29287;// level 15
assign po1933 = w29290;// level 15
assign po1934 = w29293;// level 15
assign po1935 = w29296;// level 15
assign po1936 = w29299;// level 15
assign po1937 = w29302;// level 15
assign po1938 = w29310;// level 14
assign po1939 = w29314;// level 12
assign po1940 = w29317;// level 12
assign po1941 = w29320;// level 12
assign po1942 = w29323;// level 12
assign po1943 = w29327;// level 13
assign po1944 = w29330;// level 12
assign po1945 = w29333;// level 13
assign po1946 = w29336;// level 13
assign po1947 = w29339;// level 13
assign po1948 = w29342;// level 13
assign po1949 = ~w29346;// level 11
assign po1950 = pi1875;// level 0
assign po1951 = w29347;// level 1
assign po1952 = ~w29353;// level 14
assign po1953 = w29356;// level 6
assign po1954 = w29363;// level 14
assign po1955 = w29365;// level 9
assign po1956 = w29366;// level 6
assign po1957 = ~w29369;// level 11
assign po1958 = w29376;// level 14
assign po1959 = w29379;// level 9
assign po1960 = w29382;// level 13
assign po1961 = w29385;// level 13
assign po1962 = w29388;// level 13
assign po1963 = w29391;// level 13
assign po1964 = w29394;// level 13
assign po1965 = w29397;// level 13
assign po1966 = w29400;// level 13
assign po1967 = w29403;// level 13
assign po1968 = w29406;// level 12
assign po1969 = w29409;// level 12
assign po1970 = w29412;// level 12
assign po1971 = w29415;// level 12
assign po1972 = w29418;// level 12
assign po1973 = w29421;// level 12
assign po1974 = w29424;// level 12
assign po1975 = w29427;// level 12
assign po1976 = ~w29431;// level 11
assign po1977 = ~w29434;// level 11
assign po1978 = w29436;// level 9
assign po1979 = w29438;// level 17
assign po1980 = w29440;// level 8
assign po1981 = w29442;// level 20
assign po1982 = w29444;// level 25
assign po1983 = w29446;// level 24
assign po1984 = ~w29449;// level 10
assign po1985 = w29451;// level 10
assign po1986 = w29454;// level 11
assign po1987 = w29456;// level 12
assign po1988 = w29458;// level 13
assign po1989 = w29460;// level 14
assign po1990 = w29462;// level 15
assign po1991 = w29467;// level 7
assign po1992 = ~w29472;// level 15
assign po1993 = w29476;// level 15
assign po1994 = w29482;// level 14
assign po1995 = w29483;// level 9
assign po1996 = ~w29487;// level 14
assign po1997 = w29492;// level 14
assign po1998 = w29493;// level 9
assign po1999 = w29496;// level 11
assign po2000 = w29499;// level 10
assign po2001 = w29502;// level 7
assign po2002 = w29505;// level 6
assign po2003 = w29508;// level 8
assign po2004 = w29511;// level 6
assign po2005 = w29513;// level 8
assign po2006 = w29515;// level 16
assign po2007 = w29517;// level 12
assign po2008 = w29519;// level 21
assign po2009 = w29521;// level 18
assign po2010 = w29526;// level 14
assign po2011 = w29531;// level 14
assign po2012 = w29536;// level 7
assign po2013 = ~w29540;// level 16
assign po2014 = ~w29545;// level 16
assign po2015 = w29548;// level 14
assign po2016 = w29551;// level 14
assign po2017 = w29554;// level 12
assign po2018 = w29558;// level 12
assign po2019 = w29561;// level 12
assign po2020 = w29564;// level 12
assign po2021 = ~w29582;// level 16
assign po2022 = ~w29588;// level 17
assign po2023 = w29591;// level 15
assign po2024 = ~w29594;// level 16
assign po2025 = ~w29597;// level 16
assign po2026 = ~w29600;// level 16
assign po2027 = ~w29603;// level 16
assign po2028 = ~w29606;// level 16
assign po2029 = ~w29609;// level 16
assign po2030 = ~w29612;// level 15
assign po2031 = ~w29615;// level 15
assign po2032 = ~w29618;// level 16
assign po2033 = ~w29621;// level 16
assign po2034 = ~w29624;// level 16
assign po2035 = ~w29629;// level 16
assign po2036 = ~w29632;// level 16
assign po2037 = ~w29635;// level 16
assign po2038 = ~w29638;// level 16
assign po2039 = ~w29641;// level 16
assign po2040 = ~w29644;// level 16
assign po2041 = ~w29647;// level 16
assign po2042 = ~w29650;// level 16
assign po2043 = ~w29653;// level 16
assign po2044 = ~w29656;// level 16
assign po2045 = ~w29659;// level 16
assign po2046 = ~w29662;// level 16
assign po2047 = w29665;// level 9
assign po2048 = w29668;// level 9
assign po2049 = ~w29673;// level 17
assign po2050 = ~w29678;// level 17
assign po2051 = ~w29683;// level 17
assign po2052 = ~w29688;// level 17
assign po2053 = ~w29693;// level 17
assign po2054 = w29696;// level 9
assign po2055 = w29699;// level 15
assign po2056 = w29702;// level 9
assign po2057 = ~w29708;// level 16
assign po2058 = ~w29711;// level 16
assign po2059 = ~w29714;// level 16
assign po2060 = ~w29717;// level 16
assign po2061 = ~w29720;// level 16
assign po2062 = ~w29723;// level 16
assign po2063 = ~w29726;// level 16
assign po2064 = ~w29729;// level 16
assign po2065 = ~w29732;// level 16
assign po2066 = ~w29735;// level 15
assign po2067 = ~w29738;// level 15
assign po2068 = ~w29741;// level 16
assign po2069 = ~w29745;// level 16
assign po2070 = ~w29748;// level 16
assign po2071 = ~w29751;// level 16
assign po2072 = ~w29754;// level 16
assign po2073 = ~w29757;// level 16
assign po2074 = ~w29760;// level 16
assign po2075 = ~w29763;// level 16
assign po2076 = ~w29766;// level 15
assign po2077 = ~w29769;// level 16
assign po2078 = w29780;// level 9
assign po2079 = w29784;// level 7
assign po2080 = pi3557;// level 0
assign po2081 = ~w29789;// level 16
assign po2082 = ~w29792;// level 16
assign po2083 = ~w29795;// level 16
assign po2084 = ~w29798;// level 16
assign po2085 = ~w29801;// level 16
assign po2086 = ~w29804;// level 16
assign po2087 = ~w29807;// level 16
assign po2088 = ~w29810;// level 16
assign po2089 = ~w29813;// level 16
assign po2090 = ~w29816;// level 15
assign po2091 = ~w29819;// level 16
assign po2092 = ~w29822;// level 16
assign po2093 = ~w29825;// level 16
assign po2094 = ~w29828;// level 16
assign po2095 = ~w29831;// level 16
assign po2096 = ~w29838;// level 14
assign po2097 = w29840;// level 11
assign po2098 = w29842;// level 10
assign po2099 = w29850;// level 20
assign po2100 = w29858;// level 19
assign po2101 = ~w29861;// level 16
assign po2102 = ~w29874;// level 12
assign po2103 = ~w29878;// level 12
assign po2104 = ~w29886;// level 12
assign po2105 = ~w29890;// level 12
assign po2106 = ~w29893;// level 16
assign po2107 = w29896;// level 15
assign po2108 = ~w29900;// level 13
assign po2109 = ~w29904;// level 12
assign po2110 = w29907;// level 12
assign po2111 = w29910;// level 12
assign po2112 = w29913;// level 12
assign po2113 = w29916;// level 12
assign po2114 = w29919;// level 12
assign po2115 = w29922;// level 12
assign po2116 = w29925;// level 12
assign po2117 = w29928;// level 12
assign po2118 = w29931;// level 12
assign po2119 = w29934;// level 12
assign po2120 = w29937;// level 13
assign po2121 = w29940;// level 14
assign po2122 = w29943;// level 14
assign po2123 = w29946;// level 14
assign po2124 = w29949;// level 14
assign po2125 = w29952;// level 14
assign po2126 = w29955;// level 14
assign po2127 = w29958;// level 14
assign po2128 = w29961;// level 14
assign po2129 = w29964;// level 14
assign po2130 = w29967;// level 14
assign po2131 = w29973;// level 7
assign po2132 = w29977;// level 13
assign po2133 = w29986;// level 11
assign po2134 = w29992;// level 12
assign po2135 = w29996;// level 12
assign po2136 = w30000;// level 12
assign po2137 = ~w30003;// level 16
assign po2138 = ~w30006;// level 16
assign po2139 = ~w30009;// level 16
assign po2140 = ~w30012;// level 16
assign po2141 = ~w30015;// level 16
assign po2142 = ~w30018;// level 16
assign po2143 = ~w30021;// level 16
assign po2144 = ~w30024;// level 16
assign po2145 = ~w30027;// level 16
assign po2146 = ~w30030;// level 16
assign po2147 = ~w30033;// level 16
assign po2148 = ~w30036;// level 16
assign po2149 = ~w30043;// level 11
assign po2150 = ~w30048;// level 16
assign po2151 = ~w30059;// level 12
assign po2152 = ~w30063;// level 12
assign po2153 = ~w30072;// level 12
assign po2154 = ~w30076;// level 12
assign po2155 = w30081;// level 14
assign po2156 = w30086;// level 14
assign po2157 = w30091;// level 14
assign po2158 = w30096;// level 14
assign po2159 = w30099;// level 6
assign po2160 = w30101;// level 6
assign po2161 = ~w30104;// level 16
assign po2162 = ~w30107;// level 16
assign po2163 = ~w30110;// level 15
assign po2164 = w30115;// level 8
assign po2165 = ~w30121;// level 13
assign po2166 = ~w30124;// level 16
assign po2167 = ~w30127;// level 16
assign po2168 = w30130;// level 14
assign po2169 = w30131;// level 1
assign po2170 = ~w30136;// level 9
assign po2171 = ~w30140;// level 10
assign po2172 = ~w30144;// level 16
assign po2173 = w30147;// level 11
assign po2174 = w30150;// level 14
assign po2175 = w30153;// level 12
assign po2176 = ~w30158;// level 16
assign po2177 = ~w30163;// level 17
assign po2178 = w30166;// level 8
assign po2179 = ~w30169;// level 15
assign po2180 = w30172;// level 8
assign po2181 = w30175;// level 8
assign po2182 = w30178;// level 11
assign po2183 = ~w30181;// level 16
assign po2184 = ~w30184;// level 16
assign po2185 = w30188;// level 5
assign po2186 = w30189;// level 8
assign po2187 = ~w30192;// level 16
assign po2188 = ~w30195;// level 16
assign po2189 = ~w30198;// level 16
assign po2190 = ~w30201;// level 16
assign po2191 = w30205;// level 16
assign po2192 = w30206;// level 3
assign po2193 = ~w30207;// level 1
assign po2194 = ~w30210;// level 16
assign po2195 = ~w30213;// level 16
assign po2196 = ~w30216;// level 16
assign po2197 = ~w30219;// level 16
assign po2198 = ~w30222;// level 16
assign po2199 = ~w30225;// level 16
assign po2200 = ~w30228;// level 15
assign po2201 = ~w30231;// level 16
assign po2202 = ~w30234;// level 16
assign po2203 = ~w30237;// level 16
assign po2204 = w30240;// level 8
assign po2205 = w30243;// level 8
assign po2206 = w30246;// level 8
assign po2207 = w30247;// level 8
assign po2208 = ~w30252;// level 16
assign po2209 = ~w30256;// level 16
assign po2210 = ~w30259;// level 16
assign po2211 = ~w30262;// level 16
assign po2212 = ~w30265;// level 16
assign po2213 = ~w30268;// level 16
assign po2214 = ~w30271;// level 15
assign po2215 = ~w30274;// level 15
assign po2216 = ~w30277;// level 16
assign po2217 = ~w30280;// level 16
assign po2218 = ~w30283;// level 16
assign po2219 = ~w30287;// level 15
assign po2220 = ~w30290;// level 16
assign po2221 = w30293;// level 8
assign po2222 = w30296;// level 8
assign po2223 = w30299;// level 8
assign po2224 = w30302;// level 8
assign po2225 = w30305;// level 8
assign po2226 = w30308;// level 11
assign po2227 = w30311;// level 8
assign po2228 = ~w30314;// level 15
assign po2229 = ~w30318;// level 16
assign po2230 = ~w30321;// level 16
assign po2231 = ~w30324;// level 16
assign po2232 = ~w30327;// level 16
assign po2233 = ~w30330;// level 16
assign po2234 = ~w30333;// level 16
assign po2235 = ~w30336;// level 16
assign po2236 = ~w30339;// level 16
assign po2237 = ~w30342;// level 16
assign po2238 = ~w30345;// level 16
assign po2239 = ~w30348;// level 15
assign po2240 = ~w30351;// level 15
assign po2241 = ~w30354;// level 16
assign po2242 = ~w30357;// level 16
assign po2243 = ~w30360;// level 16
assign po2244 = ~w30363;// level 16
assign po2245 = ~w30369;// level 32
assign po2246 = ~w30381;// level 6
assign po2247 = ~w30387;// level 5
assign po2248 = w30393;// level 9
assign po2249 = ~w30397;// level 16
assign po2250 = ~w30400;// level 16
assign po2251 = ~w30403;// level 16
assign po2252 = ~w30406;// level 16
assign po2253 = ~w30409;// level 16
assign po2254 = ~w30412;// level 16
assign po2255 = ~w30415;// level 16
assign po2256 = ~w30418;// level 16
assign po2257 = ~w30424;// level 12
assign po2258 = ~w30427;// level 12
assign po2259 = ~w30430;// level 12
assign po2260 = ~w30433;// level 12
assign po2261 = ~w30436;// level 12
assign po2262 = ~w30439;// level 12
assign po2263 = ~w30442;// level 16
assign po2264 = ~w30447;// level 12
assign po2265 = w30450;// level 11
assign po2266 = w30458;// level 20
assign po2267 = w30466;// level 20
assign po2268 = w30474;// level 20
assign po2269 = w30482;// level 20
assign po2270 = w30490;// level 20
assign po2271 = w30498;// level 20
assign po2272 = w30506;// level 20
assign po2273 = w30514;// level 20
assign po2274 = w30522;// level 19
assign po2275 = w30530;// level 20
assign po2276 = w30538;// level 20
assign po2277 = w30546;// level 20
assign po2278 = w30554;// level 20
assign po2279 = w30557;// level 11
assign po2280 = w30560;// level 11
assign po2281 = w30563;// level 11
assign po2282 = ~w30570;// level 13
assign po2283 = ~w30574;// level 14
assign po2284 = ~w30577;// level 14
assign po2285 = ~w30580;// level 14
assign po2286 = ~w30583;// level 14
assign po2287 = w30586;// level 28
assign po2288 = ~w30589;// level 26
assign po2289 = w30592;// level 27
assign po2290 = ~w30594;// level 26
assign po2291 = ~w30596;// level 27
assign po2292 = ~w30599;// level 26
assign po2293 = ~w30602;// level 27
assign po2294 = w30605;// level 28
assign po2295 = ~w30607;// level 28
assign po2296 = w30610;// level 28
assign po2297 = ~w30613;// level 13
assign po2298 = ~w30616;// level 13
assign po2299 = ~w30619;// level 13
assign po2300 = ~w30622;// level 13
assign po2301 = w30625;// level 13
assign po2302 = ~w30628;// level 13
assign po2303 = ~w30631;// level 13
assign po2304 = ~w30634;// level 13
assign po2305 = ~w30637;// level 13
assign po2306 = ~w30640;// level 13
assign po2307 = ~w30643;// level 12
assign po2308 = ~w30646;// level 12
assign po2309 = ~w30649;// level 12
assign po2310 = ~w30652;// level 12
assign po2311 = ~w30655;// level 12
assign po2312 = w30658;// level 12
assign po2313 = ~w30661;// level 12
assign po2314 = ~w30664;// level 12
assign po2315 = ~w30667;// level 12
assign po2316 = ~w30670;// level 12
assign po2317 = ~w30673;// level 12
assign po2318 = ~w30676;// level 12
assign po2319 = ~w30681;// level 13
assign po2320 = ~w30684;// level 13
assign po2321 = w30692;// level 31
assign po2322 = w30700;// level 30
assign po2323 = w30708;// level 29
assign po2324 = ~w30717;// level 29
assign po2325 = w30725;// level 29
assign po2326 = w30733;// level 30
assign po2327 = ~w30742;// level 30
assign po2328 = ~w30746;// level 11
assign po2329 = ~w30750;// level 11
assign po2330 = ~w30754;// level 11
assign po2331 = ~w30757;// level 12
assign po2332 = ~w30763;// level 11
assign po2333 = w30766;// level 11
assign po2334 = w30769;// level 11
assign po2335 = w30772;// level 11
assign po2336 = w30775;// level 11
assign po2337 = w30778;// level 11
assign po2338 = w30781;// level 11
assign po2339 = w30784;// level 11
assign po2340 = w30789;// level 11
assign po2341 = w30794;// level 11
assign po2342 = w30797;// level 11
assign po2343 = w30800;// level 11
assign po2344 = w30803;// level 11
assign po2345 = w30806;// level 11
assign po2346 = w30809;// level 11
assign po2347 = w30812;// level 11
assign po2348 = w30815;// level 11
assign po2349 = w30818;// level 11
assign po2350 = w30821;// level 11
assign po2351 = w30824;// level 11
assign po2352 = w30827;// level 11
assign po2353 = w30830;// level 11
assign po2354 = w30833;// level 11
assign po2355 = w30836;// level 11
assign po2356 = w30839;// level 11
assign po2357 = w30843;// level 11
assign po2358 = w30847;// level 11
assign po2359 = ~w30851;// level 10
assign po2360 = w30862;// level 14
assign po2361 = w30865;// level 11
assign po2362 = ~w30868;// level 16
assign po2363 = ~w30871;// level 16
assign po2364 = ~w30874;// level 16
assign po2365 = ~w30877;// level 16
assign po2366 = ~w30880;// level 16
assign po2367 = w30885;// level 6
assign po2368 = ~w30888;// level 16
assign po2369 = ~w30893;// level 16
assign po2370 = ~w30899;// level 16
assign po2371 = w30902;// level 11
assign po2372 = ~w30907;// level 16
assign po2373 = w30910;// level 11
assign po2374 = w30913;// level 11
assign po2375 = w30916;// level 11
assign po2376 = w30919;// level 11
assign po2377 = w30922;// level 11
assign po2378 = ~w30925;// level 16
assign po2379 = ~w30928;// level 16
assign po2380 = ~w30931;// level 13
assign po2381 = ~w30934;// level 12
assign po2382 = ~w30937;// level 12
assign po2383 = ~w30940;// level 13
assign po2384 = ~w30943;// level 12
assign po2385 = ~w30946;// level 13
assign po2386 = ~w30949;// level 13
assign po2387 = ~w30952;// level 13
assign po2388 = ~w30955;// level 13
assign po2389 = ~w30958;// level 12
assign po2390 = w30966;// level 11
assign po2391 = w30975;// level 11
assign po2392 = w30980;// level 11
assign po2393 = w30996;// level 15
assign po2394 = w31005;// level 11
assign po2395 = ~w31008;// level 16
assign po2396 = ~w31012;// level 18
assign po2397 = w31020;// level 11
assign po2398 = ~w31023;// level 16
assign po2399 = ~w31026;// level 16
assign po2400 = ~w31029;// level 16
assign po2401 = w31032;// level 16
assign po2402 = w31035;// level 16
assign po2403 = w31038;// level 16
assign po2404 = w31041;// level 16
assign po2405 = w31044;// level 16
assign po2406 = w31047;// level 15
assign po2407 = w31050;// level 16
assign po2408 = w31053;// level 16
assign po2409 = w31056;// level 16
assign po2410 = w31057;// level 3
assign po2411 = ~w31058;// level 1
assign po2412 = w31059;// level 15
assign po2413 = w31069;// level 16
assign po2414 = w31078;// level 16
assign po2415 = w31087;// level 16
assign po2416 = w31096;// level 16
assign po2417 = w31105;// level 16
assign po2418 = w31114;// level 16
assign po2419 = w31123;// level 16
assign po2420 = w31132;// level 16
assign po2421 = w31141;// level 15
assign po2422 = w31150;// level 16
assign po2423 = ~w31153;// level 16
assign po2424 = ~w31157;// level 32
assign po2425 = w31161;// level 15
assign po2426 = ~w31168;// level 13
assign po2427 = ~w31171;// level 12
assign po2428 = ~w31174;// level 12
assign po2429 = ~w31177;// level 12
assign po2430 = ~w31180;// level 12
assign po2431 = ~w31183;// level 12
assign po2432 = ~w31186;// level 12
assign po2433 = ~w31189;// level 12
assign po2434 = ~w31192;// level 16
assign po2435 = w31201;// level 15
assign po2436 = ~w31205;// level 17
assign po2437 = ~w31208;// level 17
assign po2438 = ~w31211;// level 17
assign po2439 = ~w31214;// level 16
assign po2440 = ~w31217;// level 16
assign po2441 = ~w31220;// level 17
assign po2442 = ~w31223;// level 17
assign po2443 = ~w31226;// level 16
assign po2444 = ~w31229;// level 17
assign po2445 = ~w31232;// level 15
assign po2446 = ~w31235;// level 16
assign po2447 = ~w31238;// level 16
assign po2448 = ~w31241;// level 16
assign po2449 = ~w31244;// level 16
assign po2450 = ~w31247;// level 17
assign po2451 = ~w31250;// level 17
assign po2452 = ~w31253;// level 12
assign po2453 = w31262;// level 16
assign po2454 = ~w31264;// level 11
assign po2455 = w31266;// level 7
assign po2456 = ~w31267;// level 12
assign po2457 = ~w31270;// level 18
assign po2458 = ~w31273;// level 18
assign po2459 = ~w31276;// level 18
assign po2460 = ~w31279;// level 18
assign po2461 = ~w31282;// level 18
assign po2462 = ~w31285;// level 18
assign po2463 = ~w31288;// level 18
assign po2464 = ~w31291;// level 18
assign po2465 = ~w31294;// level 17
assign po2466 = ~w31297;// level 17
assign po2467 = ~w31300;// level 18
assign po2468 = ~w31303;// level 18
assign po2469 = ~w31306;// level 18
assign po2470 = ~w31309;// level 18
assign po2471 = ~w31312;// level 16
assign po2472 = w31315;// level 20
assign po2473 = w31318;// level 19
assign po2474 = ~w31322;// level 17
assign po2475 = ~w31325;// level 17
assign po2476 = ~w31328;// level 17
assign po2477 = ~w31331;// level 16
assign po2478 = ~w31334;// level 16
assign po2479 = ~w31337;// level 17
assign po2480 = ~w31340;// level 17
assign po2481 = ~w31343;// level 16
assign po2482 = ~w31346;// level 17
assign po2483 = ~w31349;// level 15
assign po2484 = ~w31352;// level 16
assign po2485 = ~w31355;// level 16
assign po2486 = ~w31358;// level 16
assign po2487 = ~w31361;// level 16
assign po2488 = ~w31364;// level 17
assign po2489 = ~w31367;// level 17
assign po2490 = ~w31371;// level 17
assign po2491 = ~w31374;// level 17
assign po2492 = ~w31377;// level 17
assign po2493 = ~w31380;// level 16
assign po2494 = ~w31383;// level 16
assign po2495 = ~w31386;// level 17
assign po2496 = ~w31389;// level 17
assign po2497 = ~w31392;// level 16
assign po2498 = ~w31395;// level 17
assign po2499 = ~w31398;// level 15
assign po2500 = ~w31401;// level 16
assign po2501 = ~w31404;// level 16
assign po2502 = ~w31407;// level 16
assign po2503 = ~w31410;// level 16
assign po2504 = ~w31413;// level 17
assign po2505 = ~w31416;// level 17
assign po2506 = w31420;// level 11
assign po2507 = w31425;// level 11
assign po2508 = w31433;// level 11
assign po2509 = w31438;// level 11
assign po2510 = w31443;// level 11
assign po2511 = w31451;// level 11
assign po2512 = w31456;// level 11
assign po2513 = w31461;// level 11
assign po2514 = ~w31464;// level 16
assign po2515 = ~w31467;// level 16
assign po2516 = ~w31470;// level 16
assign po2517 = ~w31473;// level 16
assign po2518 = ~w31476;// level 16
assign po2519 = ~w31479;// level 16
assign po2520 = ~w31482;// level 16
assign po2521 = ~w31485;// level 16
assign po2522 = ~w31488;// level 16
assign po2523 = ~w31491;// level 16
assign po2524 = ~w31494;// level 16
assign po2525 = ~w31497;// level 16
assign po2526 = ~w31500;// level 16
assign po2527 = ~w31503;// level 16
assign po2528 = ~w31505;// level 16
assign po2529 = ~w31508;// level 16
assign po2530 = ~w31511;// level 16
assign po2531 = ~w31514;// level 16
assign po2532 = ~w31517;// level 16
assign po2533 = ~w31520;// level 16
assign po2534 = ~w31523;// level 16
assign po2535 = ~w31526;// level 16
assign po2536 = ~w31529;// level 16
assign po2537 = ~w31532;// level 16
assign po2538 = ~w31535;// level 16
assign po2539 = ~w31538;// level 16
assign po2540 = ~w31541;// level 16
assign po2541 = ~w31544;// level 16
assign po2542 = ~w31547;// level 16
assign po2543 = ~w31550;// level 16
assign po2544 = ~w31552;// level 16
assign po2545 = ~w31555;// level 16
assign po2546 = ~w31557;// level 16
assign po2547 = ~w31559;// level 16
assign po2548 = ~w31562;// level 16
assign po2549 = ~w31564;// level 16
assign po2550 = ~w31567;// level 16
assign po2551 = ~w31570;// level 16
assign po2552 = ~w31573;// level 16
assign po2553 = ~w31575;// level 16
assign po2554 = ~w31578;// level 16
assign po2555 = ~w31580;// level 16
assign po2556 = ~w31583;// level 16
assign po2557 = ~w31586;// level 16
assign po2558 = ~w31589;// level 16
assign po2559 = ~w31592;// level 16
assign po2560 = ~w31595;// level 16
assign po2561 = ~w31598;// level 16
assign po2562 = ~w31601;// level 16
assign po2563 = ~w31604;// level 16
assign po2564 = ~w31607;// level 16
assign po2565 = ~w31610;// level 16
assign po2566 = ~w31613;// level 16
assign po2567 = ~w31616;// level 16
assign po2568 = ~w31619;// level 16
assign po2569 = ~w31622;// level 16
assign po2570 = ~w31624;// level 28
assign po2571 = w31627;// level 26
assign po2572 = ~w31630;// level 26
assign po2573 = ~w31632;// level 27
assign po2574 = ~w31634;// level 28
assign po2575 = ~w31637;// level 26
assign po2576 = w31640;// level 27
assign po2577 = w31643;// level 26
assign po2578 = w31646;// level 27
assign po2579 = ~w31648;// level 26
assign po2580 = ~w31650;// level 27
assign po2581 = ~w31652;// level 28
assign po2582 = ~w31655;// level 28
assign po2583 = w31658;// level 28
assign po2584 = w31661;// level 28
assign po2585 = ~w31663;// level 26
assign po2586 = ~w31665;// level 26
assign po2587 = ~w31668;// level 26
assign po2588 = ~w31670;// level 27
assign po2589 = w31673;// level 28
assign po2590 = w31676;// level 28
assign po2591 = ~w31679;// level 28
assign po2592 = ~w31682;// level 16
assign po2593 = ~w31685;// level 16
assign po2594 = ~w31688;// level 16
assign po2595 = ~w31691;// level 16
assign po2596 = ~w31694;// level 16
assign po2597 = ~w31697;// level 16
assign po2598 = ~w31700;// level 16
assign po2599 = ~w31703;// level 16
assign po2600 = ~w31706;// level 16
assign po2601 = ~w31709;// level 16
assign po2602 = ~w31712;// level 16
assign po2603 = ~w31715;// level 16
assign po2604 = ~w31718;// level 16
assign po2605 = ~w31721;// level 16
assign po2606 = ~w31724;// level 16
assign po2607 = ~w31727;// level 16
assign po2608 = ~w31730;// level 16
assign po2609 = ~w31733;// level 16
assign po2610 = ~w31736;// level 16
assign po2611 = ~w31739;// level 16
assign po2612 = ~w31742;// level 16
assign po2613 = ~w31745;// level 16
assign po2614 = ~w31748;// level 16
assign po2615 = ~w31751;// level 16
assign po2616 = ~w31753;// level 16
assign po2617 = ~w31756;// level 16
assign po2618 = ~w31759;// level 16
assign po2619 = ~w31762;// level 16
assign po2620 = ~w31765;// level 16
assign po2621 = ~w31767;// level 16
assign po2622 = ~w31769;// level 16
assign po2623 = ~w31771;// level 16
assign po2624 = ~w31774;// level 16
assign po2625 = ~w31777;// level 16
assign po2626 = ~w31780;// level 16
assign po2627 = ~w31783;// level 16
assign po2628 = ~w31786;// level 16
assign po2629 = ~w31789;// level 16
assign po2630 = ~w31792;// level 16
assign po2631 = ~w31795;// level 16
assign po2632 = ~w31798;// level 16
assign po2633 = ~w31801;// level 16
assign po2634 = ~w31803;// level 16
assign po2635 = ~w31806;// level 16
assign po2636 = ~w31809;// level 16
assign po2637 = ~w31811;// level 16
assign po2638 = ~w31814;// level 16
assign po2639 = ~w31817;// level 16
assign po2640 = ~w31819;// level 16
assign po2641 = w31822;// level 13
assign po2642 = w31825;// level 13
assign po2643 = ~w31828;// level 13
assign po2644 = ~w31831;// level 13
assign po2645 = ~w31834;// level 13
assign po2646 = ~w31837;// level 13
assign po2647 = ~w31840;// level 13
assign po2648 = w31843;// level 13
assign po2649 = ~w31846;// level 12
assign po2650 = ~w31849;// level 12
assign po2651 = w31852;// level 12
assign po2652 = ~w31855;// level 12
assign po2653 = w31858;// level 12
assign po2654 = ~w31861;// level 12
assign po2655 = ~w31864;// level 12
assign po2656 = ~w31867;// level 12
assign po2657 = ~w31870;// level 12
assign po2658 = ~w31873;// level 12
assign po2659 = ~w31876;// level 12
assign po2660 = ~w31879;// level 12
assign po2661 = ~w31882;// level 12
assign po2662 = ~w31885;// level 12
assign po2663 = ~w31888;// level 12
assign po2664 = ~w31891;// level 12
assign po2665 = ~w31894;// level 12
assign po2666 = w31897;// level 12
assign po2667 = w31900;// level 12
assign po2668 = ~w31903;// level 12
assign po2669 = ~w31906;// level 12
assign po2670 = ~w31909;// level 12
assign po2671 = w31912;// level 12
assign po2672 = ~w31915;// level 13
assign po2673 = ~w31918;// level 13
assign po2674 = ~w31921;// level 13
assign po2675 = w31924;// level 13
assign po2676 = ~w31927;// level 13
assign po2677 = w31930;// level 13
assign po2678 = ~w31933;// level 13
assign po2679 = ~w31936;// level 13
assign po2680 = ~w31939;// level 13
assign po2681 = ~w31942;// level 13
assign po2682 = ~w31945;// level 13
assign po2683 = ~w31948;// level 13
assign po2684 = ~w31951;// level 13
assign po2685 = ~w31954;// level 13
assign po2686 = w31962;// level 30
assign po2687 = w31970;// level 29
assign po2688 = w31976;// level 31
assign po2689 = w31984;// level 31
assign po2690 = w31992;// level 31
assign po2691 = w32000;// level 31
assign po2692 = ~w32002;// level 14
assign po2693 = ~w32006;// level 13
assign po2694 = ~w32015;// level 8
assign po2695 = ~w32018;// level 12
assign po2696 = ~w32023;// level 22
assign po2697 = ~w32025;// level 10
assign po2698 = ~w32031;// level 5
assign po2699 = ~w32032;// level 6
assign po2700 = ~w32062;// level 8
assign po2701 = w20920;// level 8
assign po2702 = ~w32065;// level 12
assign po2703 = ~w32068;// level 13
assign po2704 = ~w32071;// level 12
assign po2705 = ~w32074;// level 12
assign po2706 = w32082;// level 31
assign po2707 = w32085;// level 16
assign po2708 = w32088;// level 15
assign po2709 = w32091;// level 16
assign po2710 = w32094;// level 16
assign po2711 = w32097;// level 16
assign po2712 = w32100;// level 16
assign po2713 = w21419;// level 8
assign po2714 = w32109;// level 18
assign po2715 = ~w32117;// level 9
assign po2716 = w32122;// level 7
assign po2717 = ~w32130;// level 9
assign po2718 = w32138;// level 18
assign po2719 = w32141;// level 18
assign po2720 = w32144;// level 12
assign po2721 = w32147;// level 13
assign po2722 = w32151;// level 18
assign po2723 = w32155;// level 18
assign po2724 = ~w32157;// level 28
assign po2725 = ~w32159;// level 28
assign po2726 = ~w32161;// level 28
assign po2727 = ~w32163;// level 28
assign po2728 = ~w32166;// level 12
assign po2729 = ~w32173;// level 11
assign po2730 = w32175;// level 7
assign po2731 = ~w32177;// level 10
assign po2732 = ~w32180;// level 12
assign po2733 = ~w32184;// level 13
assign po2734 = w32187;// level 20
assign po2735 = w32190;// level 20
assign po2736 = w32193;// level 20
assign po2737 = w32196;// level 20
assign po2738 = w32199;// level 20
assign po2739 = w32202;// level 20
assign po2740 = w32205;// level 20
assign po2741 = w32208;// level 20
assign po2742 = w32211;// level 19
assign po2743 = w32214;// level 20
assign po2744 = w32217;// level 20
assign po2745 = w32220;// level 20
assign po2746 = ~w32222;// level 27
assign po2747 = ~w32224;// level 26
assign po2748 = ~w32226;// level 27
assign po2749 = ~w32228;// level 28
assign po2750 = ~w32231;// level 28
assign po2751 = ~w32233;// level 28
assign po2752 = w32236;// level 27
assign po2753 = w32239;// level 28
assign po2754 = ~w32241;// level 28
assign po2755 = ~w32244;// level 28
assign po2756 = ~w32246;// level 27
assign po2757 = ~w32248;// level 27
assign po2758 = ~w32251;// level 27
assign po2759 = w32254;// level 28
assign po2760 = ~w32257;// level 28
assign po2761 = w32260;// level 28
assign po2762 = ~w32266;// level 11
assign po2763 = ~w32272;// level 11
assign po2764 = ~w32278;// level 11
assign po2765 = ~w32284;// level 11
assign po2766 = ~w32286;// level 28
assign po2767 = ~w32288;// level 28
assign po2768 = ~w32290;// level 28
assign po2769 = ~w32292;// level 28
assign po2770 = ~w32294;// level 27
assign po2771 = ~w32296;// level 28
assign po2772 = ~w32298;// level 28
assign po2773 = ~w32300;// level 28
assign po2774 = ~w32302;// level 28
assign po2775 = ~w32304;// level 28
assign po2776 = ~w32306;// level 28
assign po2777 = ~w32308;// level 28
assign po2778 = ~w32310;// level 28
assign po2779 = ~w32312;// level 27
assign po2780 = ~w32315;// level 28
assign po2781 = ~w32317;// level 28
assign po2782 = ~w32319;// level 28
assign po2783 = ~w32321;// level 28
assign po2784 = ~w32323;// level 27
assign po2785 = w32326;// level 13
assign po2786 = w32329;// level 18
assign po2787 = w32332;// level 18
assign po2788 = ~w32336;// level 11
assign po2789 = ~w32339;// level 10
assign po2790 = ~w32342;// level 10
assign po2791 = ~w32345;// level 10
assign po2792 = ~w32348;// level 10
assign po2793 = ~w32351;// level 10
assign po2794 = ~w32354;// level 10
assign po2795 = ~w32357;// level 10
assign po2796 = ~w32360;// level 10
assign po2797 = ~w32363;// level 10
assign po2798 = ~w32366;// level 10
assign po2799 = ~w32369;// level 10
assign po2800 = ~w32373;// level 11
assign po2801 = ~w32375;// level 21
assign po2802 = ~w32378;// level 11
assign po2803 = ~w32383;// level 21
assign po2804 = ~w32387;// level 21
assign po2805 = ~w32391;// level 21
assign po2806 = w32396;// level 4
assign po2807 = ~w32400;// level 4
assign po2808 = ~w32404;// level 16
assign po2809 = ~w32407;// level 16
assign po2810 = ~w32410;// level 16
assign po2811 = ~w32413;// level 16
assign po2812 = ~w32416;// level 16
assign po2813 = ~w32419;// level 16
assign po2814 = ~w32422;// level 16
assign po2815 = ~w32425;// level 16
assign po2816 = ~w32428;// level 16
assign po2817 = ~w32431;// level 16
assign po2818 = w32439;// level 19
assign po2819 = w32443;// level 19
assign po2820 = w32447;// level 19
assign po2821 = w32452;// level 7
assign po2822 = w32458;// level 7
assign po2823 = w27425;// level 12
assign po2824 = w28384;// level 12
assign po2825 = w32462;// level 7
assign po2826 = w32465;// level 20
assign po2827 = ~w32468;// level 16
assign po2828 = ~w32471;// level 16
assign po2829 = w32474;// level 18
assign po2830 = ~w32476;// level 6
assign po2831 = ~w32479;// level 10
assign po2832 = ~w32482;// level 10
assign po2833 = ~w32485;// level 10
assign po2834 = w32488;// level 12
assign po2835 = ~w32490;// level 28
assign po2836 = w21451;// level 6
assign po2837 = w32494;// level 18
assign po2838 = w32495;// level 6
assign po2839 = ~w32497;// level 27
assign po2840 = ~w32499;// level 28
assign po2841 = ~w32501;// level 28
assign po2842 = ~w32503;// level 28
assign po2843 = ~w32505;// level 16
assign po2844 = ~w32508;// level 30
assign po2845 = ~w32510;// level 28
assign po2846 = ~w32512;// level 16
assign po2847 = ~w32514;// level 16
assign po2848 = ~w32516;// level 28
assign po2849 = ~w32518;// level 16
assign po2850 = ~w32520;// level 28
assign po2851 = ~w32522;// level 16
assign po2852 = ~w32526;// level 17
assign po2853 = ~w32529;// level 16
assign po2854 = ~w32532;// level 28
assign po2855 = ~w32535;// level 30
assign po2856 = ~w32538;// level 17
assign po2857 = ~w32541;// level 16
assign po2858 = ~w32544;// level 16
assign po2859 = ~w32546;// level 28
assign po2860 = ~w32549;// level 16
assign po2861 = ~w32551;// level 16
assign po2862 = ~w32554;// level 16
assign po2863 = ~w32556;// level 16
assign po2864 = ~w32559;// level 29
assign po2865 = ~w32561;// level 16
assign po2866 = ~w32564;// level 29
assign po2867 = ~w32566;// level 16
assign po2868 = ~w32569;// level 28
assign po2869 = ~w32575;// level 11
assign po2870 = w32576;// level 1
assign po2871 = ~w32582;// level 11
assign po2872 = ~w32588;// level 11
assign po2873 = ~w32594;// level 11
assign po2874 = ~w32600;// level 11
assign po2875 = ~w32602;// level 16
assign po2876 = ~w32604;// level 16
assign po2877 = ~w32606;// level 16
assign po2878 = ~w32608;// level 16
assign po2879 = pi3137;// level 0
assign po2880 = ~w32610;// level 16
assign po2881 = ~w32612;// level 16
assign po2882 = pi3142;// level 0
assign po2883 = ~w32617;// level 16
assign po2884 = ~w32620;// level 16
assign po2885 = ~w32623;// level 16
assign po2886 = ~w32626;// level 16
assign po2887 = ~w32629;// level 16
assign po2888 = ~w32632;// level 16
assign po2889 = ~w32635;// level 16
assign po2890 = ~w32638;// level 16
assign po2891 = ~w32641;// level 15
assign po2892 = ~w32644;// level 15
assign po2893 = ~w32647;// level 16
assign po2894 = ~w32650;// level 16
assign po2895 = ~w32653;// level 16
assign po2896 = ~w32656;// level 16
assign po2897 = ~w32659;// level 16
assign po2898 = w32668;// level 16
assign po2899 = w32673;// level 16
assign po2900 = w32678;// level 16
assign po2901 = w32683;// level 16
assign po2902 = w32688;// level 16
assign po2903 = w32693;// level 16
assign po2904 = w32698;// level 16
assign po2905 = w32703;// level 16
assign po2906 = w32708;// level 15
assign po2907 = w32713;// level 15
assign po2908 = w32718;// level 16
assign po2909 = w32723;// level 16
assign po2910 = w32728;// level 16
assign po2911 = w32733;// level 16
assign po2912 = w32738;// level 16
assign po2913 = w32739;// level 1
assign po2914 = ~w32742;// level 12
assign po2915 = pi3129;// level 0
assign po2916 = w32745;// level 15
assign po2917 = w32746;// level 1
assign po2918 = ~w32751;// level 4
assign po2919 = ~w32753;// level 16
assign po2920 = ~w32756;// level 16
assign po2921 = w32757;// level 3
assign po2922 = ~w32759;// level 2
assign po2923 = ~w32763;// level 18
assign po2924 = ~w32766;// level 18
assign po2925 = ~w32769;// level 18
assign po2926 = ~w32772;// level 18
assign po2927 = ~w32775;// level 18
assign po2928 = ~w32778;// level 18
assign po2929 = ~w32782;// level 18
assign po2930 = ~w32785;// level 18
assign po2931 = ~w32788;// level 18
assign po2932 = ~w32791;// level 18
assign po2933 = ~w32794;// level 16
assign po2934 = ~w32797;// level 18
assign po2935 = ~w32800;// level 18
assign po2936 = ~w32804;// level 18
assign po2937 = ~w32807;// level 18
assign po2938 = ~w32810;// level 18
assign po2939 = ~w32813;// level 18
assign po2940 = ~w32816;// level 18
assign po2941 = ~w32819;// level 18
assign po2942 = ~w32823;// level 18
assign po2943 = ~w32826;// level 18
assign po2944 = ~w32829;// level 18
assign po2945 = ~w32832;// level 18
assign po2946 = ~w32835;// level 18
assign po2947 = ~w32838;// level 18
assign po2948 = ~w32841;// level 17
assign po2949 = ~w32844;// level 17
assign po2950 = ~w32847;// level 17
assign po2951 = ~w32850;// level 16
assign po2952 = ~w32853;// level 16
assign po2953 = ~w32856;// level 17
assign po2954 = ~w32859;// level 16
assign po2955 = ~w32862;// level 17
assign po2956 = ~w32865;// level 15
assign po2957 = ~w32868;// level 16
assign po2958 = ~w32871;// level 16
assign po2959 = ~w32874;// level 16
assign po2960 = ~w32877;// level 17
assign po2961 = w32881;// level 5
assign po2962 = ~w32884;// level 30
assign po2963 = ~w32887;// level 29
assign po2964 = ~w32890;// level 28
assign po2965 = ~w32893;// level 30
assign po2966 = ~w32895;// level 16
assign po2967 = ~w32897;// level 16
assign po2968 = ~w32899;// level 16
assign po2969 = ~w32901;// level 16
assign po2970 = ~w32903;// level 16
assign po2971 = ~w32905;// level 16
assign po2972 = ~w32907;// level 16
assign po2973 = ~w32909;// level 16
assign po2974 = ~w32911;// level 16
assign po2975 = ~w32913;// level 16
assign po2976 = ~w32915;// level 16
assign po2977 = ~w32917;// level 16
assign po2978 = ~w32919;// level 16
assign po2979 = ~w32921;// level 16
assign po2980 = ~w32923;// level 16
assign po2981 = ~w32925;// level 16
assign po2982 = ~w32927;// level 16
assign po2983 = ~w32929;// level 16
assign po2984 = ~w32931;// level 16
assign po2985 = ~w32933;// level 16
assign po2986 = ~w32935;// level 16
assign po2987 = ~w32937;// level 16
assign po2988 = ~w32939;// level 16
assign po2989 = ~w32941;// level 16
assign po2990 = ~w32943;// level 16
assign po2991 = ~w32945;// level 16
assign po2992 = ~w32947;// level 16
assign po2993 = ~w32950;// level 16
assign po2994 = ~w32952;// level 16
assign po2995 = ~w32954;// level 16
assign po2996 = ~w32957;// level 16
assign po2997 = ~w32960;// level 16
assign po2998 = ~w32963;// level 16
assign po2999 = ~w32965;// level 16
assign po3000 = ~w32968;// level 16
assign po3001 = ~w32971;// level 16
assign po3002 = ~w32974;// level 16
assign po3003 = ~w32977;// level 16
assign po3004 = ~w32980;// level 16
assign po3005 = ~w32982;// level 16
assign po3006 = ~w32984;// level 16
assign po3007 = ~w32986;// level 16
assign po3008 = ~w32988;// level 16
assign po3009 = ~w32990;// level 16
assign po3010 = ~w32992;// level 16
assign po3011 = ~w32994;// level 16
assign po3012 = ~w32996;// level 16
assign po3013 = ~w32998;// level 16
assign po3014 = ~w33000;// level 16
assign po3015 = ~w33002;// level 16
assign po3016 = ~w33005;// level 27
assign po3017 = ~w33007;// level 28
assign po3018 = ~w33009;// level 28
assign po3019 = w33012;// level 27
assign po3020 = ~w33014;// level 28
assign po3021 = ~w33016;// level 28
assign po3022 = ~w33022;// level 11
assign po3023 = ~w33028;// level 11
assign po3024 = ~w33034;// level 11
assign po3025 = ~w33040;// level 11
assign po3026 = ~w33042;// level 16
assign po3027 = ~w33044;// level 16
assign po3028 = ~w33046;// level 16
assign po3029 = ~w33048;// level 16
assign po3030 = ~w33050;// level 16
assign po3031 = ~w33052;// level 16
assign po3032 = ~w33054;// level 16
assign po3033 = ~w33056;// level 16
assign po3034 = ~w33058;// level 16
assign po3035 = ~w33060;// level 16
assign po3036 = ~w33062;// level 16
assign po3037 = ~w33064;// level 16
assign po3038 = ~w33066;// level 16
assign po3039 = ~w33068;// level 16
assign po3040 = ~w33070;// level 16
assign po3041 = ~w33072;// level 16
assign po3042 = ~w33074;// level 16
assign po3043 = ~w33076;// level 16
assign po3044 = ~w33078;// level 16
assign po3045 = ~w33080;// level 16
assign po3046 = ~w33082;// level 16
assign po3047 = ~w33085;// level 16
assign po3048 = ~w33087;// level 16
assign po3049 = ~w33089;// level 16
assign po3050 = ~w33092;// level 16
assign po3051 = ~w33095;// level 16
assign po3052 = ~w33097;// level 16
assign po3053 = ~w33099;// level 16
assign po3054 = ~w33101;// level 16
assign po3055 = ~w33104;// level 16
assign po3056 = ~w33107;// level 16
assign po3057 = ~w33110;// level 16
assign po3058 = ~w33113;// level 16
assign po3059 = ~w33116;// level 16
assign po3060 = ~w33119;// level 16
assign po3061 = ~w33122;// level 16
assign po3062 = ~w33125;// level 16
assign po3063 = ~w33127;// level 16
assign po3064 = w33130;// level 28
assign po3065 = ~w33132;// level 28
assign po3066 = ~w33134;// level 28
assign po3067 = ~w33137;// level 28
assign po3068 = ~w33140;// level 28
assign po3069 = ~w33142;// level 28
assign po3070 = ~w33144;// level 28
assign po3071 = ~w33146;// level 28
assign po3072 = ~w33148;// level 28
assign po3073 = ~w33150;// level 28
assign po3074 = ~w33152;// level 28
assign po3075 = ~w33156;// level 11
assign po3076 = w33159;// level 12
assign po3077 = w33162;// level 14
assign po3078 = w33165;// level 7
assign po3079 = w33168;// level 5
assign po3080 = w33171;// level 5
assign po3081 = ~w33173;// level 20
assign po3082 = w33178;// level 16
assign po3083 = w21365;// level 6
assign po3084 = ~w33180;// level 13
assign po3085 = w33184;// level 14
assign po3086 = ~w33187;// level 16
assign po3087 = ~w33189;// level 6
assign po3088 = w33193;// level 8
assign po3089 = w33196;// level 7
assign po3090 = w33199;// level 7
assign po3091 = ~w33201;// level 16
assign po3092 = ~w33203;// level 16
assign po3093 = w33207;// level 5
assign po3094 = ~w33209;// level 28
assign po3095 = ~w33213;// level 11
assign po3096 = ~w33217;// level 18
assign po3097 = ~w33220;// level 20
assign po3098 = w33223;// level 27
assign po3099 = ~w33226;// level 18
assign po3100 = ~w33229;// level 18
assign po3101 = ~w33233;// level 17
assign po3102 = ~w33236;// level 17
assign po3103 = ~w33240;// level 12
assign po3104 = w33244;// level 5
assign po3105 = ~w33247;// level 18
assign po3106 = ~w33250;// level 30
assign po3107 = ~w33253;// level 19
assign po3108 = w33257;// level 5
assign po3109 = w33261;// level 5
assign po3110 = w33265;// level 5
assign po3111 = ~w33269;// level 17
assign po3112 = ~w33272;// level 30
assign po3113 = w33273;// level 9
assign po3114 = ~w33276;// level 29
assign po3115 = ~w33279;// level 28
assign po3116 = w33282;// level 15
assign po3117 = w33285;// level 15
assign po3118 = w33287;// level 6
assign po3119 = ~w33290;// level 16
assign po3120 = ~w33292;// level 10
assign po3121 = ~w33295;// level 16
assign po3122 = ~w33298;// level 16
assign po3123 = ~w33301;// level 15
assign po3124 = w33304;// level 5
assign po3125 = ~w33307;// level 16
assign po3126 = ~w33310;// level 16
assign po3127 = ~w33313;// level 17
assign po3128 = ~w33315;// level 27
assign po3129 = w33318;// level 5
assign po3130 = w33322;// level 11
assign po3131 = w33335;// level 15
assign po3132 = w33336;// level 12
assign po3133 = w33339;// level 5
assign po3134 = ~w33346;// level 17
assign po3135 = ~w33349;// level 17
assign po3136 = w33352;// level 5
assign po3137 = ~w33355;// level 17
assign po3138 = w33358;// level 4
assign po3139 = w33362;// level 5
assign po3140 = w33365;// level 5
assign po3141 = w33368;// level 5
assign po3142 = w33370;// level 6
assign po3143 = w33373;// level 15
assign po3144 = ~w33376;// level 17
assign po3145 = ~w33379;// level 17
assign po3146 = ~w33382;// level 17
assign po3147 = ~w33385;// level 17
assign po3148 = ~w33388;// level 17
assign po3149 = ~w33391;// level 17
assign po3150 = ~w33394;// level 17
assign po3151 = ~w33397;// level 17
assign po3152 = ~w33400;// level 17
assign po3153 = ~w33403;// level 17
assign po3154 = ~w33406;// level 17
assign po3155 = w33409;// level 5
assign po3156 = w33412;// level 5
assign po3157 = w33415;// level 5
assign po3158 = ~w33419;// level 17
assign po3159 = ~w33423;// level 17
assign po3160 = ~w33426;// level 17
assign po3161 = ~w33429;// level 17
assign po3162 = ~w33432;// level 16
assign po3163 = ~w33435;// level 16
assign po3164 = ~w33438;// level 17
assign po3165 = ~w33441;// level 17
assign po3166 = ~w33444;// level 16
assign po3167 = ~w33447;// level 17
assign po3168 = ~w33450;// level 15
assign po3169 = ~w33453;// level 16
assign po3170 = ~w33456;// level 16
assign po3171 = ~w33459;// level 16
assign po3172 = ~w33462;// level 16
assign po3173 = ~w33465;// level 17
assign po3174 = ~w33468;// level 17
assign po3175 = w33471;// level 5
assign po3176 = w33474;// level 5
assign po3177 = w33478;// level 5
assign po3178 = w33482;// level 5
assign po3179 = ~w33485;// level 17
assign po3180 = ~w33488;// level 18
assign po3181 = ~w33491;// level 18
assign po3182 = ~w33494;// level 18
assign po3183 = ~w33497;// level 18
assign po3184 = ~w33500;// level 18
assign po3185 = ~w33503;// level 17
assign po3186 = ~w33506;// level 17
assign po3187 = ~w33509;// level 17
assign po3188 = ~w33512;// level 18
assign po3189 = ~w33515;// level 18
assign po3190 = ~w33518;// level 18
assign po3191 = ~w33521;// level 18
assign po3192 = ~w33524;// level 18
assign po3193 = ~w33527;// level 18
assign po3194 = ~w33530;// level 18
assign po3195 = ~w33533;// level 17
assign po3196 = ~w33536;// level 17
assign po3197 = ~w33539;// level 16
assign po3198 = w33542;// level 5
assign po3199 = w33545;// level 5
assign po3200 = w33548;// level 5
assign po3201 = w33551;// level 5
assign po3202 = w33554;// level 5
assign po3203 = w33557;// level 5
assign po3204 = w33560;// level 5
assign po3205 = w33564;// level 5
assign po3206 = ~w33567;// level 17
assign po3207 = ~w33570;// level 17
assign po3208 = ~w33573;// level 16
assign po3209 = ~w33576;// level 17
assign po3210 = ~w33579;// level 16
assign po3211 = ~w33582;// level 17
assign po3212 = ~w33585;// level 15
assign po3213 = ~w33588;// level 16
assign po3214 = ~w33591;// level 16
assign po3215 = ~w33594;// level 17
assign po3216 = w33597;// level 5
assign po3217 = w33600;// level 5
assign po3218 = w33603;// level 5
assign po3219 = w33606;// level 5
assign po3220 = w33609;// level 5
assign po3221 = w33612;// level 5
assign po3222 = w33615;// level 5
assign po3223 = w33618;// level 5
assign po3224 = w33621;// level 5
assign po3225 = w33624;// level 5
assign po3226 = w33627;// level 5
assign po3227 = w33630;// level 5
assign po3228 = w33633;// level 5
assign po3229 = w33637;// level 11
assign po3230 = w33641;// level 11
assign po3231 = w33645;// level 11
assign po3232 = ~w33648;// level 16
assign po3233 = w33651;// level 5
assign po3234 = ~w33654;// level 18
assign po3235 = ~w33657;// level 18
assign po3236 = ~w33660;// level 18
assign po3237 = ~w33663;// level 18
assign po3238 = ~w33666;// level 18
assign po3239 = ~w33669;// level 18
assign po3240 = ~w33672;// level 18
assign po3241 = ~w33675;// level 18
assign po3242 = ~w33678;// level 17
assign po3243 = ~w33681;// level 17
assign po3244 = ~w33684;// level 18
assign po3245 = ~w33687;// level 18
assign po3246 = ~w33690;// level 18
assign po3247 = ~w33693;// level 16
assign po3248 = w33696;// level 5
assign po3249 = ~w33699;// level 17
assign po3250 = ~w33702;// level 17
assign po3251 = ~w33705;// level 17
assign po3252 = ~w33708;// level 16
assign po3253 = ~w33711;// level 17
assign po3254 = ~w33714;// level 16
assign po3255 = ~w33717;// level 17
assign po3256 = ~w33720;// level 17
assign po3257 = ~w33723;// level 17
assign po3258 = ~w33726;// level 17
assign po3259 = ~w33729;// level 16
assign po3260 = ~w33732;// level 16
assign po3261 = ~w33735;// level 17
assign po3262 = ~w33738;// level 17
assign po3263 = ~w33741;// level 16
assign po3264 = ~w33744;// level 15
assign po3265 = ~w33747;// level 16
assign po3266 = ~w33750;// level 16
assign po3267 = ~w33753;// level 16
assign po3268 = ~w33756;// level 17
assign po3269 = w33761;// level 12
assign po3270 = w33765;// level 12
assign po3271 = ~w33768;// level 30
assign po3272 = w33771;// level 5
assign po3273 = w33774;// level 5
assign po3274 = w33777;// level 5
assign po3275 = w33780;// level 5
assign po3276 = w33783;// level 5
assign po3277 = w33786;// level 5
assign po3278 = ~w33788;// level 28
assign po3279 = ~w33790;// level 28
assign po3280 = ~w33792;// level 28
assign po3281 = ~w33794;// level 28
assign po3282 = ~w33796;// level 27
assign po3283 = ~w33798;// level 28
assign po3284 = w33801;// level 28
assign po3285 = ~w33803;// level 28
assign po3286 = ~w33805;// level 27
assign po3287 = ~w33808;// level 16
assign po3288 = w33811;// level 5
assign po3289 = w33814;// level 5
assign po3290 = w33817;// level 5
assign po3291 = w33820;// level 5
assign po3292 = ~w33825;// level 16
assign po3293 = ~w33829;// level 16
assign po3294 = ~w33833;// level 16
assign po3295 = w33836;// level 5
assign po3296 = ~w33840;// level 16
assign po3297 = ~w33843;// level 16
assign po3298 = ~w33846;// level 16
assign po3299 = ~w33849;// level 16
assign po3300 = w33852;// level 11
assign po3301 = ~w33856;// level 11
assign po3302 = w33859;// level 5
assign po3303 = ~w33863;// level 8
assign po3304 = ~w33866;// level 16
assign po3305 = ~w33869;// level 15
assign po3306 = ~w33872;// level 16
assign po3307 = ~w33875;// level 16
assign po3308 = ~w33878;// level 16
assign po3309 = w33881;// level 5
assign po3310 = w27429;// level 5
assign po3311 = w28388;// level 6
assign po3312 = w33884;// level 5
assign po3313 = w33887;// level 5
assign po3314 = w33890;// level 5
assign po3315 = w33893;// level 5
assign po3316 = w33896;// level 5
assign po3317 = w33899;// level 5
assign po3318 = w33902;// level 5
assign po3319 = w33905;// level 5
assign po3320 = w33908;// level 5
assign po3321 = w33911;// level 5
assign po3322 = w33914;// level 5
assign po3323 = w33917;// level 5
assign po3324 = w33920;// level 5
assign po3325 = w33923;// level 5
assign po3326 = w33926;// level 5
assign po3327 = w33929;// level 5
assign po3328 = w33932;// level 5
assign po3329 = w33935;// level 5
assign po3330 = w33938;// level 5
assign po3331 = w33941;// level 5
assign po3332 = w33944;// level 5
assign po3333 = w33947;// level 5
assign po3334 = w33950;// level 5
assign po3335 = w33953;// level 5
assign po3336 = w33956;// level 5
assign po3337 = w33959;// level 5
assign po3338 = w33962;// level 5
assign po3339 = w33965;// level 5
assign po3340 = w33968;// level 5
assign po3341 = w33971;// level 5
assign po3342 = w33974;// level 5
assign po3343 = w33977;// level 5
assign po3344 = w33980;// level 5
assign po3345 = w33983;// level 5
assign po3346 = w33986;// level 5
assign po3347 = w33989;// level 5
assign po3348 = w33992;// level 5
assign po3349 = w33995;// level 5
assign po3350 = w33998;// level 5
assign po3351 = w34001;// level 5
assign po3352 = w34004;// level 5
assign po3353 = w34007;// level 5
assign po3354 = w34010;// level 5
assign po3355 = w34013;// level 5
assign po3356 = w34016;// level 5
assign po3357 = w34019;// level 5
assign po3358 = w34022;// level 5
assign po3359 = w34025;// level 5
assign po3360 = w34028;// level 5
assign po3361 = w34031;// level 5
assign po3362 = w34034;// level 5
assign po3363 = w34037;// level 5
assign po3364 = w34040;// level 5
assign po3365 = w34043;// level 5
assign po3366 = w34046;// level 5
assign po3367 = w34049;// level 5
assign po3368 = w34052;// level 5
assign po3369 = w34055;// level 5
assign po3370 = w34058;// level 5
assign po3371 = w34061;// level 5
assign po3372 = w34064;// level 5
assign po3373 = ~w34067;// level 5
assign po3374 = w34070;// level 5
assign po3375 = w34073;// level 5
assign po3376 = w34076;// level 5
assign po3377 = ~w34079;// level 17
assign po3378 = w34082;// level 5
assign po3379 = w34085;// level 5
assign po3380 = w34088;// level 5
assign po3381 = ~w34091;// level 16
assign po3382 = w34094;// level 5
assign po3383 = w34097;// level 11
assign po3384 = w34100;// level 5
assign po3385 = w34103;// level 5
assign po3386 = ~w34107;// level 16
assign po3387 = w34110;// level 5
assign po3388 = w34113;// level 5
assign po3389 = w34116;// level 5
assign po3390 = w34119;// level 5
assign po3391 = w34122;// level 5
assign po3392 = ~w34125;// level 16
assign po3393 = ~w34128;// level 17
assign po3394 = w34132;// level 12
assign po3395 = w34135;// level 5
assign po3396 = w34138;// level 5
assign po3397 = ~w34141;// level 16
assign po3398 = w34144;// level 5
assign po3399 = w34147;// level 5
assign po3400 = w34150;// level 5
assign po3401 = w34153;// level 5
assign po3402 = ~w34156;// level 16
assign po3403 = w34159;// level 5
assign po3404 = w34162;// level 4
assign po3405 = w34165;// level 5
assign po3406 = w34168;// level 5
assign po3407 = w34171;// level 5
assign po3408 = w34174;// level 5
assign po3409 = ~w34177;// level 16
assign po3410 = w34180;// level 5
assign po3411 = ~w34182;// level 28
assign po3412 = w34185;// level 5
assign po3413 = w34188;// level 5
assign po3414 = ~w34190;// level 28
assign po3415 = ~w34193;// level 15
assign po3416 = pi3527;// level 0
assign po3417 = w34196;// level 5
assign po3418 = ~w34199;// level 16
assign po3419 = ~w34202;// level 16
assign po3420 = ~w34205;// level 16
assign po3421 = ~w34208;// level 8
assign po3422 = w34211;// level 5
assign po3423 = ~w34214;// level 8
assign po3424 = ~w34217;// level 8
assign po3425 = ~w34220;// level 8
assign po3426 = ~w34223;// level 16
assign po3427 = w34226;// level 5
assign po3428 = ~w34229;// level 8
assign po3429 = w34232;// level 5
assign po3430 = ~w34235;// level 8
assign po3431 = ~w34238;// level 8
assign po3432 = ~w34241;// level 17
assign po3433 = ~w34248;// level 11
assign po3434 = ~w34252;// level 11
assign po3435 = ~w34256;// level 11
assign po3436 = ~w34260;// level 11
assign po3437 = ~w34266;// level 11
assign po3438 = ~w34270;// level 16
assign po3439 = ~w34274;// level 20
assign po3440 = ~w34276;// level 21
assign po3441 = ~w34279;// level 16
assign po3442 = ~w34282;// level 17
assign po3443 = ~w34286;// level 11
assign po3444 = ~w34289;// level 17
assign po3445 = ~w34292;// level 17
assign po3446 = ~w34296;// level 17
assign po3447 = ~w34299;// level 17
assign po3448 = ~w29348;// level 10
assign po3449 = ~w34302;// level 10
assign po3450 = ~w34305;// level 17
assign po3451 = ~w34308;// level 17
assign po3452 = ~w34311;// level 16
assign po3453 = ~w34314;// level 16
assign po3454 = ~w34318;// level 11
assign po3455 = w34319;// level 12
assign po3456 = ~w34342;// level 5
assign po3457 = ~w34344;// level 11
assign po3458 = ~w34348;// level 11
assign po3459 = ~w34351;// level 17
assign po3460 = ~pi3300;// level 0
assign po3461 = pi3254;// level 0
assign po3462 = ~w34354;// level 16
assign po3463 = ~pi3303;// level 0
assign po3464 = pi3205;// level 0
assign po3465 = ~w34357;// level 11
assign po3466 = ~w34359;// level 20
assign po3467 = w34360;// level 4
assign po3468 = ~w34366;// level 10
assign po3469 = ~w34369;// level 17
assign po3470 = ~w34372;// level 17
assign po3471 = ~w34375;// level 18
assign po3472 = ~w34378;// level 18
assign po3473 = ~w34381;// level 18
assign po3474 = ~w34384;// level 18
assign po3475 = ~w34387;// level 18
assign po3476 = ~w34390;// level 18
assign po3477 = ~w34393;// level 18
assign po3478 = ~w34396;// level 17
assign po3479 = ~w34399;// level 16
assign po3480 = ~w34402;// level 18
assign po3481 = ~w34405;// level 18
assign po3482 = ~w34408;// level 18
assign po3483 = ~w34411;// level 18
assign po3484 = ~w34414;// level 18
assign po3485 = ~w34417;// level 18
assign po3486 = ~w34420;// level 16
assign po3487 = ~w34423;// level 17
assign po3488 = ~w34426;// level 17
assign po3489 = ~w34429;// level 17
assign po3490 = ~w34432;// level 16
assign po3491 = ~w34435;// level 15
assign po3492 = ~w34438;// level 16
assign po3493 = ~w34441;// level 16
assign po3494 = ~w34444;// level 16
assign po3495 = ~w34447;// level 16
assign po3496 = ~w34450;// level 17
assign po3497 = ~w34453;// level 17
assign po3498 = ~w34456;// level 16
assign po3499 = ~w34459;// level 16
assign po3500 = ~w34462;// level 17
assign po3501 = ~w34465;// level 17
assign po3502 = ~w34468;// level 15
assign po3503 = ~w34471;// level 16
assign po3504 = ~w34474;// level 16
assign po3505 = ~w34477;// level 17
assign po3506 = ~w34481;// level 16
assign po3507 = ~w34485;// level 11
assign po3508 = w34487;// level 4
assign po3509 = ~w34491;// level 16
assign po3510 = ~w34494;// level 21
assign po3511 = ~w34497;// level 20
assign po3512 = ~w34501;// level 11
assign po3513 = ~w34505;// level 11
assign po3514 = ~w34509;// level 11
assign po3515 = ~w34513;// level 11
assign po3516 = ~w34517;// level 11
assign po3517 = ~w34521;// level 11
assign po3518 = ~w34525;// level 11
assign po3519 = w34528;// level 14
assign po3520 = w34530;// level 4
assign po3521 = ~w34533;// level 18
assign po3522 = ~w34536;// level 17
assign po3523 = ~w34540;// level 12
assign po3524 = ~w34542;// level 13
assign po3525 = w34544;// level 4
assign po3526 = ~w34550;// level 11
assign po3527 = ~w34556;// level 11
assign po3528 = ~w34562;// level 11
assign po3529 = ~w34568;// level 11
assign po3530 = ~w34571;// level 21
assign po3531 = ~w34573;// level 20
assign po3532 = ~w34577;// level 3
assign po3533 = ~w34581;// level 3
assign po3534 = ~w34585;// level 3
assign po3535 = ~w34592;// level 22
assign po3536 = ~w34595;// level 20
assign po3537 = ~w34599;// level 16
assign po3538 = w34605;// level 6
assign po3539 = w34611;// level 6
assign po3540 = w34617;// level 6
assign po3541 = w34623;// level 6
assign po3542 = w34629;// level 6
assign po3543 = w34635;// level 6
assign po3544 = w34641;// level 6
assign po3545 = w34647;// level 6
assign po3546 = ~w34651;// level 16
assign po3547 = ~w34655;// level 16
assign po3548 = ~w34661;// level 11
assign po3549 = ~w34667;// level 11
assign po3550 = ~w34673;// level 11
assign po3551 = ~w34679;// level 11
assign po3552 = ~w34683;// level 3
assign po3553 = w34685;// level 10
assign po3554 = ~w34691;// level 11
assign po3555 = ~w34697;// level 11
assign po3556 = ~w34701;// level 11
assign po3557 = ~w34705;// level 16
assign po3558 = ~w34709;// level 16
assign po3559 = ~w34713;// level 16
assign po3560 = w34719;// level 6
assign po3561 = w34725;// level 6
assign po3562 = w34731;// level 6
assign po3563 = w34737;// level 6
assign po3564 = ~w34740;// level 10
assign po3565 = ~w34743;// level 11
assign po3566 = ~w34748;// level 4
assign po3567 = w34750;// level 5
assign po3568 = w34754;// level 11
assign po3569 = w20918;// level 7
assign po3570 = ~w15388;// level 9
assign po3571 = w21417;// level 7
assign po3572 = w34759;// level 3
assign po3573 = w34762;// level 14
assign po3574 = w32027;// level 2
assign po3575 = ~w34765;// level 4
assign po3576 = ~w34766;// level 20
assign po3577 = ~w34767;// level 20
assign po3578 = w34770;// level 14
assign po3579 = w34773;// level 14
assign po3580 = w34776;// level 14
assign po3581 = w34779;// level 14
assign po3582 = w34782;// level 14
assign po3583 = w34785;// level 14
assign po3584 = w34788;// level 14
assign po3585 = w34791;// level 14
assign po3586 = ~w34794;// level 4
assign po3587 = w34798;// level 11
assign po3588 = ~w34801;// level 11
assign po3589 = ~w34804;// level 11
assign po3590 = w34805;// level 1
assign po3591 = ~w34809;// level 15
assign po3592 = ~w34812;// level 4
assign po3593 = w34815;// level 14
assign po3594 = w34818;// level 14
assign po3595 = w34821;// level 14
assign po3596 = w34824;// level 14
assign po3597 = w34827;// level 14
assign po3598 = w34830;// level 14
assign po3599 = w34831;// level 1
assign po3600 = ~w34835;// level 15
assign po3601 = w34838;// level 14
assign po3602 = w34841;// level 14
assign po3603 = w34845;// level 14
assign po3604 = w34848;// level 14
assign po3605 = w34851;// level 14
assign po3606 = w34854;// level 14
assign po3607 = ~w34857;// level 11
assign po3608 = w34860;// level 14
assign po3609 = w34863;// level 14
assign po3610 = w34866;// level 14
assign po3611 = w34869;// level 14
assign po3612 = w34871;// level 4
assign po3613 = ~w34875;// level 20
assign po3614 = ~w34878;// level 10
assign po3615 = ~w34882;// level 16
assign po3616 = ~w165;// level 11
assign po3617 = w34889;// level 15
assign po3618 = w34895;// level 15
assign po3619 = w34901;// level 15
assign po3620 = w34907;// level 15
assign po3621 = w34911;// level 11
assign po3622 = pi3418;// level 0
assign po3623 = ~w34913;// level 4
assign po3624 = w34914;// level 2
assign po3625 = pi3431;// level 0
assign po3626 = ~w34917;// level 3
assign po3627 = w6682;// level 5
assign po3628 = ~w34920;// level 10
assign po3629 = w34926;// level 15
assign po3630 = w34932;// level 15
assign po3631 = w34938;// level 15
assign po3632 = ~w34946;// level 16
assign po3633 = w34952;// level 15
assign po3634 = w34958;// level 15
assign po3635 = w34964;// level 15
assign po3636 = ~w34970;// level 14
assign po3637 = ~w34976;// level 14
assign po3638 = w34982;// level 15
assign po3639 = w34988;// level 15
assign po3640 = w34991;// level 4
assign po3641 = w34994;// level 4
assign po3642 = w34997;// level 4
assign po3643 = w35000;// level 4
assign po3644 = w35003;// level 4
assign po3645 = ~w113;// level 6
assign po3646 = ~w177;// level 6
assign po3647 = ~w33326;// level 10
assign po3648 = ~w35005;// level 4
assign po3649 = w35009;// level 11
assign po3650 = ~w35011;// level 4
assign po3651 = ~w35014;// level 16
assign po3652 = ~w35018;// level 11
assign po3653 = ~w35020;// level 10
assign po3654 = ~w35024;// level 11
assign po3655 = ~w35027;// level 11
assign po3656 = ~w35029;// level 4
assign po3657 = ~w35031;// level 4
assign po3658 = ~w35033;// level 4
assign po3659 = ~w35035;// level 4
assign po3660 = ~w35036;// level 1
assign po3661 = ~w35038;// level 4
assign po3662 = ~w35040;// level 4
assign po3663 = w35043;// level 4
assign po3664 = ~w35045;// level 4
assign po3665 = ~w35047;// level 4
assign po3666 = w35050;// level 14
assign po3667 = ~w35052;// level 11
assign po3668 = w35055;// level 4
assign po3669 = w35058;// level 4
assign po3670 = ~w35061;// level 11
assign po3671 = w35064;// level 4
assign po3672 = w35067;// level 4
assign po3673 = ~w35073;// level 14
assign po3674 = w35076;// level 4
assign po3675 = ~w35079;// level 11
assign po3676 = ~w35082;// level 11
assign po3677 = ~w35085;// level 11
assign po3678 = ~w35088;// level 11
assign po3679 = ~w35090;// level 4
assign po3680 = w35093;// level 4
assign po3681 = w35099;// level 15
assign po3682 = w35101;// level 29
assign po3683 = ~w35104;// level 16
assign po3684 = ~w35107;// level 16
assign po3685 = ~w19953;// level 4
assign po3686 = w35109;// level 30
assign po3687 = w35110;// level 30
assign po3688 = w35111;// level 29
assign po3689 = w35114;// level 28
assign po3690 = ~w35117;// level 10
assign po3691 = w35119;// level 28
assign po3692 = w35121;// level 28
assign po3693 = ~w35124;// level 10
assign po3694 = w35128;// level 11
assign po3695 = w35129;// level 14
assign po3696 = w35130;// level 15
assign po3697 = w35131;// level 15
assign po3698 = w35132;// level 14
assign po3699 = ~w35135;// level 3
assign po3700 = ~w35138;// level 3
assign po3701 = ~w35141;// level 10
assign po3702 = w35142;// level 28
assign po3703 = w35144;// level 28
assign po3704 = w35145;// level 28
assign po3705 = w35146;// level 3
assign po3706 = w35148;// level 2
assign po3707 = w35149;// level 28
assign po3708 = w35150;// level 28
assign po3709 = w35151;// level 29
assign po3710 = w35152;// level 29
assign po3711 = w35153;// level 29
assign po3712 = w35155;// level 32
assign po3713 = ~w35156;// level 1
assign po3714 = ~w35158;// level 10
assign po3715 = ~w35161;// level 10
assign po3716 = w35163;// level 10
assign po3717 = ~w35165;// level 10
assign po3718 = ~w35167;// level 10
assign po3719 = pi3555;// level 0
assign po3720 = w35168;// level 9
assign po3721 = ~w35171;// level 10
assign po3722 = ~w35173;// level 4
assign po3723 = ~w35175;// level 10
assign po3724 = w35176;// level 29
assign po3725 = ~w35179;// level 9
assign po3726 = ~w35182;// level 9
assign po3727 = ~w35185;// level 9
assign po3728 = ~w35188;// level 9
assign po3729 = ~w35191;// level 9
assign po3730 = ~w35194;// level 9
assign po3731 = ~w35197;// level 9
assign po3732 = w35198;// level 10
assign po3733 = ~w35201;// level 18
assign po3734 = ~w35203;// level 7
assign po3735 = pi1609;// level 0
assign po3736 = ~pi3382;// level 0
assign po3737 = ~w35206;// level 9
assign po3738 = w35210;// level 10
assign po3739 = ~w35213;// level 9
assign po3740 = ~w35216;// level 9
assign po3741 = ~w9;// level 4
assign po3742 = ~w35219;// level 2
assign po3743 = w32393;// level 2
assign po3744 = ~w35223;// level 4
assign po3745 = ~w25373;// level 1
assign po3746 = w34833;// level 13
assign po3747 = w35225;// level 8
assign po3748 = ~w35228;// level 9
assign po3749 = ~w35231;// level 9
assign po3750 = ~w35234;// level 9
assign po3751 = w35238;// level 12
assign po3752 = w35240;// level 9
assign po3753 = w35241;// level 5
assign po3754 = w35243;// level 19
assign po3755 = w35245;// level 9
assign po3756 = w35248;// level 9
assign po3757 = w35249;// level 9
assign po3758 = ~w35252;// level 9
assign po3759 = w34807;// level 13
assign po3760 = w35255;// level 23
assign po3761 = w9807;// level 23
assign po3762 = w35258;// level 23
assign po3763 = ~w35261;// level 10
assign po3764 = ~w35264;// level 10
assign po3765 = w9804;// level 23
assign po3766 = ~pi3472;// level 0
assign po3767 = ~pi3469;// level 0
assign po3768 = pi3507;// level 0
assign po3769 = w35266;// level 2
assign po3770 = ~pi3537;// level 0
assign po3771 = ~pi3536;// level 0
assign po3772 = pi0827;// level 0
assign po3773 = ~w35269;// level 2
assign po3774 = ~w35272;// level 2
assign po3775 = ~w35275;// level 2
assign po3776 = ~w35278;// level 2
assign po3777 = ~w35281;// level 24
assign po3778 = w35284;// level 23
assign po3779 = ~w35287;// level 10
assign po3780 = w35288;// level 8
assign po3781 = w35291;// level 23
assign po3782 = w35294;// level 23
assign po3783 = w35297;// level 23
assign po3784 = w9813;// level 23
assign po3785 = w9810;// level 23
assign po3786 = w35300;// level 23
assign po3787 = w35303;// level 23
assign po3788 = w9801;// level 23
assign po3789 = ~w35306;// level 15
assign po3790 = ~w35309;// level 2
assign po3791 = ~w35312;// level 2
assign po3792 = ~w35315;// level 2
assign po3793 = ~w35318;// level 2
assign po3794 = ~w35321;// level 2
assign po3795 = ~w35324;// level 2
assign po3796 = ~w35327;// level 2
assign po3797 = ~pi1882;// level 0
assign po3798 = ~w35330;// level 2
assign po3799 = ~w35333;// level 15
assign po3800 = ~pi2099;// level 0
assign po3801 = ~w35336;// level 15
assign po3802 = ~w35339;// level 2
assign po3803 = ~w35342;// level 2
assign po3804 = ~w35345;// level 2
assign po3805 = ~w35348;// level 2
assign po3806 = w35351;// level 23
assign po3807 = ~w35352;// level 6
assign po3808 = pi3549;// level 0
assign po3809 = w35354;// level 2
assign po3810 = ~pi3571;// level 0
assign po3811 = pi3531;// level 0
assign po3812 = pi3532;// level 0
assign po3813 = pi3533;// level 0
assign po3814 = pi3534;// level 0
assign po3815 = ~w35357;// level 24
assign po3816 = pi3544;// level 0
assign po3817 = ~w35360;// level 24
assign po3818 = ~w35363;// level 24
assign po3819 = pi3550;// level 0
assign po3820 = ~w35366;// level 24
assign po3821 = ~w35369;// level 24
assign po3822 = ~w35372;// level 24
assign po3823 = ~w35375;// level 24
assign po3824 = ~w35378;// level 24
assign po3825 = ~w35381;// level 24
assign po3826 = ~w35384;// level 24
assign po3827 = ~w35387;// level 24
assign po3828 = w35389;// level 8
assign po3829 = ~w35392;// level 24
assign po3830 = ~w9609;// level 9
assign po3831 = ~w342;// level 7
assign po3832 = w35393;// level 7
assign po3833 = w35394;// level 1
assign po3834 = ~w9352;// level 9
assign po3835 = ~w9304;// level 9
assign po3836 = ~w9186;// level 9
assign po3837 = ~w9126;// level 9
assign po3838 = ~w7101;// level 9
assign po3839 = ~w9669;// level 9
assign po3840 = ~w9556;// level 9
assign po3841 = w358;// level 8
assign po3842 = ~w9448;// level 9
assign po3843 = ~w9397;// level 9
assign po3844 = ~w9510;// level 9
assign po3845 = ~w7162;// level 9
assign po3846 = ~w9068;// level 9
assign po3847 = ~w9243;// level 9
assign po3848 = ~w932;// level 2
assign po3849 = ~w7173;// level 5
assign po3850 = w6677;// level 3
assign po3851 = ~w0;// level 1
assign po3852 = ~w28741;// level 7
assign po3853 = w10;// level 5
assign po3854 = pi3551;// level 0
assign po3855 = ~w926;// level 2
assign po3856 = ~pi0582;// level 0
assign po3857 = ~pi3660;// level 0
assign po3858 = ~pi3657;// level 0
assign po3859 = ~pi3658;// level 0
assign po3860 = ~pi3659;// level 0
assign po3861 = ~pi0581;// level 0
assign po3862 = ~pi3661;// level 0
assign po3863 = ~pi3656;// level 0
assign po3864 = ~pi3214;// level 0
assign po3865 = ~pi1596;// level 0
assign po3866 = ~pi3200;// level 0
assign po3867 = ~pi3213;// level 0
assign po3868 = ~pi3232;// level 0
assign po3869 = ~pi3212;// level 0
assign po3870 = ~pi3662;// level 0
assign po3871 = w941;// level 2
assign po3872 = w923;// level 4
assign po3873 = ~w323;// level 2
assign po3874 = ~w915;// level 5
assign po3875 = ~pi2399;// level 0
assign po3876 = ~pi2387;// level 0
assign po3877 = ~pi3098;// level 0
assign po3878 = ~w919;// level 3
assign po3879 = w28389;// level 13
assign po3880 = ~w10741;// level 1
assign po3881 = pi2385;// level 0
assign po3882 = w17480;// level 2
assign po3883 = pi1931;// level 0
assign po3884 = pi2111;// level 0
assign po3885 = pi0939;// level 0
assign po3886 = pi3645;// level 0
assign po3887 = pi3679;// level 0
assign po3888 = pi3674;// level 0
assign po3889 = pi3675;// level 0
assign po3890 = pi3673;// level 0
assign po3891 = pi3672;// level 0
assign po3892 = pi0565;// level 0
assign po3893 = w7177;// level 1
assign po3894 = w35395;// level 7
assign po3895 = pi3591;// level 0
assign po3896 = w27430;// level 13
assign po3897 = ~w17481;// level 3
assign po3898 = pi3585;// level 0
assign po3899 = pi0936;// level 0
assign po3900 = ~w35398;// level 15
assign po3901 = ~w35401;// level 15
assign po3902 = ~w35404;// level 15
assign po3903 = ~w35407;// level 15
assign po3904 = ~w35410;// level 15
assign po3905 = ~w35413;// level 15
assign po3906 = ~w35416;// level 15
assign po3907 = ~w35419;// level 15
assign po3908 = ~w35422;// level 15
assign po3909 = ~w35425;// level 15
assign po3910 = ~w35428;// level 15
assign po3911 = ~w35431;// level 15
assign po3912 = ~w35434;// level 15
assign po3913 = ~w35437;// level 15
assign po3914 = ~w35440;// level 15
assign po3915 = ~w35443;// level 15
assign po3916 = ~w35446;// level 15
assign po3917 = ~w35449;// level 15
assign po3918 = ~w35452;// level 15
assign po3919 = ~w35455;// level 15
assign po3920 = ~w35458;// level 15
assign po3921 = ~w35461;// level 15
assign po3922 = ~w35464;// level 15
assign po3923 = ~w35467;// level 15
assign po3924 = ~w35470;// level 15
assign po3925 = ~w35473;// level 15
assign po3926 = w35474;// level 14
assign po3927 = ~w35477;// level 15
assign po3928 = ~w35490;// level 16
assign po3929 = w35498;// level 16
assign po3930 = w35502;// level 15
assign po3931 = w35503;// level 14
assign po3932 = w35483;// level 14
assign po3933 = ~w35488;// level 14
assign po3934 = ~w35069;// level 13
assign po3935 = pi3629;// level 0
assign po3936 = pi3630;// level 0
assign po3937 = w28372;// level 8
assign po3938 = w35510;// level 11
assign po3939 = w24175;// level 5
assign po3940 = ~w35511;// level 4
assign po3941 = w35531;// level 8
assign po3942 = pi3637;// level 0
assign po3943 = w28370;// level 7
assign po3944 = pi3640;// level 0
assign po3945 = w27413;// level 8
assign po3946 = ~w341;// level 7
assign po3947 = ~w35506;// level 2
assign po3948 = ~w6681;// level 4
assign po3949 = w35532;// level 1
assign po3950 = w27411;// level 7
assign po3951 = ~pi3676;// level 0
assign po3952 = pi0853;// level 0
endmodule
