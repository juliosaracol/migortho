module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129, po130, po131, po132, po133, po134, po135, po136, po137, po138, po139, po140, po141, po142, po143, po144, po145, po146, po147, po148, po149, po150, po151, po152, po153, po154, po155, po156, po157, po158, po159, po160, po161, po162, po163, po164, po165, po166, po167, po168, po169, po170, po171, po172, po173, po174, po175, po176, po177, po178, po179, po180, po181, po182, po183, po184, po185, po186, po187, po188, po189, po190, po191, po192, po193, po194, po195, po196, po197, po198, po199, po200, po201, po202, po203, po204, po205, po206, po207, po208, po209, po210, po211, po212, po213, po214, po215, po216, po217, po218, po219, po220, po221, po222, po223, po224, po225, po226, po227, po228, po229, po230, po231, po232, po233, po234, po235, po236, po237, po238, po239, po240, po241, po242, po243, po244, po245, po246, po247, po248, po249, po250, po251, po252, po253, po254, po255, po256, po257;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452;
assign w0 = pi066 & pi081;
assign w1 = pi068 & w0;
assign w2 = w0 & w2073;
assign w3 = ~pi066 & ~pi068;
assign w4 = pi069 & pi081;
assign w5 = w3 & ~w4;
assign w6 = ~w2 & ~w5;
assign w7 = ~pi069 & ~pi081;
assign w8 = w3 & w7;
assign w9 = pi192 & w8;
assign w10 = w8 & w2074;
assign w11 = (pi064 & ~w8) | (pi064 & w2201) | (~w8 & w2201);
assign w12 = ~w10 & ~w11;
assign w13 = w6 & ~w12;
assign w14 = (pi037 & ~w8) | (pi037 & w2075) | (~w8 & w2075);
assign w15 = w8 & w2076;
assign w16 = ~w14 & ~w15;
assign w17 = ~w6 & ~w16;
assign w18 = ~w13 & ~w17;
assign w19 = ~pi193 & ~w18;
assign w20 = ~w6 & ~w7;
assign w21 = (pi048 & ~w8) | (pi048 & w2077) | (~w8 & w2077);
assign w22 = w8 & w2078;
assign w23 = ~w21 & ~w22;
assign w24 = w20 & ~w23;
assign w25 = (pi065 & ~w8) | (pi065 & w2079) | (~w8 & w2079);
assign w26 = w8 & w2080;
assign w27 = ~w25 & ~w26;
assign w28 = w8 & ~w27;
assign w29 = (pi045 & ~w8) | (pi045 & w2081) | (~w8 & w2081);
assign w30 = w8 & w2082;
assign w31 = ~w29 & ~w30;
assign w32 = ~w24 & ~w28;
assign w33 = (pi193 & ~w32) | (pi193 & w2220) | (~w32 & w2220);
assign w34 = ~w19 & ~w33;
assign w35 = pi021 & ~w9;
assign w36 = pi219 & w9;
assign w37 = ~w35 & ~w36;
assign w38 = ~w34 & w37;
assign w39 = w34 & ~w37;
assign w40 = ~w38 & ~w39;
assign w41 = w8 & w2083;
assign w42 = (pi078 & ~w8) | (pi078 & w2084) | (~w8 & w2084);
assign w43 = ~w41 & ~w42;
assign w44 = w6 & ~w43;
assign w45 = w8 & w2085;
assign w46 = ~pi192 & w8;
assign w47 = w8 & w2175;
assign w48 = (pi039 & ~w8) | (pi039 & w2086) | (~w8 & w2086);
assign w49 = w8 & w2087;
assign w50 = ~w48 & ~w49;
assign w51 = w20 & ~w50;
assign w52 = (pi193 & ~w8) | (pi193 & w2221) | (~w8 & w2221);
assign w53 = ~w47 & w52;
assign w54 = ~w44 & w53;
assign w55 = ~w51 & w54;
assign w56 = w8 & w2088;
assign w57 = (pi083 & ~w8) | (pi083 & w2089) | (~w8 & w2089);
assign w58 = ~w56 & ~w57;
assign w59 = w6 & ~w58;
assign w60 = (pi059 & ~w8) | (pi059 & w2090) | (~w8 & w2090);
assign w61 = w8 & w2091;
assign w62 = ~w60 & ~w61;
assign w63 = ~w6 & ~w62;
assign w64 = (~pi193 & w58) | (~pi193 & w2178) | (w58 & w2178);
assign w65 = ~w63 & w64;
assign w66 = ~w55 & ~w65;
assign w67 = pi007 & ~w9;
assign w68 = pi253 & w9;
assign w69 = ~w67 & ~w68;
assign w70 = ~w55 & w2222;
assign w71 = (~w69 & w55) | (~w69 & w2223) | (w55 & w2223);
assign w72 = ~w70 & ~w71;
assign w73 = w8 & w2092;
assign w74 = (pi074 & ~w8) | (pi074 & w2093) | (~w8 & w2093);
assign w75 = ~w73 & ~w74;
assign w76 = w6 & ~w75;
assign w77 = w8 & w2094;
assign w78 = w8 & w2171;
assign w79 = (pi041 & ~w8) | (pi041 & w2095) | (~w8 & w2095);
assign w80 = w8 & w2096;
assign w81 = ~w79 & ~w80;
assign w82 = w20 & ~w81;
assign w83 = (pi193 & ~w8) | (pi193 & w2224) | (~w8 & w2224);
assign w84 = ~w78 & w83;
assign w85 = ~w76 & w84;
assign w86 = ~w82 & w85;
assign w87 = w8 & w2097;
assign w88 = (pi076 & ~w8) | (pi076 & w2098) | (~w8 & w2098);
assign w89 = ~w87 & ~w88;
assign w90 = w6 & ~w89;
assign w91 = w8 & w2099;
assign w92 = (pi091 & ~w8) | (pi091 & w2100) | (~w8 & w2100);
assign w93 = ~w91 & ~w92;
assign w94 = ~w6 & ~w93;
assign w95 = (~pi193 & w89) | (~pi193 & w2178) | (w89 & w2178);
assign w96 = ~w94 & w95;
assign w97 = ~w86 & ~w96;
assign w98 = pi026 & ~w9;
assign w99 = pi203 & w9;
assign w100 = ~w98 & ~w99;
assign w101 = ~w86 & w2225;
assign w102 = (~w100 & w86) | (~w100 & w2226) | (w86 & w2226);
assign w103 = ~w101 & ~w102;
assign w104 = ~w72 & w103;
assign w105 = w72 & ~w103;
assign w106 = ~w104 & ~w105;
assign w107 = (pi047 & ~w8) | (pi047 & w2101) | (~w8 & w2101);
assign w108 = w8 & w2102;
assign w109 = ~w107 & ~w108;
assign w110 = w20 & ~w109;
assign w111 = (pi061 & ~w8) | (pi061 & w2103) | (~w8 & w2103);
assign w112 = w8 & w2104;
assign w113 = ~w111 & ~w112;
assign w114 = ~w6 & ~w113;
assign w115 = w7 & w114;
assign w116 = (pi035 & ~w8) | (pi035 & w2105) | (~w8 & w2105);
assign w117 = w8 & w2106;
assign w118 = ~w116 & ~w117;
assign w119 = w6 & ~w118;
assign w120 = pi193 & ~w110;
assign w121 = ~w119 & w120;
assign w122 = ~w115 & w121;
assign w123 = w8 & w2107;
assign w124 = (pi075 & ~w8) | (pi075 & w2181) | (~w8 & w2181);
assign w125 = ~w123 & ~w124;
assign w126 = w6 & ~w125;
assign w127 = (pi053 & ~w8) | (pi053 & w2108) | (~w8 & w2108);
assign w128 = w8 & w2109;
assign w129 = ~w127 & ~w128;
assign w130 = ~w6 & ~w129;
assign w131 = ~pi193 & ~w126;
assign w132 = ~w130 & w131;
assign w133 = ~w122 & ~w132;
assign w134 = pi029 & ~w9;
assign w135 = pi211 & w9;
assign w136 = ~w134 & ~w135;
assign w137 = ~w122 & w2227;
assign w138 = (~w136 & w122) | (~w136 & w2228) | (w122 & w2228);
assign w139 = ~w137 & ~w138;
assign w140 = ~w105 & w139;
assign w141 = (pi072 & ~w8) | (pi072 & w2110) | (~w8 & w2110);
assign w142 = w8 & w2111;
assign w143 = ~w141 & ~w142;
assign w144 = ~w6 & ~w143;
assign w145 = (pi077 & ~w8) | (pi077 & w2112) | (~w8 & w2112);
assign w146 = w8 & w2113;
assign w147 = ~w145 & ~w146;
assign w148 = w6 & ~w147;
assign w149 = ~w144 & ~w148;
assign w150 = ~pi193 & ~w149;
assign w151 = (pi092 & ~w8) | (pi092 & w2114) | (~w8 & w2114);
assign w152 = w8 & w2115;
assign w153 = ~w151 & ~w152;
assign w154 = ~w6 & ~w153;
assign w155 = ~w153 & w2229;
assign w156 = (pi054 & ~w8) | (pi054 & w2116) | (~w8 & w2116);
assign w157 = w8 & w2117;
assign w158 = ~w156 & ~w157;
assign w159 = w6 & ~w158;
assign w160 = (pi042 & ~w8) | (pi042 & w2118) | (~w8 & w2118);
assign w161 = w8 & w2119;
assign w162 = ~w160 & ~w161;
assign w163 = w20 & ~w162;
assign w164 = ~w159 & ~w163;
assign w165 = (pi193 & ~w164) | (pi193 & w2230) | (~w164 & w2230);
assign w166 = ~w150 & ~w165;
assign w167 = pi017 & ~w9;
assign w168 = pi195 & w9;
assign w169 = ~w167 & ~w168;
assign w170 = ~w166 & w169;
assign w171 = w166 & ~w169;
assign w172 = ~w170 & ~w171;
assign w173 = ~w140 & ~w172;
assign w174 = ~w106 & w173;
assign w175 = w72 & w172;
assign w176 = ~w40 & w139;
assign w177 = w175 & ~w176;
assign w178 = (~w40 & w174) | (~w40 & w2293) | (w174 & w2293);
assign w179 = ~w139 & w172;
assign w180 = ~w106 & ~w176;
assign w181 = (~w180 & w178) | (~w180 & w2378) | (w178 & w2378);
assign w182 = w6 & ~w109;
assign w183 = ~w6 & ~w118;
assign w184 = ~w182 & ~w183;
assign w185 = ~pi193 & ~w184;
assign w186 = (pi040 & ~w8) | (pi040 & w2231) | (~w8 & w2231);
assign w187 = w8 & w2232;
assign w188 = ~w186 & ~w187;
assign w189 = ~w6 & ~w188;
assign w190 = w7 & w189;
assign w191 = w8 & w2120;
assign w192 = (pi058 & ~w8) | (pi058 & w2247) | (~w8 & w2247);
assign w193 = ~w191 & ~w192;
assign w194 = w20 & ~w193;
assign w195 = ~w148 & ~w194;
assign w196 = ~w190 & w195;
assign w197 = pi193 & ~w196;
assign w198 = ~w185 & ~w197;
assign w199 = pi020 & ~w9;
assign w200 = pi227 & w9;
assign w201 = ~w199 & ~w200;
assign w202 = ~w198 & w201;
assign w203 = w198 & ~w201;
assign w204 = ~w202 & ~w203;
assign w205 = w40 & ~w204;
assign w206 = w72 & ~w172;
assign w207 = w106 & ~w206;
assign w208 = ~w172 & w207;
assign w209 = w205 & w208;
assign w210 = w72 & w103;
assign w211 = w139 & ~w172;
assign w212 = w40 & w210;
assign w213 = w211 & w212;
assign w214 = ~w72 & w172;
assign w215 = w139 & w172;
assign w216 = ~w103 & w215;
assign w217 = (~w104 & ~w215) | (~w104 & w2379) | (~w215 & w2379);
assign w218 = w40 & ~w214;
assign w219 = ~w217 & w218;
assign w220 = w40 & ~w139;
assign w221 = ~w206 & ~w214;
assign w222 = ~w221 & w2380;
assign w223 = w104 & ~w172;
assign w224 = w139 & w223;
assign w225 = w204 & ~w224;
assign w226 = ~w40 & w106;
assign w227 = ~w211 & w226;
assign w228 = w225 & ~w227;
assign w229 = w228 & w2381;
assign w230 = ~w104 & ~w211;
assign w231 = w104 & ~w215;
assign w232 = ~w230 & ~w231;
assign w233 = ~w204 & ~w232;
assign w234 = ~w178 & w233;
assign w235 = ~w229 & ~w234;
assign w236 = ~w209 & ~w213;
assign w237 = ~w181 & w236;
assign w238 = ~w235 & w237;
assign w239 = pi139 & ~w9;
assign w240 = ~pi236 & w9;
assign w241 = ~w239 & ~w240;
assign w242 = ~w238 & w241;
assign w243 = w238 & ~w241;
assign w244 = ~w242 & ~w243;
assign w245 = (pi088 & ~w8) | (pi088 & w2121) | (~w8 & w2121);
assign w246 = w8 & w2122;
assign w247 = ~w245 & ~w246;
assign w248 = (pi033 & ~w8) | (pi033 & w2123) | (~w8 & w2123);
assign w249 = w8 & w2124;
assign w250 = ~w248 & ~w249;
assign w251 = w6 & ~w250;
assign w252 = (pi036 & ~w8) | (pi036 & w2125) | (~w8 & w2125);
assign w253 = w8 & w2126;
assign w254 = ~w252 & ~w253;
assign w255 = w20 & ~w254;
assign w256 = (pi193 & w247) | (pi193 & w2233) | (w247 & w2233);
assign w257 = ~w251 & ~w255;
assign w258 = w256 & w257;
assign w259 = (pi073 & ~w8) | (pi073 & w2127) | (~w8 & w2127);
assign w260 = w8 & w2128;
assign w261 = ~w259 & ~w260;
assign w262 = (pi044 & ~w8) | (pi044 & w2129) | (~w8 & w2129);
assign w263 = w8 & w2130;
assign w264 = ~w262 & ~w263;
assign w265 = w6 & ~w264;
assign w266 = (~pi193 & w261) | (~pi193 & w2189) | (w261 & w2189);
assign w267 = ~w265 & w266;
assign w268 = ~w258 & ~w267;
assign w269 = pi019 & ~w9;
assign w270 = pi209 & w9;
assign w271 = ~w269 & ~w270;
assign w272 = ~w258 & w2234;
assign w273 = (~w271 & w258) | (~w271 & w2235) | (w258 & w2235);
assign w274 = ~w272 & ~w273;
assign w275 = (pi089 & ~w8) | (pi089 & w2131) | (~w8 & w2131);
assign w276 = w8 & w2132;
assign w277 = ~w275 & ~w276;
assign w278 = (pi079 & ~w8) | (pi079 & w2133) | (~w8 & w2133);
assign w279 = w8 & w2134;
assign w280 = ~w278 & ~w279;
assign w281 = w20 & ~w280;
assign w282 = (pi057 & ~w8) | (pi057 & w2135) | (~w8 & w2135);
assign w283 = w8 & w2136;
assign w284 = ~w282 & ~w283;
assign w285 = w6 & ~w284;
assign w286 = (pi193 & w277) | (pi193 & w2233) | (w277 & w2233);
assign w287 = ~w281 & ~w285;
assign w288 = w286 & w287;
assign w289 = (pi034 & ~w8) | (pi034 & w2137) | (~w8 & w2137);
assign w290 = w8 & w2138;
assign w291 = ~w289 & ~w290;
assign w292 = (pi055 & ~w8) | (pi055 & w2139) | (~w8 & w2139);
assign w293 = w8 & w2140;
assign w294 = ~w292 & ~w293;
assign w295 = w6 & ~w294;
assign w296 = (~pi193 & w291) | (~pi193 & w2189) | (w291 & w2189);
assign w297 = ~w295 & w296;
assign w298 = ~w288 & ~w297;
assign w299 = pi023 & ~w9;
assign w300 = pi201 & w9;
assign w301 = ~w299 & ~w300;
assign w302 = ~w288 & w2236;
assign w303 = (~w301 & w288) | (~w301 & w2237) | (w288 & w2237);
assign w304 = ~w302 & ~w303;
assign w305 = w274 & ~w304;
assign w306 = (pi085 & ~w8) | (pi085 & w2141) | (~w8 & w2141);
assign w307 = w8 & w2142;
assign w308 = ~w306 & ~w307;
assign w309 = w20 & ~w264;
assign w310 = w6 & ~w261;
assign w311 = (pi193 & w308) | (pi193 & w2233) | (w308 & w2233);
assign w312 = ~w309 & ~w310;
assign w313 = w311 & w312;
assign w314 = w6 & ~w280;
assign w315 = (~pi193 & w284) | (~pi193 & w2189) | (w284 & w2189);
assign w316 = ~w314 & w315;
assign w317 = ~w313 & ~w316;
assign w318 = pi003 & ~w9;
assign w319 = pi251 & w9;
assign w320 = ~w318 & ~w319;
assign w321 = ~w313 & w2238;
assign w322 = (~w320 & w313) | (~w320 & w2239) | (w313 & w2239);
assign w323 = ~w321 & ~w322;
assign w324 = w304 & ~w323;
assign w325 = (pi067 & ~w8) | (pi067 & w2143) | (~w8 & w2143);
assign w326 = w8 & w2144;
assign w327 = ~w325 & ~w326;
assign w328 = (pi032 & ~w8) | (pi032 & w2145) | (~w8 & w2145);
assign w329 = w8 & w2146;
assign w330 = ~w328 & ~w329;
assign w331 = w6 & ~w330;
assign w332 = (pi070 & ~w8) | (pi070 & w2147) | (~w8 & w2147);
assign w333 = w8 & w2148;
assign w334 = ~w332 & ~w333;
assign w335 = w20 & ~w334;
assign w336 = (pi193 & w327) | (pi193 & w2233) | (w327 & w2233);
assign w337 = ~w331 & ~w335;
assign w338 = w336 & w337;
assign w339 = (pi038 & ~w8) | (pi038 & w2149) | (~w8 & w2149);
assign w340 = w8 & w2150;
assign w341 = ~w339 & ~w340;
assign w342 = (pi052 & ~w8) | (pi052 & w2151) | (~w8 & w2151);
assign w343 = w8 & w2152;
assign w344 = ~w342 & ~w343;
assign w345 = w6 & ~w344;
assign w346 = (~pi193 & w341) | (~pi193 & w2189) | (w341 & w2189);
assign w347 = ~w345 & w346;
assign w348 = ~w338 & ~w347;
assign w349 = pi002 & ~w9;
assign w350 = pi217 & w9;
assign w351 = ~w349 & ~w350;
assign w352 = ~w338 & w2240;
assign w353 = (~w351 & w338) | (~w351 & w2241) | (w338 & w2241);
assign w354 = ~w352 & ~w353;
assign w355 = ~w324 & ~w354;
assign w356 = w304 & w323;
assign w357 = w354 & ~w356;
assign w358 = ~w355 & ~w357;
assign w359 = (pi046 & ~w8) | (pi046 & w2153) | (~w8 & w2153);
assign w360 = w8 & w2154;
assign w361 = ~w359 & ~w360;
assign w362 = (pi051 & ~w8) | (pi051 & w2155) | (~w8 & w2155);
assign w363 = w8 & w2156;
assign w364 = ~w362 & ~w363;
assign w365 = w6 & ~w364;
assign w366 = (pi084 & ~w8) | (pi084 & w2157) | (~w8 & w2157);
assign w367 = w8 & w2158;
assign w368 = ~w366 & ~w367;
assign w369 = w20 & ~w368;
assign w370 = (pi193 & w361) | (pi193 & w2233) | (w361 & w2233);
assign w371 = ~w365 & ~w369;
assign w372 = w370 & w371;
assign w373 = (pi043 & ~w8) | (pi043 & w2159) | (~w8 & w2159);
assign w374 = w8 & w2160;
assign w375 = ~w373 & ~w374;
assign w376 = (pi086 & ~w8) | (pi086 & w2161) | (~w8 & w2161);
assign w377 = w8 & w2162;
assign w378 = ~w376 & ~w377;
assign w379 = w6 & ~w378;
assign w380 = (~pi193 & w375) | (~pi193 & w2189) | (w375 & w2189);
assign w381 = ~w379 & w380;
assign w382 = ~w372 & ~w381;
assign w383 = pi028 & ~w9;
assign w384 = pi225 & w9;
assign w385 = ~w383 & ~w384;
assign w386 = ~w372 & w2242;
assign w387 = (~w385 & w372) | (~w385 & w2243) | (w372 & w2243);
assign w388 = ~w386 & ~w387;
assign w389 = (~w388 & w358) | (~w388 & w923) | (w358 & w923);
assign w390 = ~w323 & w354;
assign w391 = w274 & w390;
assign w392 = w390 & w2294;
assign w393 = w304 & w392;
assign w394 = w274 & w323;
assign w395 = w304 & ~w394;
assign w396 = ~w354 & w388;
assign w397 = ~w305 & w396;
assign w398 = ~w395 & w397;
assign w399 = (pi087 & ~w8) | (pi087 & w2163) | (~w8 & w2163);
assign w400 = w8 & w2164;
assign w401 = ~w399 & ~w400;
assign w402 = w6 & ~w401;
assign w403 = (pi063 & ~w8) | (pi063 & w2165) | (~w8 & w2165);
assign w404 = w8 & w2166;
assign w405 = ~w403 & ~w404;
assign w406 = ~w6 & ~w405;
assign w407 = ~w402 & ~w406;
assign w408 = ~pi193 & ~w407;
assign w409 = (pi049 & ~w8) | (pi049 & w2167) | (~w8 & w2167);
assign w410 = w8 & w2168;
assign w411 = ~w409 & ~w410;
assign w412 = w8 & ~w411;
assign w413 = (pi062 & ~w8) | (pi062 & w2169) | (~w8 & w2169);
assign w414 = w8 & w2170;
assign w415 = ~w413 & ~w414;
assign w416 = ~w415 & w20;
assign w417 = ~w379 & ~w412;
assign w418 = (pi193 & ~w417) | (pi193 & w2295) | (~w417 & w2295);
assign w419 = ~w408 & ~w418;
assign w420 = pi030 & ~w9;
assign w421 = pi233 & w9;
assign w422 = ~w420 & ~w421;
assign w423 = ~w419 & w422;
assign w424 = w419 & ~w422;
assign w425 = ~w423 & ~w424;
assign w426 = ~w398 & ~w425;
assign w427 = ~w393 & w426;
assign w428 = ~w388 & w425;
assign w429 = ~w304 & w323;
assign w430 = ~w324 & ~w429;
assign w431 = ~w304 & w354;
assign w432 = ~w274 & ~w431;
assign w433 = ~w430 & w432;
assign w434 = w428 & ~w433;
assign w435 = (~w434 & ~w427) | (~w434 & w2296) | (~w427 & w2296);
assign w436 = w305 & ~w323;
assign w437 = ~w354 & w436;
assign w438 = w274 & w304;
assign w439 = ~w356 & ~w394;
assign w440 = ~w438 & ~w439;
assign w441 = w354 & w440;
assign w442 = ~w437 & ~w441;
assign w443 = w324 & w354;
assign w444 = ~w355 & ~w443;
assign w445 = ~w429 & w444;
assign w446 = w388 & w425;
assign w447 = ~w440 & w446;
assign w448 = ~w445 & w447;
assign w449 = (~w448 & w435) | (~w448 & w2382) | (w435 & w2382);
assign w450 = ~w388 & ~w425;
assign w451 = ~w274 & ~w323;
assign w452 = w431 & w451;
assign w453 = ~w450 & w452;
assign w454 = ~w449 & ~w453;
assign w455 = pi145 & ~w9;
assign w456 = ~pi244 & w9;
assign w457 = ~w455 & ~w456;
assign w458 = w454 & ~w457;
assign w459 = ~w454 & w457;
assign w460 = ~w458 & ~w459;
assign w461 = (pi090 & ~w8) | (pi090 & w2171) | (~w8 & w2171);
assign w462 = ~w77 & ~w461;
assign w463 = w6 & ~w462;
assign w464 = w8 & w2098;
assign w465 = w20 & ~w93;
assign w466 = (pi193 & ~w8) | (pi193 & w2244) | (~w8 & w2244);
assign w467 = ~w464 & w466;
assign w468 = ~w463 & w467;
assign w469 = ~w465 & w468;
assign w470 = w6 & ~w50;
assign w471 = ~w6 & ~w43;
assign w472 = (~pi193 & w50) | (~pi193 & w2178) | (w50 & w2178);
assign w473 = ~w471 & w472;
assign w474 = ~w469 & ~w473;
assign w475 = pi014 & ~w9;
assign w476 = pi255 & w9;
assign w477 = ~w475 & ~w476;
assign w478 = ~w469 & w2245;
assign w479 = (~w477 & w469) | (~w477 & w2246) | (w469 & w2246);
assign w480 = ~w478 & ~w479;
assign w481 = w6 & ~w143;
assign w482 = w8 & w2247;
assign w483 = w20 & ~w147;
assign w484 = (pi193 & ~w8) | (pi193 & w2248) | (~w8 & w2248);
assign w485 = ~w482 & w484;
assign w486 = ~w481 & w485;
assign w487 = ~w483 & w486;
assign w488 = (~pi193 & w118) | (~pi193 & w2178) | (w118 & w2178);
assign w489 = ~w189 & w488;
assign w490 = ~w487 & ~w489;
assign w491 = pi013 & ~w9;
assign w492 = pi197 & w9;
assign w493 = ~w491 & ~w492;
assign w494 = ~w487 & w2249;
assign w495 = (~w493 & w487) | (~w493 & w2250) | (w487 & w2250);
assign w496 = ~w494 & ~w495;
assign w497 = w6 & ~w129;
assign w498 = w8 & w2172;
assign w499 = w8 & w2183;
assign w500 = w20 & ~w125;
assign w501 = (pi193 & ~w8) | (pi193 & w2251) | (~w8 & w2251);
assign w502 = ~w499 & w501;
assign w503 = ~w497 & w502;
assign w504 = ~w500 & w503;
assign w505 = w6 & ~w23;
assign w506 = ~w6 & ~w31;
assign w507 = (~pi193 & w23) | (~pi193 & w2178) | (w23 & w2178);
assign w508 = ~w506 & w507;
assign w509 = ~w504 & ~w508;
assign w510 = pi027 & ~w9;
assign w511 = pi205 & w9;
assign w512 = ~w510 & ~w511;
assign w513 = ~w504 & w2252;
assign w514 = (~w512 & w504) | (~w512 & w2253) | (w504 & w2253);
assign w515 = ~w513 & ~w514;
assign w516 = ~w496 & w515;
assign w517 = ~w480 & w516;
assign w518 = ~w6 & ~w162;
assign w519 = w6 & ~w153;
assign w520 = ~w518 & ~w519;
assign w521 = ~pi193 & ~w520;
assign w522 = w6 & ~w62;
assign w523 = w8 & ~w158;
assign w524 = ~w6 & ~w58;
assign w525 = ~w58 & w20;
assign w526 = ~w522 & ~w523;
assign w527 = (pi193 & ~w526) | (pi193 & w2297) | (~w526 & w2297);
assign w528 = ~w521 & ~w527;
assign w529 = pi012 & ~w9;
assign w530 = pi221 & w9;
assign w531 = ~w529 & ~w530;
assign w532 = ~w528 & w531;
assign w533 = w528 & ~w531;
assign w534 = ~w532 & ~w533;
assign w535 = ~w517 & ~w534;
assign w536 = w480 & ~w496;
assign w537 = w6 & ~w16;
assign w538 = w8 & w2093;
assign w539 = ~w12 & w20;
assign w540 = (pi193 & ~w8) | (pi193 & w2254) | (~w8 & w2254);
assign w541 = ~w538 & w540;
assign w542 = ~w537 & w541;
assign w543 = ~w539 & w542;
assign w544 = ~w6 & ~w81;
assign w545 = (~pi193 & w462) | (~pi193 & w2178) | (w462 & w2178);
assign w546 = ~w544 & w545;
assign w547 = ~w543 & ~w546;
assign w548 = pi031 & ~w9;
assign w549 = pi213 & w9;
assign w550 = ~w548 & ~w549;
assign w551 = ~w543 & w2255;
assign w552 = (~w550 & w543) | (~w550 & w2256) | (w543 & w2256);
assign w553 = ~w551 & ~w552;
assign w554 = ~w515 & w553;
assign w555 = w536 & w554;
assign w556 = w480 & ~w516;
assign w557 = ~w480 & ~w496;
assign w558 = w496 & ~w553;
assign w559 = ~w114 & ~w497;
assign w560 = ~pi193 & ~w559;
assign w561 = w8 & ~w109;
assign w562 = w6 & ~w188;
assign w563 = w20 & ~w118;
assign w564 = ~w561 & ~w562;
assign w565 = ~w563 & w564;
assign w566 = pi193 & ~w565;
assign w567 = ~w560 & ~w566;
assign w568 = pi024 & ~w9;
assign w569 = pi229 & w9;
assign w570 = ~w568 & ~w569;
assign w571 = ~w567 & w570;
assign w572 = w567 & ~w570;
assign w573 = ~w571 & ~w572;
assign w574 = ~w558 & ~w573;
assign w575 = ~w556 & ~w557;
assign w576 = w574 & w575;
assign w577 = w480 & ~w553;
assign w578 = w516 & w577;
assign w579 = w534 & ~w555;
assign w580 = ~w578 & w579;
assign w581 = ~w576 & w580;
assign w582 = ~w535 & ~w581;
assign w583 = w517 & w553;
assign w584 = w480 & w496;
assign w585 = ~w515 & w584;
assign w586 = w534 & ~w585;
assign w587 = ~w480 & w558;
assign w588 = w586 & ~w587;
assign w589 = ~w515 & ~w536;
assign w590 = ~w553 & ~w589;
assign w591 = ~w480 & w554;
assign w592 = ~w516 & ~w534;
assign w593 = ~w591 & w592;
assign w594 = ~w590 & w593;
assign w595 = ~w588 & ~w594;
assign w596 = w573 & ~w583;
assign w597 = ~w595 & w596;
assign w598 = ~w553 & w557;
assign w599 = ~w515 & w598;
assign w600 = ~w534 & ~w553;
assign w601 = ~w534 & w2383;
assign w602 = w496 & ~w515;
assign w603 = w577 & w602;
assign w604 = w553 & w584;
assign w605 = ~w534 & w604;
assign w606 = ~w555 & ~w573;
assign w607 = ~w603 & w606;
assign w608 = ~w599 & ~w601;
assign w609 = ~w605 & w608;
assign w610 = w607 & w609;
assign w611 = ~w597 & ~w610;
assign w612 = ~w582 & ~w611;
assign w613 = pi147 & ~w9;
assign w614 = ~pi216 & w9;
assign w615 = ~w613 & ~w614;
assign w616 = w612 & ~w615;
assign w617 = ~w612 & w615;
assign w618 = ~w616 & ~w617;
assign w619 = (~w230 & w178) | (~w230 & w2384) | (w178 & w2384);
assign w620 = w40 & w175;
assign w621 = ~w176 & ~w220;
assign w622 = ~w172 & w621;
assign w623 = (~w105 & w622) | (~w105 & w2385) | (w622 & w2385);
assign w624 = ~w40 & w172;
assign w625 = ~w106 & w624;
assign w626 = ~w204 & ~w625;
assign w627 = ~w222 & w626;
assign w628 = ~w623 & w627;
assign w629 = (~w624 & w221) | (~w624 & w2298) | (w221 & w2298);
assign w630 = w210 & ~w629;
assign w631 = w207 & w2386;
assign w632 = ~w224 & ~w631;
assign w633 = w40 & ~w105;
assign w634 = w179 & ~w633;
assign w635 = w40 & w216;
assign w636 = w176 & w206;
assign w637 = w204 & ~w634;
assign w638 = ~w636 & w637;
assign w639 = ~w635 & w638;
assign w640 = w639 & w2387;
assign w641 = (~w619 & w640) | (~w619 & w2299) | (w640 & w2299);
assign w642 = pi149 & ~w9;
assign w643 = ~pi250 & w9;
assign w644 = ~w642 & ~w643;
assign w645 = w641 & ~w644;
assign w646 = ~w641 & w644;
assign w647 = ~w645 & ~w646;
assign w648 = w103 & ~w221;
assign w649 = ~w139 & w648;
assign w650 = w632 & ~w649;
assign w651 = w214 & w220;
assign w652 = w176 & ~w207;
assign w653 = (~w176 & w221) | (~w176 & w2388) | (w221 & w2388);
assign w654 = ~w652 & ~w653;
assign w655 = w105 & w621;
assign w656 = w204 & ~w651;
assign w657 = ~w655 & w656;
assign w658 = ~w654 & w657;
assign w659 = ~w103 & w214;
assign w660 = w621 & w659;
assign w661 = ~w220 & w223;
assign w662 = w177 & ~w655;
assign w663 = ~w204 & ~w661;
assign w664 = ~w652 & w663;
assign w665 = ~w660 & w664;
assign w666 = ~w662 & w665;
assign w667 = ~w658 & ~w666;
assign w668 = pi129 & ~w9;
assign w669 = ~pi248 & w9;
assign w670 = ~w668 & ~w669;
assign w671 = ~w667 & w2389;
assign w672 = (w670 & w667) | (w670 & w2390) | (w667 & w2390);
assign w673 = ~w671 & ~w672;
assign w674 = (w553 & ~w584) | (w553 & w2391) | (~w584 & w2391);
assign w675 = w496 & w515;
assign w676 = ~w480 & w675;
assign w677 = ~w553 & ~w676;
assign w678 = ~w674 & ~w677;
assign w679 = w553 & w593;
assign w680 = w480 & w515;
assign w681 = ~w558 & w680;
assign w682 = ~w598 & ~w603;
assign w683 = (~w534 & ~w682) | (~w534 & w2300) | (~w682 & w2300);
assign w684 = w586 & ~w681;
assign w685 = ~w599 & w684;
assign w686 = ~w679 & ~w683;
assign w687 = ~w685 & w686;
assign w688 = (~w573 & w687) | (~w573 & w2392) | (w687 & w2392);
assign w689 = ~w480 & w602;
assign w690 = w602 & w2393;
assign w691 = ~w534 & w690;
assign w692 = ~w516 & ~w536;
assign w693 = ~w515 & w534;
assign w694 = ~w598 & ~w693;
assign w695 = ~w692 & ~w694;
assign w696 = w534 & ~w602;
assign w697 = w553 & w696;
assign w698 = w696 & w2393;
assign w699 = ~w695 & ~w698;
assign w700 = (w573 & ~w699) | (w573 & w2394) | (~w699 & w2394);
assign w701 = w496 & w680;
assign w702 = ~w689 & ~w701;
assign w703 = (~w553 & w702) | (~w553 & w2395) | (w702 & w2395);
assign w704 = ~w517 & w674;
assign w705 = w534 & ~w704;
assign w706 = ~w703 & w705;
assign w707 = ~w691 & ~w706;
assign w708 = ~w700 & w707;
assign w709 = ~w688 & w708;
assign w710 = pi136 & ~w9;
assign w711 = ~pi238 & w9;
assign w712 = ~w710 & ~w711;
assign w713 = w709 & ~w712;
assign w714 = ~w709 & w712;
assign w715 = ~w713 & ~w714;
assign w716 = w536 & ~w553;
assign w717 = ~w601 & ~w716;
assign w718 = w696 & ~w716;
assign w719 = ~w692 & w718;
assign w720 = ~w605 & ~w690;
assign w721 = ~w719 & w720;
assign w722 = (w573 & ~w721) | (w573 & w2396) | (~w721 & w2396);
assign w723 = ~w577 & ~w602;
assign w724 = ~w556 & ~w723;
assign w725 = ~w583 & ~w724;
assign w726 = ~w534 & ~w725;
assign w727 = w577 & w693;
assign w728 = w553 & w675;
assign w729 = ~w555 & ~w701;
assign w730 = w535 & w729;
assign w731 = w554 & w557;
assign w732 = w534 & ~w676;
assign w733 = ~w731 & w732;
assign w734 = ~w730 & ~w733;
assign w735 = ~w578 & ~w728;
assign w736 = ~w734 & w735;
assign w737 = ~w573 & ~w736;
assign w738 = ~w726 & ~w727;
assign w739 = ~w722 & w738;
assign w740 = ~w737 & w739;
assign w741 = pi121 & ~w9;
assign w742 = ~pi256 & w9;
assign w743 = ~w741 & ~w742;
assign w744 = ~w740 & w743;
assign w745 = w740 & ~w743;
assign w746 = ~w744 & ~w745;
assign w747 = ~w6 & ~w364;
assign w748 = w6 & ~w368;
assign w749 = ~w747 & ~w748;
assign w750 = ~pi193 & ~w749;
assign w751 = w6 & ~w327;
assign w752 = w8 & ~w344;
assign w753 = w20 & ~w341;
assign w754 = ~w751 & ~w752;
assign w755 = (pi193 & ~w754) | (pi193 & w2257) | (~w754 & w2257);
assign w756 = ~w750 & ~w755;
assign w757 = pi025 & ~w9;
assign w758 = pi223 & w9;
assign w759 = ~w757 & ~w758;
assign w760 = ~w756 & w759;
assign w761 = w756 & ~w759;
assign w762 = ~w760 & ~w761;
assign w763 = w6 & ~w254;
assign w764 = ~w6 & ~w250;
assign w765 = ~w763 & ~w764;
assign w766 = ~pi193 & ~w765;
assign w767 = (pi050 & ~w8) | (pi050 & w2258) | (~w8 & w2258);
assign w768 = w8 & w2259;
assign w769 = ~w767 & ~w768;
assign w770 = w8 & ~w769;
assign w771 = w6 & ~w405;
assign w772 = ~w401 & w20;
assign w773 = ~w770 & ~w771;
assign w774 = (pi193 & ~w773) | (pi193 & w2301) | (~w773 & w2301);
assign w775 = ~w766 & ~w774;
assign w776 = pi010 & ~w9;
assign w777 = pi231 & w9;
assign w778 = ~w776 & ~w777;
assign w779 = ~w775 & w778;
assign w780 = w775 & ~w778;
assign w781 = ~w779 & ~w780;
assign w782 = w762 & ~w781;
assign w783 = ~w762 & w781;
assign w784 = (pi060 & ~w8) | (pi060 & w2260) | (~w8 & w2260);
assign w785 = w8 & w2261;
assign w786 = ~w784 & ~w785;
assign w787 = ~w6 & ~w786;
assign w788 = (pi056 & ~w8) | (pi056 & w2173) | (~w8 & w2173);
assign w789 = w8 & w2174;
assign w790 = ~w788 & ~w789;
assign w791 = w6 & ~w790;
assign w792 = ~w787 & ~w791;
assign w793 = ~pi193 & ~w792;
assign w794 = w20 & ~w291;
assign w795 = w8 & ~w294;
assign w796 = ~w794 & ~w795;
assign w797 = (pi193 & ~w796) | (pi193 & w2262) | (~w796 & w2262);
assign w798 = ~w793 & ~w797;
assign w799 = pi008 & ~w9;
assign w800 = pi199 & w9;
assign w801 = ~w799 & ~w800;
assign w802 = ~w798 & w801;
assign w803 = w798 & ~w801;
assign w804 = ~w802 & ~w803;
assign w805 = w6 & ~w308;
assign w806 = ~w6 & ~w264;
assign w807 = ~w805 & ~w806;
assign w808 = ~pi193 & ~w807;
assign w809 = w8 & ~w261;
assign w810 = w20 & ~w247;
assign w811 = ~w763 & ~w809;
assign w812 = (pi193 & ~w811) | (pi193 & w2263) | (~w811 & w2263);
assign w813 = ~w808 & ~w812;
assign w814 = pi016 & ~w9;
assign w815 = pi207 & w9;
assign w816 = ~w814 & ~w815;
assign w817 = ~w813 & w816;
assign w818 = w813 & ~w816;
assign w819 = ~w817 & ~w818;
assign w820 = ~w804 & w819;
assign w821 = w6 & ~w341;
assign w822 = ~w6 & ~w327;
assign w823 = ~w821 & ~w822;
assign w824 = ~pi193 & ~w823;
assign w825 = w8 & ~w334;
assign w826 = w20 & ~w330;
assign w827 = ~w791 & ~w825;
assign w828 = (pi193 & ~w827) | (pi193 & w2264) | (~w827 & w2264);
assign w829 = ~w824 & ~w828;
assign w830 = pi006 & ~w9;
assign w831 = pi257 & w9;
assign w832 = ~w830 & ~w831;
assign w833 = ~w829 & w832;
assign w834 = w829 & ~w832;
assign w835 = ~w833 & ~w834;
assign w836 = ~w804 & w835;
assign w837 = w804 & ~w835;
assign w838 = ~w836 & ~w837;
assign w839 = ~w6 & ~w411;
assign w840 = ~w771 & ~w839;
assign w841 = ~pi193 & ~w840;
assign w842 = w20 & ~w378;
assign w843 = w8 & ~w415;
assign w844 = ~w842 & ~w843;
assign w845 = (pi193 & ~w844) | (pi193 & w2265) | (~w844 & w2265);
assign w846 = ~w841 & ~w845;
assign w847 = pi011 & ~w9;
assign w848 = pi215 & w9;
assign w849 = ~w847 & ~w848;
assign w850 = ~w846 & w849;
assign w851 = w846 & ~w849;
assign w852 = ~w850 & ~w851;
assign w853 = w838 & ~w852;
assign w854 = w838 & w2302;
assign w855 = ~w835 & w852;
assign w856 = w819 & w855;
assign w857 = (~w783 & w854) | (~w783 & w2397) | (w854 & w2397);
assign w858 = ~w781 & w852;
assign w859 = ~w819 & ~w835;
assign w860 = ~w804 & w859;
assign w861 = w858 & w860;
assign w862 = ~w835 & ~w852;
assign w863 = w819 & w862;
assign w864 = w804 & ~w852;
assign w865 = ~w804 & w852;
assign w866 = ~w864 & ~w865;
assign w867 = w762 & w781;
assign w868 = ~w863 & w867;
assign w869 = ~w866 & w868;
assign w870 = ~w861 & ~w869;
assign w871 = ~w819 & w855;
assign w872 = ~w869 & w2303;
assign w873 = (~w782 & w872) | (~w782 & w2398) | (w872 & w2398);
assign w874 = w819 & w835;
assign w875 = ~w859 & ~w874;
assign w876 = ~w852 & w875;
assign w877 = w804 & ~w819;
assign w878 = w783 & ~w877;
assign w879 = w876 & w878;
assign w880 = ~w804 & w875;
assign w881 = w819 & ~w836;
assign w882 = w858 & ~w881;
assign w883 = w880 & w882;
assign w884 = ~w852 & w874;
assign w885 = w867 & w884;
assign w886 = w762 & w835;
assign w887 = ~w820 & ~w877;
assign w888 = w852 & w886;
assign w889 = w887 & w888;
assign w890 = w804 & w852;
assign w891 = ~w859 & ~w890;
assign w892 = ~w835 & w890;
assign w893 = ~w891 & ~w892;
assign w894 = ~w804 & w884;
assign w895 = w781 & w894;
assign w896 = ~w893 & w2399;
assign w897 = ~w895 & w896;
assign w898 = ~w804 & ~w819;
assign w899 = ~w862 & ~w898;
assign w900 = w782 & ~w899;
assign w901 = ~w854 & w900;
assign w902 = ~w885 & ~w889;
assign w903 = ~w879 & w902;
assign w904 = w903 & w2304;
assign w905 = ~w897 & w904;
assign w906 = pi142 & ~w9;
assign w907 = ~pi252 & w9;
assign w908 = ~w906 & ~w907;
assign w909 = w905 & w2400;
assign w910 = (w908 & ~w905) | (w908 & w2401) | (~w905 & w2401);
assign w911 = ~w909 & ~w910;
assign w912 = w304 & ~w354;
assign w913 = ~w388 & ~w912;
assign w914 = ~w431 & w913;
assign w915 = ~w441 & w914;
assign w916 = ~w274 & w388;
assign w917 = ~w443 & ~w916;
assign w918 = ~w432 & ~w917;
assign w919 = (~w425 & w915) | (~w425 & w2305) | (w915 & w2305);
assign w920 = ~w395 & ~w431;
assign w921 = w428 & ~w443;
assign w922 = ~w920 & w921;
assign w923 = w305 & ~w388;
assign w924 = ~w441 & w2306;
assign w925 = ~w439 & w2402;
assign w926 = w274 & w430;
assign w927 = w324 & w2307;
assign w928 = (w425 & w926) | (w425 & w2308) | (w926 & w2308);
assign w929 = ~w394 & ~w451;
assign w930 = w912 & w929;
assign w931 = ~w925 & ~w930;
assign w932 = ~w928 & w931;
assign w933 = w388 & ~w932;
assign w934 = ~w922 & ~w924;
assign w935 = ~w919 & w934;
assign w936 = pi154 & ~w9;
assign w937 = ~pi198 & w9;
assign w938 = ~w936 & ~w937;
assign w939 = (w938 & ~w935) | (w938 & w2403) | (~w935 & w2403);
assign w940 = w935 & w2404;
assign w941 = ~w939 & ~w940;
assign w942 = ~w305 & w929;
assign w943 = w428 & w942;
assign w944 = w323 & ~w431;
assign w945 = ~w438 & w446;
assign w946 = ~w944 & w945;
assign w947 = ~w943 & ~w946;
assign w948 = ~w912 & ~w947;
assign w949 = ~w274 & ~w388;
assign w950 = w324 & w949;
assign w951 = ~w928 & ~w950;
assign w952 = ~w354 & ~w951;
assign w953 = w323 & w912;
assign w954 = ~w436 & ~w953;
assign w955 = w388 & ~w954;
assign w956 = w929 & w2309;
assign w957 = (~w438 & w391) | (~w438 & w2405) | (w391 & w2405);
assign w958 = w914 & ~w929;
assign w959 = w429 & w916;
assign w960 = ~w950 & ~w959;
assign w961 = ~w392 & w960;
assign w962 = ~w957 & w961;
assign w963 = (~w425 & ~w962) | (~w425 & w2406) | (~w962 & w2406);
assign w964 = ~w955 & ~w956;
assign w965 = ~w948 & w964;
assign w966 = ~w952 & w965;
assign w967 = pi130 & ~w9;
assign w968 = ~pi242 & w9;
assign w969 = ~w967 & ~w968;
assign w970 = w966 & w2310;
assign w971 = (w969 & ~w966) | (w969 & w2311) | (~w966 & w2311);
assign w972 = ~w970 & ~w971;
assign w973 = w20 & ~w364;
assign w974 = w8 & ~w368;
assign w975 = (pi193 & w344) | (pi193 & w2188) | (w344 & w2188);
assign w976 = ~w973 & ~w974;
assign w977 = w975 & w976;
assign w978 = ~w6 & ~w361;
assign w979 = (~pi193 & w375) | (~pi193 & w2178) | (w375 & w2178);
assign w980 = ~w978 & w979;
assign w981 = ~w977 & ~w980;
assign w982 = ~w977 & w2266;
assign w983 = (~w422 & w977) | (~w422 & w2267) | (w977 & w2267);
assign w984 = ~w982 & ~w983;
assign w985 = w8 & ~w284;
assign w986 = w20 & ~w308;
assign w987 = (pi193 & w264) | (pi193 & w2188) | (w264 & w2188);
assign w988 = ~w985 & ~w986;
assign w989 = w987 & w988;
assign w990 = ~w6 & ~w280;
assign w991 = (~pi193 & w277) | (~pi193 & w2178) | (w277 & w2178);
assign w992 = ~w990 & w991;
assign w993 = ~w989 & ~w992;
assign w994 = pi022 & ~w9;
assign w995 = pi241 & w9;
assign w996 = ~w994 & ~w995;
assign w997 = ~w989 & w2268;
assign w998 = (~w996 & w989) | (~w996 & w2269) | (w989 & w2269);
assign w999 = ~w997 & ~w998;
assign w1000 = w6 & ~w415;
assign w1001 = w20 & ~w411;
assign w1002 = w8 & ~w405;
assign w1003 = (pi193 & w415) | (pi193 & w2188) | (w415 & w2188);
assign w1004 = ~w1001 & ~w1002;
assign w1005 = w1003 & w1004;
assign w1006 = w6 & ~w769;
assign w1007 = (~pi193 & w401) | (~pi193 & w2189) | (w401 & w2189);
assign w1008 = ~w1006 & w1007;
assign w1009 = ~w1005 & ~w1008;
assign w1010 = pi004 & ~w9;
assign w1011 = pi249 & w9;
assign w1012 = ~w1010 & ~w1011;
assign w1013 = ~w1005 & w2270;
assign w1014 = (~w1012 & w1005) | (~w1012 & w2271) | (w1005 & w2271);
assign w1015 = ~w1013 & ~w1014;
assign w1016 = w999 & w1015;
assign w1017 = ~w999 & ~w1015;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = ~w984 & w1018;
assign w1020 = w984 & ~w999;
assign w1021 = w20 & ~w375;
assign w1022 = w6 & ~w361;
assign w1023 = w8 & ~w378;
assign w1024 = pi193 & ~w1021;
assign w1025 = ~w1022 & ~w1023;
assign w1026 = w1024 & w1025;
assign w1027 = w6 & ~w411;
assign w1028 = (~pi193 & w415) | (~pi193 & w2189) | (w415 & w2189);
assign w1029 = ~w1027 & w1028;
assign w1030 = ~w1026 & ~w1029;
assign w1031 = ~w1026 & w2272;
assign w1032 = (~w385 & w1026) | (~w385 & w2273) | (w1026 & w2273);
assign w1033 = ~w1031 & ~w1032;
assign w1034 = w999 & w1033;
assign w1035 = ~w1020 & ~w1034;
assign w1036 = ~w1015 & ~w1033;
assign w1037 = w1015 & w1033;
assign w1038 = ~w1036 & ~w1037;
assign w1039 = ~w984 & ~w1033;
assign w1040 = ~w999 & w1033;
assign w1041 = ~w1039 & ~w1040;
assign w1042 = w1038 & ~w1041;
assign w1043 = ~w1035 & ~w1042;
assign w1044 = ~w1019 & ~w1043;
assign w1045 = w984 & w1015;
assign w1046 = ~w1015 & w1039;
assign w1047 = ~w1045 & ~w1046;
assign w1048 = (~w1033 & w1046) | (~w1033 & w2312) | (w1046 & w2312);
assign w1049 = w6 & ~w334;
assign w1050 = ~w6 & ~w330;
assign w1051 = ~w1049 & ~w1050;
assign w1052 = ~pi193 & ~w1051;
assign w1053 = w8 & ~w790;
assign w1054 = w20 & ~w786;
assign w1055 = ~w295 & ~w1053;
assign w1056 = (pi193 & ~w1055) | (pi193 & w2313) | (~w1055 & w2313);
assign w1057 = ~w1052 & ~w1056;
assign w1058 = w832 & ~w1057;
assign w1059 = ~w832 & w1057;
assign w1060 = ~w1058 & ~w1059;
assign w1061 = ~w1048 & ~w1060;
assign w1062 = w984 & ~w1038;
assign w1063 = (w1060 & w1038) | (w1060 & w2314) | (w1038 & w2314);
assign w1064 = ~w1061 & ~w1063;
assign w1065 = ~w1020 & ~w1033;
assign w1066 = ~w1016 & ~w1065;
assign w1067 = w984 & w1034;
assign w1068 = ~w1042 & ~w1067;
assign w1069 = ~w984 & ~w999;
assign w1070 = ~w1037 & w1069;
assign w1071 = ~w1060 & ~w1070;
assign w1072 = (w1071 & ~w1068) | (w1071 & w2274) | (~w1068 & w2274);
assign w1073 = w984 & w1040;
assign w1074 = w1060 & ~w1073;
assign w1075 = ~w1015 & w1060;
assign w1076 = w1060 & w2407;
assign w1077 = w1034 & w1076;
assign w1078 = (~w1077 & w1072) | (~w1077 & w2315) | (w1072 & w2315);
assign w1079 = ~w1044 & ~w1064;
assign w1080 = ~w1078 & w1079;
assign w1081 = ~w6 & ~w247;
assign w1082 = ~w310 & ~w1081;
assign w1083 = ~pi193 & ~w1082;
assign w1084 = w8 & ~w254;
assign w1085 = w20 & ~w250;
assign w1086 = ~w1006 & ~w1084;
assign w1087 = ~w1085 & w1086;
assign w1088 = pi193 & ~w1087;
assign w1089 = ~w1083 & ~w1088;
assign w1090 = w801 & ~w1089;
assign w1091 = ~w801 & w1089;
assign w1092 = ~w1090 & ~w1091;
assign w1093 = (w1074 & w1043) | (w1074 & w2316) | (w1043 & w2316);
assign w1094 = ~w1020 & w1037;
assign w1095 = ~w1060 & ~w1094;
assign w1096 = w1020 & ~w1037;
assign w1097 = w999 & w1039;
assign w1098 = w1039 & w2408;
assign w1099 = w1095 & ~w1096;
assign w1100 = (w1092 & ~w1099) | (w1092 & w2317) | (~w1099 & w2317);
assign w1101 = ~w1093 & w1100;
assign w1102 = w1033 & ~w1070;
assign w1103 = w1047 & ~w1102;
assign w1104 = w984 & w1033;
assign w1105 = (~w1060 & ~w1018) | (~w1060 & w2318) | (~w1018 & w2318);
assign w1106 = w1020 & ~w1033;
assign w1107 = w1060 & ~w1067;
assign w1108 = ~w1106 & w1107;
assign w1109 = ~w1019 & w1108;
assign w1110 = (~w1092 & w1103) | (~w1092 & w2319) | (w1103 & w2319);
assign w1111 = ~w1109 & w1110;
assign w1112 = ~w1101 & ~w1111;
assign w1113 = ~w1080 & w1112;
assign w1114 = pi148 & ~w9;
assign w1115 = ~pi230 & w9;
assign w1116 = ~w1114 & ~w1115;
assign w1117 = w1113 & ~w1116;
assign w1118 = ~w1113 & w1116;
assign w1119 = ~w1117 & ~w1118;
assign w1120 = (~w6 & w192) | (~w6 & w2275) | (w192 & w2275);
assign w1121 = ~w562 & ~w1120;
assign w1122 = ~pi193 & ~w1121;
assign w1123 = w8 & ~w147;
assign w1124 = w20 & ~w143;
assign w1125 = ~w519 & ~w1123;
assign w1126 = (pi193 & ~w1125) | (pi193 & w2276) | (~w1125 & w2276);
assign w1127 = ~w1122 & ~w1126;
assign w1128 = pi000 & ~w9;
assign w1129 = pi237 & w9;
assign w1130 = ~w1128 & ~w1129;
assign w1131 = ~w1127 & w1130;
assign w1132 = w1127 & ~w1130;
assign w1133 = ~w1131 & ~w1132;
assign w1134 = ~w159 & ~w524;
assign w1135 = ~pi193 & ~w1134;
assign w1136 = w8 & ~w62;
assign w1137 = (pi080 & ~w8) | (pi080 & w2175) | (~w8 & w2175);
assign w1138 = ~w45 & ~w1137;
assign w1139 = w20 & ~w1138;
assign w1140 = ~w470 & ~w1136;
assign w1141 = (pi193 & ~w1140) | (pi193 & w2176) | (~w1140 & w2176);
assign w1142 = ~w1135 & ~w1141;
assign w1143 = pi001 & ~w9;
assign w1144 = pi245 & w9;
assign w1145 = ~w1143 & ~w1144;
assign w1146 = ~w1142 & w1145;
assign w1147 = w1142 & ~w1145;
assign w1148 = ~w1146 & ~w1147;
assign w1149 = ~w1133 & ~w1148;
assign w1150 = w6 & ~w81;
assign w1151 = w8 & w2100;
assign w1152 = w20 & ~w462;
assign w1153 = (pi193 & ~w8) | (pi193 & w2177) | (~w8 & w2177);
assign w1154 = ~w1151 & w1153;
assign w1155 = ~w1150 & w1154;
assign w1156 = ~w1152 & w1155;
assign w1157 = ~w6 & ~w89;
assign w1158 = (~pi193 & w43) | (~pi193 & w2178) | (w43 & w2178);
assign w1159 = ~w1157 & w1158;
assign w1160 = ~w1156 & ~w1159;
assign w1161 = ~w1156 & w2179;
assign w1162 = (~w570 & w1156) | (~w570 & w2180) | (w1156 & w2180);
assign w1163 = ~w1161 & ~w1162;
assign w1164 = w6 & ~w113;
assign w1165 = w8 & w2181;
assign w1166 = w20 & ~w129;
assign w1167 = (pi193 & ~w8) | (pi193 & w2182) | (~w8 & w2182);
assign w1168 = ~w1165 & w1167;
assign w1169 = ~w1164 & w1168;
assign w1170 = ~w1166 & w1169;
assign w1171 = (pi071 & ~w8) | (pi071 & w2183) | (~w8 & w2183);
assign w1172 = ~w498 & ~w1171;
assign w1173 = ~w6 & ~w1172;
assign w1174 = (~pi193 & w31) | (~pi193 & w2178) | (w31 & w2178);
assign w1175 = ~w1173 & w1174;
assign w1176 = ~w1170 & ~w1175;
assign w1177 = ~w1170 & w2184;
assign w1178 = (~w531 & w1170) | (~w531 & w2185) | (w1170 & w2185);
assign w1179 = ~w1177 & ~w1178;
assign w1180 = w1163 & w1179;
assign w1181 = ~w1163 & ~w1179;
assign w1182 = ~w1180 & ~w1181;
assign w1183 = w1149 & w1182;
assign w1184 = w1148 & w1179;
assign w1185 = w1148 & w1180;
assign w1186 = ~w1183 & ~w1185;
assign w1187 = ~w6 & ~w27;
assign w1188 = ~w537 & ~w1187;
assign w1189 = ~pi193 & ~w1188;
assign w1190 = w8 & ~w23;
assign w1191 = w6 & ~w1172;
assign w1192 = w20 & ~w31;
assign w1193 = ~w1190 & ~w1191;
assign w1194 = (pi193 & ~w1193) | (pi193 & w2277) | (~w1193 & w2277);
assign w1195 = ~w1189 & ~w1194;
assign w1196 = w69 & ~w1195;
assign w1197 = ~w69 & w1195;
assign w1198 = ~w1196 & ~w1197;
assign w1199 = (w1198 & w1183) | (w1198 & w2186) | (w1183 & w2186);
assign w1200 = w1133 & w1179;
assign w1201 = ~w1133 & ~w1179;
assign w1202 = ~w1200 & ~w1201;
assign w1203 = ~w1133 & w1163;
assign w1204 = ~w1202 & w2187;
assign w1205 = ~w1199 & ~w1204;
assign w1206 = ~w1133 & w1179;
assign w1207 = w1148 & ~w1163;
assign w1208 = w1206 & ~w1207;
assign w1209 = w1205 & w1208;
assign w1210 = ~w1148 & w1163;
assign w1211 = (~w1179 & w1148) | (~w1179 & w1181) | (w1148 & w1181);
assign w1212 = ~w1207 & w1211;
assign w1213 = ~w1133 & w1212;
assign w1214 = ~w1133 & ~w1163;
assign w1215 = w1148 & ~w1214;
assign w1216 = w1179 & w1198;
assign w1217 = ~w1149 & w1216;
assign w1218 = ~w1215 & w1217;
assign w1219 = ~w1213 & ~w1218;
assign w1220 = ~w154 & ~w481;
assign w1221 = ~pi193 & ~w1220;
assign w1222 = w8 & ~w162;
assign w1223 = ~w158 & w20;
assign w1224 = ~w59 & ~w1222;
assign w1225 = (pi193 & ~w1224) | (pi193 & w2320) | (~w1224 & w2320);
assign w1226 = ~w1221 & ~w1225;
assign w1227 = w169 & ~w1226;
assign w1228 = ~w169 & w1226;
assign w1229 = ~w1227 & ~w1228;
assign w1230 = (~w1229 & w1209) | (~w1229 & w2321) | (w1209 & w2321);
assign w1231 = w1198 & ~w1212;
assign w1232 = ~w1163 & w1179;
assign w1233 = ~w1198 & ~w1232;
assign w1234 = ~w1198 & ~w1229;
assign w1235 = w1133 & ~w1233;
assign w1236 = ~w1234 & w1235;
assign w1237 = ~w1231 & w1236;
assign w1238 = ~w1205 & w1229;
assign w1239 = w1133 & w1163;
assign w1240 = ~w1202 & w2322;
assign w1241 = w1148 & w1229;
assign w1242 = w1181 & w1241;
assign w1243 = w1202 & w1210;
assign w1244 = ~w1242 & ~w1243;
assign w1245 = (~w1198 & ~w1244) | (~w1198 & w2323) | (~w1244 & w2323);
assign w1246 = ~w1237 & ~w1238;
assign w1247 = ~w1245 & w1246;
assign w1248 = pi123 & ~w9;
assign w1249 = ~pi214 & w9;
assign w1250 = ~w1248 & ~w1249;
assign w1251 = (w1250 & ~w1247) | (w1250 & w2324) | (~w1247 & w2324);
assign w1252 = w1247 & w2325;
assign w1253 = ~w1251 & ~w1252;
assign w1254 = w8 & ~w401;
assign w1255 = w20 & ~w405;
assign w1256 = (pi193 & w411) | (pi193 & w2188) | (w411 & w2188);
assign w1257 = ~w1254 & ~w1255;
assign w1258 = w1256 & w1257;
assign w1259 = ~w6 & ~w769;
assign w1260 = (~pi193 & w250) | (~pi193 & w2178) | (w250 & w2178);
assign w1261 = ~w1259 & w1260;
assign w1262 = ~w1258 & ~w1261;
assign w1263 = ~w1258 & w2278;
assign w1264 = (~w778 & w1258) | (~w778 & w2279) | (w1258 & w2279);
assign w1265 = ~w1263 & ~w1264;
assign w1266 = w8 & ~w280;
assign w1267 = w20 & ~w284;
assign w1268 = (pi193 & w308) | (pi193 & w2188) | (w308 & w2188);
assign w1269 = ~w1266 & ~w1267;
assign w1270 = w1268 & w1269;
assign w1271 = w6 & ~w291;
assign w1272 = (~pi193 & w277) | (~pi193 & w2189) | (w277 & w2189);
assign w1273 = ~w1271 & w1272;
assign w1274 = ~w1270 & ~w1273;
assign w1275 = ~w1270 & w2190;
assign w1276 = (~w759 & w1270) | (~w759 & w2191) | (w1270 & w2191);
assign w1277 = ~w1275 & ~w1276;
assign w1278 = ~w1265 & ~w1277;
assign w1279 = ~w6 & ~w790;
assign w1280 = ~w331 & ~w1279;
assign w1281 = ~pi193 & ~w1280;
assign w1282 = w8 & ~w786;
assign w1283 = ~w6 & ~w294;
assign w1284 = ~w294 & w20;
assign w1285 = ~w1271 & ~w1282;
assign w1286 = (pi193 & ~w1285) | (pi193 & w2192) | (~w1285 & w2192);
assign w1287 = ~w1281 & ~w1286;
assign w1288 = pi015 & ~w9;
assign w1289 = pi247 & w9;
assign w1290 = ~w1288 & ~w1289;
assign w1291 = ~w1287 & w1290;
assign w1292 = w1287 & ~w1290;
assign w1293 = ~w1291 & ~w1292;
assign w1294 = w1278 & ~w1293;
assign w1295 = ~w6 & ~w308;
assign w1296 = ~w285 & ~w1295;
assign w1297 = ~pi193 & ~w1296;
assign w1298 = w6 & ~w247;
assign w1299 = w8 & ~w264;
assign w1300 = w20 & ~w261;
assign w1301 = ~w1298 & ~w1299;
assign w1302 = (pi193 & ~w1301) | (pi193 & w2280) | (~w1301 & w2280);
assign w1303 = ~w1297 & ~w1302;
assign w1304 = w477 & ~w1303;
assign w1305 = ~w477 & w1303;
assign w1306 = ~w1304 & ~w1305;
assign w1307 = ~w6 & ~w368;
assign w1308 = ~w1022 & ~w1307;
assign w1309 = ~pi193 & ~w1308;
assign w1310 = w8 & ~w364;
assign w1311 = ~w6 & ~w344;
assign w1312 = ~w344 & w20;
assign w1313 = ~w821 & ~w1310;
assign w1314 = (pi193 & ~w1313) | (pi193 & w2281) | (~w1313 & w2281);
assign w1315 = ~w1309 & ~w1314;
assign w1316 = pi005 & ~w9;
assign w1317 = pi239 & w9;
assign w1318 = ~w1316 & ~w1317;
assign w1319 = ~w1315 & w1318;
assign w1320 = w1315 & ~w1318;
assign w1321 = ~w1319 & ~w1320;
assign w1322 = ~w1306 & w1321;
assign w1323 = w1294 & w1322;
assign w1324 = w1265 & w1277;
assign w1325 = w1293 & w1324;
assign w1326 = ~w1278 & ~w1324;
assign w1327 = ~w1321 & ~w1326;
assign w1328 = (~w1306 & w1325) | (~w1306 & w2326) | (w1325 & w2326);
assign w1329 = ~w1327 & w1328;
assign w1330 = ~w6 & ~w378;
assign w1331 = ~w1000 & ~w1330;
assign w1332 = ~pi193 & ~w1331;
assign w1333 = w8 & ~w375;
assign w1334 = w20 & ~w361;
assign w1335 = ~w748 & ~w1333;
assign w1336 = (pi193 & ~w1335) | (pi193 & w2282) | (~w1335 & w2282);
assign w1337 = ~w1332 & ~w1336;
assign w1338 = w493 & ~w1337;
assign w1339 = ~w493 & w1337;
assign w1340 = ~w1338 & ~w1339;
assign w1341 = w1293 & ~w1321;
assign w1342 = w1265 & ~w1277;
assign w1343 = w1341 & w1342;
assign w1344 = ~w1323 & ~w1340;
assign w1345 = ~w1343 & w1344;
assign w1346 = ~w1329 & w1345;
assign w1347 = w1294 & w1306;
assign w1348 = ~w1265 & w1277;
assign w1349 = w1321 & w1348;
assign w1350 = w1293 & w1349;
assign w1351 = ~w1347 & ~w1350;
assign w1352 = ~w1293 & w1321;
assign w1353 = w1342 & w1352;
assign w1354 = ~w1306 & ~w1326;
assign w1355 = w1277 & w1293;
assign w1356 = ~w1294 & ~w1355;
assign w1357 = w1354 & w1356;
assign w1358 = ~w1321 & w1324;
assign w1359 = w1306 & w1358;
assign w1360 = (w1340 & ~w1352) | (w1340 & w2327) | (~w1352 & w2327);
assign w1361 = ~w1359 & w1360;
assign w1362 = w1351 & ~w1357;
assign w1363 = w1361 & w1362;
assign w1364 = ~w1346 & ~w1363;
assign w1365 = w1293 & ~w1306;
assign w1366 = ~w1324 & ~w1365;
assign w1367 = ~w1321 & ~w1355;
assign w1368 = ~w1366 & w1367;
assign w1369 = w1265 & w1368;
assign w1370 = w1341 & w1348;
assign w1371 = w1294 & ~w1321;
assign w1372 = ~w1294 & w1321;
assign w1373 = (~w1324 & w1294) | (~w1324 & w2328) | (w1294 & w2328);
assign w1374 = w1321 & w1326;
assign w1375 = (w1340 & ~w1326) | (w1340 & w2193) | (~w1326 & w2193);
assign w1376 = ~w1355 & ~w1373;
assign w1377 = ~w1375 & w1376;
assign w1378 = ~w1370 & ~w1371;
assign w1379 = (w1306 & w1377) | (w1306 & w2409) | (w1377 & w2409);
assign w1380 = ~w1364 & ~w1369;
assign w1381 = pi138 & ~w9;
assign w1382 = ~pi220 & w9;
assign w1383 = ~w1381 & ~w1382;
assign w1384 = w1380 & w2329;
assign w1385 = (w1383 & ~w1380) | (w1383 & w2330) | (~w1380 & w2330);
assign w1386 = ~w1384 & ~w1385;
assign w1387 = w913 & w944;
assign w1388 = (w388 & w956) | (w388 & w2410) | (w956 & w2410);
assign w1389 = (w390 & w926) | (w390 & w2331) | (w926 & w2331);
assign w1390 = ~w1387 & ~w1389;
assign w1391 = (w425 & ~w1390) | (w425 & w2411) | (~w1390 & w2411);
assign w1392 = w914 & w926;
assign w1393 = ~w443 & w929;
assign w1394 = ~w425 & w438;
assign w1395 = (~w1394 & w1393) | (~w1394 & w2412) | (w1393 & w2412);
assign w1396 = ~w444 & ~w1395;
assign w1397 = w356 & w916;
assign w1398 = ~w431 & ~w451;
assign w1399 = ~w388 & ~w390;
assign w1400 = ~w1398 & w1399;
assign w1401 = (~w425 & w1400) | (~w425 & w2413) | (w1400 & w2413);
assign w1402 = ~w392 & ~w1392;
assign w1403 = ~w1401 & w1402;
assign w1404 = ~w1396 & w1403;
assign w1405 = pi127 & ~w9;
assign w1406 = ~pi196 & w9;
assign w1407 = ~w1405 & ~w1406;
assign w1408 = (w1407 & ~w1404) | (w1407 & w2414) | (~w1404 & w2414);
assign w1409 = w1404 & w2415;
assign w1410 = ~w1408 & ~w1409;
assign w1411 = w781 & w890;
assign w1412 = w856 & w1411;
assign w1413 = w855 & ~w887;
assign w1414 = (w762 & ~w875) | (w762 & w1425) | (~w875 & w1425);
assign w1415 = ~w1413 & w1414;
assign w1416 = (~w781 & w893) | (~w781 & w782) | (w893 & w782);
assign w1417 = ~w1415 & w1416;
assign w1418 = ~w838 & w852;
assign w1419 = ~w853 & ~w1418;
assign w1420 = w783 & ~w1419;
assign w1421 = (w819 & w781) | (w819 & w2194) | (w781 & w2194);
assign w1422 = ~w819 & ~w867;
assign w1423 = w838 & ~w1421;
assign w1424 = ~w1422 & w1423;
assign w1425 = w762 & w804;
assign w1426 = w876 & w1425;
assign w1427 = ~w894 & ~w1412;
assign w1428 = ~w1424 & w1427;
assign w1429 = ~w1426 & w1428;
assign w1430 = ~w1420 & w1429;
assign w1431 = pi146 & ~w9;
assign w1432 = ~pi254 & w9;
assign w1433 = ~w1431 & ~w1432;
assign w1434 = w1430 & w2332;
assign w1435 = (w1433 & ~w1430) | (w1433 & w2333) | (~w1430 & w2333);
assign w1436 = ~w1434 & ~w1435;
assign w1437 = w20 & ~w62;
assign w1438 = w8 & w2089;
assign w1439 = w6 & ~w1138;
assign w1440 = (pi193 & ~w8) | (pi193 & w2195) | (~w8 & w2195);
assign w1441 = ~w1438 & w1440;
assign w1442 = ~w1437 & w1441;
assign w1443 = ~w1439 & w1442;
assign w1444 = w6 & ~w162;
assign w1445 = (~pi193 & w158) | (~pi193 & w2189) | (w158 & w2189);
assign w1446 = ~w1444 & w1445;
assign w1447 = ~w1443 & ~w1446;
assign w1448 = ~w1443 & w2196;
assign w1449 = (~w37 & w1443) | (~w37 & w2197) | (w1443 & w2197);
assign w1450 = ~w1448 & ~w1449;
assign w1451 = w6 & ~w93;
assign w1452 = w8 & w2084;
assign w1453 = w20 & ~w89;
assign w1454 = (pi193 & ~w8) | (pi193 & w2198) | (~w8 & w2198);
assign w1455 = ~w1452 & w1454;
assign w1456 = ~w1451 & w1455;
assign w1457 = ~w1453 & w1456;
assign w1458 = ~w6 & ~w50;
assign w1459 = (~pi193 & w1138) | (~pi193 & w2178) | (w1138 & w2178);
assign w1460 = ~w1458 & w1459;
assign w1461 = ~w1457 & ~w1460;
assign w1462 = ~w1457 & w2199;
assign w1463 = (~w201 & w1457) | (~w201 & w2200) | (w1457 & w2200);
assign w1464 = ~w1462 & ~w1463;
assign w1465 = w1450 & ~w1464;
assign w1466 = w6 & ~w27;
assign w1467 = w8 & w2201;
assign w1468 = ~w16 & w20;
assign w1469 = (pi193 & ~w8) | (pi193 & w2202) | (~w8 & w2202);
assign w1470 = ~w1467 & w1469;
assign w1471 = ~w1466 & w1470;
assign w1472 = ~w1468 & w1471;
assign w1473 = ~w6 & ~w75;
assign w1474 = (~pi193 & w81) | (~pi193 & w2178) | (w81 & w2178);
assign w1475 = ~w1473 & w1474;
assign w1476 = ~w1472 & ~w1475;
assign w1477 = pi009 & ~w9;
assign w1478 = pi243 & w9;
assign w1479 = ~w1477 & ~w1478;
assign w1480 = ~w1472 & w2203;
assign w1481 = (~w1479 & w1472) | (~w1479 & w2204) | (w1472 & w2204);
assign w1482 = ~w1480 & ~w1481;
assign w1483 = w8 & ~w143;
assign w1484 = w20 & ~w153;
assign w1485 = (pi193 & w162) | (pi193 & w2188) | (w162 & w2188);
assign w1486 = ~w1483 & ~w1484;
assign w1487 = w1485 & w1486;
assign w1488 = (w6 & w192) | (w6 & w2205) | (w192 & w2205);
assign w1489 = (~pi193 & w147) | (~pi193 & w2189) | (w147 & w2189);
assign w1490 = ~w1488 & w1489;
assign w1491 = ~w1487 & ~w1490;
assign w1492 = pi018 & ~w9;
assign w1493 = pi235 & w9;
assign w1494 = ~w1492 & ~w1493;
assign w1495 = ~w1487 & w2206;
assign w1496 = (~w1494 & w1487) | (~w1494 & w2207) | (w1487 & w2207);
assign w1497 = ~w1495 & ~w1496;
assign w1498 = ~w1482 & w1497;
assign w1499 = ~w1450 & w1498;
assign w1500 = ~w1465 & ~w1499;
assign w1501 = w1482 & ~w1497;
assign w1502 = ~w1450 & ~w1501;
assign w1503 = ~w1501 & w1530;
assign w1504 = w1450 & w1482;
assign w1505 = w1464 & w1504;
assign w1506 = ~w6 & ~w125;
assign w1507 = ~w1191 & ~w1506;
assign w1508 = ~pi193 & ~w1507;
assign w1509 = w8 & ~w129;
assign w1510 = w20 & ~w113;
assign w1511 = ~w182 & ~w1509;
assign w1512 = (pi193 & ~w1511) | (pi193 & w2283) | (~w1511 & w2283);
assign w1513 = ~w1508 & ~w1512;
assign w1514 = w320 & ~w1513;
assign w1515 = ~w320 & w1513;
assign w1516 = ~w1514 & ~w1515;
assign w1517 = ~w1505 & w1516;
assign w1518 = ~w1464 & ~w1497;
assign w1519 = ~w1503 & ~w1518;
assign w1520 = w1517 & w1519;
assign w1521 = ~w1464 & w1482;
assign w1522 = ~w1450 & w1521;
assign w1523 = w1516 & ~w1522;
assign w1524 = w1464 & w1501;
assign w1525 = ~w1516 & ~w1524;
assign w1526 = w1450 & w1518;
assign w1527 = w1525 & ~w1526;
assign w1528 = ~w1523 & ~w1527;
assign w1529 = w1502 & w1518;
assign w1530 = ~w1450 & w1464;
assign w1531 = w1498 & w1530;
assign w1532 = ~w1529 & ~w1531;
assign w1533 = ~w1503 & ~w1522;
assign w1534 = ~w1528 & w2284;
assign w1535 = ~w6 & ~w23;
assign w1536 = ~w1466 & ~w1535;
assign w1537 = ~pi193 & ~w1536;
assign w1538 = w8 & ~w31;
assign w1539 = w20 & ~w1172;
assign w1540 = ~w126 & ~w1538;
assign w1541 = (pi193 & ~w1540) | (pi193 & w2334) | (~w1540 & w2334);
assign w1542 = ~w1537 & ~w1541;
assign w1543 = w301 & ~w1542;
assign w1544 = ~w301 & w1542;
assign w1545 = ~w1543 & ~w1544;
assign w1546 = (w1545 & w1534) | (w1545 & w2335) | (w1534 & w2335);
assign w1547 = w1482 & w1530;
assign w1548 = w1530 & w2285;
assign w1549 = w1521 & w2286;
assign w1550 = ~w1548 & ~w1549;
assign w1551 = w1450 & ~w1497;
assign w1552 = w1464 & w1551;
assign w1553 = w1550 & ~w1552;
assign w1554 = (w1516 & ~w1550) | (w1516 & w2336) | (~w1550 & w2336);
assign w1555 = (~w1545 & w1528) | (~w1545 & w2337) | (w1528 & w2337);
assign w1556 = w1465 & ~w1482;
assign w1557 = ~w1505 & ~w1556;
assign w1558 = w1465 & w1498;
assign w1559 = w1516 & ~w1558;
assign w1560 = ~w1557 & ~w1559;
assign w1561 = ~w1554 & ~w1560;
assign w1562 = ~w1555 & w1561;
assign w1563 = ~w1546 & w1562;
assign w1564 = pi125 & ~w9;
assign w1565 = ~pi246 & w9;
assign w1566 = ~w1564 & ~w1565;
assign w1567 = w1563 & ~w1566;
assign w1568 = ~w1563 & w1566;
assign w1569 = ~w1567 & ~w1568;
assign w1570 = w1293 & w1342;
assign w1571 = ~w1293 & w1348;
assign w1572 = ~w1570 & ~w1571;
assign w1573 = ~w1340 & ~w1572;
assign w1574 = ~w1327 & w1375;
assign w1575 = w1277 & ~w1293;
assign w1576 = ~w1374 & w1575;
assign w1577 = ~w1574 & ~w1576;
assign w1578 = ~w1327 & w1572;
assign w1579 = (~w1573 & w1577) | (~w1573 & w2338) | (w1577 & w2338);
assign w1580 = (~w1570 & w1374) | (~w1570 & w2208) | (w1374 & w2208);
assign w1581 = w1340 & ~w1580;
assign w1582 = w1278 & w1341;
assign w1583 = ~w1350 & ~w1358;
assign w1584 = ~w1582 & w1583;
assign w1585 = ~w1581 & w1584;
assign w1586 = ~w1306 & ~w1585;
assign w1587 = w1322 & w1342;
assign w1588 = w1348 & w1365;
assign w1589 = w1293 & w1358;
assign w1590 = ~w1371 & ~w1587;
assign w1591 = ~w1588 & ~w1589;
assign w1592 = w1590 & w1591;
assign w1593 = w1321 & w1570;
assign w1594 = ~w1323 & ~w1593;
assign w1595 = (w1594 & w1592) | (w1594 & w2339) | (w1592 & w2339);
assign w1596 = ~w1586 & w1595;
assign w1597 = pi135 & ~w9;
assign w1598 = ~pi206 & w9;
assign w1599 = ~w1597 & ~w1598;
assign w1600 = (w1599 & ~w1596) | (w1599 & w2340) | (~w1596 & w2340);
assign w1601 = w1596 & w2341;
assign w1602 = ~w1600 & ~w1601;
assign w1603 = w553 & w557;
assign w1604 = ~w604 & ~w689;
assign w1605 = ~w554 & ~w1604;
assign w1606 = w534 & ~w1603;
assign w1607 = ~w1605 & w1606;
assign w1608 = w574 & ~w723;
assign w1609 = (~w534 & ~w598) | (~w534 & w2416) | (~w598 & w2416);
assign w1610 = ~w1608 & w1609;
assign w1611 = ~w1607 & ~w1610;
assign w1612 = ~w600 & w701;
assign w1613 = ~w680 & w697;
assign w1614 = ~w573 & ~w583;
assign w1615 = ~w1612 & w1614;
assign w1616 = ~w1613 & w1615;
assign w1617 = ~w534 & ~w676;
assign w1618 = ~w718 & ~w1617;
assign w1619 = w573 & ~w585;
assign w1620 = ~w731 & w1619;
assign w1621 = ~w1618 & w1620;
assign w1622 = ~w1616 & ~w1621;
assign w1623 = w600 & w676;
assign w1624 = ~w578 & ~w1623;
assign w1625 = ~w1611 & w1624;
assign w1626 = ~w1622 & w1625;
assign w1627 = pi152 & ~w9;
assign w1628 = ~pi194 & w9;
assign w1629 = ~w1627 & ~w1628;
assign w1630 = w1626 & ~w1629;
assign w1631 = ~w1626 & w1629;
assign w1632 = ~w1630 & ~w1631;
assign w1633 = ~w860 & ~w884;
assign w1634 = (w781 & ~w1633) | (w781 & w2209) | (~w1633 & w2209);
assign w1635 = ~w864 & w881;
assign w1636 = ~w819 & w864;
assign w1637 = (~w781 & w1635) | (~w781 & w2342) | (w1635 & w2342);
assign w1638 = ~w883 & ~w894;
assign w1639 = ~w1634 & w1638;
assign w1640 = (~w762 & ~w1639) | (~w762 & w2210) | (~w1639 & w2210);
assign w1641 = ~w819 & w835;
assign w1642 = ~w886 & ~w1641;
assign w1643 = w1411 & ~w1642;
assign w1644 = ~w881 & w2343;
assign w1645 = ~w837 & ~w865;
assign w1646 = ~w874 & w1645;
assign w1647 = ~w1644 & ~w1646;
assign w1648 = pi128 & ~w9;
assign w1649 = ~pi234 & w9;
assign w1650 = ~w1648 & ~w1649;
assign w1651 = (w1650 & w1640) | (w1650 & w2346) | (w1640 & w2346);
assign w1652 = ~w1640 & w2347;
assign w1653 = ~w1651 & ~w1652;
assign w1654 = (~w1072 & w2417) | (~w1072 & w2418) | (w2417 & w2418);
assign w1655 = ~w999 & ~w1047;
assign w1656 = w1075 & w1106;
assign w1657 = ~w1063 & ~w1656;
assign w1658 = ~w1655 & ~w1657;
assign w1659 = ~w1105 & ~w1658;
assign w1660 = ~w1040 & ~w1097;
assign w1661 = w1074 & ~w1660;
assign w1662 = ~w1035 & w1095;
assign w1663 = w1016 & w1039;
assign w1664 = ~w1661 & ~w1663;
assign w1665 = (~w1092 & ~w1664) | (~w1092 & w2348) | (~w1664 & w2348);
assign w1666 = ~w1659 & ~w1665;
assign w1667 = pi151 & ~w9;
assign w1668 = ~pi208 & w9;
assign w1669 = ~w1667 & ~w1668;
assign w1670 = (w1669 & ~w1666) | (w1669 & w2419) | (~w1666 & w2419);
assign w1671 = w1666 & w2420;
assign w1672 = ~w1670 & ~w1671;
assign w1673 = ~w1183 & ~w1229;
assign w1674 = ~w1214 & ~w1239;
assign w1675 = ~w1232 & w1674;
assign w1676 = w1186 & ~w1675;
assign w1677 = w1215 & ~w1676;
assign w1678 = ~w1148 & ~w1182;
assign w1679 = ~w1148 & ~w1180;
assign w1680 = (w2214 & w2349) | (w2214 & w2350) | (w2349 & w2350);
assign w1681 = ~w1677 & w1680;
assign w1682 = (~w1198 & w1681) | (~w1198 & w2215) | (w1681 & w2215);
assign w1683 = ~w1200 & ~w1211;
assign w1684 = w1133 & ~w1182;
assign w1685 = ~w1210 & w1684;
assign w1686 = w1229 & ~w1683;
assign w1687 = ~w1685 & w1686;
assign w1688 = (w1198 & w1687) | (w1198 & w2351) | (w1687 & w2351);
assign w1689 = w1684 & w2287;
assign w1690 = ~w1148 & w1198;
assign w1691 = ~w1232 & ~w1690;
assign w1692 = w1202 & ~w1691;
assign w1693 = ~w1689 & ~w1692;
assign w1694 = w1203 & w1241;
assign w1695 = (~w1694 & w1693) | (~w1694 & w2352) | (w1693 & w2352);
assign w1696 = ~w1688 & w1695;
assign w1697 = pi155 & ~w9;
assign w1698 = ~pi226 & w9;
assign w1699 = ~w1697 & ~w1698;
assign w1700 = (w1699 & w1682) | (w1699 & w2353) | (w1682 & w2353);
assign w1701 = ~w1682 & w2354;
assign w1702 = ~w1700 & ~w1701;
assign w1703 = w1015 & w1060;
assign w1704 = ~w1020 & w1703;
assign w1705 = w1068 & ~w1704;
assign w1706 = (w1060 & ~w1018) | (w1060 & w2216) | (~w1018 & w2216);
assign w1707 = ~w1068 & w1706;
assign w1708 = ~w1705 & ~w1707;
assign w1709 = w1046 & w1060;
assign w1710 = (~w1092 & w1708) | (~w1092 & w2217) | (w1708 & w2217);
assign w1711 = ~w984 & w1034;
assign w1712 = ~w1060 & w1711;
assign w1713 = ~w1661 & ~w1712;
assign w1714 = ~w1064 & w1713;
assign w1715 = (w1015 & w1070) | (w1015 & w2218) | (w1070 & w2218);
assign w1716 = w1062 & ~w1703;
assign w1717 = ~w1712 & ~w1715;
assign w1718 = ~w1716 & w1717;
assign w1719 = w1662 & w1718;
assign w1720 = w1040 & w1703;
assign w1721 = ~w1098 & ~w1656;
assign w1722 = ~w1720 & w1721;
assign w1723 = ~w1719 & w1722;
assign w1724 = ~w1710 & w1723;
assign w1725 = pi150 & ~w9;
assign w1726 = ~pi218 & w9;
assign w1727 = ~w1725 & ~w1726;
assign w1728 = (w1727 & ~w1724) | (w1727 & w2355) | (~w1724 & w2355);
assign w1729 = w1724 & w2356;
assign w1730 = ~w1728 & ~w1729;
assign w1731 = w856 & w1425;
assign w1732 = w804 & ~w875;
assign w1733 = ~w880 & ~w1732;
assign w1734 = w781 & ~w855;
assign w1735 = w1733 & ~w1734;
assign w1736 = (~w762 & w1733) | (~w762 & w2357) | (w1733 & w2357);
assign w1737 = ~w1735 & w1736;
assign w1738 = w782 & ~w859;
assign w1739 = ~w865 & w1738;
assign w1740 = ~w853 & w1739;
assign w1741 = ~w1731 & ~w1740;
assign w1742 = w870 & w1741;
assign w1743 = ~w1737 & w1742;
assign w1744 = pi137 & ~w9;
assign w1745 = ~pi240 & w9;
assign w1746 = ~w1744 & ~w1745;
assign w1747 = w1743 & ~w1746;
assign w1748 = ~w1743 & w1746;
assign w1749 = ~w1747 & ~w1748;
assign w1750 = (~w1340 & w1327) | (~w1340 & w2358) | (w1327 & w2358);
assign w1751 = ~w1341 & ~w1348;
assign w1752 = ~w1265 & w1293;
assign w1753 = ~w1751 & ~w1752;
assign w1754 = ~w1750 & ~w1753;
assign w1755 = w1306 & ~w1754;
assign w1756 = ~w1293 & ~w1342;
assign w1757 = ~w1340 & ~w1570;
assign w1758 = ~w1756 & w1757;
assign w1759 = w1751 & w1758;
assign w1760 = ~w1353 & ~w1370;
assign w1761 = (~w1306 & w1759) | (~w1306 & w2421) | (w1759 & w2421);
assign w1762 = ~w1326 & ~w1340;
assign w1763 = w1277 & w1306;
assign w1764 = w1340 & ~w1763;
assign w1765 = w1352 & ~w1762;
assign w1766 = w1354 & ~w1372;
assign w1767 = ~w1588 & ~w1593;
assign w1768 = ~w1766 & w1767;
assign w1769 = w1340 & ~w1768;
assign w1770 = (~w1371 & ~w1765) | (~w1371 & w2359) | (~w1765 & w2359);
assign w1771 = ~w1769 & w1770;
assign w1772 = ~w1755 & w1771;
assign w1773 = pi131 & ~w9;
assign w1774 = ~pi200 & w9;
assign w1775 = ~w1773 & ~w1774;
assign w1776 = (w1775 & ~w1772) | (w1775 & w2360) | (~w1772 & w2360);
assign w1777 = w1772 & w2361;
assign w1778 = ~w1776 & ~w1777;
assign w1779 = ~w1517 & ~w1554;
assign w1780 = w1518 & ~w1556;
assign w1781 = ~w1482 & w1551;
assign w1782 = w1551 & w2288;
assign w1783 = w1545 & ~w1547;
assign w1784 = ~w1558 & w1783;
assign w1785 = ~w1780 & ~w1782;
assign w1786 = w1784 & w1785;
assign w1787 = w1497 & ~w1530;
assign w1788 = ~w1465 & w1787;
assign w1789 = ~w1545 & ~w1781;
assign w1790 = ~w1788 & w1789;
assign w1791 = ~w1786 & ~w1790;
assign w1792 = ~w1779 & ~w1791;
assign w1793 = ~w1482 & ~w1530;
assign w1794 = ~w1499 & ~w1552;
assign w1795 = (~w1793 & ~w1794) | (~w1793 & w2362) | (~w1794 & w2362);
assign w1796 = w1464 & w1482;
assign w1797 = w1788 & ~w1796;
assign w1798 = ~w1545 & ~w1551;
assign w1799 = ~w1547 & w1798;
assign w1800 = ~w1797 & w1799;
assign w1801 = w1450 & w1497;
assign w1802 = w1521 & w1801;
assign w1803 = ~w1499 & ~w1781;
assign w1804 = w1545 & ~w1803;
assign w1805 = ~w1516 & ~w1802;
assign w1806 = ~w1804 & w1805;
assign w1807 = ~w1795 & w1806;
assign w1808 = ~w1800 & w1807;
assign w1809 = ~w1792 & ~w1808;
assign w1810 = pi140 & ~w9;
assign w1811 = ~pi228 & w9;
assign w1812 = ~w1810 & ~w1811;
assign w1813 = ~w1809 & w2363;
assign w1814 = (w1812 & w1809) | (w1812 & w2364) | (w1809 & w2364);
assign w1815 = ~w1813 & ~w1814;
assign w1816 = (~w620 & ~w208) | (~w620 & w2365) | (~w208 & w2365);
assign w1817 = w139 & ~w1816;
assign w1818 = ~w173 & ~w223;
assign w1819 = ~w225 & ~w1818;
assign w1820 = ~w139 & w210;
assign w1821 = (~w40 & w1819) | (~w40 & w2366) | (w1819 & w2366);
assign w1822 = ~w40 & w204;
assign w1823 = ~w205 & ~w1822;
assign w1824 = ~w659 & w1823;
assign w1825 = ~w174 & w1824;
assign w1826 = ~w179 & ~w211;
assign w1827 = w204 & ~w206;
assign w1828 = ~w1826 & w1827;
assign w1829 = ~w648 & ~w1823;
assign w1830 = ~w1828 & w1829;
assign w1831 = ~w1825 & ~w1830;
assign w1832 = ~w1817 & ~w1821;
assign w1833 = ~w1831 & w1832;
assign w1834 = pi141 & ~w9;
assign w1835 = ~pi222 & w9;
assign w1836 = ~w1834 & ~w1835;
assign w1837 = ~w1833 & w1836;
assign w1838 = w1833 & ~w1836;
assign w1839 = ~w1837 & ~w1838;
assign w1840 = ~w1294 & ~w1348;
assign w1841 = w1265 & ~w1352;
assign w1842 = w1840 & ~w1841;
assign w1843 = (~w1842 & ~w1577) | (~w1842 & w2367) | (~w1577 & w2367);
assign w1844 = ~w1374 & w1840;
assign w1845 = (w1306 & w1374) | (w1306 & w2219) | (w1374 & w2219);
assign w1846 = ~w1844 & w1845;
assign w1847 = (~w1340 & w1846) | (~w1340 & w2368) | (w1846 & w2368);
assign w1848 = w1321 & ~w1351;
assign w1849 = (~w1340 & ~w1358) | (~w1340 & w2369) | (~w1358 & w2369);
assign w1850 = ~w1293 & ~w1321;
assign w1851 = w1326 & w1850;
assign w1852 = ~w1325 & ~w1582;
assign w1853 = ~w1851 & w1852;
assign w1854 = w1306 & ~w1849;
assign w1855 = ~w1853 & w1854;
assign w1856 = ~w1848 & ~w1855;
assign w1857 = ~w1847 & w1856;
assign w1858 = pi157 & ~w9;
assign w1859 = ~pi202 & w9;
assign w1860 = ~w1858 & ~w1859;
assign w1861 = (w1860 & ~w1857) | (w1860 & w2370) | (~w1857 & w2370);
assign w1862 = w1857 & w2371;
assign w1863 = ~w1861 & ~w1862;
assign w1864 = ~w1067 & ~w1069;
assign w1865 = ~w1092 & ~w1864;
assign w1866 = ~w1045 & ~w1097;
assign w1867 = w1065 & w1866;
assign w1868 = ~w1865 & ~w1867;
assign w1869 = ~w1060 & ~w1868;
assign w1870 = ~w1076 & ~w1106;
assign w1871 = w1038 & ~w1870;
assign w1872 = (w1060 & w1097) | (w1060 & w2422) | (w1097 & w2422);
assign w1873 = ~w1092 & ~w1872;
assign w1874 = ~w1871 & w1873;
assign w1875 = (w1092 & w1068) | (w1092 & w2372) | (w1068 & w2372);
assign w1876 = w1718 & w1875;
assign w1877 = ~w1874 & ~w1876;
assign w1878 = pi143 & ~w9;
assign w1879 = ~pi204 & w9;
assign w1880 = ~w1878 & ~w1879;
assign w1881 = (w1880 & w1877) | (w1880 & w2423) | (w1877 & w2423);
assign w1882 = ~w1877 & w2424;
assign w1883 = ~w1881 & ~w1882;
assign w1884 = ~w1180 & w1683;
assign w1885 = w1149 & w1232;
assign w1886 = ~w1185 & ~w1229;
assign w1887 = ~w1885 & w1886;
assign w1888 = ~w1884 & w1887;
assign w1889 = ~w1201 & w1678;
assign w1890 = ~w1240 & ~w1889;
assign w1891 = (w1229 & ~w1149) | (w1229 & w2373) | (~w1149 & w2373);
assign w1892 = w1890 & w1891;
assign w1893 = ~w1198 & ~w1888;
assign w1894 = ~w1892 & w1893;
assign w1895 = w1201 & w1690;
assign w1896 = ~w1184 & ~w1229;
assign w1897 = w1198 & w1203;
assign w1898 = w1896 & w1897;
assign w1899 = ~w1216 & ~w1239;
assign w1900 = ~w1200 & w1241;
assign w1901 = ~w1899 & w1900;
assign w1902 = w1198 & w1239;
assign w1903 = ~w1896 & w1902;
assign w1904 = ~w1206 & ~w1229;
assign w1905 = ~w1239 & w1904;
assign w1906 = w1890 & w1905;
assign w1907 = ~w1895 & ~w1898;
assign w1908 = ~w1901 & ~w1903;
assign w1909 = w1907 & w1908;
assign w1910 = ~w1906 & w1909;
assign w1911 = ~w1894 & w1910;
assign w1912 = pi126 & ~w9;
assign w1913 = ~pi224 & w9;
assign w1914 = ~w1912 & ~w1913;
assign w1915 = ~w1911 & w1914;
assign w1916 = w1911 & ~w1914;
assign w1917 = ~w1915 & ~w1916;
assign w1918 = w1516 & ~w1532;
assign w1919 = ~w1502 & w1517;
assign w1920 = ~w1521 & ~w1782;
assign w1921 = (~w1518 & w1919) | (~w1518 & w2289) | (w1919 & w2289);
assign w1922 = w1796 & ~w1801;
assign w1923 = ~w1516 & ~w1793;
assign w1924 = ~w1922 & w1923;
assign w1925 = (~w1545 & w1921) | (~w1545 & w2374) | (w1921 & w2374);
assign w1926 = ~w1504 & w1787;
assign w1927 = w1525 & ~w1926;
assign w1928 = ~w1520 & ~w1927;
assign w1929 = ~w1464 & w1781;
assign w1930 = (w1545 & w1928) | (w1545 & w2425) | (w1928 & w2425);
assign w1931 = ~w1918 & ~w1925;
assign w1932 = pi144 & ~w9;
assign w1933 = ~pi210 & w9;
assign w1934 = ~w1932 & ~w1933;
assign w1935 = (w1934 & ~w1931) | (w1934 & w2426) | (~w1931 & w2426);
assign w1936 = w1931 & w2427;
assign w1937 = ~w1935 & ~w1936;
assign w1938 = w1553 & w1780;
assign w1939 = ~w1548 & w1559;
assign w1940 = ~w1516 & ~w1781;
assign w1941 = ~w1549 & w1940;
assign w1942 = (~w1941 & w1938) | (~w1941 & w2428) | (w1938 & w2428);
assign w1943 = w1464 & ~w1516;
assign w1944 = w1450 & w1501;
assign w1945 = ~w1943 & ~w1944;
assign w1946 = w1796 & w1945;
assign w1947 = (~w1516 & ~w1794) | (~w1516 & w2429) | (~w1794 & w2429);
assign w1948 = ~w1545 & ~w1782;
assign w1949 = w1550 & w1948;
assign w1950 = ~w1946 & w1949;
assign w1951 = ~w1947 & w1950;
assign w1952 = ~w1516 & w1922;
assign w1953 = ~w1945 & ~w1952;
assign w1954 = w1497 & w1522;
assign w1955 = ~w1531 & w1545;
assign w1956 = ~w1954 & w1955;
assign w1957 = ~w1953 & w1956;
assign w1958 = ~w1951 & ~w1957;
assign w1959 = pi156 & ~w9;
assign w1960 = ~pi232 & w9;
assign w1961 = ~w1959 & ~w1960;
assign w1962 = ~w1958 & w2430;
assign w1963 = (w1961 & w1958) | (w1961 & w2431) | (w1958 & w2431);
assign w1964 = ~w1962 & ~w1963;
assign w1965 = w1241 & w2432;
assign w1966 = (w2214 & w2375) | (w2214 & w2376) | (w2375 & w2376);
assign w1967 = ~w1206 & w1233;
assign w1968 = ~w1211 & w1967;
assign w1969 = ~w1179 & w1198;
assign w1970 = ~w1674 & w1969;
assign w1971 = w1891 & ~w1968;
assign w1972 = ~w1970 & w1971;
assign w1973 = ~w1966 & ~w1972;
assign w1974 = w1184 & ~w1203;
assign w1975 = w1212 & ~w1229;
assign w1976 = (~w1198 & w1975) | (~w1198 & w2433) | (w1975 & w2433);
assign w1977 = w1232 & w1690;
assign w1978 = w1202 & w1691;
assign w1979 = w1231 & w1978;
assign w1980 = ~w1965 & ~w1977;
assign w1981 = ~w1979 & w1980;
assign w1982 = ~w1973 & w2377;
assign w1983 = pi153 & ~w9;
assign w1984 = ~pi212 & w9;
assign w1985 = ~w1983 & ~w1984;
assign w1986 = ~w1982 & w1985;
assign w1987 = w1982 & ~w1985;
assign w1988 = ~w1986 & ~w1987;
assign w1989 = ~w6 & ~w334;
assign w1990 = ~w751 & ~w1989;
assign w1991 = ~pi193 & ~w1990;
assign w1992 = w8 & ~w330;
assign w1993 = w6 & ~w786;
assign w1994 = w20 & ~w790;
assign w1995 = ~w1992 & ~w1993;
assign w1996 = ~w1994 & w1995;
assign w1997 = pi193 & ~w1996;
assign w1998 = ~w1991 & ~w1997;
assign w1999 = ~w6 & ~w254;
assign w2000 = ~w1298 & ~w1999;
assign w2001 = ~pi193 & ~w2000;
assign w2002 = w8 & ~w250;
assign w2003 = w20 & ~w769;
assign w2004 = ~w402 & ~w2002;
assign w2005 = ~w2003 & w2004;
assign w2006 = pi193 & ~w2005;
assign w2007 = ~w2001 & ~w2006;
assign w2008 = ~w1283 & ~w1993;
assign w2009 = ~pi193 & ~w2008;
assign w2010 = w8 & ~w291;
assign w2011 = w20 & ~w277;
assign w2012 = ~w314 & ~w2010;
assign w2013 = ~w2011 & w2012;
assign w2014 = pi193 & ~w2013;
assign w2015 = ~w2009 & ~w2014;
assign w2016 = ~w6 & ~w109;
assign w2017 = ~w1164 & ~w2016;
assign w2018 = ~pi193 & ~w2017;
assign w2019 = w8 & ~w118;
assign w2020 = w20 & ~w188;
assign w2021 = ~w1488 & ~w2019;
assign w2022 = ~w2020 & w2021;
assign w2023 = pi193 & ~w2022;
assign w2024 = ~w2018 & ~w2023;
assign w2025 = ~w6 & ~w12;
assign w2026 = ~w76 & ~w2025;
assign w2027 = ~pi193 & ~w2026;
assign w2028 = w8 & ~w16;
assign w2029 = w20 & ~w27;
assign w2030 = ~w505 & ~w2028;
assign w2031 = ~w2029 & w2030;
assign w2032 = pi193 & ~w2031;
assign w2033 = ~w2027 & ~w2032;
assign w2034 = ~w365 & ~w1311;
assign w2035 = ~pi193 & ~w2034;
assign w2036 = w8 & ~w341;
assign w2037 = w20 & ~w327;
assign w2038 = ~w1049 & ~w2036;
assign w2039 = ~w2037 & w2038;
assign w2040 = pi193 & ~w2039;
assign w2041 = ~w2035 & ~w2040;
assign w2042 = ~w6 & ~w1138;
assign w2043 = ~w522 & ~w2042;
assign w2044 = ~pi193 & ~w2043;
assign w2045 = w8 & ~w50;
assign w2046 = w20 & ~w43;
assign w2047 = ~w90 & ~w2045;
assign w2048 = ~w2046 & w2047;
assign w2049 = pi193 & ~w2048;
assign w2050 = ~w2044 & ~w2049;
assign w2051 = ~w6 & ~w462;
assign w2052 = ~w1451 & ~w2051;
assign w2053 = ~pi193 & ~w2052;
assign w2054 = w8 & ~w81;
assign w2055 = w20 & ~w75;
assign w2056 = ~w13 & ~w2054;
assign w2057 = ~w2055 & w2056;
assign w2058 = pi193 & ~w2057;
assign w2059 = ~w2053 & ~w2058;
assign w2060 = ~pi066 & ~pi081;
assign w2061 = ~w0 & ~w2060;
assign w2062 = ~pi068 & ~w0;
assign w2063 = ~w1 & ~w8;
assign w2064 = ~w2062 & w2063;
assign w2065 = ~pi069 & ~w1;
assign w2066 = ~w2 & ~w8;
assign w2067 = ~w2065 & w2066;
assign w2068 = ~pi081 & w2066;
assign w2069 = ~w9 & ~w2068;
assign w2070 = pi082 & ~w8;
assign w2071 = ~w46 & ~w2070;
assign w2072 = ~pi082 & w46;
assign w2073 = pi068 & pi069;
assign w2074 = pi192 & pi307;
assign w2075 = ~pi192 & pi037;
assign w2076 = pi192 & pi300;
assign w2077 = ~pi192 & pi048;
assign w2078 = pi192 & pi286;
assign w2079 = ~pi192 & pi065;
assign w2080 = pi192 & pi293;
assign w2081 = ~pi192 & pi045;
assign w2082 = pi192 & pi279;
assign w2083 = pi192 & pi294;
assign w2084 = ~pi192 & pi078;
assign w2085 = pi192 & pi308;
assign w2086 = ~pi192 & pi039;
assign w2087 = pi192 & pi301;
assign w2088 = pi192 & pi267;
assign w2089 = ~pi192 & pi083;
assign w2090 = ~pi192 & pi059;
assign w2091 = pi192 & pi260;
assign w2092 = pi192 & pi259;
assign w2093 = ~pi192 & pi074;
assign w2094 = pi192 & pi273;
assign w2095 = ~pi192 & pi041;
assign w2096 = pi192 & pi266;
assign w2097 = pi192 & pi287;
assign w2098 = ~pi192 & pi076;
assign w2099 = pi192 & pi280;
assign w2100 = ~pi192 & pi091;
assign w2101 = ~pi192 & pi047;
assign w2102 = pi192 & pi303;
assign w2103 = ~pi192 & pi061;
assign w2104 = pi192 & pi310;
assign w2105 = ~pi192 & pi035;
assign w2106 = pi192 & pi296;
assign w2107 = pi192 & pi265;
assign w2108 = ~pi192 & pi053;
assign w2109 = pi192 & pi258;
assign w2110 = ~pi192 & pi072;
assign w2111 = pi192 & pi295;
assign w2112 = ~pi192 & pi077;
assign w2113 = pi192 & pi302;
assign w2114 = ~pi192 & pi092;
assign w2115 = pi192 & pi288;
assign w2116 = ~pi192 & pi054;
assign w2117 = pi192 & pi274;
assign w2118 = ~pi192 & pi042;
assign w2119 = pi192 & pi281;
assign w2120 = pi192 & pi309;
assign w2121 = ~pi192 & pi088;
assign w2122 = pi192 & pi277;
assign w2123 = ~pi192 & pi033;
assign w2124 = pi192 & pi263;
assign w2125 = ~pi192 & pi036;
assign w2126 = pi192 & pi270;
assign w2127 = ~pi192 & pi073;
assign w2128 = pi192 & pi284;
assign w2129 = ~pi192 & pi044;
assign w2130 = pi192 & pi291;
assign w2131 = ~pi192 & pi089;
assign w2132 = pi192 & pi262;
assign w2133 = ~pi192 & pi079;
assign w2134 = pi192 & pi312;
assign w2135 = ~pi192 & pi057;
assign w2136 = pi192 & pi305;
assign w2137 = ~pi192 & pi034;
assign w2138 = pi192 & pi269;
assign w2139 = ~pi192 & pi055;
assign w2140 = pi192 & pi276;
assign w2141 = ~pi192 & pi085;
assign w2142 = pi192 & pi298;
assign w2143 = ~pi192 & pi067;
assign w2144 = pi192 & pi311;
assign w2145 = ~pi192 & pi032;
assign w2146 = pi192 & pi297;
assign w2147 = ~pi192 & pi070;
assign w2148 = pi192 & pi304;
assign w2149 = ~pi192 & pi038;
assign w2150 = pi192 & pi261;
assign w2151 = ~pi192 & pi052;
assign w2152 = pi192 & pi268;
assign w2153 = ~pi192 & pi046;
assign w2154 = pi192 & pi264;
assign w2155 = ~pi192 & pi051;
assign w2156 = pi192 & pi275;
assign w2157 = ~pi192 & pi084;
assign w2158 = pi192 & pi282;
assign w2159 = ~pi192 & pi043;
assign w2160 = pi192 & pi271;
assign w2161 = ~pi192 & pi086;
assign w2162 = pi192 & pi278;
assign w2163 = ~pi192 & pi087;
assign w2164 = pi192 & pi306;
assign w2165 = ~pi192 & pi063;
assign w2166 = pi192 & pi299;
assign w2167 = ~pi192 & pi049;
assign w2168 = pi192 & pi292;
assign w2169 = ~pi192 & pi062;
assign w2170 = pi192 & pi285;
assign w2171 = ~pi192 & pi090;
assign w2172 = pi192 & pi272;
assign w2173 = ~pi192 & pi056;
assign w2174 = pi192 & pi290;
assign w2175 = ~pi192 & pi080;
assign w2176 = w1139 & pi193;
assign w2177 = ~w2099 & pi193;
assign w2178 = ~w6 & ~pi193;
assign w2179 = ~w1159 & w570;
assign w2180 = w1159 & ~w570;
assign w2181 = ~pi192 & pi075;
assign w2182 = ~w2107 & pi193;
assign w2183 = ~pi192 & pi071;
assign w2184 = ~w1175 & w531;
assign w2185 = w1175 & ~w531;
assign w2186 = w1185 & w1198;
assign w2187 = w1148 & ~w1203;
assign w2188 = ~w6 & pi193;
assign w2189 = w6 & ~pi193;
assign w2190 = ~w1273 & w759;
assign w2191 = w1273 & ~w759;
assign w2192 = w1284 & pi193;
assign w2193 = ~w1321 & w1340;
assign w2194 = ~w852 & w819;
assign w2195 = ~w2088 & pi193;
assign w2196 = ~w1446 & w37;
assign w2197 = w1446 & ~w37;
assign w2198 = ~w2083 & pi193;
assign w2199 = ~w1460 & w201;
assign w2200 = w1460 & ~w201;
assign w2201 = ~pi192 & pi064;
assign w2202 = ~w2074 & pi193;
assign w2203 = ~w1475 & w1479;
assign w2204 = w1475 & ~w1479;
assign w2205 = w191 & w6;
assign w2206 = ~w1490 & w1494;
assign w2207 = w1490 & ~w1494;
assign w2208 = ~w1575 & ~w1570;
assign w2209 = w892 & w781;
assign w2210 = w1637 & ~w762;
assign w2211 = w864 & w2434;
assign w2212 = (w880 & w867) | (w880 & w2435) | (w867 & w2435);
assign w2213 = w1077 & w1092;
assign w2214 = ~w1678 & ~w1229;
assign w2215 = ~w1676 & w2436;
assign w2216 = ~w1104 & w1060;
assign w2217 = w1709 & ~w1092;
assign w2218 = w1034 & w1015;
assign w2219 = ~w1575 & w1306;
assign w2220 = ~w31 & w2290;
assign w2221 = ~w2085 & pi193;
assign w2222 = ~w65 & w69;
assign w2223 = w65 & ~w69;
assign w2224 = ~w2094 & pi193;
assign w2225 = ~w96 & w100;
assign w2226 = w96 & ~w100;
assign w2227 = (w136 & ~w131) | (w136 & w2291) | (~w131 & w2291);
assign w2228 = w131 & w2292;
assign w2229 = ~w6 & w7;
assign w2230 = w155 & pi193;
assign w2231 = ~pi192 & pi040;
assign w2232 = pi192 & pi289;
assign w2233 = ~w8 & pi193;
assign w2234 = ~w267 & w271;
assign w2235 = w267 & ~w271;
assign w2236 = ~w297 & w301;
assign w2237 = w297 & ~w301;
assign w2238 = ~w316 & w320;
assign w2239 = w316 & ~w320;
assign w2240 = ~w347 & w351;
assign w2241 = w347 & ~w351;
assign w2242 = ~w381 & w385;
assign w2243 = w381 & ~w385;
assign w2244 = ~w2097 & pi193;
assign w2245 = ~w473 & w477;
assign w2246 = w473 & ~w477;
assign w2247 = ~pi192 & pi058;
assign w2248 = ~w2120 & pi193;
assign w2249 = ~w489 & w493;
assign w2250 = w489 & ~w493;
assign w2251 = ~w2172 & pi193;
assign w2252 = ~w508 & w512;
assign w2253 = w508 & ~w512;
assign w2254 = ~w2092 & pi193;
assign w2255 = ~w546 & w550;
assign w2256 = w546 & ~w550;
assign w2257 = w753 & pi193;
assign w2258 = ~pi192 & pi050;
assign w2259 = pi192 & pi313;
assign w2260 = ~pi192 & pi060;
assign w2261 = pi192 & pi283;
assign w2262 = ~w277 & w2290;
assign w2263 = w810 & pi193;
assign w2264 = w826 & pi193;
assign w2265 = ~w375 & w2290;
assign w2266 = ~w980 & w422;
assign w2267 = w980 & ~w422;
assign w2268 = ~w992 & w996;
assign w2269 = w992 & ~w996;
assign w2270 = ~w1008 & w1012;
assign w2271 = w1008 & ~w1012;
assign w2272 = ~w1029 & w385;
assign w2273 = w1029 & ~w385;
assign w2274 = w1066 & w1071;
assign w2275 = w191 & ~w6;
assign w2276 = w1124 & pi193;
assign w2277 = w1192 & pi193;
assign w2278 = ~w1261 & w778;
assign w2279 = w1261 & ~w778;
assign w2280 = w1300 & pi193;
assign w2281 = w1312 & pi193;
assign w2282 = w1334 & pi193;
assign w2283 = w1510 & pi193;
assign w2284 = w1532 & ~w1533;
assign w2285 = w1482 & w1497;
assign w2286 = ~w1450 & ~w1497;
assign w2287 = ~w1210 & w1198;
assign w2288 = ~w1482 & w1464;
assign w2289 = ~w1920 & ~w1518;
assign w2290 = w6 & pi193;
assign w2291 = w130 & w136;
assign w2292 = ~w130 & ~w136;
assign w2293 = w177 & ~w40;
assign w2294 = w274 & w388;
assign w2295 = w416 & pi193;
assign w2296 = w389 & ~w434;
assign w2297 = w525 & pi193;
assign w2298 = ~w220 & ~w624;
assign w2299 = w628 & ~w619;
assign w2300 = w681 & ~w534;
assign w2301 = w772 & pi193;
assign w2302 = ~w852 & ~w820;
assign w2303 = ~w861 & w871;
assign w2304 = ~w883 & ~w901;
assign w2305 = w918 & ~w425;
assign w2306 = ~w437 & w923;
assign w2307 = w354 & ~w274;
assign w2308 = w927 & w425;
assign w2309 = ~w305 & w431;
assign w2310 = ~w963 & ~w969;
assign w2311 = w963 & w969;
assign w2312 = w1045 & ~w1033;
assign w2313 = w1054 & pi193;
assign w2314 = ~w984 & w1060;
assign w2315 = w1074 & ~w1077;
assign w2316 = w1019 & w1074;
assign w2317 = w1098 & w1092;
assign w2318 = ~w1104 & ~w1060;
assign w2319 = ~w1105 & ~w1092;
assign w2320 = w1223 & pi193;
assign w2321 = ~w1219 & ~w1229;
assign w2322 = w1148 & ~w1239;
assign w2323 = w1240 & ~w1198;
assign w2324 = w1230 & w1250;
assign w2325 = ~w1230 & ~w1250;
assign w2326 = ~w1321 & ~w1306;
assign w2327 = ~w1342 & w1340;
assign w2328 = ~w1321 & ~w1324;
assign w2329 = ~w1379 & ~w1383;
assign w2330 = w1379 & w1383;
assign w2331 = w927 & w390;
assign w2332 = ~w1417 & ~w1433;
assign w2333 = w1417 & w1433;
assign w2334 = w1539 & pi193;
assign w2335 = w1520 & w2437;
assign w2336 = w1552 & w1516;
assign w2337 = (~w1545 & w1529) | (~w1545 & w2438) | (w1529 & w2438);
assign w2338 = ~w1578 & ~w1573;
assign w2339 = w1340 & w1594;
assign w2340 = ~w1579 & w2439;
assign w2341 = (~w1599 & w1579) | (~w1599 & w2440) | (w1579 & w2440);
assign w2342 = w1636 & ~w781;
assign w2343 = w858 & ~w1641;
assign w2344 = ~w1643 & ~w762;
assign w2345 = ~w1643 & w1647;
assign w2346 = (~w2345 & w2441) | (~w2345 & w2442) | (w2441 & w2442);
assign w2347 = (w2345 & w2443) | (w2345 & w2444) | (w2443 & w2444);
assign w2348 = w1662 & ~w1092;
assign w2349 = ~w1679 & ~w1229;
assign w2350 = ~w1679 & ~w1202;
assign w2351 = w1212 & w2445;
assign w2352 = w1229 & ~w1694;
assign w2353 = ~w1696 & w1699;
assign w2354 = w1696 & ~w1699;
assign w2355 = ~w1714 & w2446;
assign w2356 = (~w1727 & w1714) | (~w1727 & w2447) | (w1714 & w2447);
assign w2357 = ~w1734 & ~w762;
assign w2358 = w1349 & ~w1340;
assign w2359 = w1764 & ~w1371;
assign w2360 = w1761 & w1775;
assign w2361 = ~w1761 & ~w1775;
assign w2362 = w1548 & ~w1793;
assign w2363 = ~w1549 & ~w1812;
assign w2364 = w1549 & w1812;
assign w2365 = ~w205 & ~w620;
assign w2366 = w1820 & ~w40;
assign w2367 = ~w1340 & ~w1842;
assign w2368 = w1368 & ~w1340;
assign w2369 = ~w1293 & ~w1340;
assign w2370 = ~w1843 & w2448;
assign w2371 = (~w1860 & w1843) | (~w1860 & w2449) | (w1843 & w2449);
assign w2372 = ~w1706 & w1092;
assign w2373 = ~w1232 & w1229;
assign w2374 = w1924 & ~w1545;
assign w2375 = ~w1897 & ~w1229;
assign w2376 = ~w1897 & ~w1202;
assign w2377 = w1981 & ~w1976;
assign w2378 = w179 & ~w180;
assign w2379 = w103 & ~w104;
assign w2380 = w220 & ~w210;
assign w2381 = ~w219 & ~w222;
assign w2382 = ~w442 & ~w448;
assign w2383 = ~w553 & ~w480;
assign w2384 = w179 & ~w230;
assign w2385 = w175 & w633;
assign w2386 = ~w172 & w220;
assign w2387 = ~w630 & w632;
assign w2388 = ~w103 & ~w176;
assign w2389 = (~w670 & w650) | (~w670 & w2450) | (w650 & w2450);
assign w2390 = ~w650 & w2451;
assign w2391 = w515 & w553;
assign w2392 = w678 & ~w573;
assign w2393 = ~w480 & w553;
assign w2394 = w683 & w573;
assign w2395 = ~w573 & ~w553;
assign w2396 = ~w717 & w2452;
assign w2397 = w856 & ~w783;
assign w2398 = w857 & ~w782;
assign w2399 = ~w762 & w874;
assign w2400 = ~w873 & ~w908;
assign w2401 = w873 & w908;
assign w2402 = ~w438 & ~w425;
assign w2403 = w933 & w938;
assign w2404 = ~w933 & ~w938;
assign w2405 = w912 & ~w438;
assign w2406 = w958 & ~w425;
assign w2407 = ~w1015 & ~w984;
assign w2408 = w999 & ~w1015;
assign w2409 = ~w1378 & w1306;
assign w2410 = w438 & w388;
assign w2411 = w1388 & w425;
assign w2412 = ~w388 & ~w1394;
assign w2413 = w1397 & ~w425;
assign w2414 = w1391 & w1407;
assign w2415 = ~w1391 & ~w1407;
assign w2416 = w515 & ~w534;
assign w2417 = w2213 & w1092;
assign w2418 = (w1092 & w2213) | (w1092 & ~w1074) | (w2213 & ~w1074);
assign w2419 = w1654 & w1669;
assign w2420 = ~w1654 & ~w1669;
assign w2421 = ~w1760 & ~w1306;
assign w2422 = w1045 & w1060;
assign w2423 = w1869 & w1880;
assign w2424 = ~w1869 & ~w1880;
assign w2425 = w1929 & w1545;
assign w2426 = w1930 & w1934;
assign w2427 = ~w1930 & ~w1934;
assign w2428 = ~w1939 & ~w1941;
assign w2429 = w1802 & ~w1516;
assign w2430 = ~w1942 & ~w1961;
assign w2431 = w1942 & w1961;
assign w2432 = w1181 & ~w1133;
assign w2433 = w1974 & ~w1198;
assign w2434 = ~w819 & w781;
assign w2435 = w762 & w2211;
assign w2436 = ~w1673 & ~w1198;
assign w2437 = ~w1500 & w1545;
assign w2438 = w1531 & ~w1545;
assign w2439 = w1306 & w1599;
assign w2440 = ~w1306 & ~w1599;
assign w2441 = w1650 & w2212;
assign w2442 = w1650 & ~w2344;
assign w2443 = ~w1650 & ~w2212;
assign w2444 = ~w1650 & w2344;
assign w2445 = ~w1133 & w1198;
assign w2446 = w1092 & w1727;
assign w2447 = ~w1092 & ~w1727;
assign w2448 = ~w1306 & w1860;
assign w2449 = w1306 & ~w1860;
assign w2450 = w621 & ~w670;
assign w2451 = ~w621 & w670;
assign w2452 = ~w516 & w573;
assign one = 1;
assign po000 = pi170;// level 0
assign po001 = pi119;// level 0
assign po002 = pi186;// level 0
assign po003 = pi098;// level 0
assign po004 = pi165;// level 0
assign po005 = pi120;// level 0
assign po006 = pi184;// level 0
assign po007 = pi096;// level 0
assign po008 = pi174;// level 0
assign po009 = pi134;// level 0
assign po010 = pi162;// level 0
assign po011 = pi106;// level 0
assign po012 = pi183;// level 0
assign po013 = pi112;// level 0
assign po014 = pi163;// level 0
assign po015 = pi133;// level 0
assign po016 = pi168;// level 0
assign po017 = pi105;// level 0
assign po018 = pi158;// level 0
assign po019 = pi122;// level 0
assign po020 = pi181;// level 0
assign po021 = pi102;// level 0
assign po022 = pi173;// level 0
assign po023 = pi117;// level 0
assign po024 = pi175;// level 0
assign po025 = pi124;// level 0
assign po026 = pi189;// level 0
assign po027 = pi110;// level 0
assign po028 = pi160;// level 0
assign po029 = pi103;// level 0
assign po030 = pi188;// level 0
assign po031 = pi095;// level 0
assign po032 = pi172;// level 0
assign po033 = pi115;// level 0
assign po034 = pi171;// level 0
assign po035 = pi107;// level 0
assign po036 = pi166;// level 0
assign po037 = pi116;// level 0
assign po038 = pi169;// level 0
assign po039 = pi132;// level 0
assign po040 = pi182;// level 0
assign po041 = pi101;// level 0
assign po042 = pi159;// level 0
assign po043 = pi104;// level 0
assign po044 = pi161;// level 0
assign po045 = pi111;// level 0
assign po046 = pi167;// level 0
assign po047 = pi109;// level 0
assign po048 = pi179;// level 0
assign po049 = pi094;// level 0
assign po050 = pi164;// level 0
assign po051 = pi113;// level 0
assign po052 = pi176;// level 0
assign po053 = pi100;// level 0
assign po054 = pi185;// level 0
assign po055 = pi097;// level 0
assign po056 = pi178;// level 0
assign po057 = pi118;// level 0
assign po058 = pi187;// level 0
assign po059 = pi108;// level 0
assign po060 = pi177;// level 0
assign po061 = pi114;// level 0
assign po062 = pi180;// level 0
assign po063 = pi099;// level 0
assign po064 = pi093;// level 0
assign po065 = pi191;// level 0
assign po066 = one;// level 0
assign po067 = pi190;// level 0
assign po068 = w244;// level 19
assign po069 = w460;// level 19
assign po070 = w618;// level 19
assign po071 = w647;// level 19
assign po072 = w673;// level 19
assign po073 = w715;// level 19
assign po074 = w746;// level 19
assign po075 = w911;// level 19
assign po076 = w941;// level 18
assign po077 = w972;// level 19
assign po078 = ~w1119;// level 19
assign po079 = ~w1253;// level 19
assign po080 = ~w1386;// level 19
assign po081 = w1410;// level 18
assign po082 = w1436;// level 19
assign po083 = w1569;// level 19
assign po084 = w1602;// level 19
assign po085 = w1632;// level 19
assign po086 = w1653;// level 19
assign po087 = w1672;// level 18
assign po088 = ~w1702;// level 19
assign po089 = w1730;// level 19
assign po090 = w1749;// level 19
assign po091 = ~w1778;// level 19
assign po092 = w1815;// level 19
assign po093 = w1839;// level 19
assign po094 = ~w1863;// level 19
assign po095 = w1883;// level 18
assign po096 = w1917;// level 19
assign po097 = w1937;// level 18
assign po098 = ~w1964;// level 18
assign po099 = w1988;// level 19
assign po100 = ~w1998;// level 9
assign po101 = ~w2007;// level 9
assign po102 = ~w2015;// level 9
assign po103 = ~w2024;// level 9
assign po104 = ~w1089;// level 9
assign po105 = ~w2033;// level 9
assign po106 = ~w2041;// level 9
assign po107 = ~w2050;// level 9
assign po108 = ~w198;// level 9
assign po109 = ~w2059;// level 9
assign po110 = ~w1226;// level 8
assign po111 = ~w1337;// level 8
assign po112 = ~w1303;// level 8
assign po113 = ~w1542;// level 8
assign po114 = w382;// level 8
assign po115 = ~w567;// level 9
assign po116 = ~w1195;// level 8
assign po117 = ~w419;// level 8
assign po118 = ~w775;// level 8
assign po119 = ~w1315;// level 8
assign po120 = ~w756;// level 8
assign po121 = ~w1513;// level 8
assign po122 = ~w528;// level 8
assign po123 = ~w798;// level 8
assign po124 = ~w1057;// level 8
assign po125 = w993;// level 8
assign po126 = w490;// level 8
assign po127 = ~w1142;// level 8
assign po128 = ~w1287;// level 8
assign po129 = w133;// level 9
assign po130 = ~w846;// level 8
assign po131 = w1009;// level 8
assign po132 = w1476;// level 8
assign po133 = ~w34;// level 8
assign po134 = w2061;// level 2
assign po135 = w348;// level 8
assign po136 = w2064;// level 4
assign po137 = w2067;// level 4
assign po138 = ~w829;// level 8
assign po139 = w509;// level 8
assign po140 = w1491;// level 8
assign po141 = ~w813;// level 8
assign po142 = w547;// level 8
assign po143 = w1176;// level 8
assign po144 = w474;// level 8
assign po145 = ~w1127;// level 8
assign po146 = w1461;// level 8
assign po147 = w1274;// level 8
assign po148 = w66;// level 8
assign po149 = ~w2069;// level 5
assign po150 = ~w2071;// level 4
assign po151 = w1447;// level 8
assign po152 = w981;// level 8
assign po153 = w317;// level 8
assign po154 = w1030;// level 8
assign po155 = w1262;// level 8
assign po156 = w268;// level 8
assign po157 = w298;// level 8
assign po158 = w97;// level 8
assign po159 = w1160;// level 8
assign po160 = ~w166;// level 8
assign po161 = w2072;// level 4
assign po162 = ~pi130;// level 0
assign po163 = ~pi126;// level 0
assign po164 = ~pi131;// level 0
assign po165 = ~pi129;// level 0
assign po166 = ~pi127;// level 0
assign po167 = ~pi121;// level 0
assign po168 = ~pi125;// level 0
assign po169 = ~pi128;// level 0
assign po170 = ~pi123;// level 0
assign po171 = ~pi141;// level 0
assign po172 = ~pi139;// level 0
assign po173 = ~pi144;// level 0
assign po174 = ~pi143;// level 0
assign po175 = ~pi140;// level 0
assign po176 = ~pi142;// level 0
assign po177 = ~pi137;// level 0
assign po178 = ~pi138;// level 0
assign po179 = ~pi136;// level 0
assign po180 = ~pi135;// level 0
assign po181 = ~pi145;// level 0
assign po182 = ~pi146;// level 0
assign po183 = ~pi155;// level 0
assign po184 = ~pi148;// level 0
assign po185 = ~pi147;// level 0
assign po186 = ~pi149;// level 0
assign po187 = ~pi152;// level 0
assign po188 = ~pi154;// level 0
assign po189 = ~w832;// level 5
assign po190 = ~pi153;// level 0
assign po191 = ~w849;// level 5
assign po192 = ~pi150;// level 0
assign po193 = ~w1290;// level 5
assign po194 = ~w385;// level 5
assign po195 = ~w493;// level 5
assign po196 = ~w1494;// level 5
assign po197 = ~w1012;// level 5
assign po198 = ~w1479;// level 5
assign po199 = ~w301;// level 5
assign po200 = ~pi156;// level 0
assign po201 = ~pi151;// level 0
assign po202 = ~pi157;// level 0
assign po203 = ~w816;// level 5
assign po204 = ~w1318;// level 5
assign po205 = ~w996;// level 5
assign po206 = ~w531;// level 5
assign po207 = ~w1130;// level 5
assign po208 = ~w570;// level 5
assign po209 = ~w759;// level 5
assign po210 = ~w69;// level 5
assign po211 = ~w512;// level 5
assign po212 = ~w136;// level 5
assign po213 = ~w1145;// level 5
assign po214 = ~w477;// level 5
assign po215 = ~w351;// level 5
assign po216 = ~w778;// level 5
assign po217 = ~w320;// level 5
assign po218 = ~w37;// level 5
assign po219 = ~w271;// level 5
assign po220 = ~w169;// level 5
assign po221 = ~w550;// level 5
assign po222 = ~w801;// level 5
assign po223 = ~w201;// level 5
assign po224 = ~w422;// level 5
assign po225 = ~w100;// level 5
assign po226 = pi031;// level 0
assign po227 = pi000;// level 0
assign po228 = pi025;// level 0
assign po229 = pi005;// level 0
assign po230 = pi027;// level 0
assign po231 = pi019;// level 0
assign po232 = pi001;// level 0
assign po233 = pi008;// level 0
assign po234 = pi010;// level 0
assign po235 = pi022;// level 0
assign po236 = pi029;// level 0
assign po237 = pi030;// level 0
assign po238 = pi017;// level 0
assign po239 = pi024;// level 0
assign po240 = pi020;// level 0
assign po241 = pi002;// level 0
assign po242 = pi026;// level 0
assign po243 = pi021;// level 0
assign po244 = pi015;// level 0
assign po245 = pi014;// level 0
assign po246 = pi003;// level 0
assign po247 = pi009;// level 0
assign po248 = pi006;// level 0
assign po249 = pi011;// level 0
assign po250 = pi018;// level 0
assign po251 = pi016;// level 0
assign po252 = pi023;// level 0
assign po253 = pi004;// level 0
assign po254 = pi013;// level 0
assign po255 = pi007;// level 0
assign po256 = pi028;// level 0
assign po257 = pi012;// level 0
endmodule
