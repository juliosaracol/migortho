module top (
            pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518, 
            po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142, w7143, w7144, w7145, w7146, w7147, w7148, w7149, w7150, w7151, w7152, w7153, w7154, w7155, w7156, w7157, w7158, w7159, w7160, w7161, w7162, w7163, w7164, w7165, w7166, w7167, w7168, w7169, w7170, w7171, w7172, w7173, w7174, w7175, w7176, w7177, w7178, w7179, w7180, w7181, w7182, w7183, w7184, w7185, w7186, w7187, w7188, w7189, w7190, w7191, w7192, w7193, w7194, w7195, w7196, w7197, w7198, w7199, w7200, w7201, w7202, w7203, w7204, w7205, w7206, w7207, w7208, w7209, w7210, w7211, w7212, w7213, w7214, w7215, w7216, w7217, w7218, w7219, w7220, w7221, w7222, w7223, w7224, w7225, w7226, w7227, w7228, w7229, w7230, w7231, w7232, w7233, w7234, w7235, w7236, w7237, w7238, w7239, w7240, w7241, w7242, w7243, w7244, w7245, w7246, w7247, w7248, w7249, w7250, w7251, w7252, w7253, w7254, w7255, w7256, w7257, w7258, w7259, w7260, w7261, w7262, w7263, w7264, w7265, w7266, w7267, w7268, w7269, w7270, w7271, w7272, w7273, w7274, w7275, w7276, w7277, w7278, w7279, w7280, w7281, w7282, w7283, w7284, w7285, w7286, w7287, w7288, w7289, w7290, w7291, w7292, w7293, w7294, w7295, w7296, w7297, w7298, w7299, w7300, w7301, w7302, w7303, w7304, w7305, w7306, w7307, w7308, w7309, w7310, w7311, w7312, w7313, w7314, w7315, w7316, w7317, w7318, w7319, w7320, w7321, w7322, w7323, w7324, w7325, w7326, w7327, w7328, w7329, w7330, w7331, w7332, w7333, w7334, w7335, w7336, w7337, w7338, w7339, w7340, w7341, w7342, w7343, w7344, w7345, w7346, w7347, w7348, w7349, w7350, w7351, w7352, w7353, w7354, w7355, w7356, w7357, w7358, w7359, w7360, w7361, w7362, w7363, w7364, w7365, w7366, w7367, w7368, w7369, w7370, w7371, w7372, w7373, w7374, w7375, w7376, w7377, w7378, w7379, w7380, w7381, w7382, w7383, w7384, w7385, w7386, w7387, w7388, w7389, w7390, w7391, w7392, w7393, w7394, w7395, w7396, w7397, w7398, w7399, w7400, w7401, w7402, w7403, w7404, w7405, w7406, w7407, w7408, w7409, w7410, w7411, w7412, w7413, w7414, w7415, w7416, w7417, w7418, w7419, w7420, w7421, w7422, w7423, w7424, w7425, w7426, w7427, w7428, w7429, w7430, w7431, w7432, w7433, w7434, w7435, w7436, w7437, w7438, w7439, w7440, w7441, w7442, w7443, w7444, w7445, w7446, w7447, w7448, w7449, w7450, w7451, w7452, w7453, w7454, w7455, w7456, w7457, w7458, w7459, w7460, w7461, w7462, w7463, w7464, w7465, w7466, w7467, w7468, w7469, w7470, w7471, w7472, w7473, w7474, w7475, w7476, w7477, w7478, w7479, w7480, w7481, w7482, w7483, w7484, w7485, w7486, w7487, w7488, w7489, w7490, w7491, w7492, w7493, w7494, w7495, w7496, w7497, w7498, w7499, w7500, w7501, w7502, w7503, w7504, w7505, w7506, w7507, w7508, w7509, w7510, w7511, w7512, w7513, w7514, w7515, w7516, w7517, w7518, w7519, w7520, w7521, w7522, w7523, w7524, w7525, w7526, w7527, w7528, w7529, w7530, w7531, w7532, w7533, w7534, w7535, w7536, w7537, w7538, w7539, w7540, w7541, w7542, w7543, w7544, w7545, w7546, w7547, w7548, w7549, w7550, w7551, w7552, w7553, w7554, w7555, w7556, w7557, w7558, w7559, w7560, w7561, w7562, w7563, w7564, w7565, w7566, w7567, w7568, w7569, w7570, w7571, w7572, w7573, w7574, w7575, w7576, w7577, w7578, w7579, w7580, w7581, w7582, w7583, w7584, w7585, w7586, w7587, w7588, w7589, w7590, w7591, w7592, w7593, w7594, w7595, w7596, w7597, w7598, w7599, w7600, w7601, w7602, w7603, w7604, w7605, w7606, w7607, w7608, w7609, w7610, w7611, w7612, w7613, w7614, w7615, w7616, w7617, w7618, w7619, w7620, w7621, w7622, w7623, w7624, w7625, w7626, w7627, w7628, w7629, w7630, w7631, w7632, w7633, w7634, w7635, w7636, w7637, w7638, w7639, w7640, w7641, w7642, w7643, w7644, w7645, w7646, w7647, w7648, w7649, w7650, w7651, w7652, w7653, w7654, w7655, w7656, w7657, w7658, w7659, w7660, w7661, w7662, w7663, w7664, w7665, w7666, w7667, w7668, w7669, w7670, w7671, w7672, w7673, w7674, w7675, w7676, w7677, w7678, w7679, w7680, w7681, w7682, w7683, w7684, w7685, w7686, w7687, w7688, w7689, w7690, w7691, w7692, w7693, w7694, w7695, w7696, w7697, w7698, w7699, w7700, w7701, w7702, w7703, w7704, w7705, w7706, w7707, w7708, w7709, w7710, w7711, w7712, w7713, w7714, w7715, w7716, w7717, w7718, w7719, w7720, w7721, w7722, w7723, w7724, w7725, w7726, w7727, w7728, w7729, w7730, w7731, w7732, w7733, w7734, w7735, w7736, w7737, w7738, w7739, w7740, w7741, w7742, w7743, w7744, w7745, w7746, w7747, w7748, w7749, w7750, w7751, w7752, w7753, w7754, w7755, w7756, w7757, w7758, w7759, w7760, w7761, w7762, w7763, w7764, w7765, w7766, w7767, w7768, w7769, w7770, w7771, w7772, w7773, w7774, w7775, w7776, w7777, w7778, w7779, w7780, w7781, w7782, w7783, w7784, w7785, w7786, w7787, w7788, w7789, w7790, w7791, w7792, w7793, w7794, w7795, w7796, w7797, w7798, w7799, w7800, w7801, w7802, w7803, w7804, w7805, w7806, w7807, w7808, w7809, w7810, w7811, w7812, w7813, w7814, w7815, w7816, w7817, w7818, w7819, w7820, w7821, w7822, w7823, w7824, w7825, w7826, w7827, w7828, w7829, w7830, w7831, w7832, w7833, w7834, w7835, w7836, w7837, w7838, w7839, w7840, w7841, w7842, w7843, w7844, w7845, w7846, w7847, w7848, w7849, w7850, w7851, w7852, w7853, w7854, w7855, w7856, w7857, w7858, w7859, w7860, w7861, w7862, w7863, w7864, w7865, w7866, w7867, w7868, w7869, w7870, w7871, w7872, w7873, w7874, w7875, w7876, w7877, w7878, w7879, w7880, w7881, w7882, w7883, w7884, w7885, w7886, w7887, w7888, w7889, w7890, w7891, w7892, w7893, w7894, w7895, w7896, w7897, w7898, w7899, w7900, w7901, w7902, w7903, w7904, w7905, w7906, w7907, w7908, w7909, w7910, w7911, w7912, w7913, w7914, w7915, w7916, w7917, w7918, w7919, w7920, w7921, w7922, w7923, w7924, w7925, w7926, w7927, w7928, w7929, w7930, w7931, w7932, w7933, w7934, w7935, w7936, w7937, w7938, w7939, w7940, w7941, w7942, w7943, w7944, w7945, w7946, w7947, w7948, w7949, w7950, w7951, w7952, w7953, w7954, w7955, w7956, w7957, w7958, w7959, w7960, w7961, w7962, w7963, w7964, w7965, w7966, w7967, w7968, w7969, w7970, w7971, w7972, w7973, w7974, w7975, w7976, w7977, w7978, w7979, w7980, w7981, w7982, w7983, w7984, w7985, w7986, w7987, w7988, w7989, w7990, w7991, w7992, w7993, w7994, w7995, w7996, w7997, w7998, w7999, w8000, w8001, w8002, w8003, w8004, w8005, w8006, w8007, w8008, w8009, w8010, w8011, w8012, w8013, w8014, w8015, w8016, w8017, w8018, w8019, w8020, w8021, w8022, w8023, w8024, w8025, w8026, w8027, w8028, w8029, w8030, w8031, w8032, w8033, w8034, w8035, w8036, w8037, w8038, w8039, w8040, w8041, w8042, w8043, w8044, w8045, w8046, w8047, w8048, w8049, w8050, w8051, w8052, w8053, w8054, w8055, w8056, w8057, w8058, w8059, w8060, w8061, w8062, w8063, w8064, w8065, w8066, w8067, w8068, w8069, w8070, w8071, w8072, w8073, w8074, w8075, w8076, w8077, w8078, w8079, w8080, w8081, w8082, w8083, w8084, w8085, w8086, w8087, w8088, w8089, w8090, w8091, w8092, w8093, w8094, w8095, w8096, w8097, w8098, w8099, w8100, w8101, w8102, w8103, w8104, w8105, w8106, w8107, w8108, w8109, w8110, w8111, w8112, w8113, w8114, w8115, w8116, w8117, w8118, w8119, w8120, w8121, w8122, w8123, w8124, w8125, w8126, w8127, w8128, w8129, w8130, w8131, w8132, w8133, w8134, w8135, w8136, w8137, w8138, w8139, w8140, w8141, w8142, w8143, w8144, w8145, w8146, w8147, w8148, w8149, w8150, w8151, w8152, w8153, w8154, w8155, w8156, w8157, w8158, w8159, w8160, w8161, w8162, w8163, w8164, w8165, w8166, w8167, w8168, w8169, w8170, w8171, w8172, w8173, w8174, w8175, w8176, w8177, w8178, w8179, w8180, w8181, w8182, w8183, w8184, w8185, w8186, w8187, w8188, w8189, w8190, w8191, w8192, w8193, w8194, w8195, w8196, w8197, w8198, w8199, w8200, w8201, w8202, w8203, w8204, w8205, w8206, w8207, w8208, w8209, w8210, w8211, w8212, w8213, w8214, w8215, w8216, w8217, w8218, w8219, w8220, w8221, w8222, w8223, w8224, w8225, w8226, w8227, w8228, w8229, w8230, w8231, w8232, w8233, w8234, w8235, w8236, w8237, w8238, w8239, w8240, w8241, w8242, w8243, w8244, w8245, w8246, w8247, w8248, w8249, w8250, w8251, w8252, w8253, w8254, w8255, w8256, w8257, w8258, w8259, w8260, w8261, w8262, w8263, w8264, w8265, w8266, w8267, w8268, w8269, w8270, w8271, w8272, w8273, w8274, w8275, w8276, w8277, w8278, w8279, w8280, w8281, w8282, w8283, w8284, w8285, w8286, w8287, w8288, w8289, w8290, w8291, w8292, w8293, w8294, w8295, w8296, w8297, w8298, w8299, w8300, w8301, w8302, w8303, w8304, w8305, w8306, w8307, w8308, w8309, w8310, w8311, w8312, w8313, w8314, w8315, w8316, w8317, w8318, w8319, w8320, w8321, w8322, w8323, w8324, w8325, w8326, w8327, w8328, w8329, w8330, w8331, w8332, w8333, w8334, w8335, w8336, w8337, w8338, w8339, w8340, w8341, w8342, w8343, w8344, w8345, w8346, w8347, w8348, w8349, w8350, w8351, w8352, w8353, w8354, w8355, w8356, w8357, w8358, w8359, w8360, w8361, w8362, w8363, w8364, w8365, w8366, w8367, w8368, w8369, w8370, w8371, w8372, w8373, w8374, w8375, w8376, w8377, w8378, w8379, w8380, w8381, w8382, w8383, w8384, w8385, w8386, w8387, w8388, w8389, w8390, w8391, w8392, w8393, w8394, w8395, w8396, w8397, w8398, w8399, w8400, w8401, w8402, w8403, w8404, w8405, w8406, w8407, w8408, w8409, w8410, w8411, w8412, w8413, w8414, w8415, w8416, w8417, w8418, w8419, w8420, w8421, w8422, w8423, w8424, w8425, w8426, w8427, w8428, w8429, w8430, w8431, w8432, w8433, w8434, w8435, w8436, w8437, w8438, w8439, w8440, w8441, w8442, w8443, w8444, w8445, w8446, w8447, w8448, w8449, w8450, w8451, w8452, w8453, w8454, w8455, w8456, w8457, w8458, w8459, w8460, w8461, w8462, w8463, w8464, w8465, w8466, w8467, w8468, w8469, w8470, w8471, w8472, w8473, w8474, w8475, w8476, w8477, w8478, w8479, w8480, w8481, w8482, w8483, w8484, w8485, w8486, w8487, w8488, w8489, w8490, w8491, w8492, w8493, w8494, w8495, w8496, w8497, w8498, w8499, w8500, w8501, w8502, w8503, w8504, w8505, w8506, w8507, w8508, w8509, w8510, w8511, w8512, w8513, w8514, w8515, w8516, w8517, w8518, w8519, w8520, w8521, w8522, w8523, w8524, w8525, w8526, w8527, w8528, w8529, w8530, w8531, w8532, w8533, w8534, w8535, w8536, w8537, w8538, w8539, w8540, w8541, w8542, w8543, w8544, w8545, w8546, w8547, w8548, w8549, w8550, w8551, w8552, w8553, w8554, w8555, w8556, w8557, w8558, w8559, w8560, w8561, w8562, w8563, w8564, w8565, w8566, w8567, w8568, w8569, w8570, w8571, w8572, w8573, w8574, w8575, w8576, w8577, w8578, w8579, w8580, w8581, w8582, w8583, w8584, w8585, w8586, w8587, w8588, w8589, w8590, w8591, w8592, w8593, w8594, w8595, w8596, w8597, w8598, w8599, w8600, w8601, w8602, w8603, w8604, w8605, w8606, w8607, w8608, w8609, w8610, w8611, w8612, w8613, w8614, w8615, w8616, w8617, w8618, w8619, w8620, w8621, w8622, w8623, w8624, w8625, w8626, w8627, w8628, w8629, w8630, w8631, w8632, w8633, w8634, w8635, w8636, w8637, w8638, w8639, w8640, w8641, w8642, w8643, w8644, w8645, w8646, w8647, w8648, w8649, w8650, w8651, w8652, w8653, w8654, w8655, w8656, w8657, w8658, w8659, w8660, w8661, w8662, w8663, w8664, w8665, w8666, w8667, w8668, w8669, w8670, w8671, w8672, w8673, w8674, w8675, w8676, w8677, w8678, w8679, w8680, w8681, w8682, w8683, w8684, w8685, w8686, w8687, w8688, w8689, w8690, w8691, w8692, w8693, w8694, w8695, w8696, w8697, w8698, w8699, w8700, w8701, w8702, w8703, w8704, w8705, w8706, w8707, w8708, w8709, w8710, w8711, w8712, w8713, w8714, w8715, w8716, w8717, w8718, w8719, w8720, w8721, w8722, w8723, w8724, w8725, w8726, w8727, w8728, w8729, w8730, w8731, w8732, w8733, w8734, w8735, w8736, w8737, w8738, w8739, w8740, w8741, w8742, w8743, w8744, w8745, w8746, w8747, w8748, w8749, w8750, w8751, w8752, w8753, w8754, w8755, w8756, w8757, w8758, w8759, w8760, w8761, w8762, w8763, w8764, w8765, w8766, w8767, w8768, w8769, w8770, w8771, w8772, w8773, w8774, w8775, w8776, w8777, w8778, w8779, w8780, w8781, w8782, w8783, w8784, w8785, w8786, w8787, w8788, w8789, w8790, w8791, w8792, w8793, w8794, w8795, w8796, w8797, w8798, w8799, w8800, w8801, w8802, w8803, w8804, w8805, w8806, w8807, w8808, w8809, w8810, w8811, w8812, w8813, w8814, w8815, w8816, w8817, w8818, w8819, w8820, w8821, w8822, w8823, w8824, w8825, w8826, w8827, w8828, w8829, w8830, w8831, w8832, w8833, w8834, w8835, w8836, w8837, w8838, w8839, w8840, w8841, w8842, w8843, w8844, w8845, w8846, w8847, w8848, w8849, w8850, w8851, w8852, w8853, w8854, w8855, w8856, w8857, w8858, w8859, w8860, w8861, w8862, w8863, w8864, w8865, w8866, w8867, w8868, w8869, w8870, w8871, w8872, w8873, w8874, w8875, w8876, w8877, w8878, w8879, w8880, w8881, w8882, w8883, w8884, w8885, w8886, w8887, w8888, w8889, w8890, w8891, w8892, w8893, w8894, w8895, w8896, w8897, w8898, w8899, w8900, w8901, w8902, w8903, w8904, w8905, w8906, w8907, w8908, w8909, w8910, w8911, w8912, w8913, w8914, w8915, w8916, w8917, w8918, w8919, w8920, w8921, w8922, w8923, w8924, w8925, w8926, w8927, w8928, w8929, w8930, w8931, w8932, w8933, w8934, w8935, w8936, w8937, w8938, w8939, w8940, w8941, w8942, w8943, w8944, w8945, w8946, w8947, w8948, w8949, w8950, w8951, w8952, w8953, w8954, w8955, w8956, w8957, w8958, w8959, w8960, w8961, w8962, w8963, w8964, w8965, w8966, w8967, w8968, w8969, w8970, w8971, w8972, w8973, w8974, w8975, w8976, w8977, w8978, w8979, w8980, w8981, w8982, w8983, w8984, w8985, w8986, w8987, w8988, w8989, w8990, w8991, w8992, w8993, w8994, w8995, w8996, w8997, w8998, w8999, w9000, w9001, w9002, w9003, w9004, w9005, w9006, w9007, w9008, w9009, w9010, w9011, w9012, w9013, w9014, w9015, w9016, w9017, w9018, w9019, w9020, w9021, w9022, w9023, w9024, w9025, w9026, w9027, w9028, w9029, w9030, w9031, w9032, w9033, w9034, w9035, w9036, w9037, w9038, w9039, w9040, w9041, w9042, w9043, w9044, w9045, w9046, w9047, w9048, w9049, w9050, w9051, w9052, w9053, w9054, w9055, w9056, w9057, w9058, w9059, w9060, w9061, w9062, w9063, w9064, w9065, w9066, w9067, w9068, w9069, w9070, w9071, w9072, w9073, w9074, w9075, w9076, w9077, w9078, w9079, w9080, w9081, w9082, w9083, w9084, w9085, w9086, w9087, w9088, w9089, w9090, w9091, w9092, w9093, w9094, w9095, w9096, w9097, w9098, w9099, w9100, w9101, w9102, w9103, w9104, w9105, w9106, w9107, w9108, w9109, w9110, w9111, w9112, w9113, w9114, w9115, w9116, w9117, w9118, w9119, w9120, w9121, w9122, w9123, w9124, w9125, w9126, w9127, w9128, w9129, w9130, w9131, w9132, w9133, w9134, w9135, w9136, w9137, w9138, w9139, w9140, w9141, w9142, w9143, w9144, w9145, w9146, w9147, w9148, w9149, w9150, w9151, w9152, w9153, w9154, w9155, w9156, w9157, w9158, w9159, w9160, w9161, w9162, w9163, w9164, w9165, w9166, w9167, w9168, w9169, w9170, w9171, w9172, w9173, w9174, w9175, w9176, w9177, w9178, w9179, w9180, w9181, w9182, w9183, w9184, w9185, w9186, w9187, w9188, w9189, w9190, w9191, w9192, w9193, w9194, w9195, w9196, w9197, w9198, w9199, w9200, w9201, w9202, w9203, w9204, w9205, w9206, w9207, w9208, w9209, w9210, w9211, w9212, w9213, w9214, w9215, w9216, w9217, w9218, w9219, w9220, w9221, w9222, w9223, w9224, w9225, w9226, w9227, w9228, w9229, w9230, w9231, w9232, w9233, w9234, w9235, w9236, w9237, w9238, w9239, w9240, w9241, w9242, w9243, w9244, w9245, w9246, w9247, w9248, w9249, w9250, w9251, w9252, w9253, w9254, w9255, w9256, w9257, w9258, w9259, w9260, w9261, w9262, w9263, w9264, w9265, w9266, w9267, w9268, w9269, w9270, w9271, w9272, w9273, w9274, w9275, w9276, w9277, w9278, w9279, w9280, w9281, w9282, w9283, w9284, w9285, w9286, w9287, w9288, w9289, w9290, w9291, w9292, w9293, w9294, w9295, w9296, w9297, w9298, w9299, w9300, w9301, w9302, w9303, w9304, w9305, w9306, w9307, w9308, w9309, w9310, w9311, w9312, w9313, w9314, w9315, w9316, w9317, w9318, w9319, w9320, w9321, w9322, w9323, w9324, w9325, w9326, w9327, w9328, w9329, w9330, w9331, w9332, w9333, w9334, w9335, w9336, w9337, w9338, w9339, w9340, w9341, w9342, w9343, w9344, w9345, w9346, w9347, w9348, w9349, w9350, w9351, w9352, w9353, w9354, w9355, w9356, w9357, w9358, w9359, w9360, w9361, w9362, w9363, w9364, w9365, w9366, w9367, w9368, w9369, w9370, w9371, w9372, w9373, w9374, w9375, w9376, w9377, w9378, w9379, w9380, w9381, w9382, w9383, w9384, w9385, w9386, w9387, w9388, w9389, w9390, w9391, w9392, w9393, w9394, w9395, w9396, w9397, w9398, w9399, w9400, w9401, w9402, w9403, w9404, w9405, w9406, w9407, w9408, w9409, w9410, w9411, w9412, w9413, w9414, w9415, w9416, w9417, w9418, w9419, w9420, w9421, w9422, w9423, w9424, w9425, w9426, w9427, w9428, w9429, w9430, w9431, w9432, w9433, w9434, w9435, w9436, w9437, w9438, w9439, w9440, w9441, w9442, w9443, w9444, w9445, w9446, w9447, w9448, w9449, w9450, w9451, w9452, w9453, w9454, w9455, w9456, w9457, w9458, w9459, w9460, w9461, w9462, w9463, w9464, w9465, w9466, w9467, w9468, w9469, w9470, w9471, w9472, w9473, w9474, w9475, w9476, w9477, w9478, w9479, w9480, w9481, w9482, w9483, w9484, w9485, w9486, w9487, w9488, w9489, w9490, w9491, w9492, w9493, w9494, w9495, w9496, w9497, w9498, w9499, w9500, w9501, w9502, w9503, w9504, w9505, w9506, w9507, w9508, w9509, w9510, w9511, w9512, w9513, w9514, w9515, w9516, w9517, w9518, w9519, w9520, w9521, w9522, w9523, w9524, w9525, w9526, w9527, w9528, w9529, w9530, w9531, w9532, w9533, w9534, w9535, w9536, w9537, w9538, w9539, w9540, w9541, w9542, w9543, w9544, w9545, w9546, w9547, w9548, w9549, w9550, w9551, w9552, w9553, w9554, w9555, w9556, w9557, w9558, w9559, w9560, w9561, w9562, w9563, w9564, w9565, w9566, w9567, w9568, w9569, w9570, w9571, w9572, w9573, w9574, w9575, w9576, w9577, w9578, w9579, w9580, w9581, w9582, w9583, w9584, w9585, w9586, w9587, w9588, w9589, w9590, w9591, w9592, w9593, w9594, w9595, w9596, w9597, w9598, w9599, w9600, w9601, w9602, w9603, w9604, w9605, w9606, w9607, w9608, w9609, w9610, w9611, w9612, w9613, w9614, w9615, w9616, w9617, w9618, w9619, w9620, w9621, w9622, w9623, w9624, w9625, w9626, w9627, w9628, w9629, w9630, w9631, w9632, w9633, w9634, w9635, w9636, w9637, w9638, w9639, w9640, w9641, w9642, w9643, w9644, w9645, w9646, w9647, w9648, w9649, w9650, w9651, w9652, w9653, w9654, w9655, w9656, w9657, w9658, w9659, w9660, w9661, w9662, w9663, w9664, w9665, w9666, w9667, w9668, w9669, w9670, w9671, w9672, w9673, w9674, w9675, w9676, w9677, w9678, w9679, w9680, w9681, w9682, w9683, w9684, w9685, w9686, w9687, w9688, w9689, w9690, w9691, w9692, w9693, w9694, w9695, w9696, w9697, w9698, w9699, w9700, w9701, w9702, w9703, w9704, w9705, w9706, w9707, w9708, w9709, w9710, w9711, w9712, w9713, w9714, w9715, w9716, w9717, w9718, w9719, w9720, w9721, w9722, w9723, w9724, w9725, w9726, w9727, w9728, w9729, w9730, w9731, w9732, w9733, w9734, w9735, w9736, w9737, w9738, w9739, w9740, w9741, w9742, w9743, w9744, w9745, w9746, w9747, w9748, w9749, w9750, w9751, w9752, w9753, w9754, w9755, w9756, w9757, w9758, w9759, w9760, w9761, w9762, w9763, w9764, w9765, w9766, w9767, w9768, w9769, w9770, w9771, w9772, w9773, w9774, w9775, w9776, w9777, w9778, w9779, w9780, w9781, w9782, w9783, w9784, w9785, w9786, w9787, w9788, w9789, w9790, w9791, w9792, w9793, w9794, w9795, w9796, w9797, w9798, w9799, w9800, w9801, w9802, w9803, w9804, w9805, w9806, w9807, w9808, w9809, w9810, w9811, w9812, w9813, w9814, w9815, w9816, w9817, w9818, w9819, w9820, w9821, w9822, w9823, w9824, w9825, w9826, w9827, w9828, w9829, w9830, w9831, w9832, w9833, w9834, w9835, w9836, w9837, w9838, w9839, w9840, w9841, w9842, w9843, w9844, w9845, w9846, w9847, w9848, w9849, w9850, w9851, w9852, w9853, w9854, w9855, w9856, w9857, w9858, w9859, w9860, w9861, w9862, w9863, w9864, w9865, w9866, w9867, w9868, w9869, w9870, w9871, w9872, w9873, w9874, w9875, w9876, w9877, w9878, w9879, w9880, w9881, w9882, w9883, w9884, w9885, w9886, w9887, w9888, w9889, w9890, w9891, w9892, w9893, w9894, w9895, w9896, w9897, w9898, w9899, w9900, w9901, w9902, w9903, w9904, w9905, w9906, w9907, w9908, w9909, w9910, w9911, w9912, w9913, w9914, w9915, w9916, w9917, w9918, w9919, w9920, w9921, w9922, w9923, w9924, w9925, w9926, w9927, w9928, w9929, w9930, w9931, w9932, w9933, w9934, w9935, w9936, w9937, w9938, w9939, w9940, w9941, w9942, w9943, w9944, w9945, w9946, w9947, w9948, w9949, w9950, w9951, w9952, w9953, w9954, w9955, w9956, w9957, w9958, w9959, w9960, w9961, w9962, w9963, w9964, w9965, w9966, w9967, w9968, w9969, w9970, w9971, w9972, w9973, w9974, w9975, w9976, w9977, w9978, w9979, w9980, w9981, w9982, w9983, w9984, w9985, w9986, w9987, w9988, w9989, w9990, w9991, w9992, w9993, w9994, w9995, w9996, w9997, w9998, w9999, w10000, w10001, w10002, w10003, w10004, w10005, w10006, w10007, w10008, w10009, w10010, w10011, w10012, w10013, w10014, w10015, w10016, w10017, w10018, w10019, w10020, w10021, w10022, w10023, w10024, w10025, w10026, w10027, w10028, w10029, w10030, w10031, w10032, w10033, w10034, w10035, w10036, w10037, w10038, w10039, w10040, w10041, w10042, w10043, w10044, w10045, w10046, w10047, w10048, w10049, w10050, w10051, w10052, w10053, w10054, w10055, w10056, w10057, w10058, w10059, w10060, w10061, w10062, w10063, w10064, w10065, w10066, w10067, w10068, w10069, w10070, w10071, w10072, w10073, w10074, w10075, w10076, w10077, w10078, w10079, w10080, w10081, w10082, w10083, w10084, w10085, w10086, w10087, w10088, w10089, w10090, w10091, w10092, w10093, w10094, w10095, w10096, w10097, w10098, w10099, w10100, w10101, w10102, w10103, w10104, w10105, w10106, w10107, w10108, w10109, w10110, w10111, w10112, w10113, w10114, w10115, w10116, w10117, w10118, w10119, w10120, w10121, w10122, w10123, w10124, w10125, w10126, w10127, w10128, w10129, w10130, w10131, w10132, w10133, w10134, w10135, w10136, w10137, w10138, w10139, w10140, w10141, w10142, w10143, w10144, w10145, w10146, w10147, w10148, w10149, w10150, w10151, w10152, w10153, w10154, w10155, w10156, w10157, w10158, w10159, w10160, w10161, w10162, w10163, w10164, w10165, w10166, w10167, w10168, w10169, w10170, w10171, w10172, w10173, w10174, w10175, w10176, w10177, w10178, w10179, w10180, w10181, w10182, w10183, w10184, w10185, w10186, w10187, w10188, w10189, w10190, w10191, w10192, w10193, w10194, w10195, w10196, w10197, w10198, w10199, w10200, w10201, w10202, w10203, w10204, w10205, w10206, w10207, w10208, w10209, w10210, w10211, w10212, w10213, w10214, w10215, w10216, w10217, w10218, w10219, w10220, w10221, w10222, w10223, w10224, w10225, w10226, w10227, w10228, w10229, w10230, w10231, w10232, w10233, w10234, w10235, w10236, w10237, w10238, w10239, w10240, w10241, w10242, w10243, w10244, w10245, w10246, w10247, w10248, w10249, w10250, w10251, w10252, w10253, w10254, w10255, w10256, w10257, w10258, w10259, w10260, w10261, w10262, w10263, w10264, w10265, w10266, w10267, w10268, w10269, w10270, w10271, w10272, w10273, w10274, w10275, w10276, w10277, w10278, w10279, w10280, w10281, w10282, w10283, w10284, w10285, w10286, w10287, w10288, w10289, w10290, w10291, w10292, w10293, w10294, w10295, w10296, w10297, w10298, w10299, w10300, w10301, w10302, w10303, w10304, w10305, w10306, w10307, w10308, w10309, w10310, w10311, w10312, w10313, w10314, w10315, w10316, w10317, w10318, w10319, w10320, w10321, w10322, w10323, w10324, w10325, w10326, w10327, w10328, w10329, w10330, w10331, w10332, w10333, w10334, w10335, w10336, w10337, w10338, w10339, w10340, w10341, w10342, w10343, w10344, w10345, w10346, w10347, w10348, w10349, w10350, w10351, w10352, w10353, w10354, w10355, w10356, w10357, w10358, w10359, w10360, w10361, w10362, w10363, w10364, w10365, w10366, w10367, w10368, w10369, w10370, w10371, w10372, w10373, w10374, w10375, w10376, w10377, w10378, w10379, w10380, w10381, w10382, w10383, w10384, w10385, w10386, w10387, w10388, w10389, w10390, w10391, w10392, w10393, w10394, w10395, w10396, w10397, w10398, w10399, w10400, w10401, w10402, w10403, w10404, w10405, w10406, w10407, w10408, w10409, w10410, w10411, w10412, w10413, w10414, w10415, w10416, w10417, w10418, w10419, w10420, w10421, w10422, w10423, w10424, w10425, w10426, w10427, w10428, w10429, w10430, w10431, w10432, w10433, w10434, w10435, w10436, w10437, w10438, w10439, w10440, w10441, w10442, w10443, w10444, w10445, w10446, w10447, w10448, w10449, w10450, w10451, w10452, w10453, w10454, w10455, w10456, w10457, w10458, w10459, w10460, w10461, w10462, w10463, w10464, w10465, w10466, w10467, w10468, w10469, w10470, w10471, w10472, w10473, w10474, w10475, w10476, w10477, w10478, w10479, w10480, w10481, w10482, w10483, w10484, w10485, w10486, w10487, w10488, w10489, w10490, w10491, w10492, w10493, w10494, w10495, w10496, w10497, w10498, w10499, w10500, w10501, w10502, w10503, w10504, w10505, w10506, w10507, w10508, w10509, w10510, w10511, w10512, w10513, w10514, w10515, w10516, w10517, w10518, w10519, w10520, w10521, w10522, w10523, w10524, w10525, w10526, w10527, w10528, w10529, w10530, w10531, w10532, w10533, w10534, w10535, w10536, w10537, w10538, w10539, w10540, w10541, w10542, w10543, w10544, w10545, w10546, w10547, w10548, w10549, w10550, w10551, w10552, w10553, w10554, w10555, w10556, w10557, w10558, w10559, w10560, w10561, w10562, w10563, w10564, w10565, w10566, w10567, w10568, w10569, w10570, w10571, w10572, w10573, w10574, w10575, w10576, w10577, w10578, w10579, w10580, w10581, w10582, w10583, w10584, w10585, w10586, w10587, w10588, w10589, w10590, w10591, w10592, w10593, w10594, w10595, w10596, w10597, w10598, w10599, w10600, w10601, w10602, w10603, w10604, w10605, w10606, w10607, w10608, w10609, w10610, w10611, w10612, w10613, w10614, w10615, w10616, w10617, w10618, w10619, w10620, w10621, w10622, w10623, w10624, w10625, w10626, w10627, w10628, w10629, w10630, w10631, w10632, w10633, w10634, w10635, w10636, w10637, w10638, w10639, w10640, w10641, w10642, w10643, w10644, w10645, w10646, w10647, w10648, w10649, w10650, w10651, w10652, w10653, w10654, w10655, w10656, w10657, w10658, w10659, w10660, w10661, w10662, w10663, w10664, w10665, w10666, w10667, w10668, w10669, w10670, w10671, w10672, w10673, w10674, w10675, w10676, w10677, w10678, w10679, w10680, w10681, w10682, w10683, w10684, w10685, w10686, w10687, w10688, w10689, w10690, w10691, w10692, w10693, w10694, w10695, w10696, w10697, w10698, w10699, w10700, w10701, w10702, w10703, w10704, w10705, w10706, w10707, w10708, w10709, w10710, w10711, w10712, w10713, w10714, w10715, w10716, w10717, w10718, w10719, w10720, w10721, w10722, w10723, w10724, w10725, w10726, w10727, w10728, w10729, w10730, w10731, w10732, w10733, w10734, w10735, w10736, w10737, w10738, w10739, w10740, w10741, w10742, w10743, w10744, w10745, w10746, w10747, w10748, w10749, w10750, w10751, w10752, w10753, w10754, w10755, w10756, w10757, w10758, w10759, w10760, w10761, w10762, w10763, w10764, w10765, w10766, w10767, w10768, w10769, w10770, w10771, w10772, w10773, w10774, w10775, w10776, w10777, w10778, w10779, w10780, w10781, w10782, w10783, w10784, w10785, w10786, w10787, w10788, w10789, w10790, w10791, w10792, w10793, w10794, w10795, w10796, w10797, w10798, w10799, w10800, w10801, w10802, w10803, w10804, w10805, w10806, w10807, w10808, w10809, w10810, w10811, w10812, w10813, w10814, w10815, w10816, w10817, w10818, w10819, w10820, w10821, w10822, w10823, w10824, w10825, w10826, w10827, w10828, w10829, w10830, w10831, w10832, w10833, w10834, w10835, w10836, w10837, w10838, w10839, w10840, w10841, w10842, w10843, w10844, w10845, w10846, w10847, w10848, w10849, w10850, w10851, w10852, w10853, w10854, w10855, w10856, w10857, w10858, w10859, w10860, w10861, w10862, w10863, w10864, w10865, w10866, w10867, w10868, w10869, w10870, w10871, w10872, w10873, w10874, w10875, w10876, w10877, w10878, w10879, w10880, w10881, w10882, w10883, w10884, w10885, w10886, w10887, w10888, w10889, w10890, w10891, w10892, w10893, w10894, w10895, w10896, w10897, w10898, w10899, w10900, w10901, w10902, w10903, w10904, w10905, w10906, w10907, w10908, w10909, w10910, w10911, w10912, w10913, w10914, w10915, w10916, w10917, w10918, w10919, w10920, w10921, w10922, w10923, w10924, w10925, w10926, w10927, w10928, w10929, w10930, w10931, w10932, w10933, w10934, w10935, w10936, w10937, w10938, w10939, w10940, w10941, w10942, w10943, w10944, w10945, w10946, w10947, w10948, w10949, w10950, w10951, w10952, w10953, w10954, w10955, w10956, w10957, w10958, w10959, w10960, w10961, w10962, w10963, w10964, w10965, w10966, w10967, w10968, w10969, w10970, w10971, w10972, w10973, w10974, w10975, w10976, w10977, w10978, w10979, w10980, w10981, w10982, w10983, w10984, w10985, w10986, w10987, w10988, w10989, w10990, w10991, w10992, w10993, w10994, w10995, w10996, w10997, w10998, w10999, w11000, w11001, w11002, w11003, w11004, w11005, w11006, w11007, w11008, w11009, w11010, w11011, w11012, w11013, w11014, w11015, w11016, w11017, w11018, w11019, w11020, w11021, w11022, w11023, w11024, w11025, w11026, w11027, w11028, w11029, w11030, w11031, w11032, w11033, w11034, w11035, w11036, w11037, w11038, w11039, w11040, w11041, w11042, w11043, w11044, w11045, w11046, w11047, w11048, w11049, w11050, w11051, w11052, w11053, w11054, w11055, w11056, w11057, w11058, w11059, w11060, w11061, w11062, w11063, w11064, w11065, w11066, w11067, w11068, w11069, w11070, w11071, w11072, w11073, w11074, w11075, w11076, w11077, w11078, w11079, w11080, w11081, w11082, w11083, w11084, w11085, w11086, w11087, w11088, w11089, w11090, w11091, w11092, w11093, w11094, w11095, w11096, w11097, w11098, w11099, w11100, w11101, w11102, w11103, w11104, w11105, w11106, w11107, w11108, w11109, w11110, w11111, w11112, w11113, w11114, w11115, w11116, w11117, w11118, w11119, w11120, w11121, w11122, w11123, w11124, w11125, w11126, w11127, w11128, w11129, w11130, w11131, w11132, w11133, w11134, w11135, w11136, w11137, w11138, w11139, w11140, w11141, w11142, w11143, w11144, w11145, w11146, w11147, w11148, w11149, w11150, w11151, w11152, w11153, w11154, w11155, w11156, w11157, w11158, w11159, w11160, w11161, w11162, w11163, w11164, w11165, w11166, w11167, w11168, w11169, w11170, w11171, w11172, w11173, w11174, w11175, w11176, w11177, w11178, w11179, w11180, w11181, w11182, w11183, w11184, w11185, w11186, w11187, w11188, w11189, w11190, w11191, w11192, w11193, w11194, w11195, w11196, w11197, w11198, w11199, w11200, w11201, w11202, w11203, w11204, w11205, w11206, w11207, w11208, w11209, w11210, w11211, w11212, w11213, w11214, w11215, w11216, w11217, w11218, w11219, w11220, w11221, w11222, w11223, w11224, w11225, w11226, w11227, w11228, w11229, w11230, w11231, w11232, w11233, w11234, w11235, w11236, w11237, w11238, w11239, w11240, w11241, w11242, w11243, w11244, w11245, w11246, w11247, w11248, w11249, w11250, w11251, w11252, w11253, w11254, w11255, w11256, w11257, w11258, w11259, w11260, w11261, w11262, w11263, w11264, w11265, w11266, w11267, w11268, w11269, w11270, w11271, w11272, w11273, w11274, w11275, w11276, w11277, w11278, w11279, w11280, w11281, w11282, w11283, w11284, w11285, w11286, w11287, w11288, w11289, w11290, w11291, w11292, w11293, w11294, w11295, w11296, w11297, w11298, w11299, w11300, w11301, w11302, w11303, w11304, w11305, w11306, w11307, w11308, w11309, w11310, w11311, w11312, w11313, w11314, w11315, w11316, w11317, w11318, w11319, w11320, w11321, w11322, w11323, w11324, w11325, w11326, w11327, w11328, w11329, w11330, w11331, w11332, w11333, w11334, w11335, w11336, w11337, w11338, w11339, w11340, w11341, w11342, w11343, w11344, w11345, w11346, w11347, w11348, w11349, w11350, w11351, w11352, w11353, w11354, w11355, w11356, w11357, w11358, w11359, w11360, w11361, w11362, w11363, w11364, w11365, w11366, w11367, w11368, w11369, w11370, w11371, w11372, w11373, w11374, w11375, w11376, w11377, w11378, w11379, w11380, w11381, w11382, w11383, w11384, w11385, w11386, w11387, w11388, w11389, w11390, w11391, w11392, w11393, w11394, w11395, w11396, w11397, w11398, w11399, w11400, w11401, w11402, w11403, w11404, w11405, w11406, w11407, w11408, w11409, w11410, w11411, w11412, w11413, w11414, w11415, w11416, w11417, w11418, w11419, w11420, w11421, w11422, w11423, w11424, w11425, w11426, w11427, w11428, w11429, w11430, w11431, w11432, w11433, w11434, w11435, w11436, w11437, w11438, w11439, w11440, w11441, w11442, w11443, w11444, w11445, w11446, w11447, w11448, w11449, w11450, w11451, w11452, w11453, w11454, w11455, w11456, w11457, w11458, w11459, w11460, w11461, w11462, w11463, w11464, w11465, w11466, w11467, w11468, w11469, w11470, w11471, w11472, w11473, w11474, w11475, w11476, w11477, w11478, w11479, w11480, w11481, w11482, w11483, w11484, w11485, w11486, w11487, w11488, w11489, w11490, w11491, w11492, w11493, w11494, w11495, w11496, w11497, w11498, w11499, w11500, w11501, w11502, w11503, w11504, w11505, w11506, w11507, w11508, w11509, w11510, w11511, w11512, w11513, w11514, w11515, w11516, w11517, w11518, w11519, w11520, w11521, w11522, w11523, w11524, w11525, w11526, w11527, w11528, w11529, w11530, w11531, w11532, w11533, w11534, w11535, w11536, w11537, w11538, w11539, w11540, w11541, w11542, w11543, w11544, w11545, w11546, w11547, w11548, w11549, w11550, w11551, w11552, w11553, w11554, w11555, w11556, w11557, w11558, w11559, w11560, w11561, w11562, w11563, w11564, w11565, w11566, w11567, w11568, w11569, w11570, w11571, w11572, w11573, w11574, w11575, w11576, w11577, w11578, w11579, w11580, w11581, w11582, w11583, w11584, w11585, w11586, w11587, w11588, w11589, w11590, w11591, w11592, w11593, w11594, w11595, w11596, w11597, w11598, w11599, w11600, w11601, w11602, w11603, w11604, w11605, w11606, w11607, w11608, w11609, w11610, w11611, w11612, w11613, w11614, w11615, w11616, w11617, w11618, w11619, w11620, w11621, w11622, w11623, w11624, w11625, w11626, w11627, w11628, w11629, w11630, w11631, w11632, w11633, w11634, w11635, w11636, w11637, w11638, w11639, w11640, w11641, w11642, w11643, w11644, w11645, w11646, w11647, w11648, w11649, w11650, w11651, w11652, w11653, w11654, w11655, w11656, w11657, w11658, w11659, w11660, w11661, w11662, w11663, w11664, w11665, w11666, w11667, w11668, w11669, w11670, w11671, w11672, w11673, w11674, w11675, w11676, w11677, w11678, w11679, w11680, w11681, w11682, w11683, w11684, w11685, w11686, w11687, w11688, w11689, w11690, w11691, w11692, w11693, w11694, w11695, w11696, w11697, w11698, w11699, w11700, w11701, w11702, w11703, w11704, w11705, w11706, w11707, w11708, w11709, w11710, w11711, w11712, w11713, w11714, w11715, w11716, w11717, w11718, w11719, w11720, w11721, w11722, w11723, w11724, w11725, w11726, w11727, w11728, w11729, w11730, w11731, w11732, w11733, w11734, w11735, w11736, w11737, w11738, w11739, w11740, w11741, w11742, w11743, w11744, w11745, w11746, w11747, w11748, w11749, w11750, w11751, w11752, w11753, w11754, w11755, w11756, w11757, w11758, w11759, w11760, w11761, w11762, w11763, w11764, w11765, w11766, w11767, w11768, w11769, w11770, w11771, w11772, w11773, w11774, w11775, w11776, w11777, w11778, w11779, w11780, w11781, w11782, w11783, w11784, w11785, w11786, w11787, w11788, w11789, w11790, w11791, w11792, w11793, w11794, w11795, w11796, w11797, w11798, w11799, w11800, w11801, w11802, w11803, w11804, w11805, w11806, w11807, w11808, w11809, w11810, w11811, w11812, w11813, w11814, w11815, w11816, w11817, w11818, w11819, w11820, w11821, w11822, w11823, w11824, w11825, w11826, w11827, w11828, w11829, w11830, w11831, w11832, w11833, w11834, w11835, w11836, w11837, w11838, w11839, w11840, w11841, w11842, w11843, w11844, w11845, w11846, w11847, w11848, w11849, w11850, w11851, w11852, w11853, w11854, w11855, w11856, w11857, w11858, w11859, w11860, w11861, w11862, w11863, w11864, w11865, w11866, w11867, w11868, w11869, w11870, w11871, w11872, w11873, w11874, w11875, w11876, w11877, w11878, w11879, w11880, w11881, w11882, w11883, w11884, w11885, w11886, w11887, w11888, w11889, w11890, w11891, w11892, w11893, w11894, w11895, w11896, w11897, w11898, w11899, w11900, w11901, w11902, w11903, w11904, w11905, w11906, w11907, w11908, w11909, w11910, w11911, w11912, w11913, w11914, w11915, w11916, w11917, w11918, w11919, w11920, w11921, w11922, w11923, w11924, w11925, w11926, w11927, w11928, w11929, w11930, w11931, w11932, w11933, w11934, w11935, w11936, w11937, w11938, w11939, w11940, w11941, w11942, w11943, w11944, w11945, w11946, w11947, w11948, w11949, w11950, w11951, w11952, w11953, w11954, w11955, w11956, w11957, w11958, w11959, w11960, w11961, w11962, w11963, w11964, w11965, w11966, w11967, w11968, w11969, w11970, w11971, w11972, w11973, w11974, w11975, w11976, w11977, w11978, w11979, w11980, w11981, w11982, w11983, w11984, w11985, w11986, w11987, w11988, w11989, w11990, w11991, w11992, w11993, w11994, w11995, w11996, w11997, w11998, w11999, w12000, w12001, w12002, w12003, w12004, w12005, w12006, w12007, w12008, w12009, w12010, w12011, w12012, w12013, w12014, w12015, w12016, w12017, w12018, w12019, w12020, w12021, w12022, w12023, w12024, w12025, w12026, w12027, w12028, w12029, w12030, w12031, w12032, w12033, w12034, w12035, w12036, w12037, w12038, w12039, w12040, w12041, w12042, w12043, w12044, w12045, w12046, w12047, w12048, w12049, w12050, w12051, w12052, w12053, w12054, w12055, w12056, w12057, w12058, w12059, w12060, w12061, w12062, w12063, w12064, w12065, w12066, w12067, w12068, w12069, w12070, w12071, w12072, w12073, w12074, w12075, w12076, w12077, w12078, w12079, w12080, w12081, w12082, w12083, w12084, w12085, w12086, w12087, w12088, w12089, w12090, w12091, w12092, w12093, w12094, w12095, w12096, w12097, w12098, w12099, w12100, w12101, w12102, w12103, w12104, w12105, w12106, w12107, w12108, w12109, w12110, w12111, w12112, w12113, w12114, w12115, w12116, w12117, w12118, w12119, w12120, w12121, w12122, w12123, w12124, w12125, w12126, w12127, w12128, w12129, w12130, w12131, w12132, w12133, w12134, w12135, w12136, w12137, w12138, w12139, w12140, w12141, w12142, w12143, w12144, w12145, w12146, w12147, w12148, w12149, w12150, w12151, w12152, w12153, w12154, w12155, w12156, w12157, w12158, w12159, w12160, w12161, w12162, w12163, w12164, w12165, w12166, w12167, w12168, w12169, w12170, w12171, w12172, w12173, w12174, w12175, w12176, w12177, w12178, w12179, w12180, w12181, w12182, w12183, w12184, w12185, w12186, w12187, w12188, w12189, w12190, w12191, w12192, w12193, w12194, w12195, w12196, w12197, w12198, w12199, w12200, w12201, w12202, w12203, w12204, w12205, w12206, w12207, w12208, w12209, w12210, w12211, w12212, w12213, w12214, w12215, w12216, w12217, w12218, w12219, w12220, w12221, w12222, w12223, w12224, w12225, w12226, w12227, w12228, w12229, w12230, w12231, w12232, w12233, w12234, w12235, w12236, w12237, w12238, w12239, w12240, w12241, w12242, w12243, w12244, w12245, w12246, w12247, w12248, w12249, w12250, w12251, w12252, w12253, w12254, w12255, w12256, w12257, w12258, w12259, w12260, w12261, w12262, w12263, w12264, w12265, w12266, w12267, w12268, w12269, w12270, w12271, w12272, w12273, w12274, w12275, w12276, w12277, w12278, w12279, w12280, w12281, w12282, w12283, w12284, w12285, w12286, w12287, w12288, w12289, w12290, w12291, w12292, w12293, w12294, w12295, w12296, w12297, w12298, w12299, w12300, w12301, w12302, w12303, w12304, w12305, w12306, w12307, w12308, w12309, w12310, w12311, w12312, w12313, w12314, w12315, w12316, w12317, w12318, w12319, w12320, w12321, w12322, w12323, w12324, w12325, w12326, w12327, w12328, w12329, w12330, w12331, w12332, w12333, w12334, w12335, w12336, w12337, w12338, w12339, w12340, w12341, w12342, w12343, w12344, w12345, w12346, w12347, w12348, w12349, w12350, w12351, w12352, w12353, w12354, w12355, w12356, w12357, w12358, w12359, w12360, w12361, w12362, w12363, w12364, w12365, w12366, w12367, w12368, w12369, w12370, w12371, w12372, w12373, w12374, w12375, w12376, w12377, w12378, w12379, w12380, w12381, w12382, w12383, w12384, w12385, w12386, w12387, w12388, w12389, w12390, w12391, w12392, w12393, w12394, w12395, w12396, w12397, w12398, w12399, w12400, w12401, w12402, w12403, w12404, w12405, w12406, w12407, w12408, w12409, w12410, w12411, w12412, w12413, w12414, w12415, w12416, w12417, w12418, w12419, w12420, w12421, w12422, w12423, w12424, w12425, w12426, w12427, w12428, w12429, w12430, w12431, w12432, w12433, w12434, w12435, w12436, w12437, w12438, w12439, w12440, w12441, w12442, w12443, w12444, w12445, w12446, w12447, w12448, w12449, w12450, w12451, w12452, w12453, w12454, w12455, w12456, w12457, w12458, w12459, w12460, w12461, w12462, w12463, w12464, w12465, w12466, w12467, w12468, w12469, w12470, w12471, w12472, w12473, w12474, w12475, w12476, w12477, w12478, w12479, w12480, w12481, w12482, w12483, w12484, w12485, w12486, w12487, w12488, w12489, w12490, w12491, w12492, w12493, w12494, w12495, w12496, w12497, w12498, w12499, w12500, w12501, w12502, w12503, w12504, w12505, w12506, w12507, w12508, w12509, w12510, w12511, w12512, w12513, w12514, w12515, w12516, w12517, w12518, w12519, w12520, w12521, w12522, w12523, w12524, w12525, w12526, w12527, w12528, w12529, w12530, w12531, w12532, w12533, w12534, w12535, w12536, w12537, w12538, w12539, w12540, w12541, w12542, w12543, w12544, w12545, w12546, w12547, w12548, w12549, w12550, w12551, w12552, w12553, w12554, w12555, w12556, w12557, w12558, w12559, w12560, w12561, w12562, w12563, w12564, w12565, w12566, w12567, w12568, w12569, w12570, w12571, w12572, w12573, w12574, w12575, w12576, w12577, w12578, w12579, w12580, w12581, w12582, w12583, w12584, w12585, w12586, w12587, w12588, w12589, w12590, w12591, w12592, w12593, w12594, w12595, w12596, w12597, w12598, w12599, w12600, w12601, w12602, w12603, w12604, w12605, w12606, w12607, w12608, w12609, w12610, w12611, w12612, w12613, w12614, w12615, w12616, w12617, w12618, w12619, w12620, w12621, w12622, w12623, w12624, w12625, w12626, w12627, w12628, w12629, w12630, w12631, w12632, w12633, w12634, w12635, w12636, w12637, w12638, w12639, w12640, w12641, w12642, w12643, w12644, w12645, w12646, w12647, w12648, w12649, w12650, w12651, w12652, w12653, w12654, w12655, w12656, w12657, w12658, w12659, w12660, w12661, w12662, w12663, w12664, w12665, w12666, w12667, w12668, w12669, w12670, w12671, w12672, w12673, w12674, w12675, w12676, w12677, w12678, w12679, w12680, w12681, w12682, w12683, w12684, w12685, w12686, w12687, w12688, w12689, w12690, w12691, w12692, w12693, w12694, w12695, w12696, w12697, w12698, w12699, w12700, w12701, w12702, w12703, w12704, w12705, w12706, w12707, w12708, w12709, w12710, w12711, w12712, w12713, w12714, w12715, w12716, w12717, w12718, w12719, w12720, w12721, w12722, w12723, w12724, w12725, w12726, w12727, w12728, w12729, w12730, w12731, w12732, w12733, w12734, w12735, w12736, w12737, w12738, w12739, w12740, w12741, w12742, w12743, w12744, w12745, w12746, w12747, w12748, w12749, w12750, w12751, w12752, w12753, w12754, w12755, w12756, w12757, w12758, w12759, w12760, w12761, w12762, w12763, w12764, w12765, w12766, w12767, w12768, w12769, w12770, w12771, w12772, w12773, w12774, w12775, w12776, w12777, w12778, w12779, w12780, w12781, w12782, w12783, w12784, w12785, w12786, w12787, w12788, w12789, w12790, w12791, w12792, w12793, w12794, w12795, w12796, w12797, w12798, w12799, w12800, w12801, w12802, w12803, w12804, w12805, w12806, w12807, w12808, w12809, w12810, w12811, w12812, w12813, w12814, w12815, w12816, w12817, w12818, w12819, w12820, w12821, w12822, w12823, w12824, w12825, w12826, w12827, w12828, w12829, w12830, w12831, w12832, w12833, w12834, w12835, w12836, w12837, w12838, w12839, w12840, w12841, w12842, w12843, w12844, w12845, w12846, w12847, w12848, w12849, w12850, w12851, w12852, w12853, w12854, w12855, w12856, w12857, w12858, w12859, w12860, w12861, w12862, w12863, w12864, w12865, w12866, w12867, w12868, w12869, w12870, w12871, w12872, w12873, w12874, w12875, w12876, w12877, w12878, w12879, w12880, w12881, w12882, w12883, w12884, w12885, w12886, w12887, w12888, w12889, w12890, w12891, w12892, w12893, w12894, w12895, w12896, w12897, w12898, w12899, w12900, w12901, w12902, w12903, w12904, w12905, w12906, w12907, w12908, w12909, w12910, w12911, w12912, w12913, w12914, w12915, w12916, w12917, w12918, w12919, w12920, w12921, w12922, w12923, w12924, w12925, w12926, w12927, w12928, w12929, w12930, w12931, w12932, w12933, w12934, w12935, w12936, w12937, w12938, w12939, w12940, w12941, w12942, w12943, w12944, w12945, w12946, w12947, w12948, w12949, w12950, w12951, w12952, w12953, w12954, w12955, w12956, w12957, w12958, w12959, w12960, w12961, w12962, w12963, w12964, w12965, w12966, w12967, w12968, w12969, w12970, w12971, w12972, w12973, w12974, w12975, w12976, w12977, w12978, w12979, w12980, w12981, w12982, w12983, w12984, w12985, w12986, w12987, w12988, w12989, w12990, w12991, w12992, w12993, w12994, w12995, w12996, w12997, w12998, w12999, w13000, w13001, w13002, w13003, w13004, w13005, w13006, w13007, w13008, w13009, w13010, w13011, w13012, w13013, w13014, w13015, w13016, w13017, w13018, w13019, w13020, w13021, w13022, w13023, w13024, w13025, w13026, w13027, w13028, w13029, w13030, w13031, w13032, w13033, w13034, w13035, w13036, w13037, w13038, w13039, w13040, w13041, w13042, w13043, w13044, w13045, w13046, w13047, w13048, w13049, w13050, w13051, w13052, w13053, w13054, w13055, w13056, w13057, w13058, w13059, w13060, w13061, w13062, w13063, w13064, w13065, w13066, w13067, w13068, w13069, w13070, w13071, w13072, w13073, w13074, w13075, w13076, w13077, w13078, w13079, w13080, w13081, w13082, w13083, w13084, w13085, w13086, w13087, w13088, w13089, w13090, w13091, w13092, w13093, w13094, w13095, w13096, w13097, w13098, w13099, w13100, w13101, w13102, w13103, w13104, w13105, w13106, w13107, w13108, w13109, w13110, w13111, w13112, w13113, w13114, w13115, w13116, w13117, w13118, w13119, w13120, w13121, w13122, w13123, w13124, w13125, w13126, w13127, w13128, w13129, w13130, w13131, w13132, w13133, w13134, w13135, w13136, w13137, w13138, w13139, w13140, w13141, w13142, w13143, w13144, w13145, w13146, w13147, w13148, w13149, w13150, w13151, w13152, w13153, w13154, w13155, w13156, w13157, w13158, w13159, w13160, w13161, w13162, w13163, w13164, w13165, w13166, w13167, w13168, w13169, w13170, w13171, w13172, w13173, w13174, w13175, w13176, w13177, w13178, w13179, w13180, w13181, w13182, w13183, w13184, w13185, w13186, w13187, w13188, w13189, w13190, w13191, w13192, w13193, w13194, w13195, w13196, w13197, w13198, w13199, w13200, w13201, w13202, w13203, w13204, w13205, w13206, w13207, w13208, w13209, w13210, w13211, w13212, w13213, w13214, w13215, w13216, w13217, w13218, w13219, w13220, w13221, w13222, w13223, w13224, w13225, w13226, w13227, w13228, w13229, w13230, w13231, w13232, w13233, w13234, w13235, w13236, w13237, w13238, w13239, w13240, w13241, w13242, w13243, w13244, w13245, w13246, w13247, w13248, w13249, w13250, w13251, w13252, w13253, w13254, w13255, w13256, w13257, w13258, w13259, w13260, w13261, w13262, w13263, w13264, w13265, w13266, w13267, w13268, w13269, w13270, w13271, w13272, w13273, w13274, w13275, w13276, w13277, w13278, w13279, w13280, w13281, w13282, w13283, w13284, w13285, w13286, w13287, w13288, w13289, w13290, w13291, w13292, w13293, w13294, w13295, w13296, w13297, w13298, w13299, w13300, w13301, w13302, w13303, w13304, w13305, w13306, w13307, w13308, w13309, w13310, w13311, w13312, w13313, w13314, w13315, w13316, w13317, w13318, w13319, w13320, w13321, w13322, w13323, w13324, w13325, w13326, w13327, w13328, w13329, w13330, w13331, w13332, w13333, w13334, w13335, w13336, w13337, w13338, w13339, w13340, w13341, w13342, w13343, w13344, w13345, w13346, w13347, w13348, w13349, w13350, w13351, w13352, w13353, w13354, w13355, w13356, w13357, w13358, w13359, w13360, w13361, w13362, w13363, w13364, w13365, w13366, w13367, w13368, w13369, w13370, w13371, w13372, w13373, w13374, w13375, w13376, w13377, w13378, w13379, w13380, w13381, w13382, w13383, w13384, w13385, w13386, w13387, w13388, w13389, w13390, w13391, w13392, w13393, w13394, w13395, w13396, w13397, w13398, w13399, w13400, w13401, w13402, w13403, w13404, w13405, w13406, w13407, w13408, w13409, w13410, w13411, w13412, w13413, w13414, w13415, w13416, w13417, w13418, w13419, w13420, w13421, w13422, w13423, w13424, w13425, w13426, w13427, w13428, w13429, w13430, w13431, w13432, w13433, w13434, w13435, w13436, w13437, w13438, w13439, w13440, w13441, w13442, w13443, w13444, w13445, w13446, w13447, w13448, w13449, w13450, w13451, w13452, w13453, w13454, w13455, w13456, w13457, w13458, w13459, w13460, w13461, w13462, w13463, w13464, w13465, w13466, w13467, w13468, w13469, w13470, w13471, w13472, w13473, w13474, w13475, w13476, w13477, w13478, w13479, w13480, w13481, w13482, w13483, w13484, w13485, w13486, w13487, w13488, w13489, w13490, w13491, w13492, w13493, w13494, w13495, w13496, w13497, w13498, w13499, w13500, w13501, w13502, w13503, w13504, w13505, w13506, w13507, w13508, w13509, w13510, w13511, w13512, w13513, w13514, w13515, w13516, w13517, w13518, w13519, w13520, w13521, w13522, w13523, w13524, w13525, w13526, w13527, w13528, w13529, w13530, w13531, w13532, w13533, w13534, w13535, w13536, w13537, w13538, w13539, w13540, w13541, w13542, w13543, w13544, w13545, w13546, w13547, w13548, w13549, w13550, w13551, w13552, w13553, w13554, w13555, w13556, w13557, w13558, w13559, w13560, w13561, w13562, w13563, w13564, w13565, w13566, w13567, w13568, w13569, w13570, w13571, w13572, w13573, w13574, w13575, w13576, w13577, w13578, w13579, w13580, w13581, w13582, w13583, w13584, w13585, w13586, w13587, w13588, w13589, w13590, w13591, w13592, w13593, w13594, w13595, w13596, w13597, w13598, w13599, w13600, w13601, w13602, w13603, w13604, w13605, w13606, w13607, w13608, w13609, w13610, w13611, w13612, w13613, w13614, w13615, w13616, w13617, w13618, w13619, w13620, w13621, w13622, w13623, w13624, w13625, w13626, w13627, w13628, w13629, w13630, w13631, w13632, w13633, w13634, w13635, w13636, w13637, w13638, w13639, w13640, w13641, w13642, w13643, w13644, w13645, w13646, w13647, w13648, w13649, w13650, w13651, w13652, w13653, w13654, w13655, w13656, w13657, w13658, w13659, w13660, w13661, w13662, w13663, w13664, w13665, w13666, w13667, w13668, w13669, w13670, w13671, w13672, w13673, w13674, w13675, w13676, w13677, w13678, w13679, w13680, w13681, w13682, w13683, w13684, w13685, w13686, w13687, w13688, w13689, w13690, w13691, w13692, w13693, w13694, w13695, w13696, w13697, w13698, w13699, w13700, w13701, w13702, w13703, w13704, w13705, w13706, w13707, w13708, w13709, w13710, w13711, w13712, w13713, w13714, w13715, w13716, w13717, w13718, w13719, w13720, w13721, w13722, w13723, w13724, w13725, w13726, w13727, w13728, w13729, w13730, w13731, w13732, w13733, w13734, w13735, w13736, w13737, w13738, w13739, w13740, w13741, w13742, w13743, w13744, w13745, w13746, w13747, w13748, w13749, w13750, w13751, w13752, w13753, w13754, w13755, w13756, w13757, w13758, w13759, w13760, w13761, w13762, w13763, w13764, w13765, w13766, w13767, w13768, w13769, w13770, w13771, w13772, w13773, w13774, w13775, w13776, w13777, w13778, w13779, w13780, w13781, w13782, w13783, w13784, w13785, w13786, w13787, w13788, w13789, w13790, w13791, w13792, w13793, w13794, w13795, w13796, w13797, w13798, w13799, w13800, w13801, w13802, w13803, w13804, w13805, w13806, w13807, w13808, w13809, w13810, w13811, w13812, w13813, w13814, w13815, w13816, w13817, w13818, w13819, w13820, w13821, w13822, w13823, w13824, w13825, w13826, w13827, w13828, w13829, w13830, w13831, w13832, w13833, w13834, w13835, w13836, w13837, w13838, w13839, w13840, w13841, w13842, w13843, w13844, w13845, w13846, w13847, w13848, w13849, w13850, w13851, w13852, w13853, w13854, w13855, w13856, w13857, w13858, w13859, w13860, w13861, w13862, w13863, w13864, w13865, w13866, w13867, w13868, w13869, w13870, w13871, w13872, w13873, w13874, w13875, w13876, w13877, w13878, w13879, w13880, w13881, w13882, w13883, w13884, w13885, w13886, w13887, w13888, w13889, w13890, w13891, w13892, w13893, w13894, w13895, w13896, w13897, w13898, w13899, w13900, w13901, w13902, w13903, w13904, w13905, w13906, w13907, w13908, w13909, w13910, w13911, w13912, w13913, w13914, w13915, w13916, w13917, w13918, w13919, w13920, w13921, w13922, w13923, w13924, w13925, w13926, w13927, w13928, w13929, w13930, w13931, w13932, w13933, w13934, w13935, w13936, w13937, w13938, w13939, w13940, w13941, w13942, w13943, w13944, w13945, w13946, w13947, w13948, w13949, w13950, w13951, w13952, w13953, w13954, w13955, w13956, w13957, w13958, w13959, w13960, w13961, w13962, w13963, w13964, w13965, w13966, w13967, w13968, w13969, w13970, w13971, w13972, w13973, w13974, w13975, w13976, w13977, w13978, w13979, w13980, w13981, w13982, w13983, w13984, w13985, w13986, w13987, w13988, w13989, w13990, w13991, w13992, w13993, w13994, w13995, w13996, w13997, w13998, w13999, w14000, w14001, w14002, w14003, w14004, w14005, w14006, w14007, w14008, w14009, w14010, w14011, w14012, w14013, w14014, w14015, w14016, w14017, w14018, w14019, w14020, w14021, w14022, w14023, w14024, w14025, w14026, w14027, w14028, w14029, w14030, w14031, w14032, w14033, w14034, w14035, w14036, w14037, w14038, w14039, w14040, w14041, w14042, w14043, w14044, w14045, w14046, w14047, w14048, w14049, w14050, w14051, w14052, w14053, w14054, w14055, w14056, w14057, w14058, w14059, w14060, w14061, w14062, w14063, w14064, w14065, w14066, w14067, w14068, w14069, w14070, w14071, w14072, w14073, w14074, w14075, w14076, w14077, w14078, w14079, w14080, w14081, w14082, w14083, w14084, w14085, w14086, w14087, w14088, w14089, w14090, w14091, w14092, w14093, w14094, w14095, w14096, w14097, w14098, w14099, w14100, w14101, w14102, w14103, w14104, w14105, w14106, w14107, w14108, w14109, w14110, w14111, w14112, w14113, w14114, w14115, w14116, w14117, w14118, w14119, w14120, w14121, w14122, w14123, w14124, w14125, w14126, w14127, w14128, w14129, w14130, w14131, w14132, w14133, w14134, w14135, w14136, w14137, w14138, w14139, w14140, w14141, w14142, w14143, w14144, w14145, w14146, w14147, w14148, w14149, w14150, w14151, w14152, w14153, w14154, w14155, w14156, w14157, w14158, w14159, w14160, w14161, w14162, w14163, w14164, w14165, w14166, w14167, w14168, w14169, w14170, w14171, w14172, w14173, w14174, w14175, w14176, w14177, w14178, w14179, w14180, w14181, w14182, w14183, w14184, w14185, w14186, w14187, w14188, w14189, w14190, w14191, w14192, w14193, w14194, w14195, w14196, w14197, w14198, w14199, w14200, w14201, w14202, w14203, w14204, w14205, w14206, w14207, w14208, w14209, w14210, w14211, w14212, w14213, w14214, w14215, w14216, w14217, w14218, w14219, w14220, w14221, w14222, w14223, w14224, w14225, w14226, w14227, w14228, w14229, w14230, w14231, w14232, w14233, w14234, w14235, w14236, w14237, w14238, w14239, w14240, w14241, w14242, w14243, w14244, w14245, w14246, w14247, w14248, w14249, w14250, w14251, w14252, w14253, w14254, w14255, w14256, w14257, w14258, w14259, w14260, w14261, w14262, w14263, w14264, w14265, w14266, w14267, w14268, w14269, w14270, w14271, w14272, w14273, w14274, w14275, w14276, w14277, w14278, w14279, w14280, w14281, w14282, w14283, w14284, w14285, w14286, w14287, w14288, w14289, w14290, w14291, w14292, w14293, w14294, w14295, w14296, w14297, w14298, w14299, w14300, w14301, w14302, w14303, w14304, w14305, w14306, w14307, w14308, w14309, w14310, w14311, w14312, w14313, w14314, w14315, w14316, w14317, w14318, w14319, w14320, w14321, w14322, w14323, w14324, w14325, w14326, w14327, w14328, w14329, w14330, w14331, w14332, w14333, w14334, w14335, w14336, w14337, w14338, w14339, w14340, w14341, w14342, w14343, w14344, w14345, w14346, w14347, w14348, w14349, w14350, w14351, w14352, w14353, w14354, w14355, w14356, w14357, w14358, w14359, w14360, w14361, w14362, w14363, w14364, w14365, w14366, w14367, w14368, w14369, w14370, w14371, w14372, w14373, w14374, w14375, w14376, w14377, w14378, w14379, w14380, w14381, w14382, w14383, w14384, w14385, w14386, w14387, w14388, w14389, w14390, w14391, w14392, w14393, w14394, w14395, w14396, w14397, w14398, w14399, w14400, w14401, w14402, w14403, w14404, w14405, w14406, w14407, w14408, w14409, w14410, w14411, w14412, w14413, w14414, w14415, w14416, w14417, w14418, w14419, w14420, w14421, w14422, w14423, w14424, w14425, w14426, w14427, w14428, w14429, w14430, w14431, w14432, w14433, w14434, w14435, w14436, w14437, w14438, w14439, w14440, w14441, w14442, w14443, w14444, w14445, w14446, w14447, w14448, w14449, w14450, w14451, w14452, w14453, w14454, w14455, w14456, w14457, w14458, w14459, w14460, w14461, w14462, w14463, w14464, w14465, w14466, w14467, w14468, w14469, w14470, w14471, w14472, w14473, w14474, w14475, w14476, w14477, w14478, w14479, w14480, w14481, w14482, w14483, w14484, w14485, w14486, w14487, w14488, w14489, w14490, w14491, w14492, w14493, w14494, w14495, w14496, w14497, w14498, w14499, w14500, w14501, w14502, w14503, w14504, w14505, w14506, w14507, w14508, w14509, w14510, w14511, w14512, w14513, w14514, w14515, w14516, w14517, w14518, w14519, w14520, w14521, w14522, w14523, w14524, w14525, w14526, w14527, w14528, w14529, w14530, w14531, w14532, w14533, w14534, w14535, w14536, w14537, w14538, w14539, w14540, w14541, w14542, w14543, w14544, w14545, w14546, w14547, w14548, w14549, w14550, w14551, w14552, w14553, w14554, w14555, w14556, w14557, w14558, w14559, w14560, w14561, w14562, w14563, w14564, w14565, w14566, w14567, w14568, w14569, w14570, w14571, w14572, w14573, w14574, w14575, w14576, w14577, w14578, w14579, w14580, w14581, w14582, w14583, w14584, w14585, w14586, w14587, w14588, w14589, w14590, w14591, w14592, w14593, w14594, w14595, w14596, w14597, w14598, w14599, w14600, w14601, w14602, w14603, w14604, w14605, w14606, w14607, w14608, w14609, w14610, w14611, w14612, w14613, w14614, w14615, w14616, w14617, w14618, w14619, w14620, w14621, w14622, w14623, w14624, w14625, w14626, w14627, w14628, w14629, w14630, w14631, w14632, w14633, w14634, w14635, w14636, w14637, w14638, w14639, w14640, w14641, w14642, w14643, w14644, w14645, w14646, w14647, w14648, w14649, w14650, w14651, w14652, w14653, w14654, w14655, w14656, w14657, w14658, w14659, w14660, w14661, w14662, w14663, w14664, w14665, w14666, w14667, w14668, w14669, w14670, w14671, w14672, w14673, w14674, w14675, w14676, w14677, w14678, w14679, w14680, w14681, w14682, w14683, w14684, w14685, w14686, w14687, w14688, w14689, w14690, w14691, w14692, w14693, w14694, w14695, w14696, w14697, w14698, w14699, w14700, w14701, w14702, w14703, w14704, w14705, w14706, w14707, w14708, w14709, w14710, w14711, w14712, w14713, w14714, w14715, w14716, w14717, w14718, w14719, w14720, w14721, w14722, w14723, w14724, w14725, w14726, w14727, w14728, w14729, w14730, w14731, w14732, w14733, w14734, w14735, w14736, w14737, w14738, w14739, w14740, w14741, w14742, w14743, w14744, w14745, w14746, w14747, w14748, w14749, w14750, w14751, w14752, w14753, w14754, w14755, w14756, w14757, w14758, w14759, w14760, w14761, w14762, w14763, w14764, w14765, w14766, w14767, w14768, w14769, w14770, w14771, w14772, w14773, w14774, w14775, w14776, w14777, w14778, w14779, w14780, w14781, w14782, w14783, w14784, w14785, w14786, w14787, w14788, w14789, w14790, w14791, w14792, w14793, w14794, w14795, w14796, w14797, w14798, w14799, w14800, w14801, w14802, w14803, w14804, w14805, w14806, w14807, w14808, w14809, w14810, w14811, w14812, w14813, w14814, w14815, w14816, w14817, w14818, w14819, w14820, w14821, w14822, w14823, w14824, w14825, w14826, w14827, w14828, w14829, w14830, w14831, w14832, w14833, w14834, w14835, w14836, w14837, w14838, w14839, w14840, w14841, w14842, w14843, w14844, w14845, w14846, w14847, w14848, w14849, w14850, w14851, w14852, w14853, w14854, w14855, w14856, w14857, w14858, w14859, w14860, w14861, w14862, w14863, w14864, w14865, w14866, w14867, w14868, w14869, w14870, w14871, w14872, w14873, w14874, w14875, w14876, w14877, w14878, w14879, w14880, w14881, w14882, w14883, w14884, w14885, w14886, w14887, w14888, w14889, w14890, w14891, w14892, w14893, w14894, w14895, w14896, w14897, w14898, w14899, w14900, w14901, w14902, w14903, w14904, w14905, w14906, w14907, w14908, w14909, w14910, w14911, w14912, w14913, w14914, w14915, w14916, w14917, w14918, w14919, w14920, w14921, w14922, w14923, w14924, w14925, w14926, w14927, w14928, w14929, w14930, w14931, w14932, w14933, w14934, w14935, w14936, w14937, w14938, w14939, w14940, w14941, w14942, w14943, w14944, w14945, w14946, w14947, w14948, w14949, w14950, w14951, w14952, w14953, w14954, w14955, w14956, w14957, w14958, w14959, w14960, w14961, w14962, w14963, w14964, w14965, w14966, w14967, w14968, w14969, w14970, w14971, w14972, w14973, w14974, w14975, w14976, w14977, w14978, w14979, w14980, w14981, w14982, w14983, w14984, w14985, w14986, w14987, w14988, w14989, w14990, w14991, w14992, w14993, w14994, w14995, w14996, w14997, w14998, w14999, w15000, w15001, w15002, w15003, w15004, w15005, w15006, w15007, w15008, w15009, w15010, w15011, w15012, w15013, w15014, w15015, w15016, w15017, w15018, w15019, w15020, w15021, w15022, w15023, w15024, w15025, w15026, w15027, w15028, w15029, w15030, w15031, w15032, w15033, w15034, w15035, w15036, w15037, w15038, w15039, w15040, w15041, w15042, w15043, w15044, w15045, w15046, w15047, w15048, w15049, w15050, w15051, w15052, w15053, w15054, w15055, w15056, w15057, w15058, w15059, w15060, w15061, w15062, w15063, w15064, w15065, w15066, w15067, w15068, w15069, w15070, w15071, w15072, w15073, w15074, w15075, w15076, w15077, w15078, w15079, w15080, w15081, w15082, w15083, w15084, w15085, w15086, w15087, w15088, w15089, w15090, w15091, w15092, w15093, w15094, w15095, w15096, w15097, w15098, w15099, w15100, w15101, w15102, w15103, w15104, w15105, w15106, w15107, w15108, w15109, w15110, w15111, w15112, w15113, w15114, w15115, w15116, w15117, w15118, w15119, w15120, w15121, w15122, w15123, w15124, w15125, w15126, w15127, w15128, w15129, w15130, w15131, w15132, w15133, w15134, w15135, w15136, w15137, w15138, w15139, w15140, w15141, w15142, w15143, w15144, w15145, w15146, w15147, w15148, w15149, w15150, w15151, w15152, w15153, w15154, w15155, w15156, w15157, w15158, w15159, w15160, w15161, w15162, w15163, w15164, w15165, w15166, w15167, w15168, w15169, w15170, w15171, w15172, w15173, w15174, w15175, w15176, w15177, w15178, w15179, w15180, w15181, w15182, w15183, w15184, w15185, w15186, w15187, w15188, w15189, w15190, w15191, w15192, w15193, w15194, w15195, w15196, w15197, w15198, w15199, w15200, w15201, w15202, w15203, w15204, w15205, w15206, w15207, w15208, w15209, w15210, w15211, w15212, w15213, w15214, w15215, w15216, w15217, w15218, w15219, w15220, w15221, w15222, w15223, w15224, w15225, w15226, w15227, w15228, w15229, w15230, w15231, w15232, w15233, w15234, w15235, w15236, w15237, w15238, w15239, w15240, w15241, w15242, w15243, w15244, w15245, w15246, w15247, w15248, w15249, w15250, w15251, w15252, w15253, w15254, w15255, w15256, w15257, w15258, w15259, w15260, w15261, w15262, w15263, w15264, w15265, w15266, w15267, w15268, w15269, w15270, w15271, w15272, w15273, w15274, w15275, w15276, w15277, w15278, w15279, w15280, w15281, w15282, w15283, w15284, w15285, w15286, w15287, w15288, w15289, w15290, w15291, w15292, w15293, w15294, w15295, w15296, w15297, w15298, w15299, w15300, w15301, w15302, w15303, w15304, w15305, w15306, w15307, w15308, w15309, w15310, w15311, w15312, w15313, w15314, w15315, w15316, w15317, w15318, w15319, w15320, w15321, w15322, w15323, w15324, w15325, w15326, w15327, w15328, w15329, w15330, w15331, w15332, w15333, w15334, w15335, w15336, w15337, w15338, w15339, w15340, w15341, w15342, w15343, w15344, w15345, w15346, w15347, w15348, w15349, w15350, w15351, w15352, w15353, w15354, w15355, w15356, w15357, w15358, w15359, w15360, w15361, w15362, w15363, w15364, w15365, w15366, w15367, w15368, w15369, w15370, w15371, w15372, w15373, w15374, w15375, w15376, w15377, w15378, w15379, w15380, w15381, w15382, w15383, w15384, w15385, w15386, w15387, w15388, w15389, w15390, w15391, w15392, w15393, w15394, w15395, w15396, w15397, w15398, w15399, w15400, w15401, w15402, w15403, w15404, w15405, w15406, w15407, w15408, w15409, w15410, w15411, w15412, w15413, w15414, w15415, w15416, w15417, w15418, w15419, w15420, w15421, w15422, w15423, w15424, w15425, w15426, w15427, w15428, w15429, w15430, w15431, w15432, w15433, w15434, w15435, w15436, w15437, w15438, w15439, w15440, w15441, w15442, w15443, w15444, w15445, w15446, w15447, w15448, w15449, w15450, w15451, w15452, w15453, w15454, w15455, w15456, w15457, w15458, w15459, w15460, w15461, w15462, w15463, w15464, w15465, w15466, w15467, w15468, w15469, w15470, w15471, w15472, w15473, w15474, w15475, w15476, w15477, w15478, w15479, w15480, w15481, w15482, w15483, w15484, w15485, w15486, w15487, w15488, w15489, w15490, w15491, w15492, w15493, w15494, w15495, w15496, w15497, w15498, w15499, w15500, w15501, w15502, w15503, w15504, w15505, w15506, w15507, w15508, w15509, w15510, w15511, w15512, w15513, w15514, w15515, w15516, w15517, w15518, w15519, w15520, w15521, w15522, w15523, w15524, w15525, w15526, w15527, w15528, w15529, w15530, w15531, w15532, w15533, w15534, w15535, w15536, w15537, w15538, w15539, w15540, w15541, w15542, w15543, w15544, w15545, w15546, w15547, w15548, w15549, w15550, w15551, w15552, w15553, w15554, w15555, w15556, w15557, w15558, w15559, w15560, w15561, w15562, w15563, w15564, w15565, w15566, w15567, w15568, w15569, w15570, w15571, w15572, w15573, w15574, w15575, w15576, w15577, w15578, w15579, w15580, w15581, w15582, w15583, w15584, w15585, w15586, w15587, w15588, w15589, w15590, w15591, w15592, w15593, w15594, w15595, w15596, w15597, w15598, w15599, w15600, w15601, w15602, w15603, w15604, w15605, w15606, w15607, w15608, w15609, w15610, w15611, w15612, w15613, w15614, w15615, w15616, w15617, w15618, w15619, w15620, w15621, w15622, w15623, w15624, w15625, w15626, w15627, w15628, w15629, w15630, w15631, w15632, w15633, w15634, w15635, w15636, w15637, w15638, w15639, w15640, w15641, w15642, w15643, w15644, w15645, w15646, w15647, w15648, w15649, w15650, w15651, w15652, w15653, w15654, w15655, w15656, w15657, w15658, w15659, w15660, w15661, w15662, w15663, w15664, w15665, w15666, w15667, w15668, w15669, w15670, w15671, w15672, w15673, w15674, w15675, w15676, w15677, w15678, w15679, w15680, w15681, w15682, w15683, w15684, w15685, w15686, w15687, w15688, w15689, w15690, w15691, w15692, w15693, w15694, w15695, w15696, w15697, w15698, w15699, w15700, w15701, w15702, w15703, w15704, w15705, w15706, w15707, w15708, w15709, w15710, w15711, w15712, w15713, w15714, w15715, w15716, w15717, w15718, w15719, w15720, w15721, w15722, w15723, w15724, w15725, w15726, w15727, w15728, w15729, w15730, w15731, w15732, w15733, w15734, w15735, w15736, w15737, w15738, w15739, w15740, w15741, w15742, w15743, w15744, w15745, w15746, w15747, w15748, w15749, w15750, w15751, w15752, w15753, w15754, w15755, w15756, w15757, w15758, w15759, w15760, w15761, w15762, w15763, w15764, w15765, w15766, w15767, w15768, w15769, w15770, w15771, w15772, w15773, w15774, w15775, w15776, w15777, w15778, w15779, w15780, w15781, w15782, w15783, w15784, w15785, w15786, w15787, w15788, w15789, w15790, w15791, w15792, w15793, w15794, w15795, w15796, w15797, w15798, w15799, w15800, w15801, w15802, w15803, w15804, w15805, w15806, w15807, w15808, w15809, w15810, w15811, w15812, w15813, w15814, w15815, w15816, w15817, w15818, w15819, w15820, w15821, w15822, w15823, w15824, w15825, w15826, w15827, w15828, w15829, w15830, w15831, w15832, w15833, w15834, w15835, w15836, w15837, w15838, w15839, w15840, w15841, w15842, w15843, w15844, w15845, w15846, w15847, w15848, w15849, w15850, w15851, w15852, w15853, w15854, w15855, w15856, w15857, w15858, w15859, w15860, w15861, w15862, w15863, w15864, w15865, w15866, w15867, w15868, w15869, w15870, w15871, w15872, w15873, w15874, w15875, w15876, w15877, w15878, w15879, w15880, w15881, w15882, w15883, w15884, w15885, w15886, w15887, w15888, w15889, w15890, w15891, w15892, w15893, w15894, w15895, w15896, w15897, w15898, w15899, w15900, w15901, w15902, w15903, w15904, w15905, w15906, w15907, w15908, w15909, w15910, w15911, w15912, w15913, w15914, w15915, w15916, w15917, w15918, w15919, w15920, w15921, w15922, w15923, w15924, w15925, w15926, w15927, w15928, w15929, w15930, w15931, w15932, w15933, w15934, w15935, w15936, w15937, w15938, w15939, w15940, w15941, w15942, w15943, w15944, w15945, w15946, w15947, w15948, w15949, w15950, w15951, w15952, w15953, w15954, w15955, w15956, w15957, w15958, w15959, w15960, w15961, w15962, w15963, w15964, w15965, w15966, w15967, w15968, w15969, w15970, w15971, w15972, w15973, w15974, w15975, w15976, w15977, w15978, w15979, w15980, w15981, w15982, w15983, w15984, w15985, w15986, w15987, w15988, w15989, w15990, w15991, w15992, w15993, w15994, w15995, w15996, w15997, w15998, w15999, w16000, w16001, w16002, w16003, w16004, w16005, w16006, w16007, w16008, w16009, w16010, w16011, w16012, w16013, w16014, w16015, w16016, w16017, w16018, w16019, w16020, w16021, w16022, w16023, w16024, w16025, w16026, w16027, w16028, w16029, w16030, w16031, w16032, w16033, w16034, w16035, w16036, w16037, w16038, w16039, w16040, w16041, w16042, w16043, w16044, w16045, w16046, w16047, w16048, w16049, w16050, w16051, w16052, w16053, w16054, w16055, w16056, w16057, w16058, w16059, w16060, w16061, w16062, w16063, w16064, w16065, w16066, w16067, w16068, w16069, w16070, w16071, w16072, w16073, w16074, w16075, w16076, w16077, w16078, w16079, w16080, w16081, w16082, w16083, w16084, w16085, w16086, w16087, w16088, w16089, w16090, w16091, w16092, w16093, w16094, w16095, w16096, w16097, w16098, w16099, w16100, w16101, w16102, w16103, w16104, w16105, w16106, w16107, w16108, w16109, w16110, w16111, w16112, w16113, w16114, w16115, w16116, w16117, w16118, w16119, w16120, w16121, w16122, w16123, w16124, w16125, w16126, w16127, w16128, w16129, w16130, w16131, w16132, w16133, w16134, w16135, w16136, w16137, w16138, w16139, w16140, w16141, w16142, w16143, w16144, w16145, w16146, w16147, w16148, w16149, w16150, w16151, w16152, w16153, w16154, w16155, w16156, w16157, w16158, w16159, w16160, w16161, w16162, w16163, w16164, w16165, w16166, w16167, w16168, w16169, w16170, w16171, w16172, w16173, w16174, w16175, w16176, w16177, w16178, w16179, w16180, w16181, w16182, w16183, w16184, w16185, w16186, w16187, w16188, w16189, w16190, w16191, w16192, w16193, w16194, w16195, w16196, w16197, w16198, w16199, w16200, w16201, w16202, w16203, w16204, w16205, w16206, w16207, w16208, w16209, w16210, w16211, w16212, w16213, w16214, w16215, w16216, w16217, w16218, w16219, w16220, w16221, w16222, w16223, w16224, w16225, w16226, w16227, w16228, w16229, w16230, w16231, w16232, w16233, w16234, w16235, w16236, w16237, w16238, w16239, w16240, w16241, w16242, w16243, w16244, w16245, w16246, w16247, w16248, w16249, w16250, w16251, w16252, w16253, w16254, w16255, w16256, w16257, w16258, w16259, w16260, w16261, w16262, w16263, w16264, w16265, w16266, w16267, w16268, w16269, w16270, w16271, w16272, w16273, w16274, w16275, w16276, w16277, w16278, w16279, w16280, w16281, w16282, w16283, w16284, w16285, w16286, w16287, w16288, w16289, w16290, w16291, w16292, w16293, w16294, w16295, w16296, w16297, w16298, w16299, w16300, w16301, w16302, w16303, w16304, w16305, w16306, w16307, w16308, w16309, w16310, w16311, w16312, w16313, w16314, w16315, w16316, w16317, w16318, w16319, w16320, w16321, w16322, w16323, w16324, w16325, w16326, w16327, w16328, w16329, w16330, w16331, w16332, w16333, w16334, w16335, w16336, w16337, w16338, w16339, w16340, w16341, w16342, w16343, w16344, w16345, w16346, w16347, w16348, w16349, w16350, w16351, w16352, w16353, w16354, w16355, w16356, w16357, w16358, w16359, w16360, w16361, w16362, w16363, w16364, w16365, w16366, w16367, w16368, w16369, w16370, w16371, w16372, w16373, w16374, w16375, w16376, w16377, w16378, w16379, w16380, w16381, w16382, w16383, w16384, w16385, w16386, w16387, w16388, w16389, w16390, w16391, w16392, w16393, w16394, w16395, w16396, w16397, w16398, w16399, w16400, w16401, w16402, w16403, w16404, w16405, w16406, w16407, w16408, w16409, w16410, w16411, w16412, w16413, w16414, w16415, w16416, w16417, w16418, w16419, w16420, w16421, w16422, w16423, w16424, w16425, w16426, w16427, w16428, w16429, w16430, w16431, w16432, w16433, w16434, w16435, w16436, w16437, w16438, w16439, w16440, w16441, w16442, w16443, w16444, w16445, w16446, w16447, w16448, w16449, w16450, w16451, w16452, w16453, w16454, w16455, w16456, w16457, w16458, w16459, w16460, w16461, w16462, w16463, w16464, w16465, w16466, w16467, w16468, w16469, w16470, w16471, w16472, w16473, w16474, w16475, w16476, w16477, w16478, w16479, w16480, w16481, w16482, w16483, w16484, w16485, w16486, w16487, w16488, w16489, w16490, w16491, w16492, w16493, w16494, w16495, w16496, w16497, w16498, w16499, w16500, w16501, w16502, w16503, w16504, w16505, w16506, w16507, w16508, w16509, w16510, w16511, w16512, w16513, w16514, w16515, w16516, w16517, w16518, w16519, w16520, w16521, w16522, w16523, w16524, w16525, w16526, w16527, w16528, w16529, w16530, w16531, w16532, w16533, w16534, w16535, w16536, w16537, w16538, w16539, w16540, w16541, w16542, w16543, w16544, w16545, w16546, w16547, w16548, w16549, w16550, w16551, w16552, w16553, w16554, w16555, w16556, w16557, w16558, w16559, w16560, w16561, w16562, w16563, w16564, w16565, w16566, w16567, w16568, w16569, w16570, w16571, w16572, w16573, w16574, w16575, w16576, w16577, w16578, w16579, w16580, w16581, w16582, w16583, w16584, w16585, w16586, w16587, w16588, w16589, w16590, w16591, w16592, w16593, w16594, w16595, w16596, w16597, w16598, w16599, w16600, w16601, w16602, w16603, w16604, w16605, w16606, w16607, w16608, w16609, w16610, w16611, w16612, w16613, w16614, w16615, w16616, w16617, w16618, w16619, w16620, w16621, w16622, w16623, w16624, w16625, w16626, w16627, w16628, w16629, w16630, w16631, w16632, w16633, w16634, w16635, w16636, w16637, w16638, w16639, w16640, w16641, w16642, w16643, w16644, w16645, w16646, w16647, w16648, w16649, w16650, w16651, w16652, w16653, w16654, w16655, w16656, w16657, w16658, w16659, w16660, w16661, w16662, w16663, w16664, w16665, w16666, w16667, w16668, w16669, w16670, w16671, w16672, w16673, w16674, w16675, w16676, w16677, w16678, w16679, w16680, w16681, w16682, w16683, w16684, w16685, w16686, w16687, w16688, w16689, w16690, w16691, w16692, w16693, w16694, w16695, w16696, w16697, w16698, w16699, w16700, w16701, w16702, w16703, w16704, w16705, w16706, w16707, w16708, w16709, w16710, w16711, w16712, w16713, w16714, w16715, w16716, w16717, w16718, w16719, w16720, w16721, w16722, w16723, w16724, w16725, w16726, w16727, w16728, w16729, w16730, w16731, w16732, w16733, w16734, w16735, w16736, w16737, w16738, w16739, w16740, w16741, w16742, w16743, w16744, w16745, w16746, w16747, w16748, w16749, w16750, w16751, w16752, w16753, w16754, w16755, w16756, w16757, w16758, w16759, w16760, w16761, w16762, w16763, w16764, w16765, w16766, w16767, w16768, w16769, w16770, w16771, w16772, w16773, w16774, w16775, w16776, w16777, w16778, w16779, w16780, w16781, w16782, w16783, w16784, w16785, w16786, w16787, w16788, w16789, w16790, w16791, w16792, w16793, w16794, w16795, w16796, w16797, w16798, w16799, w16800, w16801, w16802, w16803, w16804, w16805, w16806, w16807, w16808, w16809, w16810, w16811, w16812, w16813, w16814, w16815, w16816, w16817, w16818, w16819, w16820, w16821, w16822, w16823, w16824, w16825, w16826, w16827, w16828, w16829, w16830, w16831, w16832, w16833, w16834, w16835, w16836, w16837, w16838, w16839, w16840, w16841, w16842, w16843, w16844, w16845, w16846, w16847, w16848, w16849, w16850, w16851, w16852, w16853, w16854, w16855, w16856, w16857, w16858, w16859, w16860, w16861, w16862, w16863, w16864, w16865, w16866, w16867, w16868, w16869, w16870, w16871, w16872, w16873, w16874, w16875, w16876, w16877, w16878, w16879, w16880, w16881, w16882, w16883, w16884, w16885, w16886, w16887, w16888, w16889, w16890, w16891, w16892, w16893, w16894, w16895, w16896, w16897, w16898, w16899, w16900, w16901, w16902, w16903, w16904, w16905, w16906, w16907, w16908, w16909, w16910, w16911, w16912, w16913, w16914, w16915, w16916, w16917, w16918, w16919, w16920, w16921, w16922, w16923, w16924, w16925, w16926, w16927, w16928, w16929, w16930, w16931, w16932, w16933, w16934, w16935, w16936, w16937, w16938, w16939, w16940, w16941, w16942, w16943, w16944, w16945, w16946, w16947, w16948, w16949, w16950, w16951, w16952, w16953, w16954, w16955, w16956, w16957, w16958, w16959, w16960, w16961, w16962, w16963, w16964, w16965, w16966, w16967, w16968, w16969, w16970, w16971, w16972, w16973, w16974, w16975, w16976, w16977, w16978, w16979, w16980, w16981, w16982, w16983, w16984, w16985, w16986, w16987, w16988, w16989, w16990, w16991, w16992, w16993, w16994, w16995, w16996, w16997, w16998, w16999, w17000, w17001, w17002, w17003, w17004, w17005, w17006, w17007, w17008, w17009, w17010, w17011, w17012, w17013, w17014, w17015, w17016, w17017, w17018, w17019, w17020, w17021, w17022, w17023, w17024, w17025, w17026, w17027, w17028, w17029, w17030, w17031, w17032, w17033, w17034, w17035, w17036, w17037, w17038, w17039, w17040, w17041, w17042, w17043, w17044, w17045, w17046, w17047, w17048, w17049, w17050, w17051, w17052, w17053, w17054, w17055, w17056, w17057, w17058, w17059, w17060, w17061, w17062, w17063, w17064, w17065, w17066, w17067, w17068, w17069, w17070, w17071, w17072, w17073, w17074, w17075, w17076, w17077, w17078, w17079, w17080, w17081, w17082, w17083, w17084, w17085, w17086, w17087, w17088, w17089, w17090, w17091, w17092, w17093, w17094, w17095, w17096, w17097, w17098, w17099, w17100, w17101, w17102, w17103, w17104, w17105, w17106, w17107, w17108, w17109, w17110, w17111, w17112, w17113, w17114, w17115, w17116, w17117, w17118, w17119, w17120, w17121, w17122, w17123, w17124, w17125, w17126, w17127, w17128, w17129, w17130, w17131, w17132, w17133, w17134, w17135, w17136, w17137, w17138, w17139, w17140, w17141, w17142, w17143, w17144, w17145, w17146, w17147, w17148, w17149, w17150, w17151, w17152, w17153, w17154, w17155, w17156, w17157, w17158, w17159, w17160, w17161, w17162, w17163, w17164, w17165, w17166, w17167, w17168, w17169, w17170, w17171, w17172, w17173, w17174, w17175, w17176, w17177, w17178, w17179, w17180, w17181, w17182, w17183, w17184, w17185, w17186, w17187, w17188, w17189, w17190, w17191, w17192, w17193, w17194, w17195, w17196, w17197, w17198, w17199, w17200, w17201, w17202, w17203, w17204, w17205, w17206, w17207, w17208, w17209, w17210, w17211, w17212, w17213, w17214, w17215, w17216, w17217, w17218, w17219, w17220, w17221, w17222, w17223, w17224, w17225, w17226, w17227, w17228, w17229, w17230, w17231, w17232, w17233, w17234, w17235, w17236, w17237, w17238, w17239, w17240, w17241, w17242, w17243, w17244, w17245, w17246, w17247, w17248, w17249, w17250, w17251, w17252, w17253, w17254, w17255, w17256, w17257, w17258, w17259, w17260, w17261, w17262, w17263, w17264, w17265, w17266, w17267, w17268, w17269, w17270, w17271, w17272, w17273, w17274, w17275, w17276, w17277, w17278, w17279, w17280, w17281, w17282, w17283, w17284, w17285, w17286, w17287, w17288, w17289, w17290, w17291, w17292, w17293, w17294, w17295, w17296, w17297, w17298, w17299, w17300, w17301, w17302, w17303, w17304, w17305, w17306, w17307, w17308, w17309, w17310, w17311, w17312, w17313, w17314, w17315, w17316, w17317, w17318, w17319, w17320, w17321, w17322, w17323, w17324, w17325, w17326, w17327, w17328, w17329, w17330, w17331, w17332, w17333, w17334, w17335, w17336, w17337, w17338, w17339, w17340, w17341, w17342, w17343, w17344, w17345, w17346, w17347, w17348, w17349, w17350, w17351, w17352, w17353, w17354, w17355, w17356, w17357, w17358, w17359, w17360, w17361, w17362, w17363, w17364, w17365, w17366, w17367, w17368, w17369, w17370, w17371, w17372, w17373, w17374, w17375, w17376, w17377, w17378, w17379, w17380, w17381, w17382, w17383, w17384, w17385, w17386, w17387, w17388, w17389, w17390, w17391, w17392, w17393, w17394, w17395, w17396, w17397, w17398, w17399, w17400, w17401, w17402, w17403, w17404, w17405, w17406, w17407, w17408, w17409, w17410, w17411, w17412, w17413, w17414, w17415, w17416, w17417, w17418, w17419, w17420, w17421, w17422, w17423, w17424, w17425, w17426, w17427, w17428, w17429, w17430, w17431, w17432, w17433, w17434, w17435, w17436, w17437, w17438, w17439, w17440, w17441, w17442, w17443, w17444, w17445, w17446, w17447, w17448, w17449, w17450, w17451, w17452, w17453, w17454, w17455, w17456, w17457, w17458, w17459, w17460, w17461, w17462, w17463, w17464, w17465, w17466, w17467, w17468, w17469, w17470, w17471, w17472, w17473, w17474, w17475, w17476, w17477, w17478, w17479, w17480, w17481, w17482, w17483, w17484, w17485, w17486, w17487, w17488, w17489, w17490, w17491, w17492, w17493, w17494, w17495, w17496, w17497, w17498, w17499, w17500, w17501, w17502, w17503, w17504, w17505, w17506, w17507, w17508, w17509, w17510, w17511, w17512, w17513, w17514, w17515, w17516, w17517, w17518, w17519, w17520, w17521, w17522, w17523, w17524, w17525, w17526, w17527, w17528, w17529, w17530, w17531, w17532, w17533, w17534, w17535, w17536, w17537, w17538, w17539, w17540, w17541, w17542, w17543, w17544, w17545, w17546, w17547, w17548, w17549, w17550, w17551, w17552, w17553, w17554, w17555, w17556, w17557, w17558, w17559, w17560, w17561, w17562, w17563, w17564, w17565, w17566, w17567, w17568, w17569, w17570, w17571, w17572, w17573, w17574, w17575, w17576, w17577, w17578, w17579, w17580, w17581, w17582, w17583, w17584, w17585, w17586, w17587, w17588, w17589, w17590, w17591, w17592, w17593, w17594, w17595, w17596, w17597, w17598, w17599, w17600, w17601, w17602, w17603, w17604, w17605, w17606, w17607, w17608, w17609, w17610, w17611, w17612, w17613, w17614, w17615, w17616, w17617, w17618, w17619, w17620, w17621, w17622, w17623, w17624, w17625, w17626, w17627, w17628, w17629, w17630, w17631, w17632, w17633, w17634, w17635, w17636, w17637, w17638, w17639, w17640, w17641, w17642, w17643, w17644, w17645, w17646, w17647, w17648, w17649, w17650, w17651, w17652, w17653, w17654, w17655, w17656, w17657, w17658, w17659, w17660, w17661, w17662, w17663, w17664, w17665, w17666, w17667, w17668, w17669, w17670, w17671, w17672, w17673, w17674, w17675, w17676, w17677, w17678, w17679, w17680, w17681, w17682, w17683, w17684, w17685, w17686, w17687, w17688, w17689, w17690, w17691, w17692, w17693, w17694, w17695, w17696, w17697, w17698, w17699, w17700, w17701, w17702, w17703, w17704, w17705, w17706, w17707, w17708, w17709, w17710, w17711, w17712, w17713, w17714, w17715, w17716, w17717, w17718, w17719, w17720, w17721, w17722, w17723, w17724, w17725, w17726, w17727, w17728, w17729, w17730, w17731, w17732, w17733, w17734, w17735, w17736, w17737, w17738, w17739, w17740, w17741, w17742, w17743, w17744, w17745, w17746, w17747, w17748, w17749, w17750, w17751, w17752, w17753, w17754, w17755, w17756, w17757, w17758, w17759, w17760, w17761, w17762, w17763, w17764, w17765, w17766, w17767, w17768, w17769, w17770, w17771, w17772, w17773, w17774, w17775, w17776, w17777, w17778, w17779, w17780, w17781, w17782, w17783, w17784, w17785, w17786, w17787, w17788, w17789, w17790, w17791, w17792, w17793, w17794, w17795, w17796, w17797, w17798, w17799, w17800, w17801, w17802, w17803, w17804, w17805, w17806, w17807, w17808, w17809, w17810, w17811, w17812, w17813, w17814, w17815, w17816, w17817, w17818, w17819, w17820, w17821, w17822, w17823, w17824, w17825, w17826, w17827, w17828, w17829, w17830, w17831, w17832, w17833, w17834, w17835, w17836, w17837, w17838, w17839, w17840, w17841, w17842, w17843, w17844, w17845, w17846, w17847, w17848, w17849, w17850, w17851, w17852, w17853, w17854, w17855, w17856, w17857, w17858, w17859, w17860, w17861, w17862, w17863, w17864, w17865, w17866, w17867, w17868, w17869, w17870, w17871, w17872, w17873, w17874, w17875, w17876, w17877, w17878, w17879, w17880, w17881, w17882, w17883, w17884, w17885, w17886, w17887, w17888, w17889, w17890, w17891, w17892, w17893, w17894, w17895, w17896, w17897, w17898, w17899, w17900, w17901, w17902, w17903, w17904, w17905, w17906, w17907, w17908, w17909, w17910, w17911, w17912, w17913, w17914, w17915, w17916, w17917, w17918, w17919, w17920, w17921, w17922, w17923, w17924, w17925, w17926, w17927, w17928, w17929, w17930, w17931, w17932, w17933, w17934, w17935, w17936, w17937, w17938, w17939, w17940, w17941, w17942, w17943, w17944, w17945, w17946, w17947, w17948, w17949, w17950, w17951, w17952, w17953, w17954, w17955, w17956, w17957, w17958, w17959, w17960, w17961, w17962, w17963, w17964, w17965, w17966, w17967, w17968, w17969, w17970, w17971, w17972, w17973, w17974, w17975, w17976, w17977, w17978, w17979, w17980, w17981, w17982, w17983, w17984, w17985, w17986, w17987, w17988, w17989, w17990, w17991, w17992, w17993, w17994, w17995, w17996, w17997, w17998, w17999, w18000, w18001, w18002, w18003, w18004, w18005, w18006, w18007, w18008, w18009, w18010, w18011, w18012, w18013, w18014, w18015, w18016, w18017, w18018, w18019, w18020, w18021, w18022, w18023, w18024, w18025, w18026, w18027, w18028, w18029, w18030, w18031, w18032, w18033, w18034, w18035, w18036, w18037, w18038, w18039, w18040, w18041, w18042, w18043, w18044, w18045, w18046, w18047, w18048, w18049, w18050, w18051, w18052, w18053, w18054, w18055, w18056, w18057, w18058, w18059, w18060, w18061, w18062, w18063, w18064, w18065, w18066, w18067, w18068, w18069, w18070, w18071, w18072, w18073, w18074, w18075, w18076, w18077, w18078, w18079, w18080, w18081, w18082, w18083, w18084, w18085, w18086, w18087, w18088, w18089, w18090, w18091, w18092, w18093, w18094, w18095, w18096, w18097, w18098, w18099, w18100, w18101, w18102, w18103, w18104, w18105, w18106, w18107, w18108, w18109, w18110, w18111, w18112, w18113, w18114, w18115, w18116, w18117, w18118, w18119, w18120, w18121, w18122, w18123, w18124, w18125, w18126, w18127, w18128, w18129, w18130, w18131, w18132, w18133, w18134, w18135, w18136, w18137, w18138, w18139, w18140, w18141, w18142, w18143, w18144, w18145, w18146, w18147, w18148, w18149, w18150, w18151, w18152, w18153, w18154, w18155, w18156, w18157, w18158, w18159, w18160, w18161, w18162, w18163, w18164, w18165, w18166, w18167, w18168, w18169, w18170, w18171, w18172, w18173, w18174, w18175, w18176, w18177, w18178, w18179, w18180, w18181, w18182, w18183, w18184, w18185, w18186, w18187, w18188, w18189, w18190, w18191, w18192, w18193, w18194, w18195, w18196, w18197, w18198, w18199, w18200, w18201, w18202, w18203, w18204, w18205, w18206, w18207, w18208, w18209, w18210, w18211, w18212, w18213, w18214, w18215, w18216, w18217, w18218, w18219, w18220, w18221, w18222, w18223, w18224, w18225, w18226, w18227, w18228, w18229, w18230, w18231, w18232, w18233, w18234, w18235, w18236, w18237, w18238, w18239, w18240, w18241, w18242, w18243, w18244, w18245, w18246, w18247, w18248, w18249, w18250, w18251, w18252, w18253, w18254, w18255, w18256, w18257, w18258, w18259, w18260, w18261, w18262, w18263, w18264, w18265, w18266, w18267, w18268, w18269, w18270, w18271, w18272, w18273, w18274, w18275, w18276, w18277, w18278, w18279, w18280, w18281, w18282, w18283, w18284, w18285, w18286, w18287, w18288, w18289, w18290, w18291, w18292, w18293, w18294, w18295, w18296, w18297, w18298, w18299, w18300, w18301, w18302, w18303, w18304, w18305, w18306, w18307, w18308, w18309, w18310, w18311, w18312, w18313, w18314, w18315, w18316, w18317, w18318, w18319, w18320, w18321, w18322, w18323, w18324, w18325, w18326, w18327, w18328, w18329, w18330, w18331, w18332, w18333, w18334, w18335, w18336, w18337, w18338, w18339, w18340, w18341, w18342, w18343, w18344, w18345, w18346, w18347, w18348, w18349, w18350, w18351, w18352, w18353, w18354, w18355, w18356, w18357, w18358, w18359, w18360, w18361, w18362, w18363, w18364, w18365, w18366, w18367, w18368, w18369, w18370, w18371, w18372, w18373, w18374, w18375, w18376, w18377, w18378, w18379, w18380, w18381, w18382, w18383, w18384, w18385, w18386, w18387, w18388, w18389, w18390, w18391, w18392, w18393, w18394, w18395, w18396, w18397, w18398, w18399, w18400, w18401, w18402, w18403, w18404, w18405, w18406, w18407, w18408, w18409, w18410, w18411, w18412, w18413, w18414, w18415, w18416, w18417, w18418, w18419, w18420, w18421, w18422, w18423, w18424, w18425, w18426, w18427, w18428, w18429, w18430, w18431, w18432, w18433, w18434, w18435, w18436, w18437, w18438, w18439, w18440, w18441, w18442, w18443, w18444, w18445, w18446, w18447, w18448, w18449, w18450, w18451, w18452, w18453, w18454, w18455, w18456, w18457, w18458, w18459, w18460, w18461, w18462, w18463, w18464, w18465, w18466, w18467, w18468, w18469, w18470, w18471, w18472, w18473, w18474, w18475, w18476, w18477, w18478, w18479, w18480, w18481, w18482, w18483, w18484, w18485, w18486, w18487, w18488, w18489, w18490, w18491, w18492, w18493, w18494, w18495, w18496, w18497, w18498, w18499, w18500, w18501, w18502, w18503, w18504, w18505, w18506, w18507, w18508, w18509, w18510, w18511, w18512, w18513, w18514, w18515, w18516, w18517, w18518, w18519, w18520, w18521, w18522, w18523, w18524, w18525, w18526, w18527, w18528, w18529, w18530, w18531, w18532, w18533, w18534, w18535, w18536, w18537, w18538, w18539, w18540, w18541, w18542, w18543, w18544, w18545, w18546, w18547, w18548, w18549, w18550, w18551, w18552, w18553, w18554, w18555, w18556, w18557, w18558, w18559, w18560, w18561, w18562, w18563, w18564, w18565, w18566, w18567, w18568, w18569, w18570, w18571, w18572, w18573, w18574, w18575, w18576, w18577, w18578, w18579, w18580, w18581, w18582, w18583, w18584, w18585, w18586, w18587, w18588, w18589, w18590, w18591, w18592, w18593, w18594, w18595, w18596, w18597, w18598, w18599, w18600, w18601, w18602;
assign w0 = w15407 & w17892;
assign w1 = pi1379 & ~w4256;
assign w2 = (pi1192 & ~w5437) | (pi1192 & w4935) | (~w5437 & w4935);
assign w3 = pi1717 & ~w2253;
assign w4 = ~w16856 & ~w14321;
assign w5 = w11209 & ~w16110;
assign w6 = ~pi0986 & w15707;
assign w7 = ~w6895 & ~w8012;
assign w8 = w13509 & w6582;
assign w9 = pi1778 & w10335;
assign w10 = w13395 & w7112;
assign w11 = ~w18344 & ~w9205;
assign w12 = ~pi1936 & w16041;
assign w13 = ~w4288 & ~w3236;
assign w14 = ~w18145 & ~w15209;
assign w15 = ~pi1774 & pi3141;
assign w16 = w1962 & ~w7020;
assign w17 = pi1885 & ~w15036;
assign w18 = ~w14037 & ~w10757;
assign w19 = ~w1646 & ~w8544;
assign w20 = ~pi0295 & w4058;
assign w21 = ~w13451 & ~w800;
assign w22 = ~w3428 & ~w2236;
assign w23 = ~pi3092 & w16815;
assign w24 = pi1449 & ~w6448;
assign w25 = pi0043 & ~w14148;
assign w26 = pi1430 & ~w13753;
assign w27 = pi3507 & w13367;
assign w28 = ~pi1152 & pi1154;
assign w29 = ~w14046 & ~w15055;
assign w30 = ~w2341 & pi0834;
assign w31 = ~w3337 & ~w1720;
assign w32 = w4207 & w5995;
assign w33 = pi1529 & ~w14918;
assign w34 = ~pi2988 & w9504;
assign w35 = ~pi0621 & w14641;
assign w36 = pi1759 & ~w10389;
assign w37 = ~pi3053 & w6463;
assign w38 = ~w1741 & ~w2617;
assign w39 = ~w7097 & ~w3086;
assign w40 = ~pi0333 & w4058;
assign w41 = w16091 & w11248;
assign w42 = ~pi0281 & w4058;
assign w43 = pi2364 & ~w3223;
assign w44 = w13509 & w12590;
assign w45 = ~w14327 & ~w12469;
assign w46 = ~w7552 & ~w8578;
assign w47 = w3223 & w2753;
assign w48 = ~pi1764 & ~pi3171;
assign w49 = ~pi2992 & ~w3987;
assign w50 = ~w7844 & pi0608;
assign w51 = ~pi3287 & w17935;
assign w52 = ~w781 & ~w18317;
assign w53 = ~w14335 & ~w11789;
assign w54 = w14932 & w18301;
assign w55 = w8754 & w13221;
assign w56 = pi2845 & w14148;
assign w57 = ~w14228 & pi0634;
assign w58 = w14228 & ~w3374;
assign w59 = pi3082 & w16815;
assign w60 = ~pi2975 & w4508;
assign w61 = w13551 & w3796;
assign w62 = ~w8087 & w2206;
assign w63 = pi1950 & ~w14833;
assign w64 = w1368 & pi0381;
assign w65 = ~pi3164 & w1843;
assign w66 = ~w18476 & ~w12533;
assign w67 = ~w5824 & ~w16433;
assign w68 = ~pi2382 & w16041;
assign w69 = w3203 & ~w305;
assign w70 = ~pi0953 & w795;
assign w71 = ~pi3295 & w7090;
assign w72 = ~w15704 & ~w2181;
assign w73 = w10647 & ~w8099;
assign w74 = ~w14967 & ~w7103;
assign w75 = (w17562 & ~w7799) | (w17562 & w9832) | (~w7799 & w9832);
assign w76 = (pi0844 & ~w13509) | (pi0844 & w14441) | (~w13509 & w14441);
assign w77 = ~w9186 & ~w4088;
assign w78 = w16506 & ~w1340;
assign w79 = ~w4582 & ~w9597;
assign w80 = w11383 & w1072;
assign w81 = pi1494 & w13753;
assign w82 = w1391 & ~w9852;
assign w83 = ~pi3091 & w261;
assign w84 = ~w241 & ~w14928;
assign w85 = ~w1391 & pi0761;
assign w86 = ~w11483 & ~w9804;
assign w87 = pi2213 & ~w15271;
assign w88 = w7807 & w1946;
assign w89 = w10818 & ~w13091;
assign w90 = w14648 & ~pi2606;
assign w91 = w13509 & w12024;
assign w92 = ~w4163 & ~w17816;
assign w93 = ~w3381 & ~w10724;
assign w94 = pi1618 & ~w7090;
assign w95 = pi3066 & ~w16502;
assign w96 = ~w1391 & pi0777;
assign w97 = ~pi2039 & w13204;
assign w98 = ~w11469 & ~w7963;
assign w99 = pi1734 & ~w4058;
assign w100 = w10189 & pi0383;
assign w101 = (pi0381 & w5560) | (pi0381 & w64) | (w5560 & w64);
assign w102 = pi0115 & w3748;
assign w103 = ~w7844 & pi1001;
assign w104 = w10731 & w3129;
assign w105 = (pi0792 & ~w13509) | (pi0792 & w10380) | (~w13509 & w10380);
assign w106 = w6785 & ~w16498;
assign w107 = w14158 & w5547;
assign w108 = ~w1901 & w7413;
assign w109 = ~w400 & ~w6944;
assign w110 = pi3131 & ~pi3136;
assign w111 = ~w6865 & ~pi2920;
assign w112 = ~pi2026 & w7455;
assign w113 = ~pi0483 & pi3382;
assign w114 = ~pi3169 & w3982;
assign w115 = ~pi1906 & w11313;
assign w116 = (pi0772 & ~w13509) | (pi0772 & w4070) | (~w13509 & w4070);
assign w117 = ~pi0593 & w12825;
assign w118 = w11774 & w6443;
assign w119 = ~w6256 & ~w14883;
assign w120 = (pi1779 & w7215) | (pi1779 & w651) | (w7215 & w651);
assign w121 = w7959 & w1201;
assign w122 = ~w1391 & pi0764;
assign w123 = ~pi3154 & w3982;
assign w124 = ~pi0794 & w543;
assign w125 = pi2558 & ~w5274;
assign w126 = w2920 & pi0044;
assign w127 = (pi0701 & ~w13509) | (pi0701 & w5481) | (~w13509 & w5481);
assign w128 = ~w17018 & w11817;
assign w129 = w7703 & w5715;
assign w130 = ~w3470 & w11493;
assign w131 = w7842 & ~w14000;
assign w132 = ~pi1997 & w3019;
assign w133 = w15122 & ~pi2878;
assign w134 = w6575 & ~w3381;
assign w135 = w6224 & w5513;
assign w136 = w11209 & ~w13455;
assign w137 = ~pi3364 & ~pi3366;
assign w138 = ~w745 & ~w7496;
assign w139 = (pi1109 & ~w13509) | (pi1109 & w17567) | (~w13509 & w17567);
assign w140 = ~w344 & ~w11470;
assign w141 = pi2210 & ~w3223;
assign w142 = ~w7943 & ~w11038;
assign w143 = w7703 & w11837;
assign w144 = ~pi1954 & w11688;
assign w145 = ~w9507 & ~w5256;
assign w146 = ~w14560 & pi0225;
assign w147 = ~pi1322 & pi1345;
assign w148 = pi1323 & pi1345;
assign w149 = pi2440 & ~w3223;
assign w150 = ~w17427 & ~w16644;
assign w151 = ~w3069 & w14416;
assign w152 = w12460 & w16304;
assign w153 = pi1501 & ~w16922;
assign w154 = pi2414 & ~w3223;
assign w155 = (~w13367 & w17577) | (~w13367 & w6799) | (w17577 & w6799);
assign w156 = w10299 & w6320;
assign w157 = ~w18045 & ~w4759;
assign w158 = w6857 & w17933;
assign w159 = pi1451 & ~w6448;
assign w160 = ~w12857 & ~w13590;
assign w161 = pi1231 & ~pi1267;
assign w162 = w539 & ~w15223;
assign w163 = ~w8115 & ~w17082;
assign w164 = ~w10291 & ~w8458;
assign w165 = w11209 & ~w3283;
assign w166 = ~w10715 & w13435;
assign w167 = ~w9993 & ~w3653;
assign w168 = pi1596 & ~w13753;
assign w169 = w1391 & ~w2587;
assign w170 = w17477 & w5223;
assign w171 = ~w15328 & w10241;
assign w172 = (pi0367 & w6195) | (pi0367 & w8023) | (w6195 & w8023);
assign w173 = (~pi1775 & ~w7799) | (~pi1775 & w951) | (~w7799 & w951);
assign w174 = (pi0738 & ~w13509) | (pi0738 & w13375) | (~w13509 & w13375);
assign w175 = pi1182 & pi1195;
assign w176 = w7703 & w1053;
assign w177 = pi1337 & pi0261;
assign w178 = ~w2014 & w8536;
assign w179 = pi1690 & ~w15235;
assign w180 = w7703 & w11453;
assign w181 = ~pi3336 & w16922;
assign w182 = ~w10765 & ~w13452;
assign w183 = w13509 & w10752;
assign w184 = pi1711 & ~w619;
assign w185 = pi1787 & ~w8829;
assign w186 = pi2289 & ~w261;
assign w187 = pi2479 & ~w5274;
assign w188 = ~pi3145 & w15048;
assign w189 = w13509 & w8298;
assign w190 = (~pi1312 & w18092) | (~pi1312 & w8772) | (w18092 & w8772);
assign w191 = w13509 & w3226;
assign w192 = ~w12281 & ~pi0051;
assign w193 = pi1789 & ~w846;
assign w194 = ~w6030 & ~w11859;
assign w195 = ~w3686 & ~w7249;
assign w196 = pi2667 & ~w6463;
assign w197 = w13509 & w5615;
assign w198 = pi3159 & pi3207;
assign w199 = ~pi3158 & pi3207;
assign w200 = ~pi0309 & w18262;
assign w201 = w4807 & w18600;
assign w202 = ~w1368 & ~pi0455;
assign w203 = pi1964 & ~w14833;
assign w204 = ~pi2917 & ~w6045;
assign w205 = w7799 & w1219;
assign w206 = w16638 & w5156;
assign w207 = ~pi2701 & w15122;
assign w208 = ~w1277 & ~w13782;
assign w209 = w6649 & ~w15521;
assign w210 = ~w4353 & ~w10104;
assign w211 = ~w1962 & pi1119;
assign w212 = ~w7008 & ~w515;
assign w213 = pi2956 & ~w6045;
assign w214 = (~w6280 & ~w9420) | (~w6280 & w1288) | (~w9420 & w1288);
assign w215 = ~pi1316 & ~pi1301;
assign w216 = pi1854 & ~w653;
assign w217 = w11209 & ~w11029;
assign w218 = ~w6166 & ~w3281;
assign w219 = ~pi0883 & w1126;
assign w220 = ~pi2947 & ~w14417;
assign w221 = pi1758 & ~w2039;
assign w222 = pi1184 & ~w11450;
assign w223 = ~w7492 & ~w11977;
assign w224 = pi1376 & ~w11505;
assign w225 = pi3145 & w13786;
assign w226 = ~pi2922 & w11456;
assign w227 = ~w9440 & w12095;
assign w228 = ~w16575 & w6137;
assign w229 = (~pi0270 & ~w325) | (~pi0270 & w15998) | (~w325 & w15998);
assign w230 = (pi1127 & ~w13509) | (pi1127 & w8991) | (~w13509 & w8991);
assign w231 = w5437 & w13200;
assign w232 = ~w921 & ~w7061;
assign w233 = ~w1608 & ~w2573;
assign w234 = w13329 & w1858;
assign w235 = pi0111 & w9284;
assign w236 = w10335 & w9068;
assign w237 = ~pi3093 & w11406;
assign w238 = pi1442 & ~w13753;
assign w239 = ~w12996 & ~w10280;
assign w240 = pi2586 & ~w5274;
assign w241 = w7703 & w1677;
assign w242 = (pi1299 & ~w14158) | (pi1299 & w15694) | (~w14158 & w15694);
assign w243 = ~pi0836 & w93;
assign w244 = w13509 & w7169;
assign w245 = ~w3783 & ~w10240;
assign w246 = ~w18456 & ~w2073;
assign w247 = pi3021 & ~w3987;
assign w248 = pi2518 & ~w5274;
assign w249 = ~w18552 & ~w17270;
assign w250 = ~pi1268 & pi2959;
assign w251 = ~pi2680 & w13343;
assign w252 = w2341 & w4470;
assign w253 = ~pi2311 & w8617;
assign w254 = ~pi3057 & pi3207;
assign w255 = pi0250 & pi0300;
assign w256 = pi1643 & ~w13753;
assign w257 = ~pi3092 & w261;
assign w258 = ~pi3133 & w3805;
assign w259 = w4638 & w15845;
assign w260 = ~w12343 & ~w2358;
assign w261 = w6045 & w8396;
assign w262 = ~w2556 & ~w1214;
assign w263 = ~w8698 & ~w5269;
assign w264 = ~w14023 & ~w4433;
assign w265 = ~w4313 & ~w10776;
assign w266 = w922 & w10490;
assign w267 = w13509 & w13524;
assign w268 = pi2945 & w6045;
assign w269 = ~w5758 & ~w6927;
assign w270 = w6857 & w15458;
assign w271 = w8127 & w5302;
assign w272 = ~w2801 & ~w5403;
assign w273 = ~w1962 & pi1009;
assign w274 = ~w524 & ~w16129;
assign w275 = pi3157 & w9520;
assign w276 = w10189 & ~pi0472;
assign w277 = ~w7795 & ~w1361;
assign w278 = ~w10486 & ~w13416;
assign w279 = ~pi3061 & w11406;
assign w280 = pi2878 & ~w9504;
assign w281 = w10761 & w18292;
assign w282 = w11345 & w5908;
assign w283 = w4761 & w1567;
assign w284 = ~w7328 & w16393;
assign w285 = ~pi0716 & w3106;
assign w286 = ~pi0280 & w4058;
assign w287 = ~pi3043 & ~pi3207;
assign w288 = ~w12042 & ~w18125;
assign w289 = ~pi2168 & w11313;
assign w290 = ~w11974 & ~w10409;
assign w291 = ~pi0306 & pi1683;
assign w292 = pi1273 & pi1345;
assign w293 = (~pi1337 & w5855) | (~pi1337 & w14001) | (w5855 & w14001);
assign w294 = ~w7844 & pi0602;
assign w295 = ~w17157 & ~w18432;
assign w296 = w6857 & w16350;
assign w297 = ~w13250 & ~w18338;
assign w298 = ~pi2165 & w3019;
assign w299 = ~w18484 & w6275;
assign w300 = w2742 & ~w16002;
assign w301 = pi3171 & w3987;
assign w302 = ~w17534 & w12126;
assign w303 = w2764 & w14505;
assign w304 = ~pi3171 & w11132;
assign w305 = ~w2174 & ~w14402;
assign w306 = w12865 & w8631;
assign w307 = ~pi2390 & w17439;
assign w308 = ~w4820 & ~w4909;
assign w309 = (pi0777 & ~w13509) | (pi0777 & w96) | (~w13509 & w96);
assign w310 = ~w12662 & ~w17149;
assign w311 = w13509 & w14098;
assign w312 = ~w1051 & ~w1510;
assign w313 = w8337 & pi3306;
assign w314 = ~pi1828 & w7858;
assign w315 = pi0047 & w922;
assign w316 = ~w9196 & ~w2189;
assign w317 = pi1858 & ~w9021;
assign w318 = pi1394 & w13753;
assign w319 = pi1337 & ~pi0325;
assign w320 = pi1337 & pi0326;
assign w321 = w16278 & ~w2741;
assign w322 = ~w4743 & ~w11433;
assign w323 = ~pi3062 & w15235;
assign w324 = w2341 & ~w14978;
assign w325 = ~pi1858 & ~pi2911;
assign w326 = ~w6785 & pi0857;
assign w327 = w9440 & pi0186;
assign w328 = ~pi0264 & w2196;
assign w329 = pi1414 & ~w13753;
assign w330 = (pi0732 & ~w13509) | (pi0732 & w2634) | (~w13509 & w2634);
assign w331 = ~w15808 & ~pi0971;
assign w332 = ~w10558 & w11371;
assign w333 = ~pi0297 & w2196;
assign w334 = w13509 & w15384;
assign w335 = ~pi0646 & w3791;
assign w336 = ~pi0849 & w93;
assign w337 = pi0149 & ~w15479;
assign w338 = w9440 & pi0142;
assign w339 = ~w15292 & ~pi1240;
assign w340 = ~w1830 & ~w14535;
assign w341 = ~w9717 & ~w3488;
assign w342 = ~pi1375 & w5043;
assign w343 = ~w11842 & ~w17655;
assign w344 = (pi0547 & ~w13509) | (pi0547 & w13350) | (~w13509 & w13350);
assign w345 = pi1510 & ~w16922;
assign w346 = ~w3000 & ~pi2793;
assign w347 = pi3046 & ~pi3146;
assign w348 = ~w5422 & ~w5911;
assign w349 = ~w5968 & w13368;
assign w350 = w12040 & ~w1340;
assign w351 = ~pi3318 & w9781;
assign w352 = w6857 & w3364;
assign w353 = pi0135 & w5274;
assign w354 = w4019 & w8995;
assign w355 = ~pi3089 & w261;
assign w356 = ~w15145 & ~w13739;
assign w357 = w3243 & pi0311;
assign w358 = pi1467 & w13753;
assign w359 = ~w16352 & ~w16552;
assign w360 = ~w4943 & ~w5661;
assign w361 = ~w6061 & w6161;
assign w362 = w4584 & ~w8810;
assign w363 = ~w13987 & ~w6957;
assign w364 = ~w4363 & w17380;
assign w365 = pi3166 & w11272;
assign w366 = ~w1791 & w4762;
assign w367 = w16506 & ~w6680;
assign w368 = pi1395 & pi3360;
assign w369 = ~w3394 & w2845;
assign w370 = ~w1003 & ~w8469;
assign w371 = pi2313 & ~w4420;
assign w372 = pi1155 & w9420;
assign w373 = pi2510 & ~w226;
assign w374 = ~w1791 & w8819;
assign w375 = ~pi3170 & w3805;
assign w376 = pi2798 & ~w6463;
assign w377 = ~pi2973 & ~w8569;
assign w378 = w15122 & ~pi2709;
assign w379 = ~w6508 & w15029;
assign w380 = w11320 & w14069;
assign w381 = w16506 & ~w14465;
assign w382 = ~pi3094 & w15235;
assign w383 = ~w751 & w3462;
assign w384 = w15612 & w10574;
assign w385 = ~w6195 & w3687;
assign w386 = w968 & ~pi0280;
assign w387 = ~pi0657 & w12197;
assign w388 = (pi0595 & ~w13509) | (pi0595 & w1223) | (~w13509 & w1223);
assign w389 = pi1443 & ~w13753;
assign w390 = w13509 & w5498;
assign w391 = ~w9497 & w9938;
assign w392 = ~w11055 & ~w15666;
assign w393 = (~pi0486 & w17577) | (~pi0486 & w11910) | (w17577 & w11910);
assign w394 = pi0010 & ~w3748;
assign w395 = ~w6945 & ~w7174;
assign w396 = ~pi0578 & w795;
assign w397 = ~pi0413 & w17173;
assign w398 = pi0414 & w17173;
assign w399 = w6785 & ~w6680;
assign w400 = pi2754 & ~w226;
assign w401 = ~pi0517 & w14641;
assign w402 = ~pi1232 & ~pi3201;
assign w403 = ~w13850 & ~w4455;
assign w404 = w18508 & w5694;
assign w405 = pi3012 & ~w3987;
assign w406 = ~w15485 & ~w13743;
assign w407 = ~w2915 & ~w9075;
assign w408 = ~w17665 & ~w4398;
assign w409 = ~pi1995 & w3019;
assign w410 = w11813 & w4366;
assign w411 = pi0494 & pi1158;
assign w412 = w14341 & w4841;
assign w413 = ~pi3059 & w15235;
assign w414 = ~pi3029 & pi3151;
assign w415 = w13231 & ~w15173;
assign w416 = ~w94 & ~w8672;
assign w417 = ~w12601 & ~w12741;
assign w418 = ~w14574 & ~w18367;
assign w419 = ~w5473 & ~w8180;
assign w420 = ~w3976 & ~w17644;
assign w421 = pi2046 & ~w10158;
assign w422 = ~w7779 & ~w17398;
assign w423 = pi3160 & ~pi3495;
assign w424 = ~w3377 & ~w5710;
assign w425 = ~w7074 & w9241;
assign w426 = ~w17791 & ~w17054;
assign w427 = ~pi1140 & ~pi2941;
assign w428 = ~pi3020 & pi3112;
assign w429 = ~w13964 & ~w6816;
assign w430 = ~w13231 & pi1092;
assign w431 = (~pi0976 & ~w13509) | (~pi0976 & w7380) | (~w13509 & w7380);
assign w432 = w9322 & w854;
assign w433 = ~w6785 & pi0852;
assign w434 = ~w5962 & ~w8999;
assign w435 = ~w15585 & ~w14775;
assign w436 = ~pi0637 & w3791;
assign w437 = ~w3910 & w15740;
assign w438 = ~w14560 & pi0213;
assign w439 = w6649 & ~w5503;
assign w440 = (pi0315 & w3055) | (pi0315 & w5035) | (w3055 & w5035);
assign w441 = ~pi3096 & w9504;
assign w442 = ~w17665 & ~w5641;
assign w443 = ~w17665 & ~w17508;
assign w444 = ~pi0803 & w1147;
assign w445 = w13509 & w7527;
assign w446 = ~pi1761 & ~w3689;
assign w447 = pi1811 & ~pi1969;
assign w448 = ~pi0844 & w93;
assign w449 = pi1466 & w13753;
assign w450 = ~pi0806 & w1147;
assign w451 = w13825 & w10184;
assign w452 = w13509 & w16072;
assign w453 = pi1570 & ~w13753;
assign w454 = w13509 & w18085;
assign w455 = ~w14926 & ~w7562;
assign w456 = ~w3367 & w5728;
assign w457 = ~pi3072 & pi3171;
assign w458 = ~w2014 & ~w709;
assign w459 = ~w11891 & ~w13864;
assign w460 = ~pi3315 & w6448;
assign w461 = w1890 & w13945;
assign w462 = w9440 & pi0174;
assign w463 = w7799 & w2832;
assign w464 = ~pi3050 & w15235;
assign w465 = ~pi0893 & w1126;
assign w466 = pi1458 & ~w7090;
assign w467 = w14560 & pi0363;
assign w468 = ~pi2663 & w17213;
assign w469 = ~pi0783 & w543;
assign w470 = ~w4132 & ~w18227;
assign w471 = ~pi0829 & w93;
assign w472 = w7703 & w11364;
assign w473 = pi2862 & w16699;
assign w474 = ~w2464 & ~w18291;
assign w475 = ~w12806 & ~w9100;
assign w476 = (pi0755 & ~w13509) | (pi0755 & w7026) | (~w13509 & w7026);
assign w477 = ~w12568 & ~w4924;
assign w478 = ~pi0858 & w15707;
assign w479 = ~pi1014 & w12197;
assign w480 = pi3135 & w10992;
assign w481 = pi3164 & w15767;
assign w482 = w6857 & w12244;
assign w483 = ~w1368 & ~pi0458;
assign w484 = w4478 & pi0490;
assign w485 = w17495 & ~pi1315;
assign w486 = w968 & ~pi0264;
assign w487 = ~pi2967 & w5517;
assign w488 = ~w7306 & w9073;
assign w489 = ~w15071 & ~w12846;
assign w490 = ~w3505 & ~w448;
assign w491 = w13231 & ~w14597;
assign w492 = ~w9402 & w155;
assign w493 = w12040 & ~w17210;
assign w494 = ~pi2683 & w13343;
assign w495 = ~pi1959 & w11688;
assign w496 = w968 & ~pi0296;
assign w497 = w2341 & ~w9852;
assign w498 = ~pi3349 & w16922;
assign w499 = ~w12040 & pi1018;
assign w500 = pi1810 & ~w3258;
assign w501 = w9139 & w2149;
assign w502 = pi2673 & ~w226;
assign w503 = ~w9191 & ~w6686;
assign w504 = (pi3001 & ~w735) | (pi3001 & w13887) | (~w735 & w13887);
assign w505 = w13509 & w1496;
assign w506 = ~w3625 & ~w10512;
assign w507 = pi0016 & ~w14148;
assign w508 = ~pi3093 & w261;
assign w509 = w10242 & w12694;
assign w510 = (w5156 & ~w3021) | (w5156 & w206) | (~w3021 & w206);
assign w511 = ~w10628 & ~w9189;
assign w512 = w12998 & w15830;
assign w513 = w14228 & w1217;
assign w514 = pi1143 & w9420;
assign w515 = ~pi0945 & w3791;
assign w516 = ~w377 & w9882;
assign w517 = pi1888 & ~w15036;
assign w518 = ~pi1222 & ~pi3204;
assign w519 = w10912 & w7576;
assign w520 = ~w16506 & pi1133;
assign w521 = ~w12726 & ~w18505;
assign w522 = ~w15356 & ~w17200;
assign w523 = ~pi2028 & w7455;
assign w524 = ~pi3146 & w17669;
assign w525 = w3544 & pi0511;
assign w526 = ~w1319 & ~w6267;
assign w527 = ~w18315 & ~w402;
assign w528 = w13321 & ~w853;
assign w529 = ~w5560 & w202;
assign w530 = ~pi3032 & pi3135;
assign w531 = ~w12460 & w4434;
assign w532 = ~w3991 & ~w8405;
assign w533 = ~pi2921 & pi3199;
assign w534 = ~w17378 & w18569;
assign w535 = w12691 & w12929;
assign w536 = ~pi3349 & w18259;
assign w537 = w13509 & w17081;
assign w538 = ~w9317 & ~w12538;
assign w539 = w6575 & w3381;
assign w540 = w8514 & w3060;
assign w541 = pi1429 & ~w13753;
assign w542 = (~w4921 & ~w5566) | (~w4921 & w9726) | (~w5566 & w9726);
assign w543 = w134 & w12825;
assign w544 = (pi1809 & w7215) | (pi1809 & w9187) | (w7215 & w9187);
assign w545 = ~pi1973 & ~pi3117;
assign w546 = pi3155 & ~pi3166;
assign w547 = pi3116 & ~w16502;
assign w548 = w8040 & ~w4308;
assign w549 = (pi0484 & w1688) | (pi0484 & w15895) | (w1688 & w15895);
assign w550 = w9255 & w1396;
assign w551 = w11222 & w6740;
assign w552 = ~w16506 & pi1268;
assign w553 = pi1304 & ~pi1330;
assign w554 = ~pi0431 & w17173;
assign w555 = pi0432 & w17173;
assign w556 = ~w13543 & ~w14258;
assign w557 = w17562 & pi1846;
assign w558 = ~pi2187 & w2151;
assign w559 = pi0056 & w922;
assign w560 = w0 & w5983;
assign w561 = ~w4775 & w13421;
assign w562 = ~w387 & ~w8760;
assign w563 = ~w5686 & ~w14840;
assign w564 = ~pi2105 & w12724;
assign w565 = pi3136 & w4256;
assign w566 = ~pi2312 & w16041;
assign w567 = ~pi3293 & w6072;
assign w568 = ~pi2935 & pi3205;
assign w569 = ~pi0652 & w3791;
assign w570 = ~pi3059 & w16815;
assign w571 = ~w5359 & w7547;
assign w572 = ~w9462 & pi0359;
assign w573 = ~w3321 & ~w15584;
assign w574 = w17287 & w2410;
assign w575 = pi2827 & ~w3555;
assign w576 = (pi0872 & ~w13509) | (pi0872 & w2348) | (~w13509 & w2348);
assign w577 = ~w2921 & w15265;
assign w578 = pi1626 & ~w6448;
assign w579 = ~pi2093 & w12724;
assign w580 = w12040 & ~w6033;
assign w581 = (pi1183 & ~w5437) | (pi1183 & w10035) | (~w5437 & w10035);
assign w582 = pi1743 & w1924;
assign w583 = ~pi2051 & w13204;
assign w584 = ~w15808 & pi1031;
assign w585 = ~w3123 & ~w12615;
assign w586 = w934 & pi0410;
assign w587 = ~w3776 & ~w8373;
assign w588 = ~pi3133 & w4310;
assign w589 = ~w6627 & ~w8264;
assign w590 = w13509 & w3346;
assign w591 = ~w1962 & pi0644;
assign w592 = w1254 & w5046;
assign w593 = ~pi0491 & ~pi1138;
assign w594 = pi0492 & pi1139;
assign w595 = ~pi3163 & w13570;
assign w596 = ~w7736 & ~w1517;
assign w597 = ~w12460 & w1893;
assign w598 = w1451 & w17553;
assign w599 = ~w1368 & ~pi0464;
assign w600 = pi1909 & ~w14524;
assign w601 = pi3146 & w3987;
assign w602 = ~w5873 & ~w17476;
assign w603 = w16807 & w2601;
assign w604 = ~w2077 & w6250;
assign w605 = w16893 & w3858;
assign w606 = ~w10113 & w5138;
assign w607 = ~w11414 & ~w14779;
assign w608 = ~pi3158 & w11132;
assign w609 = pi2969 & w8789;
assign w610 = ~pi1696 & ~w17534;
assign w611 = ~pi3099 & w261;
assign w612 = w137 & ~w12166;
assign w613 = ~w5618 & ~w8965;
assign w614 = ~pi3136 & ~w4020;
assign w615 = ~w13849 & ~w15312;
assign w616 = ~w10510 & ~w14117;
assign w617 = ~w13362 & ~w11471;
assign w618 = ~pi0515 & ~pi1185;
assign w619 = ~w3054 & w11545;
assign w620 = ~w992 & ~w11554;
assign w621 = (~pi3369 & w18594) | (~pi3369 & w14810) | (w18594 & w14810);
assign w622 = ~pi3107 & w16502;
assign w623 = w15842 & pi2737;
assign w624 = ~w6453 & ~w17790;
assign w625 = w9543 & w7896;
assign w626 = (pi0608 & ~w13509) | (pi0608 & w50) | (~w13509 & w50);
assign w627 = ~w18459 & ~w13633;
assign w628 = pi1362 & w9653;
assign w629 = ~w2341 & pi0833;
assign w630 = pi3162 & w14951;
assign w631 = (pi0891 & ~w13509) | (pi0891 & w10204) | (~w13509 & w10204);
assign w632 = pi1309 & pi3214;
assign w633 = pi2614 & ~w261;
assign w634 = pi3160 & ~w9243;
assign w635 = ~w11461 & ~w14483;
assign w636 = (~pi0952 & ~w13509) | (~pi0952 & w8144) | (~w13509 & w8144);
assign w637 = pi1374 & ~pi3123;
assign w638 = ~w5147 & ~w5902;
assign w639 = w13509 & w1644;
assign w640 = ~pi1089 & w543;
assign w641 = ~w13098 & ~w17365;
assign w642 = ~pi1990 & w3019;
assign w643 = ~pi2925 & w6359;
assign w644 = ~pi1058 & w6200;
assign w645 = ~w16443 & w11042;
assign w646 = ~pi2550 & w5453;
assign w647 = ~w10371 & ~w13836;
assign w648 = ~pi0508 & ~pi1146;
assign w649 = pi1649 & ~w13753;
assign w650 = w7177 & w15703;
assign w651 = w8658 & pi1779;
assign w652 = pi0151 & ~w7867;
assign w653 = w1611 & w3550;
assign w654 = ~w16752 & ~w14431;
assign w655 = ~w4169 & ~w15443;
assign w656 = pi3082 & w6463;
assign w657 = w10574 & w15213;
assign w658 = pi2157 & ~w3555;
assign w659 = ~w14316 & ~w10953;
assign w660 = ~w10955 & ~w17479;
assign w661 = (w5517 & w4885) | (w5517 & w11619) | (w4885 & w11619);
assign w662 = (pi0851 & ~w13509) | (pi0851 & w1585) | (~w13509 & w1585);
assign w663 = ~w12321 & ~w16195;
assign w664 = ~w1710 & ~w14867;
assign w665 = ~pi0843 & w93;
assign w666 = ~w2182 & ~w203;
assign w667 = pi1407 & ~w1598;
assign w668 = ~w10445 & ~w15985;
assign w669 = pi2892 & ~w3555;
assign w670 = ~w2341 & pi1068;
assign w671 = ~w13361 & ~w957;
assign w672 = pi3079 & ~w3987;
assign w673 = pi1774 & ~pi3141;
assign w674 = ~pi0591 & w795;
assign w675 = ~w6195 & w146;
assign w676 = ~pi2385 & w16041;
assign w677 = w13509 & w3680;
assign w678 = pi1159 & ~pi1160;
assign w679 = pi3166 & w7946;
assign w680 = ~pi1088 & w795;
assign w681 = ~w15551 & ~w3284;
assign w682 = ~pi3160 & ~pi3171;
assign w683 = ~pi2972 & w10058;
assign w684 = w13509 & w14336;
assign w685 = ~w4259 & ~w16485;
assign w686 = ~w4769 & ~w12792;
assign w687 = w12205 & w9385;
assign w688 = w17562 & pi2559;
assign w689 = pi2045 & ~w10158;
assign w690 = w13509 & w4339;
assign w691 = w8658 & pi1789;
assign w692 = w657 & w17591;
assign w693 = w15907 & w17130;
assign w694 = ~w15808 & pi0751;
assign w695 = ~w7072 & ~w13498;
assign w696 = ~w4164 & ~w1022;
assign w697 = ~w15327 & ~pi0299;
assign w698 = w15727 & w8554;
assign w699 = w7844 & w15609;
assign w700 = w14030 & w13971;
assign w701 = ~w7033 & w932;
assign w702 = (w14755 & ~w11247) | (w14755 & w2501) | (~w11247 & w2501);
assign w703 = ~w1561 & w4222;
assign w704 = ~w4104 & ~w8906;
assign w705 = ~w18017 & ~w1246;
assign w706 = ~w1062 & ~w13632;
assign w707 = ~pi3326 & w16922;
assign w708 = pi0077 & pi0126;
assign w709 = w9323 & w7277;
assign w710 = ~w9691 & ~w15620;
assign w711 = (pi2920 & ~w384) | (pi2920 & w5287) | (~w384 & w5287);
assign w712 = w8566 & w18431;
assign w713 = ~w576 & ~w8542;
assign w714 = pi2730 & ~w3555;
assign w715 = w8611 & w12009;
assign w716 = w11345 & w8444;
assign w717 = ~pi3090 & w9504;
assign w718 = ~w2757 & ~w17562;
assign w719 = ~w280 & ~w441;
assign w720 = pi1632 & ~w13753;
assign w721 = ~w3021 & ~w1975;
assign w722 = ~w5152 & ~w9055;
assign w723 = ~pi3090 & w261;
assign w724 = pi2780 & ~w16815;
assign w725 = ~pi0717 & w3106;
assign w726 = w15951 & pi0252;
assign w727 = ~w10852 & w7290;
assign w728 = w6689 & w15289;
assign w729 = w8337 & pi3357;
assign w730 = ~w14733 & ~w60;
assign w731 = ~w595 & ~w4481;
assign w732 = ~w11297 & w16558;
assign w733 = (pi0923 & ~w13509) | (pi0923 & w14024) | (~w13509 & w14024);
assign w734 = ~w17623 & ~w12977;
assign w735 = ~pi2920 & ~pi2966;
assign w736 = ~w1052 & ~w4387;
assign w737 = ~w18325 & w14735;
assign w738 = ~pi3355 & w9781;
assign w739 = ~w14165 & ~w10674;
assign w740 = (pi1297 & ~w17477) | (pi1297 & w13901) | (~w17477 & w13901);
assign w741 = ~w5745 & w8722;
assign w742 = ~pi0781 & w543;
assign w743 = w13509 & w16663;
assign w744 = ~pi3158 & w3982;
assign w745 = (pi0644 & ~w13509) | (pi0644 & w591) | (~w13509 & w591);
assign w746 = w16888 & w11061;
assign w747 = ~pi3170 & w17387;
assign w748 = pi0005 & ~w14148;
assign w749 = ~pi2291 & w8617;
assign w750 = pi1186 & w9420;
assign w751 = ~pi1185 & w9420;
assign w752 = (~pi0499 & w17577) | (~pi0499 & w16097) | (w17577 & w16097);
assign w753 = ~w16951 & ~w1351;
assign w754 = pi2960 & pi2465;
assign w755 = ~pi0846 & w93;
assign w756 = (pi0946 & ~w13509) | (pi0946 & w7966) | (~w13509 & w7966);
assign w757 = ~w12336 & w11946;
assign w758 = ~w7479 & ~w5753;
assign w759 = pi0045 & w9240;
assign w760 = ~w11722 & ~w5925;
assign w761 = w16342 & ~w18379;
assign w762 = pi2966 & pi2588;
assign w763 = ~pi0151 & w7867;
assign w764 = ~w2829 & w7004;
assign w765 = w15808 & ~w4043;
assign w766 = ~w10901 & ~w10085;
assign w767 = ~w4177 & ~w12604;
assign w768 = w13509 & w2739;
assign w769 = w4420 & w17115;
assign w770 = pi1448 & ~w13753;
assign w771 = ~w11654 & w4410;
assign w772 = ~w14332 & ~w6874;
assign w773 = ~w10290 & ~pi1179;
assign w774 = pi1264 & ~pi2952;
assign w775 = ~pi0149 & w15479;
assign w776 = pi1293 & pi1345;
assign w777 = ~w16093 & ~w17602;
assign w778 = (~w603 & w17577) | (~w603 & w5771) | (w17577 & w5771);
assign w779 = ~pi0689 & w9110;
assign w780 = pi3080 & ~pi3141;
assign w781 = pi0075 & ~w14148;
assign w782 = ~w18404 & w12443;
assign w783 = ~pi2211 & w5075;
assign w784 = w14619 & w8069;
assign w785 = ~w13620 & w10973;
assign w786 = ~w9819 & ~w9563;
assign w787 = pi2465 & pi3362;
assign w788 = ~w3306 & ~w282;
assign w789 = ~w14228 & pi0617;
assign w790 = (pi1156 & ~w5437) | (pi1156 & w7198) | (~w5437 & w7198);
assign w791 = w15363 & w1207;
assign w792 = w11345 & w16921;
assign w793 = ~w7722 & ~w3784;
assign w794 = ~w631 & ~w15631;
assign w795 = ~w3381 & w10724;
assign w796 = ~pi0805 & w1147;
assign w797 = pi2120 & ~w412;
assign w798 = pi0298 & pi0299;
assign w799 = ~w15726 & ~w8420;
assign w800 = ~pi0505 & ~pi1192;
assign w801 = ~w17665 & ~w14887;
assign w802 = w13781 & w8540;
assign w803 = pi1902 & w9021;
assign w804 = ~w15402 & ~w15325;
assign w805 = ~w15852 & ~w12819;
assign w806 = pi1530 & w13753;
assign w807 = (pi0986 & ~w13509) | (pi0986 & w3894) | (~w13509 & w3894);
assign w808 = ~w6288 & w364;
assign w809 = ~w16278 & pi0713;
assign w810 = ~pi1878 & ~pi3512;
assign w811 = ~w8978 & ~w3666;
assign w812 = ~pi3091 & w16815;
assign w813 = ~w2735 & ~w2596;
assign w814 = ~w16712 & w5528;
assign w815 = ~pi0807 & w1147;
assign w816 = (pi0912 & ~w13509) | (pi0912 & w17471) | (~w13509 & w17471);
assign w817 = w10676 & ~w504;
assign w818 = ~pi3131 & w8515;
assign w819 = ~w9155 & w8646;
assign w820 = ~w16733 & w17878;
assign w821 = pi1419 & ~w13753;
assign w822 = w6697 & ~w7707;
assign w823 = ~pi0488 & ~pi1345;
assign w824 = ~w1863 & ~w7094;
assign w825 = pi0201 & w5274;
assign w826 = pi0018 & ~w3748;
assign w827 = ~w15555 & ~w8426;
assign w828 = ~w7750 & ~w390;
assign w829 = pi3150 & w5457;
assign w830 = pi1461 & w13753;
assign w831 = pi3169 & w7946;
assign w832 = ~w8324 & ~w2426;
assign w833 = w8268 & w8493;
assign w834 = w709 & pi1891;
assign w835 = ~pi3139 & w3982;
assign w836 = pi2460 & ~w11671;
assign w837 = pi2578 & ~w5274;
assign w838 = ~pi3318 & w17935;
assign w839 = pi1548 & ~w17935;
assign w840 = pi0444 & ~pi2911;
assign w841 = ~w15122 & ~pi1903;
assign w842 = ~w13733 & ~w13896;
assign w843 = pi2076 & ~w17683;
assign w844 = w13509 & w5471;
assign w845 = ~pi2347 & w12941;
assign w846 = ~pi1767 & ~pi3154;
assign w847 = w7621 & ~w7084;
assign w848 = ~w4153 & ~w13618;
assign w849 = ~pi3157 & w15048;
assign w850 = ~w15201 & ~w10565;
assign w851 = ~w1663 & ~w4111;
assign w852 = w16836 & pi0058;
assign w853 = pi2528 & w15191;
assign w854 = ~w950 & ~w13186;
assign w855 = ~w2771 & ~w380;
assign w856 = ~w14586 & ~w9663;
assign w857 = pi2061 & ~w4508;
assign w858 = ~w18155 & ~w7837;
assign w859 = pi1768 & ~pi3151;
assign w860 = ~w9462 & w2880;
assign w861 = ~w5928 & ~w14471;
assign w862 = ~pi3095 & w15235;
assign w863 = ~w15627 & ~w16323;
assign w864 = ~pi2472 & w5384;
assign w865 = ~pi3164 & w13730;
assign w866 = ~pi2987 & w6463;
assign w867 = ~w14228 & pi1007;
assign w868 = ~pi2410 & w5384;
assign w869 = pi2663 & ~w15235;
assign w870 = pi2955 & ~w13367;
assign w871 = w8789 & ~w16575;
assign w872 = pi1326 & pi1345;
assign w873 = ~w6323 & ~w17846;
assign w874 = ~w5167 & ~w17353;
assign w875 = ~w14648 & ~pi2694;
assign w876 = w13569 & w9941;
assign w877 = pi2831 & ~w261;
assign w878 = ~pi3313 & w17935;
assign w879 = w7703 & w9014;
assign w880 = w6179 & w4029;
assign w881 = ~w16990 & ~w13571;
assign w882 = w9108 & ~pi0444;
assign w883 = (pi0665 & ~w13509) | (pi0665 & w5816) | (~w13509 & w5816);
assign w884 = ~w15089 & ~w12110;
assign w885 = pi1373 & ~w7854;
assign w886 = ~w11110 & ~w15552;
assign w887 = ~pi1050 & w15707;
assign w888 = (pi1869 & w2014) | (pi1869 & w1287) | (w2014 & w1287);
assign w889 = pi1365 & ~w1128;
assign w890 = ~pi0082 & pi3149;
assign w891 = ~pi0483 & pi3405;
assign w892 = ~w4615 & ~w1960;
assign w893 = w14560 & pi0341;
assign w894 = w10818 & ~w12251;
assign w895 = ~w10072 & ~w11748;
assign w896 = ~w16506 & pi1263;
assign w897 = w13509 & w13124;
assign w898 = pi2309 & ~w4420;
assign w899 = ~pi3171 & w14753;
assign w900 = ~w17577 & w11161;
assign w901 = ~w17665 & ~w4649;
assign w902 = ~w5390 & w6971;
assign w903 = ~pi1827 & ~w6872;
assign w904 = ~w6745 & ~w17214;
assign w905 = ~w7844 & pi0601;
assign w906 = w14228 & ~w15296;
assign w907 = ~w11059 & w9838;
assign w908 = ~w9899 & w6890;
assign w909 = ~w18103 & ~w11549;
assign w910 = pi1877 & ~w7858;
assign w911 = ~pi0653 & w3791;
assign w912 = pi2074 & ~w17683;
assign w913 = ~pi3154 & w13730;
assign w914 = ~w5855 & w4931;
assign w915 = ~pi2145 & w13065;
assign w916 = ~pi2386 & w16041;
assign w917 = (pi1780 & w7215) | (pi1780 & w1645) | (w7215 & w1645);
assign w918 = w8356 & pi0270;
assign w919 = ~pi1102 & w17899;
assign w920 = ~w16721 & w7399;
assign w921 = pi1525 & ~w14918;
assign w922 = (~w9284 & ~w5517) | (~w9284 & w2632) | (~w5517 & w2632);
assign w923 = ~pi0723 & w17899;
assign w924 = w14812 & w8887;
assign w925 = ~pi1985 & ~w15450;
assign w926 = pi0313 & ~pi3225;
assign w927 = w2725 & ~w14465;
assign w928 = ~w601 & ~w3781;
assign w929 = w16575 & w12278;
assign w930 = ~w15670 & ~w12640;
assign w931 = ~pi3157 & w1843;
assign w932 = w9323 & ~w10384;
assign w933 = w7703 & w1023;
assign w934 = ~w968 & ~pi2486;
assign w935 = ~w5971 & ~w10547;
assign w936 = w126 & pi0040;
assign w937 = pi1337 & pi0254;
assign w938 = ~w5573 & ~w5076;
assign w939 = ~w12744 & ~w9442;
assign w940 = ~w15808 & pi0757;
assign w941 = w9440 & pi0147;
assign w942 = ~w4246 & ~w9430;
assign w943 = w17646 & w614;
assign w944 = ~w10258 & ~w4661;
assign w945 = (~pi1233 & ~w11505) | (~pi1233 & w13241) | (~w11505 & w13241);
assign w946 = ~pi3290 & w9781;
assign w947 = w16506 & ~w7707;
assign w948 = pi2400 & ~w17683;
assign w949 = ~w14648 & ~pi2781;
assign w950 = ~pi2212 & w11313;
assign w951 = ~w5453 & ~pi1775;
assign w952 = (pi1038 & ~w13509) | (pi1038 & w14758) | (~w13509 & w14758);
assign w953 = pi1644 & ~w6448;
assign w954 = ~w3055 & w8332;
assign w955 = ~w1949 & w4406;
assign w956 = ~pi2415 & w5075;
assign w957 = ~w11655 & w1731;
assign w958 = w13509 & w14367;
assign w959 = ~pi2184 & w5384;
assign w960 = pi2948 & pi2985;
assign w961 = (~pi0263 & ~w325) | (~pi0263 & w16714) | (~w325 & w16714);
assign w962 = w12460 & w17293;
assign w963 = (~w4359 & ~w5517) | (~w4359 & w8762) | (~w5517 & w8762);
assign w964 = (pi1018 & ~w13509) | (pi1018 & w499) | (~w13509 & w499);
assign w965 = ~pi0790 & w543;
assign w966 = ~w13154 & ~w23;
assign w967 = w11383 & w8045;
assign w968 = pi1692 & pi3179;
assign w969 = ~w18566 & ~w4987;
assign w970 = ~w3668 & ~w10401;
assign w971 = pi1522 & w13753;
assign w972 = w2341 & ~w3430;
assign w973 = ~pi2994 & w16922;
assign w974 = ~w2720 & ~w17330;
assign w975 = pi0250 & w5274;
assign w976 = pi0267 & pi0312;
assign w977 = w14109 & pi0439;
assign w978 = (w8789 & w4903) | (w8789 & w609) | (w4903 & w609);
assign w979 = w1009 & w16336;
assign w980 = w10818 & ~w14288;
assign w981 = pi1377 & ~w10894;
assign w982 = pi2397 & ~w10299;
assign w983 = ~w4343 & ~w1762;
assign w984 = ~w12215 & ~w16486;
assign w985 = ~w2076 & ~w3169;
assign w986 = ~w13424 & ~w2616;
assign w987 = ~pi0327 & w2196;
assign w988 = w9600 & w1392;
assign w989 = ~w4094 & ~w12659;
assign w990 = ~pi1680 & ~w7177;
assign w991 = (pi1045 & ~w13509) | (pi1045 & w16203) | (~w13509 & w16203);
assign w992 = pi3102 & ~w16502;
assign w993 = ~pi3145 & w8515;
assign w994 = pi3120 & ~w16401;
assign w995 = ~w1791 & w9222;
assign w996 = ~pi3128 & w226;
assign w997 = pi1983 & ~w4254;
assign w998 = (w2460 & ~w11232) | (w2460 & w14569) | (~w11232 & w14569);
assign w999 = w16278 & ~w6922;
assign w1000 = ~w7077 & pi0819;
assign w1001 = ~w12460 & w5681;
assign w1002 = pi1737 & w1924;
assign w1003 = pi2971 & ~w16502;
assign w1004 = ~w15536 & ~w5834;
assign w1005 = ~pi1710 & pi3143;
assign w1006 = w17248 & ~w6680;
assign w1007 = ~w17577 & w13289;
assign w1008 = ~pi1069 & w12825;
assign w1009 = ~w4641 & ~w15777;
assign w1010 = pi0067 & ~w14148;
assign w1011 = pi2945 & ~w6045;
assign w1012 = ~w968 & ~w1117;
assign w1013 = ~w6414 & w7268;
assign w1014 = ~w14262 & ~w7441;
assign w1015 = ~pi3062 & w16815;
assign w1016 = w13509 & w5321;
assign w1017 = ~w12198 & ~w7810;
assign w1018 = pi1460 & w13753;
assign w1019 = pi2854 & w15191;
assign w1020 = ~w5 & ~w9168;
assign w1021 = pi1908 & ~w3223;
assign w1022 = pi3069 & ~pi3168;
assign w1023 = w15122 & ~pi2905;
assign w1024 = ~pi2976 & w16815;
assign w1025 = pi2316 & ~w9414;
assign w1026 = ~w13480 & ~w16834;
assign w1027 = ~w487 & ~w18503;
assign w1028 = w8020 & w9253;
assign w1029 = w5985 & w18108;
assign w1030 = ~w17577 & w4936;
assign w1031 = pi2104 & ~w4420;
assign w1032 = ~w14941 & ~w18035;
assign w1033 = ~w18050 & ~w7214;
assign w1034 = ~w15542 & w2460;
assign w1035 = w5437 & w947;
assign w1036 = ~w4691 & ~w1474;
assign w1037 = pi3155 & w14951;
assign w1038 = pi1890 & ~w6463;
assign w1039 = pi2266 & ~w11671;
assign w1040 = ~w11652 & w6688;
assign w1041 = w12542 & w10716;
assign w1042 = pi2742 & ~w6463;
assign w1043 = ~pi0330 & w4058;
assign w1044 = ~w7921 & ~w15751;
assign w1045 = w8660 & w16447;
assign w1046 = ~w12588 & ~w144;
assign w1047 = (pi1142 & ~w5437) | (pi1142 & w13567) | (~w5437 & w13567);
assign w1048 = pi1335 & ~pi2553;
assign w1049 = ~pi3311 & w17935;
assign w1050 = ~pi1264 & pi2952;
assign w1051 = pi3135 & ~w15132;
assign w1052 = ~pi3131 & w15048;
assign w1053 = w15122 & ~pi1857;
assign w1054 = ~pi1159 & pi1160;
assign w1055 = ~w7077 & pi1070;
assign w1056 = ~w16575 & w4966;
assign w1057 = pi1551 & ~w17935;
assign w1058 = w4067 & w15389;
assign w1059 = ~w11536 & ~w5514;
assign w1060 = w6697 & ~w10235;
assign w1061 = w17770 & w13893;
assign w1062 = ~pi0756 & w17490;
assign w1063 = w8719 & w17849;
assign w1064 = pi1424 & ~w13753;
assign w1065 = w5437 & w14466;
assign w1066 = w10201 & w12639;
assign w1067 = ~w9614 & ~w4018;
assign w1068 = ~w8415 & ~w3110;
assign w1069 = ~pi1377 & ~pi2920;
assign w1070 = w12040 & ~w10235;
assign w1071 = w13509 & w3072;
assign w1072 = w14648 & ~pi2607;
assign w1073 = ~w7923 & ~w1397;
assign w1074 = ~w1449 & ~w8093;
assign w1075 = ~w16506 & pi1149;
assign w1076 = ~w2787 & ~w878;
assign w1077 = pi1598 & ~w16922;
assign w1078 = ~pi3158 & pi0133;
assign w1079 = ~w2725 & pi1040;
assign w1080 = ~w6794 & ~w6630;
assign w1081 = w14228 & ~w1340;
assign w1082 = (pi0800 & ~w13509) | (pi0800 & w12756) | (~w13509 & w12756);
assign w1083 = pi1587 & ~w13753;
assign w1084 = pi3141 & w8829;
assign w1085 = ~w1791 & w13912;
assign w1086 = ~w8055 & w1026;
assign w1087 = w13509 & w4876;
assign w1088 = ~w8015 & ~w18441;
assign w1089 = ~w12826 & ~w225;
assign w1090 = w10719 & ~w6918;
assign w1091 = ~w9549 & ~w611;
assign w1092 = w5236 & w12306;
assign w1093 = w5968 & pi1676;
assign w1094 = ~pi0671 & w12197;
assign w1095 = w6857 & w13194;
assign w1096 = ~w3174 & ~w14510;
assign w1097 = pi3182 & pi3320;
assign w1098 = ~w14228 & pi0622;
assign w1099 = pi1415 & ~w6072;
assign w1100 = w15188 & w12814;
assign w1101 = ~w15143 & ~w12499;
assign w1102 = ~w15667 & ~w11417;
assign w1103 = ~pi2967 & ~pi3030;
assign w1104 = ~pi2967 & pi3031;
assign w1105 = pi2951 & ~pi3199;
assign w1106 = ~w3868 & ~w6177;
assign w1107 = ~w15785 & ~w13244;
assign w1108 = pi2480 & ~w5274;
assign w1109 = pi1384 & w13753;
assign w1110 = pi2050 & ~w10158;
assign w1111 = ~w16226 & ~w3971;
assign w1112 = ~pi0483 & pi3395;
assign w1113 = w6857 & w12720;
assign w1114 = ~pi2967 & pi3035;
assign w1115 = pi1166 & w13509;
assign w1116 = pi2498 & ~w15235;
assign w1117 = ~w9960 & ~w17959;
assign w1118 = ~w1791 & w13897;
assign w1119 = ~w11911 & ~w18339;
assign w1120 = ~pi2981 & w2460;
assign w1121 = (pi0349 & w6195) | (pi0349 & w7744) | (w6195 & w7744);
assign w1122 = w5453 & pi2489;
assign w1123 = ~pi3082 & w261;
assign w1124 = pi2690 & ~w261;
assign w1125 = ~w3055 & w14855;
assign w1126 = w12543 & w3791;
assign w1127 = ~w8430 & ~w16095;
assign w1128 = w9653 & w4304;
assign w1129 = pi1613 & w13753;
assign w1130 = ~w3972 & w11825;
assign w1131 = ~w9043 & w10704;
assign w1132 = ~pi0558 & w11739;
assign w1133 = w6697 & ~w1236;
assign w1134 = ~w2725 & pi0794;
assign w1135 = ~w13554 & ~w1444;
assign w1136 = w6857 & w7637;
assign w1137 = ~w17248 & pi1055;
assign w1138 = ~pi3003 & w16502;
assign w1139 = pi3004 & w16502;
assign w1140 = w7703 & w14249;
assign w1141 = w9440 & pi0191;
assign w1142 = pi1411 & ~w13753;
assign w1143 = ~pi0592 & w795;
assign w1144 = ~w11675 & ~w1354;
assign w1145 = ~pi3150 & ~pi3160;
assign w1146 = pi3020 & ~pi3112;
assign w1147 = w12543 & w795;
assign w1148 = pi2859 & w15191;
assign w1149 = ~pi0977 & w1147;
assign w1150 = ~w1401 & ~w10883;
assign w1151 = (pi0643 & ~w13509) | (pi0643 & w15295) | (~w13509 & w15295);
assign w1152 = ~w18107 & pi0483;
assign w1153 = ~pi3154 & w13570;
assign w1154 = (pi0843 & ~w13509) | (pi0843 & w4609) | (~w13509 & w4609);
assign w1155 = ~w8662 & w5679;
assign w1156 = pi2038 & ~w17646;
assign w1157 = ~w16288 & ~w2642;
assign w1158 = ~w14073 & w16518;
assign w1159 = ~w1177 & ~w10524;
assign w1160 = ~w5490 & w2562;
assign w1161 = w15761 & w16884;
assign w1162 = w13509 & w17564;
assign w1163 = w3203 & ~w17210;
assign w1164 = ~w6829 & ~w10124;
assign w1165 = ~w128 & ~w6060;
assign w1166 = w7844 & ~w14465;
assign w1167 = ~w6697 & pi1173;
assign w1168 = ~w5453 & ~pi1777;
assign w1169 = ~pi0999 & w12825;
assign w1170 = ~w11869 & ~w4919;
assign w1171 = pi0062 & w7658;
assign w1172 = (pi0824 & ~w13509) | (pi0824 & w14577) | (~w13509 & w14577);
assign w1173 = ~pi2491 & w15122;
assign w1174 = ~w17248 & pi0948;
assign w1175 = ~w5560 & w11903;
assign w1176 = ~w5603 & ~w5392;
assign w1177 = ~pi3172 & w13570;
assign w1178 = ~w14225 & ~w3706;
assign w1179 = ~w17665 & ~w9309;
assign w1180 = pi2726 & ~w261;
assign w1181 = ~w16130 & w18033;
assign w1182 = w7703 & w2906;
assign w1183 = ~w15622 & ~w12845;
assign w1184 = ~w11239 & ~w3843;
assign w1185 = ~pi3048 & w3555;
assign w1186 = ~pi3166 & w15048;
assign w1187 = w11345 & w1922;
assign w1188 = ~w10086 & ~w12532;
assign w1189 = ~pi1844 & w9340;
assign w1190 = ~w16283 & ~w16474;
assign w1191 = pi2605 & ~w16815;
assign w1192 = pi1477 & ~w9781;
assign w1193 = ~w968 & ~w14691;
assign w1194 = w11671 & w2753;
assign w1195 = pi0096 & w3748;
assign w1196 = ~w5329 & w10944;
assign w1197 = (pi0983 & ~w13509) | (pi0983 & w6514) | (~w13509 & w6514);
assign w1198 = ~pi0284 & w4058;
assign w1199 = w16428 & w14818;
assign w1200 = ~w1934 & w5477;
assign w1201 = ~w10407 & ~w5028;
assign w1202 = ~pi1998 & w3019;
assign w1203 = ~w6466 & ~w12032;
assign w1204 = ~w2725 & pi0779;
assign w1205 = ~pi3049 & w3555;
assign w1206 = ~w5855 & w12387;
assign w1207 = w6011 & w9326;
assign w1208 = pi3147 & w18497;
assign w1209 = ~w10045 & ~w9695;
assign w1210 = ~w16371 & ~w7419;
assign w1211 = ~w11574 & ~w15844;
assign w1212 = ~pi2024 & w7455;
assign w1213 = ~pi2235 & w2151;
assign w1214 = pi2071 & ~w4508;
assign w1215 = ~w328 & ~w11666;
assign w1216 = ~pi0625 & w14641;
assign w1217 = ~w1266 & ~w147;
assign w1218 = ~w15808 & pi0921;
assign w1219 = w17562 & pi1818;
assign w1220 = ~w1862 & ~w1690;
assign w1221 = pi1350 & ~w13786;
assign w1222 = ~pi3340 & w16922;
assign w1223 = ~w7844 & pi0595;
assign w1224 = pi1609 & ~w9781;
assign w1225 = pi2960 & w3196;
assign w1226 = ~w258 & ~w12747;
assign w1227 = pi2420 & ~w10158;
assign w1228 = ~w1522 & ~w15963;
assign w1229 = ~w11366 & ~w6775;
assign w1230 = w13509 & w3566;
assign w1231 = pi2881 & ~w3555;
assign w1232 = (pi0741 & ~w13509) | (pi0741 & w2257) | (~w13509 & w2257);
assign w1233 = pi1584 & ~w16922;
assign w1234 = pi3141 & w3987;
assign w1235 = w9440 & pi0179;
assign w1236 = ~w292 & ~w18482;
assign w1237 = w11383 & w16913;
assign w1238 = w13509 & w3137;
assign w1239 = ~w16365 & ~w10134;
assign w1240 = w2341 & ~w4179;
assign w1241 = w13509 & w2264;
assign w1242 = ~pi0283 & w4058;
assign w1243 = ~pi2301 & w16041;
assign w1244 = w15195 & w3022;
assign w1245 = w3425 & w16316;
assign w1246 = w12460 & w18059;
assign w1247 = w539 & ~w18063;
assign w1248 = ~pi2009 & w11688;
assign w1249 = pi2913 & ~w3186;
assign w1250 = pi0270 & w11070;
assign w1251 = ~w13246 & ~w5300;
assign w1252 = pi1195 & w11010;
assign w1253 = ~w15928 & ~w16736;
assign w1254 = ~w3938 & ~w7252;
assign w1255 = ~pi3093 & w6463;
assign w1256 = (pi0355 & w6195) | (pi0355 & w1597) | (w6195 & w1597);
assign w1257 = ~w16747 & ~w2330;
assign w1258 = pi2930 & ~w15235;
assign w1259 = pi2361 & ~w17683;
assign w1260 = ~w14648 & ~pi2711;
assign w1261 = ~w2341 & pi0832;
assign w1262 = pi1128 & ~pi1130;
assign w1263 = ~pi3172 & w11701;
assign w1264 = w13509 & w8950;
assign w1265 = ~w16533 & ~w14919;
assign w1266 = ~pi0502 & ~pi1345;
assign w1267 = ~pi3099 & w6463;
assign w1268 = pi3142 & w13786;
assign w1269 = pi2554 & ~w5274;
assign w1270 = w1962 & ~w14143;
assign w1271 = ~w15122 & ~pi1979;
assign w1272 = w1368 & pi0382;
assign w1273 = pi1658 & ~w13753;
assign w1274 = pi1636 & ~w13753;
assign w1275 = pi3157 & w8113;
assign w1276 = w10189 & ~pi0459;
assign w1277 = ~pi0871 & w15707;
assign w1278 = pi3365 & pi0222;
assign w1279 = ~w826 & ~w14190;
assign w1280 = (~pi2920 & ~w384) | (~pi2920 & w4257) | (~w384 & w4257);
assign w1281 = ~pi2454 & w9340;
assign w1282 = (~pi0287 & ~w6857) | (~pi0287 & w10426) | (~w6857 & w10426);
assign w1283 = ~pi2267 & w3019;
assign w1284 = ~pi3060 & w16815;
assign w1285 = (pi0661 & ~w13509) | (pi0661 & w11987) | (~w13509 & w11987);
assign w1286 = (~pi1201 & ~w13509) | (~pi1201 & w3507) | (~w13509 & w3507);
assign w1287 = w709 & pi1869;
assign w1288 = pi1142 & ~w6280;
assign w1289 = (pi0818 & ~w13509) | (pi0818 & w6594) | (~w13509 & w6594);
assign w1290 = ~w11956 & ~w5612;
assign w1291 = ~w3067 & ~w17474;
assign w1292 = ~pi0978 & w543;
assign w1293 = ~w13231 & pi0567;
assign w1294 = ~w9441 & ~w17226;
assign w1295 = pi0273 & ~pi1337;
assign w1296 = w13509 & w1650;
assign w1297 = pi2542 & w14148;
assign w1298 = pi3044 & ~pi3172;
assign w1299 = ~pi3326 & w6448;
assign w1300 = (~pi0489 & w17577) | (~pi0489 & w14011) | (w17577 & w14011);
assign w1301 = w6101 & w17048;
assign w1302 = ~pi2172 & w11313;
assign w1303 = w2637 & w15466;
assign w1304 = ~w5189 & pi0925;
assign w1305 = ~w6786 & ~w8811;
assign w1306 = w9316 & w15636;
assign w1307 = w7703 & w7381;
assign w1308 = ~w16503 & ~w3802;
assign w1309 = ~w9344 & ~w15322;
assign w1310 = ~w17745 & ~w18359;
assign w1311 = w10299 & w17115;
assign w1312 = w17562 & pi2573;
assign w1313 = (~w13546 & ~w9323) | (~w13546 & w15161) | (~w9323 & w15161);
assign w1314 = (~w9834 & ~w5517) | (~w9834 & w11829) | (~w5517 & w11829);
assign w1315 = ~pi2951 & pi3199;
assign w1316 = ~w8717 & ~w3785;
assign w1317 = ~w15183 & ~w4999;
assign w1318 = w5189 & ~w11978;
assign w1319 = pi2092 & ~w4420;
assign w1320 = pi2874 & ~w2431;
assign w1321 = pi0502 & ~pi1377;
assign w1322 = (w17357 & ~w7088) | (w17357 & w10069) | (~w7088 & w10069);
assign w1323 = ~w3611 & ~w16900;
assign w1324 = w1265 & w10897;
assign w1325 = w1443 & w1925;
assign w1326 = ~w11818 & w12858;
assign w1327 = ~w6299 & ~w13406;
assign w1328 = ~w11343 & ~w13367;
assign w1329 = ~w16955 & ~w13036;
assign w1330 = w13019 & w16135;
assign w1331 = w6741 & w5209;
assign w1332 = ~w10723 & ~w11168;
assign w1333 = ~w14648 & w11383;
assign w1334 = w13231 & ~w15296;
assign w1335 = pi2019 & ~w14833;
assign w1336 = ~w11121 & ~w11565;
assign w1337 = w2341 & ~w17210;
assign w1338 = ~w5266 & ~w13769;
assign w1339 = ~w9388 & ~w14458;
assign w1340 = ~w4938 & ~w3027;
assign w1341 = ~w6812 & ~w17929;
assign w1342 = w934 & pi0424;
assign w1343 = pi0339 & ~pi3254;
assign w1344 = pi2485 & w14148;
assign w1345 = w18331 & w6429;
assign w1346 = ~w6062 & ~w1162;
assign w1347 = ~pi2994 & w6448;
assign w1348 = ~w2533 & ~w8083;
assign w1349 = w13509 & w17685;
assign w1350 = (pi0753 & ~w13509) | (pi0753 & w13130) | (~w13509 & w13130);
assign w1351 = ~w2014 & w7710;
assign w1352 = pi0004 & ~w14148;
assign w1353 = pi2895 & ~w5274;
assign w1354 = ~pi2001 & w3019;
assign w1355 = w10276 & w18098;
assign w1356 = ~w6059 & ~w8219;
assign w1357 = pi3158 & w9520;
assign w1358 = ~w9655 & ~w6610;
assign w1359 = ~w10990 & ~w2913;
assign w1360 = ~w15122 & ~pi2673;
assign w1361 = ~pi0840 & w93;
assign w1362 = ~w13367 & w1770;
assign w1363 = w13509 & w10068;
assign w1364 = ~pi1257 & ~w11505;
assign w1365 = w5453 & pi2585;
assign w1366 = ~pi3094 & w16815;
assign w1367 = w4162 & w5323;
assign w1368 = ~w14961 & ~w6468;
assign w1369 = ~pi0822 & w1147;
assign w1370 = ~w6785 & pi1051;
assign w1371 = w6649 & ~w10492;
assign w1372 = ~pi2975 & w10299;
assign w1373 = ~pi3103 & w6463;
assign w1374 = pi2897 & ~w3555;
assign w1375 = ~pi2127 & w16041;
assign w1376 = ~w7285 & ~w6727;
assign w1377 = (pi0320 & w3055) | (pi0320 & w8388) | (w3055 & w8388);
assign w1378 = pi2277 & ~w9414;
assign w1379 = ~w3007 & ~w16579;
assign w1380 = w1368 & pi0399;
assign w1381 = w14874 & w13917;
assign w1382 = ~w10640 & ~w14207;
assign w1383 = ~w12461 & ~w16982;
assign w1384 = ~w1962 & pi0649;
assign w1385 = pi3172 & w3987;
assign w1386 = pi0206 & w10959;
assign w1387 = (pi1150 & ~w5437) | (pi1150 & w4542) | (~w5437 & w4542);
assign w1388 = ~pi2970 & ~w12458;
assign w1389 = ~w1564 & ~w15906;
assign w1390 = ~w3322 & ~w14942;
assign w1391 = w7254 & w13679;
assign w1392 = w1046 & w12866;
assign w1393 = w3788 & w6197;
assign w1394 = ~w2656 & ~w11016;
assign w1395 = ~w3216 & ~w10783;
assign w1396 = ~w6158 & ~w1995;
assign w1397 = w13509 & w7990;
assign w1398 = ~w9438 & ~w4196;
assign w1399 = w17248 & ~w15173;
assign w1400 = w7703 & w5879;
assign w1401 = ~w5978 & w7732;
assign w1402 = (pi0664 & ~w13509) | (pi0664 & w11462) | (~w13509 & w11462);
assign w1403 = ~w10383 & ~w8362;
assign w1404 = ~w16677 & ~w14058;
assign w1405 = ~w8309 & ~w15961;
assign w1406 = ~pi2686 & w17213;
assign w1407 = w9720 & pi1707;
assign w1408 = (pi0632 & ~w13509) | (pi0632 & w12162) | (~w13509 & w12162);
assign w1409 = ~w5189 & pi1029;
assign w1410 = ~w14351 & ~w1139;
assign w1411 = w16278 & ~w15173;
assign w1412 = ~w12292 & ~w4106;
assign w1413 = pi0150 & w5274;
assign w1414 = (pi0689 & ~w13509) | (pi0689 & w13336) | (~w13509 & w13336);
assign w1415 = ~w12040 & pi0937;
assign w1416 = ~w8721 & ~w7616;
assign w1417 = ~pi2476 & w5384;
assign w1418 = pi1628 & ~w18259;
assign w1419 = ~w4667 & ~w11606;
assign w1420 = ~w4664 & ~w13013;
assign w1421 = w2873 & w5949;
assign w1422 = w6785 & ~w7020;
assign w1423 = pi3138 & w5457;
assign w1424 = w10158 & w3515;
assign w1425 = w7844 & ~w2776;
assign w1426 = w6857 & w11189;
assign w1427 = w12408 & w802;
assign w1428 = ~w7529 & ~w15544;
assign w1429 = ~w3457 & ~w9232;
assign w1430 = pi2489 & ~w5274;
assign w1431 = ~w16506 & pi1191;
assign w1432 = pi3160 & ~w16618;
assign w1433 = pi1849 & w7799;
assign w1434 = ~pi2069 & w8617;
assign w1435 = w15808 & ~w7020;
assign w1436 = ~w5651 & w3642;
assign w1437 = pi1459 & ~w7090;
assign w1438 = ~pi2987 & w16815;
assign w1439 = pi2969 & ~w3987;
assign w1440 = ~w7532 & ~w3635;
assign w1441 = pi1579 & w13753;
assign w1442 = ~w4991 & ~w11586;
assign w1443 = w17517 & w14182;
assign w1444 = w384 & w5462;
assign w1445 = ~w1791 & w12118;
assign w1446 = ~w6140 & ~w14726;
assign w1447 = (pi0585 & ~w13509) | (pi0585 & w7225) | (~w13509 & w7225);
assign w1448 = ~w3586 & ~w2957;
assign w1449 = pi2653 & ~w9504;
assign w1450 = (pi0737 & ~w13509) | (pi0737 & w8117) | (~w13509 & w8117);
assign w1451 = w8324 & ~w13869;
assign w1452 = ~pi0718 & w17899;
assign w1453 = w12808 & w271;
assign w1454 = (pi1198 & w4470) | (pi1198 & w6906) | (w4470 & w6906);
assign w1455 = ~w3534 & ~w6292;
assign w1456 = ~w2341 & pi1066;
assign w1457 = ~pi0546 & w3106;
assign w1458 = ~w10694 & w17640;
assign w1459 = w5189 & ~w14978;
assign w1460 = w14833 & w6320;
assign w1461 = pi1669 & w1924;
assign w1462 = pi2147 & ~w11671;
assign w1463 = (~pi3117 & w13762) | (~pi3117 & w2415) | (w13762 & w2415);
assign w1464 = w7077 & ~w305;
assign w1465 = w6187 & w3406;
assign w1466 = ~w16040 & ~w13981;
assign w1467 = ~w8026 & ~w2660;
assign w1468 = pi0053 & pi0055;
assign w1469 = (pi0897 & ~w13509) | (pi0897 & w8647) | (~w13509 & w8647);
assign w1470 = ~w139 & ~w13534;
assign w1471 = ~w14146 & ~w15200;
assign w1472 = ~w12474 & ~w16013;
assign w1473 = ~w11059 & ~w9;
assign w1474 = ~pi2835 & w13343;
assign w1475 = (w5421 & ~w9786) | (w5421 & w5664) | (~w9786 & w5664);
assign w1476 = ~w16575 & w1580;
assign w1477 = w6785 & ~w1236;
assign w1478 = w15122 & ~pi2633;
assign w1479 = ~w11230 & ~w4147;
assign w1480 = pi2969 & w11077;
assign w1481 = pi2241 & ~w4420;
assign w1482 = pi3160 & ~w17286;
assign w1483 = ~pi0305 & pi0306;
assign w1484 = pi0143 & w5274;
assign w1485 = w16873 & w14282;
assign w1486 = ~w5454 & ~w16793;
assign w1487 = pi2942 & ~pi3208;
assign w1488 = pi1423 & ~w13753;
assign w1489 = w7077 & ~w3430;
assign w1490 = w13509 & w11269;
assign w1491 = ~w4725 & ~w16964;
assign w1492 = pi3046 & ~w16502;
assign w1493 = ~pi0311 & pi0312;
assign w1494 = ~w11300 & w16211;
assign w1495 = w8789 & pi0463;
assign w1496 = w7844 & ~w9852;
assign w1497 = ~w17374 & w17232;
assign w1498 = w8324 & w1343;
assign w1499 = ~pi3058 & w16815;
assign w1500 = w7195 & w4818;
assign w1501 = (pi0593 & ~w13509) | (pi0593 & w12951) | (~w13509 & w12951);
assign w1502 = w5453 & pi2889;
assign w1503 = pi1280 & pi1345;
assign w1504 = ~w8602 & ~w1286;
assign w1505 = (~pi1219 & w907) | (~pi1219 & w15398) | (w907 & w15398);
assign w1506 = ~w17548 & ~w4012;
assign w1507 = w13509 & w17546;
assign w1508 = pi1525 & w13753;
assign w1509 = w8520 & w6194;
assign w1510 = ~pi3135 & w15132;
assign w1511 = ~w11228 & ~w1413;
assign w1512 = w2306 & w8653;
assign w1513 = w7703 & w3714;
assign w1514 = ~w7914 & ~w18055;
assign w1515 = ~pi3157 & w12427;
assign w1516 = w2579 & w17906;
assign w1517 = ~pi3005 & pi3165;
assign w1518 = pi1277 & pi1345;
assign w1519 = ~w7327 & ~w4982;
assign w1520 = pi1949 & ~w17646;
assign w1521 = ~w7695 & w17334;
assign w1522 = (pi0828 & ~w13509) | (pi0828 & w11980) | (~w13509 & w11980);
assign w1523 = pi1337 & ~pi0255;
assign w1524 = w13509 & w7002;
assign w1525 = ~pi3052 & w261;
assign w1526 = pi1395 & w12817;
assign w1527 = w13509 & w5765;
assign w1528 = w15743 & w8310;
assign w1529 = ~w11277 & ~w13075;
assign w1530 = ~w17376 & w6406;
assign w1531 = ~w3719 & ~w1436;
assign w1532 = pi2144 & ~w15883;
assign w1533 = w9440 & pi0135;
assign w1534 = pi1338 & ~w2848;
assign w1535 = ~w6195 & w3220;
assign w1536 = ~pi2015 & w11688;
assign w1537 = w15717 & ~w8345;
assign w1538 = ~pi3316 & w16922;
assign w1539 = w13509 & w15766;
assign w1540 = w8446 & w16943;
assign w1541 = ~pi0098 & w9284;
assign w1542 = pi0099 & w9284;
assign w1543 = ~w16778 & ~w13264;
assign w1544 = ~pi2910 & ~w5644;
assign w1545 = pi2487 & ~w6463;
assign w1546 = ~pi1100 & w17899;
assign w1547 = (pi1005 & ~w13509) | (pi1005 & w4078) | (~w13509 & w4078);
assign w1548 = w15271 & w14078;
assign w1549 = ~w15230 & ~w8299;
assign w1550 = (pi0801 & ~w13509) | (pi0801 & w17486) | (~w13509 & w17486);
assign w1551 = w7844 & ~w15173;
assign w1552 = ~pi3166 & w8515;
assign w1553 = w17248 & ~w12800;
assign w1554 = pi1766 & ~w14951;
assign w1555 = ~pi2115 & w12755;
assign w1556 = ~w4266 & ~w2499;
assign w1557 = ~w16541 & w16117;
assign w1558 = ~w5194 & ~w16828;
assign w1559 = pi2853 & w15191;
assign w1560 = ~pi0054 & w922;
assign w1561 = pi0055 & w922;
assign w1562 = ~pi1719 & pi3151;
assign w1563 = (pi1197 & ~w13509) | (pi1197 & w5543) | (~w13509 & w5543);
assign w1564 = w6857 & w10309;
assign w1565 = w12040 & ~w2587;
assign w1566 = w8745 & w18188;
assign w1567 = ~w7713 & ~w12148;
assign w1568 = ~pi3139 & w15048;
assign w1569 = ~pi2309 & w12724;
assign w1570 = ~w14648 & ~pi2620;
assign w1571 = ~pi1091 & w6200;
assign w1572 = pi1630 & ~w18259;
assign w1573 = pi0061 & ~w14148;
assign w1574 = ~w6785 & pi0516;
assign w1575 = ~w15309 & ~w4956;
assign w1576 = ~w11655 & w6109;
assign w1577 = pi2456 & ~w14524;
assign w1578 = ~w14571 & ~w15226;
assign w1579 = w9440 & pi0152;
assign w1580 = w10189 & pi0403;
assign w1581 = ~w16278 & pi0708;
assign w1582 = (pi0771 & ~w13509) | (pi0771 & w10270) | (~w13509 & w10270);
assign w1583 = w968 & ~pi0285;
assign w1584 = w14109 & pi0447;
assign w1585 = ~w6785 & pi0851;
assign w1586 = ~w3054 & w15596;
assign w1587 = ~w10941 & ~w13403;
assign w1588 = ~pi2928 & w15122;
assign w1589 = pi1612 & w13753;
assign w1590 = ~w1933 & ~w10513;
assign w1591 = ~pi1018 & w9110;
assign w1592 = ~w6635 & ~w14632;
assign w1593 = ~pi3313 & w6072;
assign w1594 = ~w1791 & w9883;
assign w1595 = pi0077 & pi3117;
assign w1596 = pi1337 & ~pi2989;
assign w1597 = w14560 & pi0355;
assign w1598 = pi1367 & pi1371;
assign w1599 = (~w14652 & w5855) | (~w14652 & w4660) | (w5855 & w4660);
assign w1600 = w12040 & ~w14978;
assign w1601 = pi2512 & ~w9504;
assign w1602 = ~w3000 & ~pi1747;
assign w1603 = ~pi3134 & ~pi3142;
assign w1604 = w13509 & w1240;
assign w1605 = w13367 & w18435;
assign w1606 = ~w14985 & ~w13104;
assign w1607 = w17248 & ~w14978;
assign w1608 = ~pi0683 & w9110;
assign w1609 = w384 & w4829;
assign w1610 = ~pi3061 & w3555;
assign w1611 = w17562 & w8303;
assign w1612 = pi1307 & pi3213;
assign w1613 = w6697 & ~w15296;
assign w1614 = (pi0878 & ~w13509) | (pi0878 & w7890) | (~w13509 & w7890);
assign w1615 = ~w12039 & ~w14606;
assign w1616 = w13509 & w15488;
assign w1617 = ~w13101 & ~w4430;
assign w1618 = w2946 & w15112;
assign w1619 = pi1716 & ~w619;
assign w1620 = w6282 & w6814;
assign w1621 = ~w2608 & ~w13598;
assign w1622 = (~pi0285 & ~w6857) | (~pi0285 & w1583) | (~w6857 & w1583);
assign w1623 = w2130 & ~w858;
assign w1624 = w13509 & w10436;
assign w1625 = w7077 & ~w17513;
assign w1626 = ~w5560 & w14200;
assign w1627 = ~w17248 & pi0875;
assign w1628 = ~w15746 & ~w17535;
assign w1629 = ~w7656 & pi2913;
assign w1630 = pi1591 & ~w13753;
assign w1631 = pi1437 & ~w13753;
assign w1632 = pi1329 & pi1345;
assign w1633 = pi1674 & w1924;
assign w1634 = pi1543 & w13753;
assign w1635 = w16941 & w14610;
assign w1636 = ~pi3057 & ~w18328;
assign w1637 = w2547 & w2684;
assign w1638 = ~w14269 & w17537;
assign w1639 = w6422 & w7265;
assign w1640 = pi1354 & w11685;
assign w1641 = w7582 & w1316;
assign w1642 = ~pi3088 & w11406;
assign w1643 = w14285 & w1615;
assign w1644 = w17248 & ~w7020;
assign w1645 = w8658 & pi1780;
assign w1646 = w13509 & w1435;
assign w1647 = pi1595 & ~w13786;
assign w1648 = ~w17577 & w3588;
assign w1649 = ~w4667 & ~w16721;
assign w1650 = w1391 & ~w14978;
assign w1651 = ~w10191 & ~w5749;
assign w1652 = w17248 & ~w2776;
assign w1653 = pi1629 & ~w18259;
assign w1654 = ~w5377 & ~w13405;
assign w1655 = w10189 & pi0392;
assign w1656 = ~w575 & ~w10245;
assign w1657 = ~pi2860 & w15122;
assign w1658 = ~pi3355 & w17935;
assign w1659 = pi1231 & w11655;
assign w1660 = pi0497 & pi1191;
assign w1661 = pi2669 & ~w6463;
assign w1662 = ~pi2685 & w17213;
assign w1663 = pi1749 & ~w16815;
assign w1664 = ~pi3139 & w11132;
assign w1665 = ~w13491 & ~w6298;
assign w1666 = w13509 & w16412;
assign w1667 = w2725 & ~w13195;
assign w1668 = ~pi2975 & w15271;
assign w1669 = ~w10553 & ~w17247;
assign w1670 = ~w6155 & ~w4441;
assign w1671 = ~w1791 & w4603;
assign w1672 = ~pi2006 & w11688;
assign w1673 = (pi0804 & ~w13509) | (pi0804 & w18470) | (~w13509 & w18470);
assign w1674 = ~pi3426 & w15036;
assign w1675 = ~w5371 & ~w17176;
assign w1676 = ~w10399 & ~w1424;
assign w1677 = w15122 & ~pi2700;
assign w1678 = w11383 & w10589;
assign w1679 = ~w6885 & ~w3708;
assign w1680 = w12040 & ~w14143;
assign w1681 = ~w10040 & w3866;
assign w1682 = w6352 & ~pi0444;
assign w1683 = ~pi2942 & pi3208;
assign w1684 = ~w750 & w2249;
assign w1685 = pi1351 & w14565;
assign w1686 = ~pi2322 & w12941;
assign w1687 = ~pi3008 & ~pi3207;
assign w1688 = ~w14420 & w15337;
assign w1689 = w14109 & pi0415;
assign w1690 = ~pi0890 & w1126;
assign w1691 = ~pi3159 & w3805;
assign w1692 = ~pi3158 & w17387;
assign w1693 = ~w14448 & ~w2459;
assign w1694 = ~pi2976 & w9504;
assign w1695 = ~pi3299 & w14918;
assign w1696 = pi2472 & ~w14524;
assign w1697 = ~w16601 & ~w16600;
assign w1698 = (pi0260 & ~w325) | (pi0260 & w4940) | (~w325 & w4940);
assign w1699 = w9155 & ~w8646;
assign w1700 = ~w17248 & pi0873;
assign w1701 = w14228 & w11302;
assign w1702 = ~pi3038 & ~pi3207;
assign w1703 = ~pi1109 & w12197;
assign w1704 = pi1917 & ~w15271;
assign w1705 = pi0304 & w5113;
assign w1706 = w1824 & w16938;
assign w1707 = pi2545 & w14148;
assign w1708 = w6649 & ~w6723;
assign w1709 = ~w7753 & ~w18068;
assign w1710 = ~pi1692 & ~w6857;
assign w1711 = ~w8324 & ~w2064;
assign w1712 = ~pi2967 & ~pi3105;
assign w1713 = ~w15199 & ~w15672;
assign w1714 = w16506 & ~w17513;
assign w1715 = (~pi1237 & ~w8966) | (~pi1237 & w15333) | (~w8966 & w15333);
assign w1716 = w5642 & w13318;
assign w1717 = ~w12290 & w16588;
assign w1718 = ~w8709 & ~w9418;
assign w1719 = ~w3801 & ~w17574;
assign w1720 = w13509 & w13875;
assign w1721 = pi0015 & ~w3748;
assign w1722 = w3404 & w8244;
assign w1723 = pi2243 & ~w15883;
assign w1724 = w5989 & w490;
assign w1725 = w7077 & ~w2741;
assign w1726 = ~pi3059 & w261;
assign w1727 = pi2758 & ~w3987;
assign w1728 = w13509 & w16797;
assign w1729 = ~pi1111 & w12197;
assign w1730 = (pi1007 & ~w13509) | (pi1007 & w867) | (~w13509 & w867);
assign w1731 = ~w16508 & ~w1738;
assign w1732 = ~w6189 & ~w15193;
assign w1733 = w17248 & ~w4043;
assign w1734 = ~w13714 & ~w12068;
assign w1735 = ~pi2343 & w12724;
assign w1736 = pi1592 & ~w13753;
assign w1737 = w13231 & ~w3430;
assign w1738 = ~pi1243 & pi1267;
assign w1739 = ~pi3147 & w17669;
assign w1740 = w6785 & ~w13028;
assign w1741 = pi0057 & ~w14148;
assign w1742 = pi1792 & ~w9520;
assign w1743 = ~w15861 & w9498;
assign w1744 = ~w10225 & w963;
assign w1745 = ~w4022 & ~w7644;
assign w1746 = ~pi3046 & pi3146;
assign w1747 = (~pi2966 & ~w384) | (~pi2966 & w4385) | (~w384 & w4385);
assign w1748 = w3243 & ~pi0267;
assign w1749 = pi2767 & w605;
assign w1750 = ~w9101 & ~w2048;
assign w1751 = ~w17404 & ~w12907;
assign w1752 = ~pi1171 & ~pi3209;
assign w1753 = ~w5453 & ~pi1772;
assign w1754 = w11209 & ~w1041;
assign w1755 = w16575 & w16045;
assign w1756 = ~pi3069 & pi3168;
assign w1757 = ~pi3311 & w9781;
assign w1758 = ~w24 & ~w17000;
assign w1759 = ~pi3060 & w3555;
assign w1760 = ~w4890 & ~w5555;
assign w1761 = ~w9199 & ~w11063;
assign w1762 = w10299 & w3515;
assign w1763 = ~w8024 & ~w12812;
assign w1764 = w1872 & w18174;
assign w1765 = w7307 & w13653;
assign w1766 = w11405 & ~w10843;
assign w1767 = ~w12933 & w84;
assign w1768 = w17562 & pi2562;
assign w1769 = ~pi2231 & w11313;
assign w1770 = (pi0504 & ~w6217) | (pi0504 & ~w17577) | (~w6217 & ~w17577);
assign w1771 = ~w6697 & pi0673;
assign w1772 = w13509 & w18471;
assign w1773 = ~w13748 & ~w10877;
assign w1774 = ~w312 & ~w7312;
assign w1775 = pi0514 & pi1187;
assign w1776 = ~w13822 & w10382;
assign w1777 = w11216 & w15278;
assign w1778 = w5743 & w3080;
assign w1779 = w13509 & w1006;
assign w1780 = pi3135 & w5457;
assign w1781 = ~w17248 & pi0884;
assign w1782 = ~w11820 & w13484;
assign w1783 = ~pi0707 & w3106;
assign w1784 = w15808 & ~w11978;
assign w1785 = ~w15230 & ~w2056;
assign w1786 = ~w7077 & pi0817;
assign w1787 = w17683 & w6320;
assign w1788 = ~w17338 & ~w14499;
assign w1789 = ~w8064 & ~w18370;
assign w1790 = w3243 & ~w976;
assign w1791 = ~w13695 & ~w9266;
assign w1792 = ~w15306 & w7945;
assign w1793 = ~w9997 & ~w6112;
assign w1794 = ~pi2004 & w3019;
assign w1795 = w15271 & w6320;
assign w1796 = ~w18596 & ~w4634;
assign w1797 = ~w14560 & pi0238;
assign w1798 = pi1446 & ~w13753;
assign w1799 = w13509 & w2799;
assign w1800 = ~w15917 & ~w4125;
assign w1801 = ~pi0715 & w3106;
assign w1802 = ~w1791 & w4716;
assign w1803 = ~w10487 & ~w17928;
assign w1804 = ~pi2922 & ~pi2923;
assign w1805 = ~w1715 & w224;
assign w1806 = w14228 & ~w16498;
assign w1807 = w7703 & w16845;
assign w1808 = pi3011 & w16502;
assign w1809 = w13509 & w10937;
assign w1810 = ~w6656 & ~w9428;
assign w1811 = ~w13097 & ~w7957;
assign w1812 = w13509 & w8873;
assign w1813 = w16184 & w8472;
assign w1814 = ~pi0352 & w2196;
assign w1815 = ~w16967 & w12593;
assign w1816 = ~w3812 & ~w9923;
assign w1817 = w4087 & w14273;
assign w1818 = ~pi0498 & ~w9980;
assign w1819 = ~w15122 & ~pi1883;
assign w1820 = ~w10702 & ~w8546;
assign w1821 = ~pi3138 & ~pi3160;
assign w1822 = w922 & w7952;
assign w1823 = pi1845 & ~w12558;
assign w1824 = ~w5145 & ~w2079;
assign w1825 = ~pi1035 & w6200;
assign w1826 = pi0301 & w1206;
assign w1827 = w625 & pi0496;
assign w1828 = w13509 & w1459;
assign w1829 = pi1646 & ~w6448;
assign w1830 = w12460 & w941;
assign w1831 = ~w9619 & w17714;
assign w1832 = pi1407 & ~w9781;
assign w1833 = ~w2985 & ~w342;
assign w1834 = pi0411 & w9129;
assign w1835 = ~pi2341 & w16041;
assign w1836 = ~w3947 & ~w8445;
assign w1837 = ~w4151 & ~w9018;
assign w1838 = ~w16903 & ~w5159;
assign w1839 = ~w8485 & ~w15426;
assign w1840 = ~pi2940 & pi3208;
assign w1841 = w15842 & pi2738;
assign w1842 = ~w8478 & ~w17575;
assign w1843 = ~w4020 & w3223;
assign w1844 = ~w4887 & ~w17851;
assign w1845 = w13509 & w11105;
assign w1846 = ~w4414 & ~w7484;
assign w1847 = ~w28 & ~pi1152;
assign w1848 = ~w11425 & ~w14944;
assign w1849 = ~w16575 & w2953;
assign w1850 = w7844 & ~w7707;
assign w1851 = ~w11838 & ~w1366;
assign w1852 = w17248 & ~w7707;
assign w1853 = w13549 & w12307;
assign w1854 = ~pi1337 & ~w12712;
assign w1855 = pi2630 & ~w261;
assign w1856 = ~w8351 & ~w12299;
assign w1857 = ~w7383 & ~w2972;
assign w1858 = pi0485 & pi0486;
assign w1859 = (pi0711 & ~w13509) | (pi0711 & w14353) | (~w13509 & w14353);
assign w1860 = ~w2341 & pi0831;
assign w1861 = pi1351 & ~w4324;
assign w1862 = ~pi0797 & w543;
assign w1863 = pi1314 & w11356;
assign w1864 = ~pi1209 & pi1182;
assign w1865 = w7703 & w10830;
assign w1866 = w1127 & ~w12280;
assign w1867 = w978 & ~w7161;
assign w1868 = w14648 & ~pi2734;
assign w1869 = ~w11138 & w9341;
assign w1870 = w12460 & w17754;
assign w1871 = ~w11261 & ~w17064;
assign w1872 = w16245 & w6717;
assign w1873 = ~pi1060 & w93;
assign w1874 = w13509 & w1337;
assign w1875 = pi1761 & ~pi1816;
assign w1876 = pi1570 & ~w18259;
assign w1877 = pi0090 & w9284;
assign w1878 = w14228 & ~w2587;
assign w1879 = pi1216 & ~w14583;
assign w1880 = pi2877 & ~w226;
assign w1881 = ~w3203 & pi0997;
assign w1882 = w10189 & ~pi0470;
assign w1883 = w11209 & ~w10268;
assign w1884 = ~w2461 & ~w431;
assign w1885 = ~pi3100 & w9504;
assign w1886 = ~w5855 & w4981;
assign w1887 = ~pi3162 & w11701;
assign w1888 = ~w10759 & ~w16235;
assign w1889 = ~w10055 & ~w15455;
assign w1890 = w2227 & w17379;
assign w1891 = pi1568 & ~w18259;
assign w1892 = ~pi1264 & w4880;
assign w1893 = w14109 & pi0419;
assign w1894 = ~pi2801 & w13343;
assign w1895 = (pi1792 & w5453) | (pi1792 & w7806) | (w5453 & w7806);
assign w1896 = w968 & ~pi0278;
assign w1897 = pi1549 & ~w17935;
assign w1898 = (pi0321 & w3055) | (pi0321 & w13185) | (w3055 & w13185);
assign w1899 = w11735 & w614;
assign w1900 = ~pi1984 & ~w7858;
assign w1901 = w741 & w6804;
assign w1902 = ~pi3096 & w15235;
assign w1903 = w13509 & w5791;
assign w1904 = ~w3000 & ~pi2671;
assign w1905 = (~pi1776 & ~w7799) | (~pi1776 & w10311) | (~w7799 & w10311);
assign w1906 = pi0270 & w5113;
assign w1907 = ~pi2469 & w5384;
assign w1908 = pi2995 & pi1399;
assign w1909 = w15027 & w18580;
assign w1910 = ~w4389 & ~w3760;
assign w1911 = ~pi1830 & w11313;
assign w1912 = ~w3388 & ~w4783;
assign w1913 = w14352 & w12984;
assign w1914 = (~pi0279 & ~w6857) | (~pi0279 & w14495) | (~w6857 & w14495);
assign w1915 = ~w1368 & ~pi0478;
assign w1916 = ~w3203 & pi0580;
assign w1917 = w13509 & w16615;
assign w1918 = ~pi3139 & w8515;
assign w1919 = w9720 & pi1717;
assign w1920 = ~w9264 & w5502;
assign w1921 = w934 & pi0419;
assign w1922 = ~pi0483 & pi3391;
assign w1923 = ~w13231 & pi0568;
assign w1924 = (w10959 & ~w12460) | (w10959 & w7338) | (~w12460 & w7338);
assign w1925 = ~w5536 & w11139;
assign w1926 = ~w1962 & ~pi0958;
assign w1927 = w5090 & w11720;
assign w1928 = pi3163 & w4324;
assign w1929 = ~w11021 & ~w14395;
assign w1930 = ~pi2326 & w16041;
assign w1931 = pi2286 & ~w3223;
assign w1932 = w4508 & w9407;
assign w1933 = pi1536 & ~w17935;
assign w1934 = ~w1892 & ~w13812;
assign w1935 = w5189 & ~w9852;
assign w1936 = ~w5560 & w5219;
assign w1937 = pi2707 & ~w16815;
assign w1938 = ~w17458 & ~w14966;
assign w1939 = w1453 & w7816;
assign w1940 = ~pi3340 & w9781;
assign w1941 = pi0173 & w5274;
assign w1942 = ~pi0819 & w1147;
assign w1943 = w14648 & ~pi2729;
assign w1944 = w13231 & ~w1236;
assign w1945 = w16278 & ~w12800;
assign w1946 = w17376 & pi0298;
assign w1947 = w17248 & ~w9852;
assign w1948 = ~w5453 & ~pi1774;
assign w1949 = w6857 & w2566;
assign w1950 = ~w672 & ~w13228;
assign w1951 = w16937 & w761;
assign w1952 = (pi0348 & w6195) | (pi0348 & w5211) | (w6195 & w5211);
assign w1953 = ~pi2783 & w13343;
assign w1954 = w5189 & ~w305;
assign w1955 = w14648 & ~pi2617;
assign w1956 = w9214 & w4165;
assign w1957 = (pi0859 & ~w13509) | (pi0859 & w6003) | (~w13509 & w6003);
assign w1958 = ~w16939 & pi0005;
assign w1959 = ~w14560 & pi0226;
assign w1960 = ~pi2976 & w6463;
assign w1961 = ~w6777 & ~w1021;
assign w1962 = w13867 & w6676;
assign w1963 = ~w870 & ~w8575;
assign w1964 = w11345 & w3085;
assign w1965 = w3203 & ~w9852;
assign w1966 = ~w7922 & ~w15185;
assign w1967 = w14560 & pi0373;
assign w1968 = ~pi0287 & w4058;
assign w1969 = ~w16590 & ~w6559;
assign w1970 = ~pi3333 & w9781;
assign w1971 = w6697 & ~w305;
assign w1972 = ~w5002 & ~w4834;
assign w1973 = pi2206 & ~w3223;
assign w1974 = w3988 & w17130;
assign w1975 = w10759 & w16759;
assign w1976 = w13509 & w14548;
assign w1977 = w7703 & w17678;
assign w1978 = ~w11920 & ~w10317;
assign w1979 = ~pi2243 & w12941;
assign w1980 = pi1601 & ~w9781;
assign w1981 = ~w15843 & ~w9097;
assign w1982 = ~w15064 & w13983;
assign w1983 = w8078 & w4459;
assign w1984 = ~w16506 & pi1144;
assign w1985 = w16547 & w2097;
assign w1986 = ~pi0297 & w4058;
assign w1987 = ~w17668 & ~w18448;
assign w1988 = ~w4558 & ~w7591;
assign w1989 = pi2848 & w4140;
assign w1990 = ~w9609 & ~w13317;
assign w1991 = w11383 & w4322;
assign w1992 = ~w7342 & ~w6455;
assign w1993 = pi3172 & w10992;
assign w1994 = pi3133 & w9520;
assign w1995 = ~pi0863 & w15707;
assign w1996 = w6697 & ~w6922;
assign w1997 = pi1234 & pi1376;
assign w1998 = ~w1391 & pi0765;
assign w1999 = w9440 & pi0184;
assign w2000 = pi1615 & w13753;
assign w2001 = w13509 & w69;
assign w2002 = w14524 & w9407;
assign w2003 = ~w4265 & w15695;
assign w2004 = ~w16949 & ~w2033;
assign w2005 = pi2049 & ~w10158;
assign w2006 = ~w7210 & ~w15614;
assign w2007 = pi0301 & w5274;
assign w2008 = w922 & ~w12638;
assign w2009 = ~w1292 & ~w1149;
assign w2010 = ~w17248 & pi0893;
assign w2011 = ~w5189 & ~pi0969;
assign w2012 = ~w9759 & ~w4749;
assign w2013 = ~w5724 & w14664;
assign w2014 = w9721 & w8598;
assign w2015 = (pi0669 & ~w13509) | (pi0669 & w18419) | (~w13509 & w18419);
assign w2016 = pi2299 & ~w4508;
assign w2017 = ~pi2946 & w15235;
assign w2018 = w7278 & ~w18096;
assign w2019 = ~w549 & ~w1681;
assign w2020 = ~w9164 & w16771;
assign w2021 = ~w12745 & ~w2323;
assign w2022 = ~w15064 & ~w17129;
assign w2023 = w2341 & ~w3374;
assign w2024 = w384 & w11490;
assign w2025 = ~w18473 & ~w4271;
assign w2026 = ~w2649 & ~w9567;
assign w2027 = ~w9143 & w10812;
assign w2028 = w7844 & ~w7449;
assign w2029 = w14893 & w9135;
assign w2030 = ~w3632 & ~w2451;
assign w2031 = pi2193 & ~w10299;
assign w2032 = pi3150 & w2732;
assign w2033 = pi2915 & pi2953;
assign w2034 = ~pi1960 & w11688;
assign w2035 = ~w1391 & pi1037;
assign w2036 = ~w12683 & ~w9692;
assign w2037 = w8761 & w10219;
assign w2038 = ~w10393 & ~w13199;
assign w2039 = ~pi1803 & ~pi3138;
assign w2040 = pi2113 & ~w412;
assign w2041 = ~w6891 & ~w7443;
assign w2042 = ~w8584 & w14827;
assign w2043 = ~w1 & ~w12152;
assign w2044 = (pi0996 & ~w13509) | (pi0996 & w7433) | (~w13509 & w7433);
assign w2045 = ~w1391 & pi0768;
assign w2046 = ~w13497 & w9675;
assign w2047 = w13840 & pi1365;
assign w2048 = w17302 & w10893;
assign w2049 = w12460 & w3741;
assign w2050 = ~pi0493 & ~pi1141;
assign w2051 = ~w3000 & w2263;
assign w2052 = ~w709 & pi1280;
assign w2053 = ~w6367 & ~w11249;
assign w2054 = w17248 & ~w14597;
assign w2055 = ~pi3108 & ~w3987;
assign w2056 = pi3109 & ~w3987;
assign w2057 = ~pi3313 & w18259;
assign w2058 = ~pi3416 & w15036;
assign w2059 = w13509 & w9885;
assign w2060 = pi1701 & ~w18497;
assign w2061 = w2179 & w7601;
assign w2062 = ~w10054 & ~w1264;
assign w2063 = ~w5640 & ~w16069;
assign w2064 = ~w9991 & w2354;
assign w2065 = w15244 & w2539;
assign w2066 = ~w8588 & w17683;
assign w2067 = ~w14853 & ~w996;
assign w2068 = ~pi2154 & w13065;
assign w2069 = ~pi2980 & pi3057;
assign w2070 = w13509 & w2140;
assign w2071 = w7656 & pi1211;
assign w2072 = ~w3203 & pi0590;
assign w2073 = w13509 & w513;
assign w2074 = ~pi0976 & w93;
assign w2075 = ~w12040 & pi0691;
assign w2076 = pi1951 & ~w17646;
assign w2077 = ~w7331 & ~w12463;
assign w2078 = pi3072 & ~w16502;
assign w2079 = ~pi1836 & w17439;
assign w2080 = pi0417 & w17173;
assign w2081 = w3402 & ~w16638;
assign w2082 = pi0171 & w5274;
assign w2083 = ~pi3056 & w11406;
assign w2084 = pi1251 & pi3237;
assign w2085 = ~w95 & ~w3717;
assign w2086 = ~pi2096 & w12724;
assign w2087 = pi0112 & w9284;
assign w2088 = ~w372 & ~w9779;
assign w2089 = pi2302 & ~w15883;
assign w2090 = ~pi0748 & w17490;
assign w2091 = w14228 & ~w7449;
assign w2092 = (pi1865 & w2014) | (pi1865 & w8751) | (w2014 & w8751);
assign w2093 = w4262 & w6899;
assign w2094 = ~pi3411 & w15036;
assign w2095 = (~pi0490 & w17577) | (~pi0490 & w9239) | (w17577 & w9239);
assign w2096 = ~w5189 & pi0720;
assign w2097 = ~w9193 & ~w1825;
assign w2098 = ~w9375 & ~w3764;
assign w2099 = ~w3054 & w7518;
assign w2100 = ~pi2297 & w12941;
assign w2101 = ~w16575 & w15047;
assign w2102 = ~w17212 & ~w5255;
assign w2103 = ~w11463 & ~w13407;
assign w2104 = ~w13604 & ~w13378;
assign w2105 = ~w13580 & ~w2059;
assign w2106 = w14094 & w9452;
assign w2107 = ~w16960 & ~w13474;
assign w2108 = w14109 & pi0423;
assign w2109 = ~w1274 & w6912;
assign w2110 = pi0118 & w3748;
assign w2111 = (~w4182 & ~w5517) | (~w4182 & w4471) | (~w5517 & w4471);
assign w2112 = ~pi2159 & w17439;
assign w2113 = ~w13522 & ~w6050;
assign w2114 = ~w478 & ~w4458;
assign w2115 = pi1662 & ~w4058;
assign w2116 = pi3160 & ~w10784;
assign w2117 = ~w2014 & w2983;
assign w2118 = ~w5951 & ~w17331;
assign w2119 = pi2343 & ~w4420;
assign w2120 = pi1492 & w13753;
assign w2121 = pi3008 & w16502;
assign w2122 = pi0020 & ~w3748;
assign w2123 = w7703 & w17764;
assign w2124 = ~w8538 & ~w14657;
assign w2125 = ~pi1296 & ~pi1300;
assign w2126 = ~w7826 & w7515;
assign w2127 = w1497 & w12001;
assign w2128 = (~pi1772 & ~w7799) | (~pi1772 & w1753) | (~w7799 & w1753);
assign w2129 = (pi0900 & ~w13509) | (pi0900 & w5248) | (~w13509 & w5248);
assign w2130 = ~w5843 & ~w15682;
assign w2131 = ~w394 & ~w12465;
assign w2132 = w13509 & w8104;
assign w2133 = ~w5118 & w4493;
assign w2134 = w15622 & ~w11222;
assign w2135 = ~w7102 & ~w17070;
assign w2136 = ~pi3085 & w15235;
assign w2137 = pi1137 & w9420;
assign w2138 = ~pi1136 & w9420;
assign w2139 = ~w15354 & ~w6211;
assign w2140 = w6697 & ~w2776;
assign w2141 = pi0496 & pi1143;
assign w2142 = ~w1911 & ~w1189;
assign w2143 = pi1468 & w13753;
assign w2144 = ~w5882 & ~w4926;
assign w2145 = pi2464 & ~w10299;
assign w2146 = ~w6195 & w2269;
assign w2147 = ~w16506 & pi1186;
assign w2148 = pi1655 & ~w6072;
assign w2149 = ~w10451 & ~w16944;
assign w2150 = ~pi3142 & w13570;
assign w2151 = w5767 & w17559;
assign w2152 = ~w16928 & ~w11485;
assign w2153 = w9440 & pi0172;
assign w2154 = pi2502 & ~w5274;
assign w2155 = w6857 & w2813;
assign w2156 = ~w13623 & ~w5520;
assign w2157 = ~w124 & ~w18415;
assign w2158 = ~w12775 & ~w3705;
assign w2159 = (~pi1764 & ~w7799) | (~pi1764 & w13681) | (~w7799 & w13681);
assign w2160 = pi1337 & pi0307;
assign w2161 = ~pi2178 & w5384;
assign w2162 = ~w8802 & ~w5442;
assign w2163 = pi1769 & ~w5457;
assign w2164 = w13509 & w10549;
assign w2165 = w7195 & w1206;
assign w2166 = ~pi1048 & w15707;
assign w2167 = pi3063 & w16502;
assign w2168 = w10189 & ~pi0451;
assign w2169 = ~w4294 & w5693;
assign w2170 = pi1684 & ~w7177;
assign w2171 = ~pi2375 & w12941;
assign w2172 = ~w11205 & ~w1772;
assign w2173 = w6697 & ~w3430;
assign w2174 = pi1328 & pi1345;
assign w2175 = ~w15321 & ~w2136;
assign w2176 = w12060 & w18190;
assign w2177 = ~w17466 & w11976;
assign w2178 = ~w5189 & pi0722;
assign w2179 = w5261 & w4465;
assign w2180 = w820 & w4626;
assign w2181 = w13509 & w822;
assign w2182 = ~pi3163 & w17669;
assign w2183 = ~w639 & ~w18400;
assign w2184 = pi0120 & pi2758;
assign w2185 = ~pi3165 & w17669;
assign w2186 = ~w2365 & ~w3451;
assign w2187 = (pi0678 & ~w13509) | (pi0678 & w18157) | (~w13509 & w18157);
assign w2188 = ~pi3321 & w14918;
assign w2189 = ~pi1805 & w5531;
assign w2190 = ~w6979 & ~w13989;
assign w2191 = ~w1962 & pi0654;
assign w2192 = ~w3872 & ~w13299;
assign w2193 = pi2921 & ~pi3199;
assign w2194 = w7307 & w3607;
assign w2195 = pi2801 & ~w11406;
assign w2196 = (w12095 & ~w12460) | (w12095 & w227) | (~w12460 & w227);
assign w2197 = pi2648 & ~w3555;
assign w2198 = ~pi2092 & w12724;
assign w2199 = ~w864 & ~w12044;
assign w2200 = ~w15610 & ~w15360;
assign w2201 = ~w4628 & ~w5559;
assign w2202 = w13509 & w2974;
assign w2203 = pi0021 & ~w3748;
assign w2204 = w10305 & w16659;
assign w2205 = w3243 & ~pi0313;
assign w2206 = ~w6760 & w8389;
assign w2207 = ~w16899 & ~w4744;
assign w2208 = w12460 & w1235;
assign w2209 = ~w2421 & ~w14776;
assign w2210 = ~w3778 & ~w13973;
assign w2211 = ~pi0914 & w6200;
assign w2212 = ~pi0511 & ~pi1157;
assign w2213 = ~w13418 & ~w8134;
assign w2214 = w17839 & w16414;
assign w2215 = w13509 & w10611;
assign w2216 = ~w8324 & ~w9265;
assign w2217 = pi2275 & ~w9414;
assign w2218 = w7077 & ~w10235;
assign w2219 = ~pi3117 & ~w18021;
assign w2220 = ~pi3106 & ~w3987;
assign w2221 = ~w1802 & ~w16385;
assign w2222 = w16278 & ~w9852;
assign w2223 = w9720 & pi1722;
assign w2224 = ~w5171 & ~w7980;
assign w2225 = ~w13654 & ~w2106;
assign w2226 = w9720 & pi1754;
assign w2227 = ~w9506 & ~w8240;
assign w2228 = (w13806 & ~w17173) | (w13806 & w16010) | (~w17173 & w16010);
assign w2229 = ~w472 & w4537;
assign w2230 = pi0058 & w922;
assign w2231 = ~w5785 & ~w8103;
assign w2232 = ~w3601 & ~w9929;
assign w2233 = ~pi1067 & w1147;
assign w2234 = ~w9248 & ~w1138;
assign w2235 = w17470 & w4745;
assign w2236 = pi2184 & ~w14524;
assign w2237 = ~w14716 & ~w6154;
assign w2238 = w16729 & w8885;
assign w2239 = w15122 & ~pi2467;
assign w2240 = ~w13041 & w17183;
assign w2241 = pi1539 & w13753;
assign w2242 = pi3065 & w16502;
assign w2243 = w12460 & w11148;
assign w2244 = ~w16386 & w7794;
assign w2245 = w7307 & w11153;
assign w2246 = w7681 & ~w8067;
assign w2247 = pi1984 & w14245;
assign w2248 = ~w5726 & w3098;
assign w2249 = (~w2165 & ~w17173) | (~w2165 & w14970) | (~w17173 & w14970);
assign w2250 = w16506 & pi2959;
assign w2251 = pi2927 & ~w6463;
assign w2252 = w62 & w824;
assign w2253 = w16345 & w4304;
assign w2254 = ~w18015 & ~w3502;
assign w2255 = ~w11280 & ~w1902;
assign w2256 = ~w2725 & pi0796;
assign w2257 = ~w15808 & pi0741;
assign w2258 = w5223 & ~pi1297;
assign w2259 = ~w5732 & w5496;
assign w2260 = ~w6697 & pi0670;
assign w2261 = ~w7910 & ~w7788;
assign w2262 = ~w2778 & ~w3745;
assign w2263 = ~pi2933 & w14648;
assign w2264 = w1391 & ~w10947;
assign w2265 = pi2084 & ~w17683;
assign w2266 = pi2684 & ~w11406;
assign w2267 = ~w5189 & pi0724;
assign w2268 = ~w9467 & w17273;
assign w2269 = ~w14560 & pi0214;
assign w2270 = ~w3357 & ~w175;
assign w2271 = w16278 & ~w14978;
assign w2272 = (pi0781 & ~w13509) | (pi0781 & w10452) | (~w13509 & w10452);
assign w2273 = ~w8349 & ~w5193;
assign w2274 = w16278 & ~w11978;
assign w2275 = (pi1795 & w7215) | (pi1795 & w15186) | (w7215 & w15186);
assign w2276 = pi2922 & w6045;
assign w2277 = ~w61 & w8940;
assign w2278 = ~w8523 & ~w7304;
assign w2279 = ~w17672 & ~w5875;
assign w2280 = pi0059 & pi0060;
assign w2281 = pi1440 & ~w6448;
assign w2282 = w539 & ~w7803;
assign w2283 = ~pi0483 & pi3381;
assign w2284 = pi2226 & ~w11735;
assign w2285 = w13231 & ~w4043;
assign w2286 = w2613 & w13509;
assign w2287 = (pi1025 & ~w13509) | (pi1025 & w5723) | (~w13509 & w5723);
assign w2288 = pi1702 & ~w18497;
assign w2289 = pi2819 & w605;
assign w2290 = w17562 & pi1815;
assign w2291 = w384 & w13339;
assign w2292 = ~pi2967 & pi3069;
assign w2293 = (pi1135 & ~w5437) | (pi1135 & w7542) | (~w5437 & w7542);
assign w2294 = ~w13207 & ~w6714;
assign w2295 = ~w17498 & ~w17912;
assign w2296 = ~w12291 & ~w5572;
assign w2297 = w17562 & pi1851;
assign w2298 = w16575 & w2750;
assign w2299 = ~w5135 & ~w3087;
assign w2300 = ~pi3170 & w4310;
assign w2301 = ~pi3158 & w13730;
assign w2302 = w7703 & w4778;
assign w2303 = ~w2725 & pi0785;
assign w2304 = w13509 & w1081;
assign w2305 = pi3146 & w10389;
assign w2306 = ~w7104 & ~w16284;
assign w2307 = w212 & w10193;
assign w2308 = ~w13892 & ~w7654;
assign w2309 = pi2750 & ~w226;
assign w2310 = ~w900 & w9654;
assign w2311 = pi1631 & ~w13753;
assign w2312 = ~w1859 & ~w15216;
assign w2313 = ~w10484 & ~w4883;
assign w2314 = ~pi1915 & w11313;
assign w2315 = (pi0716 & ~w13509) | (pi0716 & w5336) | (~w13509 & w5336);
assign w2316 = ~w14073 & w11639;
assign w2317 = pi2747 & ~w6463;
assign w2318 = w13321 & ~w16905;
assign w2319 = w7799 & w2290;
assign w2320 = (pi0402 & w5560) | (pi0402 & w13356) | (w5560 & w13356);
assign w2321 = ~pi1262 & pi2955;
assign w2322 = pi3517 & ~w7793;
assign w2323 = pi2982 & ~w3987;
assign w2324 = ~pi2416 & w13204;
assign w2325 = pi1296 & pi1300;
assign w2326 = w2971 & w9639;
assign w2327 = ~w15808 & pi0917;
assign w2328 = ~pi3147 & pi3168;
assign w2329 = w16506 & ~w3374;
assign w2330 = ~pi3045 & w226;
assign w2331 = ~pi2365 & w12941;
assign w2332 = w2341 & ~w305;
assign w2333 = ~pi3164 & w14753;
assign w2334 = ~pi1189 & w6200;
assign w2335 = w15122 & ~pi2500;
assign w2336 = pi1702 & w4683;
assign w2337 = pi3168 & w3987;
assign w2338 = ~w16325 & ~w13111;
assign w2339 = ~w15862 & ~w6766;
assign w2340 = w384 & w3726;
assign w2341 = w3988 & w6676;
assign w2342 = (pi0827 & ~w13509) | (pi0827 & w12613) | (~w13509 & w12613);
assign w2343 = ~w2266 & ~w12898;
assign w2344 = ~w12040 & pi1016;
assign w2345 = ~w2411 & w7858;
assign w2346 = ~w17372 & ~w1282;
assign w2347 = w17683 & w614;
assign w2348 = ~w6785 & pi0872;
assign w2349 = ~w6300 & ~w13024;
assign w2350 = ~w6550 & ~w5440;
assign w2351 = ~w13815 & ~w10017;
assign w2352 = (pi0735 & ~w13509) | (pi0735 & w8005) | (~w13509 & w8005);
assign w2353 = pi0048 & ~w14148;
assign w2354 = w16965 & ~pi3064;
assign w2355 = pi1663 & w1924;
assign w2356 = ~w5189 & pi0726;
assign w2357 = w14228 & ~w6680;
assign w2358 = pi2535 & w14148;
assign w2359 = ~w10362 & w16451;
assign w2360 = pi1337 & ~pi0248;
assign w2361 = pi1337 & pi0249;
assign w2362 = w16575 & w13377;
assign w2363 = pi2981 & ~pi2982;
assign w2364 = (~pi0327 & ~w6857) | (~pi0327 & w6923) | (~w6857 & w6923);
assign w2365 = pi2505 & ~w5274;
assign w2366 = ~pi3171 & w8515;
assign w2367 = ~w8897 & ~w2265;
assign w2368 = ~pi3028 & pi3157;
assign w2369 = pi2845 & w605;
assign w2370 = ~pi3164 & w4310;
assign w2371 = ~w8816 & w14097;
assign w2372 = ~w6846 & w15858;
assign w2373 = ~w9464 & ~w16233;
assign w2374 = ~w12847 & ~w2553;
assign w2375 = w13509 & w15829;
assign w2376 = ~w12040 & pi0683;
assign w2377 = ~w10681 & ~w15921;
assign w2378 = w14094 & w7245;
assign w2379 = ~pi0686 & w9110;
assign w2380 = ~pi1778 & w8383;
assign w2381 = (pi0635 & ~w13509) | (pi0635 & w2849) | (~w13509 & w2849);
assign w2382 = pi3158 & w18281;
assign w2383 = ~pi0291 & w4058;
assign w2384 = ~w1116 & ~w11099;
assign w2385 = w10818 & ~w12320;
assign w2386 = w7077 & ~w14597;
assign w2387 = pi0420 & w17173;
assign w2388 = (pi0305 & ~w325) | (pi0305 & w9622) | (~w325 & w9622);
assign w2389 = w6697 & ~w14597;
assign w2390 = w11320 & ~w7507;
assign w2391 = ~w6439 & ~w8734;
assign w2392 = ~pi3141 & ~pi3160;
assign w2393 = ~w9021 & w8565;
assign w2394 = ~w13231 & pi0991;
assign w2395 = w13509 & w9174;
assign w2396 = ~w10342 & ~w505;
assign w2397 = ~pi2355 & w17439;
assign w2398 = ~w12355 & ~w5322;
assign w2399 = ~pi3311 & w6448;
assign w2400 = ~w4708 & ~w3222;
assign w2401 = w13509 & w491;
assign w2402 = w10299 & w9407;
assign w2403 = ~pi3163 & w1843;
assign w2404 = ~pi1963 & w11688;
assign w2405 = ~pi0284 & w2196;
assign w2406 = w18256 & w4864;
assign w2407 = ~w8842 & ~w17233;
assign w2408 = ~w15945 & ~w2454;
assign w2409 = ~w14905 & ~w13125;
assign w2410 = ~w6493 & ~w4049;
assign w2411 = ~w14341 & ~w10635;
assign w2412 = ~pi0606 & w12825;
assign w2413 = pi1864 & ~w15036;
assign w2414 = ~w6 & ~w1729;
assign w2415 = ~w16230 & ~pi3117;
assign w2416 = ~pi3095 & w11406;
assign w2417 = ~pi2048 & w13204;
assign w2418 = (pi1076 & ~w13509) | (pi1076 & w9822) | (~w13509 & w9822);
assign w2419 = (~pi0974 & ~w13509) | (~pi0974 & w12168) | (~w13509 & w12168);
assign w2420 = w2647 & w4401;
assign w2421 = (pi0577 & ~w13509) | (pi0577 & w3370) | (~w13509 & w3370);
assign w2422 = w11383 & w10194;
assign w2423 = pi2917 & w6045;
assign w2424 = w18437 & w12719;
assign w2425 = ~w7681 & ~w8067;
assign w2426 = ~w9991 & w5810;
assign w2427 = ~w18451 & ~w8368;
assign w2428 = ~pi3419 & w15036;
assign w2429 = ~pi0516 & w15707;
assign w2430 = w2725 & ~w7449;
assign w2431 = pi1218 & w13430;
assign w2432 = ~w17042 & ~w1148;
assign w2433 = pi1465 & w13753;
assign w2434 = pi1545 & w13753;
assign w2435 = (pi0807 & ~w13509) | (pi0807 & w3675) | (~w13509 & w3675);
assign w2436 = ~w2479 & ~w14025;
assign w2437 = pi1655 & ~w13753;
assign w2438 = ~w1402 & ~w5840;
assign w2439 = ~w4175 & ~w7310;
assign w2440 = ~pi3288 & w6448;
assign w2441 = w8383 & pi0065;
assign w2442 = ~w16575 & w18517;
assign w2443 = ~pi0941 & w9110;
assign w2444 = w13329 & pi0486;
assign w2445 = ~w8126 & w13128;
assign w2446 = ~w3417 & ~w2442;
assign w2447 = ~w6402 & ~w645;
assign w2448 = ~w5189 & pi0728;
assign w2449 = w17741 & w12930;
assign w2450 = ~pi3153 & w11701;
assign w2451 = w13509 & w1334;
assign w2452 = ~w2835 & ~w8509;
assign w2453 = ~w11043 & ~w1432;
assign w2454 = w11383 & w6924;
assign w2455 = pi1421 & ~w6072;
assign w2456 = w4415 & w17493;
assign w2457 = w13509 & w5120;
assign w2458 = w5190 & pi3066;
assign w2459 = ~pi3341 & w14918;
assign w2460 = ~pi0896 & ~w8789;
assign w2461 = w13509 & w5610;
assign w2462 = pi1739 & ~w4058;
assign w2463 = w5437 & w17027;
assign w2464 = ~pi3012 & ~pi3207;
assign w2465 = ~w15330 & ~w14638;
assign w2466 = w15565 & w11843;
assign w2467 = w11735 & w17115;
assign w2468 = pi3166 & w13786;
assign w2469 = pi3207 & ~w2219;
assign w2470 = ~pi2148 & w13065;
assign w2471 = ~w15808 & pi0747;
assign w2472 = w13509 & w11370;
assign w2473 = ~pi3286 & w17935;
assign w2474 = ~w14474 & ~w15578;
assign w2475 = ~w2341 & ~pi0965;
assign w2476 = ~w3643 & ~w5378;
assign w2477 = pi1797 & pi3158;
assign w2478 = w13509 & w12467;
assign w2479 = ~pi2307 & w16041;
assign w2480 = ~w14507 & ~w3450;
assign w2481 = ~pi1881 & w17213;
assign w2482 = ~w1536 & ~w749;
assign w2483 = pi2913 & ~w16095;
assign w2484 = ~pi0857 & w15707;
assign w2485 = (pi0611 & ~w13509) | (pi0611 & w14362) | (~w13509 & w14362);
assign w2486 = pi3163 & w2848;
assign w2487 = w7307 & w13009;
assign w2488 = ~w14228 & pi1006;
assign w2489 = ~w9503 & ~w16562;
assign w2490 = ~pi0501 & ~pi1345;
assign w2491 = w14998 & w14202;
assign w2492 = pi1633 & ~w18259;
assign w2493 = ~w17638 & ~w5927;
assign w2494 = w10136 & w6997;
assign w2495 = w1368 & pi0383;
assign w2496 = ~w15656 & ~w13637;
assign w2497 = ~w11298 & ~w15357;
assign w2498 = w13509 & w4044;
assign w2499 = ~pi1983 & ~w15450;
assign w2500 = ~pi3315 & w17935;
assign w2501 = ~w918 & w14755;
assign w2502 = ~w13574 & ~w17341;
assign w2503 = (pi0850 & ~w13509) | (pi0850 & w13213) | (~w13509 & w13213);
assign w2504 = ~w9037 & ~w6344;
assign w2505 = ~w2984 & ~w16101;
assign w2506 = w7307 & w11498;
assign w2507 = ~w11344 & ~w15303;
assign w2508 = ~pi1765 & ~pi3155;
assign w2509 = w4420 & w2753;
assign w2510 = pi1283 & pi1345;
assign w2511 = (pi1807 & w5453) | (pi1807 & w9642) | (w5453 & w9642);
assign w2512 = ~w152 & ~w7995;
assign w2513 = pi1754 & ~pi3162;
assign w2514 = w3203 & ~w10235;
assign w2515 = w13509 & w13031;
assign w2516 = pi3153 & w2253;
assign w2517 = ~pi3326 & w17935;
assign w2518 = ~w13696 & ~w18253;
assign w2519 = ~pi1096 & w11739;
assign w2520 = pi2965 & ~w3987;
assign w2521 = ~w2341 & pi0830;
assign w2522 = w11383 & w16199;
assign w2523 = (~pi1801 & ~w7799) | (~pi1801 & w5283) | (~w7799 & w5283);
assign w2524 = ~w9357 & ~w3065;
assign w2525 = ~w3875 & ~w8133;
assign w2526 = ~pi3311 & w14918;
assign w2527 = ~w15316 & ~w8398;
assign w2528 = ~w5939 & w5869;
assign w2529 = pi3158 & w7705;
assign w2530 = ~pi3142 & w12427;
assign w2531 = w5453 & w8303;
assign w2532 = ~w11594 & ~w13517;
assign w2533 = ~pi1713 & ~pi3134;
assign w2534 = pi1506 & ~w16922;
assign w2535 = ~pi3328 & w9781;
assign w2536 = ~pi1232 & w5019;
assign w2537 = pi0503 & pi1155;
assign w2538 = pi2069 & ~w4508;
assign w2539 = ~w10767 & ~w8623;
assign w2540 = (pi0823 & ~w13509) | (pi0823 & w9732) | (~w13509 & w9732);
assign w2541 = ~pi1958 & w11688;
assign w2542 = pi0508 & pi1146;
assign w2543 = ~w5189 & pi0730;
assign w2544 = w6226 & w15351;
assign w2545 = ~pi3146 & w15839;
assign w2546 = ~w17329 & ~w6268;
assign w2547 = pi0496 & pi0497;
assign w2548 = ~w11427 & ~w2402;
assign w2549 = w13399 & w3616;
assign w2550 = pi1387 & w13753;
assign w2551 = pi0513 & pi1144;
assign w2552 = pi1794 & ~w9520;
assign w2553 = pi3160 & ~pi3491;
assign w2554 = pi1516 & w13753;
assign w2555 = ~w6956 & w7196;
assign w2556 = ~pi3146 & w17993;
assign w2557 = w2341 & ~w1340;
assign w2558 = ~pi1187 & w9420;
assign w2559 = ~w11247 & w3909;
assign w2560 = w2826 & w182;
assign w2561 = ~w7901 & ~w6301;
assign w2562 = w10818 & ~w9293;
assign w2563 = pi2702 & ~w16815;
assign w2564 = ~pi0956 & w12825;
assign w2565 = ~w5109 & ~w16287;
assign w2566 = w934 & pi0414;
assign w2567 = ~pi0074 & w922;
assign w2568 = pi1787 & ~w9459;
assign w2569 = pi1565 & ~w18259;
assign w2570 = w14460 & w1421;
assign w2571 = w12460 & w8281;
assign w2572 = ~pi2225 & w11313;
assign w2573 = ~pi0703 & w3106;
assign w2574 = ~pi0724 & w17899;
assign w2575 = w16506 & w5196;
assign w2576 = ~pi3086 & w261;
assign w2577 = pi1507 & ~w16922;
assign w2578 = ~w7152 & ~w18312;
assign w2579 = w17388 & w4273;
assign w2580 = ~w2170 & ~w18129;
assign w2581 = (pi0670 & ~w13509) | (pi0670 & w2260) | (~w13509 & w2260);
assign w2582 = w13509 & w17512;
assign w2583 = w12040 & ~w2776;
assign w2584 = ~w14150 & ~w7827;
assign w2585 = ~pi3045 & w261;
assign w2586 = ~w16141 & ~w9970;
assign w2587 = ~w17059 & ~w2490;
assign w2588 = (pi0763 & ~w13509) | (pi0763 & w6205) | (~w13509 & w6205);
assign w2589 = ~w3983 & ~w18272;
assign w2590 = pi1961 & ~w14833;
assign w2591 = ~w518 & ~w12616;
assign w2592 = ~pi2913 & w5292;
assign w2593 = pi1788 & ~w15767;
assign w2594 = ~w5080 & ~w7111;
assign w2595 = ~w15856 & ~w2145;
assign w2596 = w13509 & w2624;
assign w2597 = pi3136 & w13108;
assign w2598 = pi2395 & ~w18123;
assign w2599 = w16700 & w17991;
assign w2600 = w12040 & w15609;
assign w2601 = pi0988 & pi2465;
assign w2602 = (pi0873 & ~w13509) | (pi0873 & w1700) | (~w13509 & w1700);
assign w2603 = pi3078 & ~w16502;
assign w2604 = w5189 & ~w15296;
assign w2605 = w12583 & ~w778;
assign w2606 = ~w13231 & pi0569;
assign w2607 = ~w9462 & w4522;
assign w2608 = ~pi3158 & w15839;
assign w2609 = ~w4950 & ~w13074;
assign w2610 = ~w2302 & ~w1765;
assign w2611 = (w15842 & ~w384) | (w15842 & w9047) | (~w384 & w9047);
assign w2612 = ~w5288 & ~w11738;
assign w2613 = pi1152 & pi1154;
assign w2614 = w2341 & ~w14465;
assign w2615 = ~pi3160 & ~pi3169;
assign w2616 = ~w6195 & w8419;
assign w2617 = pi2865 & w14148;
assign w2618 = ~pi0329 & w2196;
assign w2619 = ~pi2102 & w12724;
assign w2620 = ~w1368 & ~pi0460;
assign w2621 = (w11186 & ~w1557) | (w11186 & w5299) | (~w1557 & w5299);
assign w2622 = w540 & w12874;
assign w2623 = (~pi0511 & w17577) | (~pi0511 & w13113) | (w17577 & w13113);
assign w2624 = w7077 & w1217;
assign w2625 = ~w3312 & ~w6435;
assign w2626 = w10823 & w11997;
assign w2627 = ~w3997 & ~w1723;
assign w2628 = pi2389 & ~w412;
assign w2629 = pi2411 & ~w17646;
assign w2630 = ~w18066 & ~w17092;
assign w2631 = pi1946 & ~w17646;
assign w2632 = pi2967 & ~w9284;
assign w2633 = w1127 & ~w7916;
assign w2634 = ~w5189 & pi0732;
assign w2635 = w1368 & pi0400;
assign w2636 = ~w10181 & ~w13202;
assign w2637 = w10721 & w1220;
assign w2638 = pi0011 & ~w3748;
assign w2639 = ~w16278 & ~pi0967;
assign w2640 = pi2923 & ~w2276;
assign w2641 = (pi1162 & w14073) | (pi1162 & w16137) | (w14073 & w16137);
assign w2642 = w13509 & w14831;
assign w2643 = ~w15808 & pi1034;
assign w2644 = ~w12836 & ~w3634;
assign w2645 = pi0178 & ~pi0190;
assign w2646 = w11383 & w16419;
assign w2647 = w10178 & w223;
assign w2648 = ~w10324 & w8101;
assign w2649 = w17741 & w9167;
assign w2650 = (~pi1766 & ~w7799) | (~pi1766 & w3399) | (~w7799 & w3399);
assign w2651 = ~w17717 & w7891;
assign w2652 = ~w1391 & pi1075;
assign w2653 = ~w8489 & ~w15878;
assign w2654 = w16575 & w2663;
assign w2655 = ~w8329 & ~w365;
assign w2656 = ~w8588 & w15271;
assign w2657 = (pi0624 & ~w13509) | (pi0624 & w7480) | (~w13509 & w7480);
assign w2658 = w13231 & ~w305;
assign w2659 = ~pi3048 & w15235;
assign w2660 = pi3147 & w10389;
assign w2661 = w14442 & w4186;
assign w2662 = pi1554 & ~w13753;
assign w2663 = w10189 & ~pi0481;
assign w2664 = ~w8963 & ~w16025;
assign w2665 = (w5517 & w235) | (w5517 & w11695) | (w235 & w11695);
assign w2666 = ~w7541 & w817;
assign w2667 = (pi0546 & ~w13509) | (pi0546 & w10938) | (~w13509 & w10938);
assign w2668 = pi2811 & ~w6463;
assign w2669 = ~w1791 & w10536;
assign w2670 = ~w8429 & ~w14904;
assign w2671 = ~pi2303 & w5075;
assign w2672 = ~w4667 & ~w18209;
assign w2673 = ~w12658 & w5814;
assign w2674 = ~pi2456 & w5384;
assign w2675 = ~pi2197 & w9340;
assign w2676 = ~w6669 & ~w3185;
assign w2677 = pi3150 & w8113;
assign w2678 = pi1214 & w5566;
assign w2679 = ~w330 & ~w18054;
assign w2680 = ~pi2797 & w17213;
assign w2681 = ~w3130 & ~w468;
assign w2682 = w8658 & pi1781;
assign w2683 = ~w6993 & ~w6046;
assign w2684 = pi0498 & pi0513;
assign w2685 = (pi0353 & w6195) | (pi0353 & w7117) | (w6195 & w7117);
assign w2686 = ~w13726 & ~w5278;
assign w2687 = ~pi3143 & pi3207;
assign w2688 = pi1490 & ~w9781;
assign w2689 = pi2731 & ~w261;
assign w2690 = pi0063 & w922;
assign w2691 = ~w4689 & ~w5519;
assign w2692 = pi2235 & ~w11735;
assign w2693 = ~pi3321 & w6072;
assign w2694 = w2725 & ~w7020;
assign w2695 = w14279 & w17045;
assign w2696 = ~w16278 & pi0717;
assign w2697 = w2626 & w16351;
assign w2698 = ~w13907 & ~w12986;
assign w2699 = (pi0385 & w5560) | (pi0385 & w13160) | (w5560 & w13160);
assign w2700 = pi1887 & ~w458;
assign w2701 = pi1659 & ~w13753;
assign w2702 = w17584 & w5228;
assign w2703 = pi1383 & ~w5043;
assign w2704 = ~w18418 & ~w5716;
assign w2705 = w7077 & ~w12800;
assign w2706 = ~pi3145 & ~pi3160;
assign w2707 = w13509 & w8334;
assign w2708 = ~w5866 & ~w5326;
assign w2709 = pi3168 & w10389;
assign w2710 = ~pi3171 & w13730;
assign w2711 = ~pi1174 & w1126;
assign w2712 = ~w5189 & pi0734;
assign w2713 = ~w247 & ~w8331;
assign w2714 = ~w14648 & ~pi2603;
assign w2715 = pi1790 & ~w18334;
assign w2716 = ~w10274 & ~w6310;
assign w2717 = ~w682 & ~w13740;
assign w2718 = ~w9494 & ~w311;
assign w2719 = ~w10079 & ~w14675;
assign w2720 = ~pi2140 & w12941;
assign w2721 = ~pi1201 & w3791;
assign w2722 = ~w18591 & ~w14015;
assign w2723 = w5275 & w4662;
assign w2724 = w9440 & pi0145;
assign w2725 = w2613 & w13679;
assign w2726 = pi0206 & ~pi0207;
assign w2727 = ~pi1992 & w3019;
assign w2728 = ~w1368 & ~pi0466;
assign w2729 = ~w7668 & ~w8497;
assign w2730 = pi2458 & ~w14524;
assign w2731 = ~pi0544 & w11739;
assign w2732 = w1611 & w17016;
assign w2733 = ~pi0590 & w795;
assign w2734 = pi3164 & w14951;
assign w2735 = (pi0820 & ~w13509) | (pi0820 & w5730) | (~w13509 & w5730);
assign w2736 = w1215 & w11991;
assign w2737 = ~pi3025 & ~pi3207;
assign w2738 = w384 & w16177;
assign w2739 = w16278 & ~w2776;
assign w2740 = (pi1193 & ~w5437) | (pi1193 & w8559) | (~w5437 & w8559);
assign w2741 = ~w3735 & ~w6886;
assign w2742 = (w2460 & ~w4084) | (w2460 & w1120) | (~w4084 & w1120);
assign w2743 = ~pi3340 & w7090;
assign w2744 = ~w1634 & w1127;
assign w2745 = w12460 & w11389;
assign w2746 = ~w16515 & ~w6925;
assign w2747 = ~w1237 & ~w16112;
assign w2748 = ~w17577 & w6095;
assign w2749 = ~pi3337 & w9781;
assign w2750 = w10189 & ~pi0462;
assign w2751 = ~w9714 & ~w3471;
assign w2752 = pi1232 & pi3027;
assign w2753 = ~pi3168 & ~w4020;
assign w2754 = ~pi3154 & w11701;
assign w2755 = pi1175 & w13509;
assign w2756 = ~pi3142 & w8515;
assign w2757 = pi2966 & pi2576;
assign w2758 = pi0024 & ~w14148;
assign w2759 = ~pi3138 & pi3207;
assign w2760 = ~w12040 & pi0690;
assign w2761 = pi2889 & ~w5274;
assign w2762 = ~pi2233 & w2151;
assign w2763 = ~w7648 & ~w10427;
assign w2764 = ~w17948 & ~w2368;
assign w2765 = ~w6697 & pi0667;
assign w2766 = ~w198 & ~w15239;
assign w2767 = w9318 & w562;
assign w2768 = ~w15233 & ~w9405;
assign w2769 = ~w14738 & w13563;
assign w2770 = ~w1907 & ~w1555;
assign w2771 = ~pi1725 & w5914;
assign w2772 = ~w1614 & ~w15512;
assign w2773 = ~pi3056 & w16815;
assign w2774 = ~w15640 & w16398;
assign w2775 = pi1669 & ~w4058;
assign w2776 = ~w12377 & ~w15211;
assign w2777 = w13509 & w14826;
assign w2778 = pi1361 & ~w4256;
assign w2779 = pi2843 & w605;
assign w2780 = ~w7656 & pi1213;
assign w2781 = (~w16158 & ~w14073) | (~w16158 & w16065) | (~w14073 & w16065);
assign w2782 = (pi1894 & w2014) | (pi1894 & w13285) | (w2014 & w13285);
assign w2783 = ~w14655 & ~w11947;
assign w2784 = ~pi1922 & w9340;
assign w2785 = pi0252 & w5113;
assign w2786 = w1500 & w14814;
assign w2787 = pi1552 & ~w17935;
assign w2788 = w13686 & w3521;
assign w2789 = ~w15335 & w14562;
assign w2790 = pi3080 & ~w16502;
assign w2791 = ~pi3171 & w11701;
assign w2792 = pi2954 & ~pi3199;
assign w2793 = w7703 & w12630;
assign w2794 = ~pi2807 & w13343;
assign w2795 = pi1800 & ~w10389;
assign w2796 = ~w11922 & ~w16395;
assign w2797 = ~pi1173 & w12197;
assign w2798 = w13509 & w15783;
assign w2799 = w5189 & w1217;
assign w2800 = w13509 & w2705;
assign w2801 = ~w16864 & w2744;
assign w2802 = (pi0761 & ~w13509) | (pi0761 & w85) | (~w13509 & w85);
assign w2803 = ~w13142 & w7166;
assign w2804 = pi2966 & pi2592;
assign w2805 = ~pi1192 & w9420;
assign w2806 = ~w1730 & ~w5260;
assign w2807 = pi3139 & w8829;
assign w2808 = w15808 & ~w10947;
assign w2809 = w3089 & w3933;
assign w2810 = ~w5812 & ~w6425;
assign w2811 = ~w5812 & ~w6426;
assign w2812 = pi2445 & ~w14524;
assign w2813 = w934 & pi0433;
assign w2814 = ~pi3154 & w17669;
assign w2815 = pi3155 & w619;
assign w2816 = ~w6119 & ~w16992;
assign w2817 = ~pi0763 & w6200;
assign w2818 = ~w16278 & pi0702;
assign w2819 = w11345 & w12096;
assign w2820 = ~w16667 & ~w5931;
assign w2821 = pi1600 & w13753;
assign w2822 = ~pi3155 & w4310;
assign w2823 = ~w9306 & ~w2171;
assign w2824 = ~w5189 & pi0736;
assign w2825 = pi0097 & w3748;
assign w2826 = w2742 & ~w4985;
assign w2827 = ~pi3290 & w17935;
assign w2828 = pi2214 & ~w11735;
assign w2829 = w291 & ~w15553;
assign w2830 = pi1860 & ~w15036;
assign w2831 = w15808 & ~w6033;
assign w2832 = w17562 & pi1823;
assign w2833 = ~w6358 & ~w14732;
assign w2834 = ~w12203 & w2051;
assign w2835 = pi0026 & ~w14148;
assign w2836 = ~w1754 & ~w9930;
assign w2837 = ~w13345 & ~w8278;
assign w2838 = ~pi3155 & w13570;
assign w2839 = w659 & w14116;
assign w2840 = ~pi3056 & w226;
assign w2841 = ~w1791 & w17123;
assign w2842 = ~w4314 & ~w14659;
assign w2843 = ~pi0816 & w1147;
assign w2844 = ~w12271 & ~w9040;
assign w2845 = ~w7236 & ~w10582;
assign w2846 = ~w3332 & ~w17336;
assign w2847 = pi2728 & ~w261;
assign w2848 = w10352 & w876;
assign w2849 = ~w1962 & pi0635;
assign w2850 = ~w18101 & ~w18243;
assign w2851 = ~w3000 & ~pi2799;
assign w2852 = ~w7077 & pi0809;
assign w2853 = w18530 & w1355;
assign w2854 = ~w14221 & ~w508;
assign w2855 = (pi0597 & ~w13509) | (pi0597 & w16260) | (~w13509 & w16260);
assign w2856 = ~w297 & ~w9180;
assign w2857 = ~w8084 & ~w1535;
assign w2858 = ~w6785 & pi0987;
assign w2859 = pi2022 & ~w17646;
assign w2860 = pi3163 & w3987;
assign w2861 = pi1337 & ~pi0271;
assign w2862 = pi0311 & ~w13184;
assign w2863 = ~w10936 & w15673;
assign w2864 = ~pi2988 & w6463;
assign w2865 = pi3172 & w8113;
assign w2866 = (pi1868 & w2014) | (pi1868 & w12991) | (w2014 & w12991);
assign w2867 = w2299 & w7999;
assign w2868 = ~w3603 & ~w7997;
assign w2869 = w539 & ~w8360;
assign w2870 = ~w14821 & ~w18090;
assign w2871 = ~w14541 & w16874;
assign w2872 = ~w9482 & ~w14849;
assign w2873 = pi0040 & pi0042;
assign w2874 = ~w5521 & w4994;
assign w2875 = ~w18275 & w15798;
assign w2876 = ~w15147 & ~w10453;
assign w2877 = ~pi0957 & w14641;
assign w2878 = w7698 & w9720;
assign w2879 = ~w2506 & ~w1865;
assign w2880 = ~w14705 & w18420;
assign w2881 = w13509 & w15980;
assign w2882 = ~pi0787 & w543;
assign w2883 = pi3031 & ~w16502;
assign w2884 = w16506 & ~w13195;
assign w2885 = ~w11279 & w3897;
assign w2886 = pi3148 & ~pi3191;
assign w2887 = pi3158 & w8113;
assign w2888 = w14648 & ~pi2748;
assign w2889 = w11383 & w8633;
assign w2890 = pi1642 & ~w13753;
assign w2891 = ~pi3120 & ~pi3160;
assign w2892 = pi0258 & pi0271;
assign w2893 = ~pi0380 & ~w6057;
assign w2894 = ~pi3057 & w16502;
assign w2895 = ~pi3131 & w4310;
assign w2896 = ~pi1023 & w3106;
assign w2897 = ~w13605 & w7189;
assign w2898 = w13509 & w15267;
assign w2899 = ~pi1045 & w93;
assign w2900 = w12205 & w16340;
assign w2901 = ~pi0124 & w9284;
assign w2902 = ~w3769 & w10183;
assign w2903 = (~pi0485 & w17577) | (~pi0485 & w5839) | (w17577 & w5839);
assign w2904 = ~w1822 & w9613;
assign w2905 = w5031 & pi1233;
assign w2906 = ~w15122 & ~pi2514;
assign w2907 = ~pi0330 & w2196;
assign w2908 = ~pi2975 & w14833;
assign w2909 = w11247 & w18238;
assign w2910 = w7307 & w346;
assign w2911 = ~pi3139 & w15839;
assign w2912 = (~pi0250 & ~w325) | (~pi0250 & w13400) | (~w325 & w13400);
assign w2913 = (pi0251 & ~w325) | (pi0251 & w13401) | (~w325 & w13401);
assign w2914 = ~pi3321 & w18259;
assign w2915 = (pi0363 & w6195) | (pi0363 & w467) | (w6195 & w467);
assign w2916 = pi0416 & w17173;
assign w2917 = ~pi0415 & w17173;
assign w2918 = ~w3075 & ~w16952;
assign w2919 = ~w14360 & ~w17395;
assign w2920 = w14460 & pi0042;
assign w2921 = (w8324 & ~w1766) | (w8324 & w9093) | (~w1766 & w9093);
assign w2922 = ~w13335 & ~w3320;
assign w2923 = pi1893 & ~w15036;
assign w2924 = ~w14731 & ~w15311;
assign w2925 = pi1348 & ~w14148;
assign w2926 = ~w9652 & ~w6149;
assign w2927 = w4420 & w3515;
assign w2928 = w13509 & w6700;
assign w2929 = ~pi3042 & pi3227;
assign w2930 = ~pi2299 & w8617;
assign w2931 = ~w4227 & ~w14698;
assign w2932 = w14228 & ~w13195;
assign w2933 = (pi0765 & ~w13509) | (pi0765 & w1998) | (~w13509 & w1998);
assign w2934 = ~pi3091 & w6463;
assign w2935 = ~w792 & ~w6921;
assign w2936 = w9440 & pi0177;
assign w2937 = w2725 & ~w2741;
assign w2938 = w3203 & ~w2776;
assign w2939 = ~w17389 & ~w6724;
assign w2940 = ~pi3049 & w11406;
assign w2941 = ~w8482 & w8123;
assign w2942 = w13509 & w6770;
assign w2943 = pi1400 & w4683;
assign w2944 = ~pi3157 & w17387;
assign w2945 = (~pi1240 & w11655) | (~pi1240 & w339) | (w11655 & w339);
assign w2946 = ~w16043 & ~w12116;
assign w2947 = pi2725 & ~w16815;
assign w2948 = ~w16750 & ~w15284;
assign w2949 = ~pi0680 & w9110;
assign w2950 = w2341 & ~w14597;
assign w2951 = ~w16506 & pi1139;
assign w2952 = pi2491 & ~w3555;
assign w2953 = w10189 & pi0395;
assign w2954 = ~pi0173 & pi0179;
assign w2955 = w5437 & w3323;
assign w2956 = pi1250 & ~w11655;
assign w2957 = pi3082 & w226;
assign w2958 = pi2765 & w14148;
assign w2959 = ~pi1852 & ~w4084;
assign w2960 = ~w6314 & ~w12236;
assign w2961 = (pi1893 & w2014) | (pi1893 & w6404) | (w2014 & w6404);
assign w2962 = ~w7504 & w12650;
assign w2963 = pi1363 & ~w11608;
assign w2964 = ~w13718 & ~w15348;
assign w2965 = ~pi2116 & w12755;
assign w2966 = pi2001 & ~w9414;
assign w2967 = ~w7218 & ~w982;
assign w2968 = ~w9324 & ~w9352;
assign w2969 = w16950 & w1416;
assign w2970 = ~pi3011 & ~pi3207;
assign w2971 = w15612 & w10676;
assign w2972 = ~pi1940 & w17439;
assign w2973 = w1225 & w14403;
assign w2974 = w7844 & ~w2587;
assign w2975 = w539 & ~w6729;
assign w2976 = ~pi1245 & w11655;
assign w2977 = ~w5350 & ~w7919;
assign w2978 = ~w17326 & ~pi0488;
assign w2979 = (pi0650 & ~w13509) | (pi0650 & w5179) | (~w13509 & w5179);
assign w2980 = w7489 & w4325;
assign w2981 = ~w14648 & ~pi2650;
assign w2982 = pi2336 & ~w412;
assign w2983 = ~w709 & ~pi1289;
assign w2984 = ~pi2101 & w12724;
assign w2985 = pi1408 & ~w5043;
assign w2986 = ~w6699 & w7906;
assign w2987 = ~w2159 & w17167;
assign w2988 = w5437 & w12335;
assign w2989 = (pi1094 & ~w13509) | (pi1094 & w3823) | (~w13509 & w3823);
assign w2990 = (pi1200 & ~w13509) | (pi1200 & w5509) | (~w13509 & w5509);
assign w2991 = ~w12567 & w14162;
assign w2992 = ~w9488 & w8541;
assign w2993 = ~pi1228 & ~pi3365;
assign w2994 = pi1626 & ~w13753;
assign w2995 = w13509 & w6994;
assign w2996 = ~pi2447 & w9340;
assign w2997 = pi2808 & ~w6463;
assign w2998 = ~w5406 & ~w1400;
assign w2999 = pi2505 & w384;
assign w3000 = ~w4295 & ~w9274;
assign w3001 = ~w17641 & ~w279;
assign w3002 = ~w16807 & w3543;
assign w3003 = w12161 & w890;
assign w3004 = ~pi2776 & w17213;
assign w3005 = ~w1791 & w18294;
assign w3006 = (pi1195 & ~w11010) | (pi1195 & w4086) | (~w11010 & w4086);
assign w3007 = pi0300 & w5113;
assign w3008 = ~w577 & ~w8525;
assign w3009 = pi0489 & pi1136;
assign w3010 = pi3143 & w8829;
assign w3011 = w7703 & w18531;
assign w3012 = pi3133 & w5457;
assign w3013 = ~w10874 & ~w16625;
assign w3014 = ~w16200 & ~w13772;
assign w3015 = ~w6195 & w11188;
assign w3016 = ~w7798 & ~w2988;
assign w3017 = ~pi0109 & w3748;
assign w3018 = (pi0636 & ~w13509) | (pi0636 & w6744) | (~w13509 & w6744);
assign w3019 = w13807 & w2425;
assign w3020 = w18377 & w10182;
assign w3021 = (~pi0085 & ~w9786) | (~pi0085 & w6532) | (~w9786 & w6532);
assign w3022 = ~w8946 & ~w6795;
assign w3023 = ~w5968 & ~pi1692;
assign w3024 = w4140 & w16318;
assign w3025 = ~w17696 & ~w7303;
assign w3026 = pi2995 & pi1595;
assign w3027 = ~pi0493 & ~pi1345;
assign w3028 = ~w9612 & ~w12969;
assign w3029 = ~w6878 & w15817;
assign w3030 = ~w8976 & ~w975;
assign w3031 = ~pi3052 & w15235;
assign w3032 = ~w12579 & ~w11647;
assign w3033 = w11383 & w8463;
assign w3034 = ~pi3159 & w15048;
assign w3035 = pi1404 & w4683;
assign w3036 = ~w7844 & ~pi0956;
assign w3037 = ~w15692 & ~w8543;
assign w3038 = pi1718 & ~w619;
assign w3039 = pi3166 & w3987;
assign w3040 = (~pi0966 & ~w13509) | (~pi0966 & w17257) | (~w13509 & w17257);
assign w3041 = w11383 & w5319;
assign w3042 = ~w15122 & ~pi2750;
assign w3043 = pi3018 & ~pi3102;
assign w3044 = pi2604 & ~w3555;
assign w3045 = ~w5036 & ~w6040;
assign w3046 = ~w15864 & ~w219;
assign w3047 = w5217 & ~w3409;
assign w3048 = ~pi0502 & pi1378;
assign w3049 = w5113 & w14503;
assign w3050 = (~pi0272 & ~w325) | (~pi0272 & w16635) | (~w325 & w16635);
assign w3051 = w3223 & w14078;
assign w3052 = w14228 & ~w14143;
assign w3053 = pi2841 & w14148;
assign w3054 = ~w18553 & ~w5386;
assign w3055 = w11924 & w13475;
assign w3056 = ~pi3089 & w226;
assign w3057 = ~pi0791 & w543;
assign w3058 = (pi0783 & ~w13509) | (pi0783 & w11602) | (~w13509 & w11602);
assign w3059 = ~pi1052 & w17490;
assign w3060 = w16672 & w13928;
assign w3061 = ~w14228 & pi0621;
assign w3062 = ~w6364 & ~w16786;
assign w3063 = w15122 & ~pi2595;
assign w3064 = w11345 & w9530;
assign w3065 = ~pi3101 & w261;
assign w3066 = ~w10725 & ~w8668;
assign w3067 = pi2991 & w8571;
assign w3068 = ~pi1084 & w795;
assign w3069 = (w8208 & ~w11247) | (w8208 & w5344) | (~w11247 & w5344);
assign w3070 = w14228 & ~w2741;
assign w3071 = ~w1368 & ~pi0469;
assign w3072 = w7077 & ~w9852;
assign w3073 = ~w837 & ~w15630;
assign w3074 = w539 & ~w4003;
assign w3075 = ~pi3147 & w3805;
assign w3076 = w15808 & ~w14143;
assign w3077 = ~w17031 & ~w6762;
assign w3078 = w5383 & ~w4004;
assign w3079 = ~w17469 & ~w3097;
assign w3080 = w6305 & w6457;
assign w3081 = ~pi1332 & pi1686;
assign w3082 = pi1678 & w14705;
assign w3083 = w13509 & w5965;
assign w3084 = ~w15364 & ~w12661;
assign w3085 = ~pi0483 & pi3404;
assign w3086 = pi3160 & ~pi3481;
assign w3087 = ~pi2119 & w12755;
assign w3088 = ~w1391 & ~pi0980;
assign w3089 = w1813 & w14832;
assign w3090 = ~w2725 & ~pi0963;
assign w3091 = ~w1099 & ~w12182;
assign w3092 = ~w10849 & ~w14485;
assign w3093 = w13509 & w15127;
assign w3094 = pi1683 & w1483;
assign w3095 = ~w8285 & ~w5210;
assign w3096 = w11735 & w6320;
assign w3097 = ~pi2523 & w14148;
assign w3098 = ~w3329 & ~w10924;
assign w3099 = ~pi0563 & w11739;
assign w3100 = (pi0726 & ~w13509) | (pi0726 & w2356) | (~w13509 & w2356);
assign w3101 = w288 & w10051;
assign w3102 = ~w3932 & ~w2463;
assign w3103 = pi2331 & ~w412;
assign w3104 = ~w7850 & w5522;
assign w3105 = ~pi3061 & w261;
assign w3106 = ~w10087 & w10724;
assign w3107 = (~w13367 & w17577) | (~w13367 & w13481) | (w17577 & w13481);
assign w3108 = ~w7070 & ~w12618;
assign w3109 = pi2553 & ~w3987;
assign w3110 = ~pi3171 & pi3207;
assign w3111 = pi3117 & pi3120;
assign w3112 = ~w658 & ~w4949;
assign w3113 = ~w14370 & w11152;
assign w3114 = w2318 & w8401;
assign w3115 = ~pi1243 & pi1256;
assign w3116 = w62 & w12357;
assign w3117 = pi2859 & w14148;
assign w3118 = ~w17679 & w1229;
assign w3119 = (w9771 & ~w2880) | (w9771 & w4611) | (~w2880 & w4611);
assign w3120 = ~w9060 & w11229;
assign w3121 = w9800 & w1910;
assign w3122 = w15842 & pi2285;
assign w3123 = pi2936 & ~w6045;
assign w3124 = ~pi2393 & w5384;
assign w3125 = w18345 & pi0359;
assign w3126 = ~pi3162 & w13570;
assign w3127 = ~w931 & ~w4782;
assign w3128 = ~pi3143 & ~pi3160;
assign w3129 = ~w17468 & ~w2774;
assign w3130 = ~w1791 & w9688;
assign w3131 = w4910 & w2142;
assign w3132 = w11833 & w6763;
assign w3133 = (pi1151 & ~w5437) | (pi1151 & w8121) | (~w5437 & w8121);
assign w3134 = ~pi2406 & w5075;
assign w3135 = ~w14128 & ~w4804;
assign w3136 = pi1333 & ~w8001;
assign w3137 = w5189 & ~w7449;
assign w3138 = w9227 & w735;
assign w3139 = ~w3751 & ~w1795;
assign w3140 = ~w10756 & ~w14208;
assign w3141 = ~w12028 & ~w3299;
assign w3142 = ~w172 & ~w7670;
assign w3143 = w968 & ~pi0283;
assign w3144 = w2725 & ~w1340;
assign w3145 = pi1641 & ~w6448;
assign w3146 = (pi0916 & ~w13509) | (pi0916 & w8191) | (~w13509 & w8191);
assign w3147 = w7307 & w12614;
assign w3148 = ~w15102 & ~w1539;
assign w3149 = w10189 & pi0384;
assign w3150 = ~w2574 & ~w14118;
assign w3151 = ~pi2315 & w12941;
assign w3152 = w13509 & w11051;
assign w3153 = ~w4241 & ~w5744;
assign w3154 = pi1469 & w13753;
assign w3155 = ~w2725 & pi0908;
assign w3156 = ~pi3164 & w11701;
assign w3157 = ~w10231 & ~w4594;
assign w3158 = pi1420 & ~w6072;
assign w3159 = ~w1146 & ~w11897;
assign w3160 = ~w3000 & ~pi1978;
assign w3161 = ~w11445 & ~w11261;
assign w3162 = ~pi2348 & w8617;
assign w3163 = ~pi0081 & ~pi1353;
assign w3164 = pi0254 & w5274;
assign w3165 = ~w1011 & ~w17083;
assign w3166 = w15590 & w406;
assign w3167 = ~pi1983 & ~pi1985;
assign w3168 = ~w2834 & w3819;
assign w3169 = w17646 & w14078;
assign w3170 = ~w13895 & ~w16060;
assign w3171 = ~pi3172 & w3805;
assign w3172 = w1391 & ~w3430;
assign w3173 = w13509 & w5541;
assign w3174 = pi2494 & ~w9504;
assign w3175 = ~pi2994 & w6072;
assign w3176 = pi0251 & w5274;
assign w3177 = w7595 & w12508;
assign w3178 = pi2377 & ~w17683;
assign w3179 = w11383 & w13439;
assign w3180 = w6649 & ~w7129;
assign w3181 = ~w12460 & w9349;
assign w3182 = ~w11172 & ~w12767;
assign w3183 = ~pi2930 & w17213;
assign w3184 = pi2152 & ~w11671;
assign w3185 = w15883 & w17115;
assign w3186 = ~pi1224 & ~pi1211;
assign w3187 = pi1944 & ~w17646;
assign w3188 = pi2399 & ~w14524;
assign w3189 = ~w13900 & ~w11410;
assign w3190 = ~pi3153 & w15839;
assign w3191 = ~w4482 & ~w12971;
assign w3192 = pi3160 & ~w8795;
assign w3193 = pi3142 & w7946;
assign w3194 = w2114 & w14093;
assign w3195 = w2725 & ~w6922;
assign w3196 = pi0483 & pi0509;
assign w3197 = pi2571 & ~w5274;
assign w3198 = ~pi0501 & pi1147;
assign w3199 = w8265 & w10;
assign w3200 = w11579 & w4989;
assign w3201 = w10647 & ~w8340;
assign w3202 = ~pi0923 & w17490;
assign w3203 = w7254 & w3988;
assign w3204 = ~w10957 & ~w9524;
assign w3205 = ~w4712 & ~w6246;
assign w3206 = ~pi2827 & w15122;
assign w3207 = ~w6524 & ~w6143;
assign w3208 = ~pi0690 & w9110;
assign w3209 = ~pi1016 & w9110;
assign w3210 = ~pi1984 & ~w15450;
assign w3211 = ~pi3135 & w15048;
assign w3212 = ~pi3048 & w226;
assign w3213 = ~w13211 & ~w6588;
assign w3214 = ~w10996 & ~w8732;
assign w3215 = ~w8764 & ~w5870;
assign w3216 = pi2160 & ~w412;
assign w3217 = pi2966 & pi2479;
assign w3218 = ~w13269 & ~w13521;
assign w3219 = ~w9468 & ~w8491;
assign w3220 = ~w14560 & pi0209;
assign w3221 = ~w3710 & ~w6882;
assign w3222 = ~w2014 & w18511;
assign w3223 = ~pi1983 & w2247;
assign w3224 = w14803 & w2853;
assign w3225 = ~pi0728 & w17899;
assign w3226 = w1391 & ~w2741;
assign w3227 = ~w5397 & ~w17195;
assign w3228 = w5756 & w3081;
assign w3229 = w15564 & w5806;
assign w3230 = w13509 & w16164;
assign w3231 = ~w2552 & ~w1994;
assign w3232 = w15122 & ~pi2722;
assign w3233 = ~w16930 & ~w15111;
assign w3234 = pi0130 & w5274;
assign w3235 = w908 & w3490;
assign w3236 = ~pi1837 & ~w4420;
assign w3237 = pi2652 & ~w16815;
assign w3238 = (~w1541 & ~w5517) | (~w1541 & w9933) | (~w5517 & w9933);
assign w3239 = w7799 & w3890;
assign w3240 = ~w17712 & ~w16696;
assign w3241 = ~w11301 & ~w13003;
assign w3242 = ~w6195 & w9225;
assign w3243 = ~w12239 & ~w1505;
assign w3244 = ~w13231 & pi0570;
assign w3245 = ~w7844 & pi0612;
assign w3246 = w7703 & w16111;
assign w3247 = ~w7969 & ~w4161;
assign w3248 = pi0038 & ~w14148;
assign w3249 = w3493 & w5703;
assign w3250 = ~w1550 & ~w6430;
assign w3251 = pi1397 & ~w6853;
assign w3252 = w13423 & w6332;
assign w3253 = pi2078 & ~w17683;
assign w3254 = ~w1791 & w17649;
assign w3255 = w17579 & w15475;
assign w3256 = ~pi2648 & w15122;
assign w3257 = ~w8341 & ~w7192;
assign w3258 = ~pi1770 & ~pi3172;
assign w3259 = pi2434 & ~w11406;
assign w3260 = ~pi2909 & w9687;
assign w3261 = ~pi3165 & w14753;
assign w3262 = ~pi2519 & ~w2431;
assign w3263 = ~pi3062 & w3555;
assign w3264 = ~w4410 & w11743;
assign w3265 = pi1178 & pi3219;
assign w3266 = pi0059 & w1171;
assign w3267 = ~pi0970 & w17899;
assign w3268 = w9353 & w988;
assign w3269 = ~pi3293 & w6448;
assign w3270 = ~pi0410 & w17173;
assign w3271 = w11735 & w2753;
assign w3272 = (~pi0280 & ~w6857) | (~pi0280 & w386) | (~w6857 & w386);
assign w3273 = (pi0564 & ~w13509) | (pi0564 & w7427) | (~w13509 & w7427);
assign w3274 = pi1337 & ~w3709;
assign w3275 = ~w1827 & ~pi0497;
assign w3276 = w7844 & ~w7020;
assign w3277 = ~pi3164 & w15048;
assign w3278 = w17562 & pi1848;
assign w3279 = ~pi3027 & ~w16550;
assign w3280 = ~w11100 & ~w12799;
assign w3281 = ~pi2123 & w11313;
assign w3282 = ~pi3150 & pi3207;
assign w3283 = w5917 & w17501;
assign w3284 = pi2394 & ~w3223;
assign w3285 = w13509 & w15701;
assign w3286 = w13509 & w17108;
assign w3287 = w5452 & w14193;
assign w3288 = ~w12079 & ~w11306;
assign w3289 = ~w8356 & w229;
assign w3290 = ~w12094 & ~w2007;
assign w3291 = ~w5419 & ~w13089;
assign w3292 = ~w15122 & ~pi2646;
assign w3293 = ~w10621 & ~w5581;
assign w3294 = w13509 & w15836;
assign w3295 = ~w2379 & ~w11431;
assign w3296 = ~w3000 & ~pi2743;
assign w3297 = ~pi0572 & w11739;
assign w3298 = w5225 & w6558;
assign w3299 = w13509 & w4624;
assign w3300 = ~w15808 & pi1030;
assign w3301 = w709 & pi1900;
assign w3302 = ~pi3138 & w11132;
assign w3303 = pi1671 & ~w4058;
assign w3304 = ~w11923 & ~w11030;
assign w3305 = w62 & ~w17477;
assign w3306 = ~w2748 & w1362;
assign w3307 = ~pi0483 & pi3394;
assign w3308 = pi2762 & w605;
assign w3309 = ~w18273 & w5649;
assign w3310 = w7307 & w18117;
assign w3311 = ~w17577 & w17619;
assign w3312 = pi0035 & ~w3748;
assign w3313 = (pi0548 & ~w13509) | (pi0548 & w16651) | (~w13509 & w16651);
assign w3314 = w1391 & ~w13195;
assign w3315 = ~w16897 & w8867;
assign w3316 = ~w1007 & w15977;
assign w3317 = w6288 & w4833;
assign w3318 = pi1759 & pi3168;
assign w3319 = ~w13519 & ~w2916;
assign w3320 = ~w5560 & w9034;
assign w3321 = (pi0580 & ~w13509) | (pi0580 & w1916) | (~w13509 & w1916);
assign w3322 = pi1613 & ~w7090;
assign w3323 = w16506 & w2042;
assign w3324 = ~w6650 & ~w1194;
assign w3325 = w17103 & w2280;
assign w3326 = w3223 & w6320;
assign w3327 = ~pi2183 & w5384;
assign w3328 = ~w14834 & ~w16275;
assign w3329 = ~w1791 & w3348;
assign w3330 = w7982 & w1486;
assign w3331 = ~pi3130 & pi1271;
assign w3332 = ~pi3518 & ~w2322;
assign w3333 = w16620 & w9084;
assign w3334 = ~pi3159 & w13570;
assign w3335 = w2280 & pi0061;
assign w3336 = ~w11134 & ~w3339;
assign w3337 = (pi0941 & ~w13509) | (pi0941 & w15983) | (~w13509 & w15983);
assign w3338 = (pi0718 & ~w13509) | (pi0718 & w10190) | (~w13509 & w10190);
assign w3339 = ~pi3311 & w16922;
assign w3340 = ~pi0041 & w922;
assign w3341 = w6697 & ~w4043;
assign w3342 = ~pi2408 & w13204;
assign w3343 = ~w14815 & ~w1658;
assign w3344 = ~w9038 & ~w9963;
assign w3345 = ~w12646 & ~w6471;
assign w3346 = w7077 & ~w4043;
assign w3347 = pi2182 & ~w14524;
assign w3348 = ~pi2647 & w15122;
assign w3349 = ~w11347 & ~w231;
assign w3350 = pi1614 & ~w7090;
assign w3351 = ~w7574 & ~w7093;
assign w3352 = ~w9067 & ~w12154;
assign w3353 = pi1337 & pi0302;
assign w3354 = ~w16278 & pi1026;
assign w3355 = w11623 & w922;
assign w3356 = w15808 & ~w7707;
assign w3357 = ~pi1182 & ~pi1195;
assign w3358 = w2971 & w14210;
assign w3359 = pi3064 & ~w16502;
assign w3360 = ~pi0712 & w3106;
assign w3361 = w709 & pi1889;
assign w3362 = ~pi3116 & pi3132;
assign w3363 = pi1169 & pi3198;
assign w3364 = w934 & pi0428;
assign w3365 = ~w9099 & ~w17137;
assign w3366 = ~pi2453 & w5384;
assign w3367 = pi1449 & ~w13753;
assign w3368 = pi2348 & ~w4508;
assign w3369 = pi3170 & w1793;
assign w3370 = ~w3203 & pi0577;
assign w3371 = ~w17723 & ~w17530;
assign w3372 = w5623 & w6563;
assign w3373 = ~pi2373 & w12755;
assign w3374 = ~w13266 & ~w13853;
assign w3375 = w14445 & w596;
assign w3376 = ~w3338 & ~w5670;
assign w3377 = ~pi3015 & ~pi3207;
assign w3378 = w13509 & w16948;
assign w3379 = w2725 & ~w14597;
assign w3380 = ~w14228 & pi0626;
assign w3381 = ~w4282 & ~w4904;
assign w3382 = ~w17665 & ~w11500;
assign w3383 = pi2271 & ~w17683;
assign w3384 = ~w810 & ~w15088;
assign w3385 = ~pi3150 & w14753;
assign w3386 = w17562 & pi1812;
assign w3387 = (pi0351 & w6195) | (pi0351 & w12642) | (w6195 & w12642);
assign w3388 = ~w11036 & w17624;
assign w3389 = ~pi1031 & w17490;
assign w3390 = w12460 & w12770;
assign w3391 = pi1824 & ~w2732;
assign w3392 = w14228 & ~w12800;
assign w3393 = w13509 & w3356;
assign w3394 = w7799 & w12186;
assign w3395 = ~pi2276 & w12724;
assign w3396 = ~w11944 & ~w5301;
assign w3397 = ~w2370 & ~w2040;
assign w3398 = ~w9493 & ~w3265;
assign w3399 = ~w5453 & ~pi1766;
assign w3400 = ~pi1367 & ~pi1371;
assign w3401 = ~w2725 & pi0798;
assign w3402 = pi1778 & w8383;
assign w3403 = w14648 & ~pi2784;
assign w3404 = ~w2793 & w11208;
assign w3405 = pi1208 & ~w11010;
assign w3406 = ~w16453 & ~w7143;
assign w3407 = ~pi1265 & ~w8804;
assign w3408 = pi3118 & w4592;
assign w3409 = ~w18153 & ~w18509;
assign w3410 = ~pi3057 & pi2980;
assign w3411 = ~pi2981 & w13584;
assign w3412 = ~w2725 & pi0787;
assign w3413 = ~w9355 & ~w12252;
assign w3414 = ~w2791 & ~w1696;
assign w3415 = w5161 & w10117;
assign w3416 = ~w18587 & pi1337;
assign w3417 = w16575 & w12455;
assign w3418 = ~w8899 & ~w10917;
assign w3419 = ~w15104 & ~w351;
assign w3420 = ~w2423 & ~w204;
assign w3421 = ~w17665 & ~w17360;
assign w3422 = (pi0881 & ~w13509) | (pi0881 & w14126) | (~w13509 & w14126);
assign w3423 = w10189 & ~pi0473;
assign w3424 = (~pi0274 & ~w6857) | (~pi0274 & w13255) | (~w6857 & w13255);
assign w3425 = ~w17288 & ~w1457;
assign w3426 = w384 & w16914;
assign w3427 = ~pi1912 & w9340;
assign w3428 = ~pi3170 & w11701;
assign w3429 = w13509 & w16376;
assign w3430 = ~w872 & ~w6021;
assign w3431 = pi1307 & ~w14094;
assign w3432 = ~pi2873 & w735;
assign w3433 = pi2830 & ~w226;
assign w3434 = (pi0992 & ~w13509) | (pi0992 & w3454) | (~w13509 & w3454);
assign w3435 = w12460 & w9329;
assign w3436 = ~pi2037 & w7455;
assign w3437 = ~pi0573 & w11739;
assign w3438 = ~w2014 & w12809;
assign w3439 = pi0389 & w12302;
assign w3440 = ~w9624 & ~w12445;
assign w3441 = w412 & w2753;
assign w3442 = w4364 & ~pi0434;
assign w3443 = ~w11234 & ~w12014;
assign w3444 = w14109 & pi0438;
assign w3445 = ~pi1197 & w11739;
assign w3446 = ~w329 & w15420;
assign w3447 = ~w16278 & pi0712;
assign w3448 = w11383 & w7723;
assign w3449 = ~w16289 & ~w3192;
assign w3450 = pi2862 & w14148;
assign w3451 = pi0145 & w5274;
assign w3452 = w2192 & w15324;
assign w3453 = ~w11335 & ~w17403;
assign w3454 = ~w13231 & pi0992;
assign w3455 = ~pi2464 & w9340;
assign w3456 = ~pi0607 & w12825;
assign w3457 = ~pi2967 & ~pi3046;
assign w3458 = w1962 & w1217;
assign w3459 = ~pi0564 & w11739;
assign w3460 = w1391 & ~w13028;
assign w3461 = pi1804 & ~pi3132;
assign w3462 = (w1599 & ~w17173) | (w1599 & w18586) | (~w17173 & w18586);
assign w3463 = ~pi0741 & w17490;
assign w3464 = ~w6464 & ~w15699;
assign w3465 = w11345 & w16068;
assign w3466 = pi1330 & ~w10296;
assign w3467 = ~pi3318 & w18259;
assign w3468 = ~w13523 & ~w3537;
assign w3469 = ~pi2478 & w5384;
assign w3470 = pi1594 & ~w13753;
assign w3471 = w5274 & w11714;
assign w3472 = ~pi3163 & w8515;
assign w3473 = ~pi3154 & pi3172;
assign w3474 = ~w6079 & w7238;
assign w3475 = pi2110 & ~w412;
assign w3476 = w13509 & w10890;
assign w3477 = pi3033 & ~w16502;
assign w3478 = ~w2393 & w13508;
assign w3479 = pi1261 & pi2553;
assign w3480 = ~w10857 & ~w13827;
assign w3481 = pi3001 & ~pi2995;
assign w3482 = ~pi0725 & w17899;
assign w3483 = ~w7844 & pi0606;
assign w3484 = pi3007 & ~pi3057;
assign w3485 = w14896 & w11130;
assign w3486 = ~w3203 & pi0587;
assign w3487 = w1962 & ~w12800;
assign w3488 = pi1158 & w9420;
assign w3489 = w13509 & w16799;
assign w3490 = w10048 & w15646;
assign w3491 = ~pi3009 & ~pi3207;
assign w3492 = ~w18097 & ~w4906;
assign w3493 = ~w11909 & ~w9050;
assign w3494 = ~w5900 & w10744;
assign w3495 = ~w10550 & ~w14829;
assign w3496 = w13509 & w5204;
assign w3497 = ~w6785 & pi0871;
assign w3498 = pi1782 & ~w10325;
assign w3499 = pi0051 & ~w14148;
assign w3500 = ~w2251 & ~w6311;
assign w3501 = w13509 & w17868;
assign w3502 = ~w18542 & w6198;
assign w3503 = pi0303 & w5274;
assign w3504 = ~w5855 & w6602;
assign w3505 = ~pi0588 & w795;
assign w3506 = w13509 & w8644;
assign w3507 = ~w1962 & ~pi1201;
assign w3508 = ~pi3440 & w15036;
assign w3509 = ~w5653 & ~w6677;
assign w3510 = ~w11355 & ~w1234;
assign w3511 = ~w11160 & ~w17106;
assign w3512 = pi3024 & ~w3987;
assign w3513 = ~w15122 & ~pi2768;
assign w3514 = (pi0893 & ~w13509) | (pi0893 & w2010) | (~w13509 & w2010);
assign w3515 = ~pi3143 & ~w4020;
assign w3516 = ~pi0487 & ~pi1345;
assign w3517 = w13509 & w6485;
assign w3518 = ~pi3298 & w6072;
assign w3519 = w535 & w4627;
assign w3520 = ~pi0628 & w14641;
assign w3521 = ~w7782 & ~w9974;
assign w3522 = ~pi3174 & w3780;
assign w3523 = w7844 & ~w10947;
assign w3524 = w539 & ~w3852;
assign w3525 = ~pi2976 & w226;
assign w3526 = ~w1501 & ~w15557;
assign w3527 = pi2058 & ~w10158;
assign w3528 = ~pi2967 & pi3051;
assign w3529 = ~w3900 & ~w42;
assign w3530 = ~w11375 & ~w11732;
assign w3531 = ~w13282 & ~w15227;
assign w3532 = w7307 & w2851;
assign w3533 = ~w16597 & ~w13755;
assign w3534 = w7703 & w13953;
assign w3535 = w13509 & w15567;
assign w3536 = pi2761 & w14148;
assign w3537 = pi3160 & ~pi3500;
assign w3538 = (pi1191 & ~w5437) | (pi1191 & w1431) | (~w5437 & w1431);
assign w3539 = pi1608 & w13753;
assign w3540 = ~w6785 & pi0866;
assign w3541 = ~w14933 & ~w12222;
assign w3542 = ~w11449 & ~w1438;
assign w3543 = w13568 & w787;
assign w3544 = w4936 & w6422;
assign w3545 = w14228 & w15609;
assign w3546 = w7620 & w6094;
assign w3547 = ~w2999 & w16377;
assign w3548 = pi2527 & w14148;
assign w3549 = w11383 & w7647;
assign w3550 = w5456 & w2878;
assign w3551 = ~w287 & ~w17520;
assign w3552 = w11350 & w2231;
assign w3553 = ~w12460 & w17725;
assign w3554 = ~w14212 & ~w6791;
assign w3555 = pi2949 & w5675;
assign w3556 = ~w16650 & ~w1929;
assign w3557 = pi2488 & ~w5274;
assign w3558 = ~pi3099 & w226;
assign w3559 = w14648 & ~pi2164;
assign w3560 = w14648 & ~pi2642;
assign w3561 = pi3134 & w653;
assign w3562 = ~w13964 & ~w2004;
assign w3563 = ~pi0294 & w4058;
assign w3564 = ~pi3098 & w16815;
assign w3565 = ~w6555 & w561;
assign w3566 = w1391 & ~w15173;
assign w3567 = w9568 & w11314;
assign w3568 = ~w17909 & ~w3083;
assign w3569 = pi3067 & ~pi3147;
assign w3570 = ~pi2081 & w17439;
assign w3571 = ~w16698 & ~w2777;
assign w3572 = w14718 & w11592;
assign w3573 = w9742 & w1764;
assign w3574 = ~pi1063 & w93;
assign w3575 = pi1390 & ~w17935;
assign w3576 = ~pi2293 & w15122;
assign w3577 = w12460 & w15931;
assign w3578 = ~pi2994 & w9781;
assign w3579 = w6009 & w16219;
assign w3580 = ~pi2427 & w5075;
assign w3581 = w5477 & ~w1341;
assign w3582 = ~pi1053 & w1126;
assign w3583 = ~w11613 & ~w910;
assign w3584 = ~w16161 & w4067;
assign w3585 = ~w17131 & w6858;
assign w3586 = pi1883 & ~w226;
assign w3587 = (pi0770 & ~w13509) | (pi0770 & w8328) | (~w13509 & w8328);
assign w3588 = w17619 & pi0508;
assign w3589 = ~pi1718 & pi3171;
assign w3590 = pi0077 & ~pi0128;
assign w3591 = ~w1962 & pi0640;
assign w3592 = pi1281 & pi1345;
assign w3593 = w12460 & w15412;
assign w3594 = ~w2673 & ~w5092;
assign w3595 = ~pi3142 & ~pi3160;
assign w3596 = w5991 & w2009;
assign w3597 = pi2876 & ~w226;
assign w3598 = ~w2003 & w16026;
assign w3599 = ~w334 & ~w13727;
assign w3600 = w8904 & w6362;
assign w3601 = pi1515 & ~w14918;
assign w3602 = ~w9080 & ~w3810;
assign w3603 = (pi0313 & w3055) | (pi0313 & w5860) | (w3055 & w5860);
assign w3604 = ~pi2122 & w12755;
assign w3605 = w13509 & w1565;
assign w3606 = pi2035 & ~w17646;
assign w3607 = ~w3000 & ~pi2487;
assign w3608 = (~pi0957 & ~w13509) | (~pi0957 & w10741) | (~w13509 & w10741);
assign w3609 = (pi1041 & ~w13509) | (pi1041 & w16448) | (~w13509 & w16448);
assign w3610 = ~w16506 & pi1155;
assign w3611 = (pi1112 & ~w13509) | (pi1112 & w8780) | (~w13509 & w8780);
assign w3612 = pi1769 & ~pi3157;
assign w3613 = ~w5012 & w13625;
assign w3614 = (pi0376 & w6195) | (pi0376 & w17628) | (w6195 & w17628);
assign w3615 = w14216 & w8671;
assign w3616 = w9552 & w3159;
assign w3617 = ~w11495 & ~w5616;
assign w3618 = ~w15429 & ~w11872;
assign w3619 = w7229 & ~w17783;
assign w3620 = ~w16572 & ~w17394;
assign w3621 = w13509 & w10657;
assign w3622 = ~w15152 & ~w12779;
assign w3623 = pi3145 & w7946;
assign w3624 = ~pi3164 & w17800;
assign w3625 = (pi1876 & w2014) | (pi1876 & w8455) | (w2014 & w8455);
assign w3626 = pi1406 & ~w3024;
assign w3627 = w14648 & ~pi2712;
assign w3628 = ~w17248 & pi1121;
assign w3629 = ~w640 & ~w17703;
assign w3630 = pi2549 & w14148;
assign w3631 = pi2818 & w605;
assign w3632 = (pi0572 & ~w13509) | (pi0572 & w15099) | (~w13509 & w15099);
assign w3633 = ~w11458 & ~w14462;
assign w3634 = w13509 & w13737;
assign w3635 = ~w10548 & w10778;
assign w3636 = ~pi0483 & pi3384;
assign w3637 = pi2018 & ~w14833;
assign w3638 = ~w5891 & ~w11759;
assign w3639 = w14648 & ~pi2613;
assign w3640 = ~w248 & ~w14965;
assign w3641 = w9989 & w18091;
assign w3642 = w1127 & ~w15802;
assign w3643 = (pi1015 & ~w13509) | (pi1015 & w9551) | (~w13509 & w9551);
assign w3644 = ~w11590 & ~w494;
assign w3645 = ~w13902 & ~w17715;
assign w3646 = ~w379 & w7877;
assign w3647 = pi2870 & w14148;
assign w3648 = w11345 & w10662;
assign w3649 = w11345 & w10663;
assign w3650 = w13509 & w2173;
assign w3651 = (~pi2969 & w10910) | (~pi2969 & w17636) | (w10910 & w17636);
assign w3652 = ~w1823 & ~w8246;
assign w3653 = w18267 & w1620;
assign w3654 = (pi1098 & ~w13509) | (pi1098 & w11601) | (~w13509 & w11601);
assign w3655 = pi3179 & ~w325;
assign w3656 = w10818 & ~w971;
assign w3657 = pi1157 & w9420;
assign w3658 = ~pi2470 & w9340;
assign w3659 = w5189 & ~w14465;
assign w3660 = ~w7721 & w11694;
assign w3661 = ~w17704 & ~w7517;
assign w3662 = w1368 & pi0394;
assign w3663 = pi1511 & ~w16922;
assign w3664 = ~pi3355 & w18259;
assign w3665 = ~w14665 & ~w13558;
assign w3666 = (~pi0273 & ~w6857) | (~pi0273 & w8825) | (~w6857 & w8825);
assign w3667 = w6665 & w1857;
assign w3668 = ~pi2214 & w2151;
assign w3669 = ~pi3158 & w17993;
assign w3670 = ~w270 & w14798;
assign w3671 = pi1372 & ~w4395;
assign w3672 = ~w6092 & w5244;
assign w3673 = w1516 & w255;
assign w3674 = ~w10813 & ~w7451;
assign w3675 = ~w7077 & pi0807;
assign w3676 = (pi1088 & ~w13509) | (pi1088 & w12279) | (~w13509 & w12279);
assign w3677 = pi3157 & w2732;
assign w3678 = ~w16161 & pi0001;
assign w3679 = ~pi3136 & pi3161;
assign w3680 = w3203 & ~w14143;
assign w3681 = ~pi3136 & ~pi3160;
assign w3682 = ~pi3172 & w15048;
assign w3683 = ~w764 & w5274;
assign w3684 = ~w15808 & pi0750;
assign w3685 = pi2108 & ~w412;
assign w3686 = (pi0739 & ~w13509) | (pi0739 & w8226) | (~w13509 & w8226);
assign w3687 = ~w14560 & pi0239;
assign w3688 = w13509 & w13258;
assign w3689 = ~pi1816 & w3709;
assign w3690 = (pi0817 & ~w13509) | (pi0817 & w1786) | (~w13509 & w1786);
assign w3691 = ~pi3286 & w6448;
assign w3692 = pi3135 & w2732;
assign w3693 = w3243 & ~pi0323;
assign w3694 = w3243 & pi0324;
assign w3695 = ~w7211 & ~w10873;
assign w3696 = ~w11734 & ~w12892;
assign w3697 = ~pi0599 & w12825;
assign w3698 = ~pi2972 & ~pi3160;
assign w3699 = ~pi0433 & w17173;
assign w3700 = pi0434 & w17173;
assign w3701 = (pi0558 & ~w13509) | (pi0558 & w11568) | (~w13509 & w11568);
assign w3702 = ~w2529 & ~w11363;
assign w3703 = ~w1976 & ~w16263;
assign w3704 = ~w5162 & ~w2395;
assign w3705 = w4009 & ~w7936;
assign w3706 = ~pi3100 & w11406;
assign w3707 = w5969 & w4345;
assign w3708 = w14524 & w6320;
assign w3709 = ~pi2525 & w13236;
assign w3710 = (pi0901 & ~w13509) | (pi0901 & w13121) | (~w13509 & w13121);
assign w3711 = ~w3761 & ~w13122;
assign w3712 = ~w11765 & ~w10259;
assign w3713 = ~pi0289 & w4058;
assign w3714 = w15122 & ~pi2638;
assign w3715 = ~w15781 & ~w3691;
assign w3716 = ~w714 & ~w6478;
assign w3717 = ~pi2990 & w16502;
assign w3718 = ~w3317 & ~w4901;
assign w3719 = ~w6490 & w15908;
assign w3720 = ~pi1257 & ~pi1238;
assign w3721 = w1368 & pi0384;
assign w3722 = w62 & ~w10359;
assign w3723 = ~w7051 & w10647;
assign w3724 = pi2849 & w7965;
assign w3725 = ~pi3098 & w226;
assign w3726 = w17562 & pi2558;
assign w3727 = ~w17248 & pi0879;
assign w3728 = pi0056 & ~w14148;
assign w3729 = pi2274 & ~w4508;
assign w3730 = ~w7568 & ~w2996;
assign w3731 = pi2918 & ~pi2943;
assign w3732 = pi1714 & ~pi3155;
assign w3733 = ~w770 & w18061;
assign w3734 = pi1650 & ~w6072;
assign w3735 = pi1325 & pi1345;
assign w3736 = w13509 & w6725;
assign w3737 = ~w12311 & ~w12470;
assign w3738 = ~w17965 & ~w16589;
assign w3739 = ~w6985 & ~w10866;
assign w3740 = w10158 & w2753;
assign w3741 = w9440 & pi0182;
assign w3742 = ~w7500 & ~w6097;
assign w3743 = ~w1391 & pi1058;
assign w3744 = ~pi0123 & w9284;
assign w3745 = pi3163 & w4256;
assign w3746 = ~w13273 & ~w11235;
assign w3747 = ~w361 & ~w16308;
assign w3748 = w1766 & w4015;
assign w3749 = (pi1268 & ~w5437) | (pi1268 & w552) | (~w5437 & w552);
assign w3750 = (pi0907 & ~w13509) | (pi0907 & w11058) | (~w13509 & w11058);
assign w3751 = pi2212 & ~w15271;
assign w3752 = ~pi1715 & pi3154;
assign w3753 = ~pi0799 & w543;
assign w3754 = ~w3422 & ~w12494;
assign w3755 = w14109 & pi0442;
assign w3756 = ~w14518 & w17168;
assign w3757 = ~pi0570 & w11739;
assign w3758 = ~w3580 & ~w11084;
assign w3759 = ~w4242 & w1708;
assign w3760 = ~pi2327 & w8617;
assign w3761 = ~pi0551 & w6200;
assign w3762 = pi2790 & ~w11406;
assign w3763 = pi2623 & ~w16815;
assign w3764 = w18123 & w6320;
assign w3765 = ~w8166 & w18382;
assign w3766 = ~pi2994 & w17935;
assign w3767 = ~w1883 & ~w18549;
assign w3768 = ~w6377 & ~w10735;
assign w3769 = ~pi2969 & w11360;
assign w3770 = (~pi0256 & ~w325) | (~pi0256 & w7040) | (~w325 & w7040);
assign w3771 = (pi0257 & ~w325) | (pi0257 & w7041) | (~w325 & w7041);
assign w3772 = (~pi0352 & ~w6857) | (~pi0352 & w16980) | (~w6857 & w16980);
assign w3773 = (pi0579 & ~w13509) | (pi0579 & w18383) | (~w13509 & w18383);
assign w3774 = w15842 & w2971;
assign w3775 = ~w5015 & ~pi0512;
assign w3776 = pi1585 & ~w14918;
assign w3777 = pi1647 & ~w6072;
assign w3778 = pi1886 & ~w15036;
assign w3779 = ~w1756 & ~w14727;
assign w3780 = pi1374 & ~pi2948;
assign w3781 = pi2997 & ~w3987;
assign w3782 = w13509 & w11749;
assign w3783 = ~pi3135 & w8515;
assign w3784 = w15883 & w9407;
assign w3785 = ~pi0278 & w2196;
assign w3786 = ~pi0492 & ~pi1345;
assign w3787 = pi3131 & w3987;
assign w3788 = ~w9807 & ~w3360;
assign w3789 = ~w9016 & ~w11181;
assign w3790 = ~w6361 & ~w2481;
assign w3791 = w3381 & ~w10724;
assign w3792 = ~pi3355 & w6448;
assign w3793 = ~w14762 & ~w16777;
assign w3794 = pi1648 & ~w17935;
assign w3795 = ~pi1800 & ~pi3146;
assign w3796 = ~w11203 & ~w10208;
assign w3797 = ~pi2194 & w9340;
assign w3798 = ~w3663 & ~w11844;
assign w3799 = ~pi2265 & w13065;
assign w3800 = w13231 & ~w6922;
assign w3801 = (pi1009 & ~w13509) | (pi1009 & w273) | (~w13509 & w273);
assign w3802 = ~pi2372 & w17439;
assign w3803 = ~w14543 & ~w16106;
assign w3804 = ~w9756 & ~w7895;
assign w3805 = ~w4020 & w9414;
assign w3806 = ~w16392 & ~w1662;
assign w3807 = ~w12140 & ~w11393;
assign w3808 = (pi1058 & ~w13509) | (pi1058 & w3743) | (~w13509 & w3743);
assign w3809 = ~pi3142 & w3982;
assign w3810 = pi2216 & ~w15271;
assign w3811 = ~w5560 & w6887;
assign w3812 = pi1168 & ~pi3194;
assign w3813 = ~w6474 & ~w8913;
assign w3814 = ~w1263 & ~w9634;
assign w3815 = ~pi2473 & w9340;
assign w3816 = w14833 & ~w8588;
assign w3817 = w7703 & w4394;
assign w3818 = (~pi0953 & ~w13509) | (~pi0953 & w10950) | (~w13509 & w10950);
assign w3819 = ~w11788 & ~w3183;
assign w3820 = ~w1563 & ~w13309;
assign w3821 = (pi0407 & w5560) | (pi0407 & w9296) | (w5560 & w9296);
assign w3822 = ~w3685 & ~w3441;
assign w3823 = ~w15808 & pi1094;
assign w3824 = w5189 & ~w10947;
assign w3825 = w13509 & w6484;
assign w3826 = ~w13364 & ~w829;
assign w3827 = ~pi0615 & w14641;
assign w3828 = ~w11839 & ~w6749;
assign w3829 = w6857 & w9269;
assign w3830 = ~pi1086 & w9110;
assign w3831 = w12067 & w16812;
assign w3832 = w11921 & w6787;
assign w3833 = ~w3043 & ~w16188;
assign w3834 = ~w12366 & ~w5358;
assign w3835 = ~w234 & ~w13367;
assign w3836 = w6617 & w5405;
assign w3837 = w13509 & w16028;
assign w3838 = ~w14560 & pi0227;
assign w3839 = ~pi3158 & w13570;
assign w3840 = ~w14516 & ~w16821;
assign w3841 = ~w10215 & ~w8468;
assign w3842 = pi1492 & ~w9781;
assign w3843 = ~pi2492 & w17213;
assign w3844 = ~pi2442 & w9340;
assign w3845 = ~pi1055 & w1126;
assign w3846 = ~pi3154 & w12427;
assign w3847 = ~pi3135 & w11132;
assign w3848 = pi1993 & ~w9414;
assign w3849 = pi1452 & ~w7090;
assign w3850 = w1391 & ~w2776;
assign w3851 = ~pi3139 & w13730;
assign w3852 = w11638 & w8021;
assign w3853 = pi1274 & pi1345;
assign w3854 = ~pi3084 & w15235;
assign w3855 = ~w4540 & ~w9768;
assign w3856 = ~w3055 & w1790;
assign w3857 = ~w18006 & ~w7426;
assign w3858 = w5383 & w5453;
assign w3859 = ~w11827 & w7460;
assign w3860 = ~w8336 & ~w4444;
assign w3861 = w16506 & ~w305;
assign w3862 = ~pi2218 & w11313;
assign w3863 = pi2174 & ~w15271;
assign w3864 = ~w17719 & ~w15035;
assign w3865 = pi0190 & w5274;
assign w3866 = ~w1688 & w4129;
assign w3867 = ~w12438 & ~w14160;
assign w3868 = w7703 & w1478;
assign w3869 = ~w2725 & pi1081;
assign w3870 = ~w978 & w11360;
assign w3871 = ~pi2940 & ~w6045;
assign w3872 = ~pi0275 & w2196;
assign w3873 = pi3160 & ~pi3478;
assign w3874 = ~w14648 & ~pi2707;
assign w3875 = ~w13250 & ~w9949;
assign w3876 = ~w3888 & ~w2537;
assign w3877 = w5063 & w13785;
assign w3878 = w10971 & w15819;
assign w3879 = w17248 & ~w14465;
assign w3880 = ~pi3097 & w3555;
assign w3881 = ~w11953 & ~w13526;
assign w3882 = w13231 & ~w14978;
assign w3883 = pi1889 & ~w15036;
assign w3884 = ~pi2164 & ~w261;
assign w3885 = ~pi3172 & w14753;
assign w3886 = ~pi1219 & ~w8198;
assign w3887 = ~pi3110 & w16502;
assign w3888 = pi0493 & pi1141;
assign w3889 = w13520 & w6035;
assign w3890 = w17562 & pi1820;
assign w3891 = ~w15459 & ~w5796;
assign w3892 = ~w2952 & ~w7579;
assign w3893 = ~pi1224 & pi2913;
assign w3894 = ~w6785 & pi0986;
assign w3895 = w13509 & w13982;
assign w3896 = ~w1350 & ~w18384;
assign w3897 = pi1337 & ~w3689;
assign w3898 = pi2103 & ~w4420;
assign w3899 = pi0027 & ~w3748;
assign w3900 = pi1730 & ~w4058;
assign w3901 = ~pi2972 & pi3057;
assign w3902 = w13509 & w7603;
assign w3903 = ~w9399 & ~w11322;
assign w3904 = ~pi3347 & w16922;
assign w3905 = ~w1368 & ~pi0451;
assign w3906 = pi1757 & ~w4630;
assign w3907 = ~w16454 & ~w16963;
assign w3908 = ~pi1378 & ~pi2920;
assign w3909 = ~w9338 & w7391;
assign w3910 = ~w3054 & w1407;
assign w3911 = ~w17248 & pi0888;
assign w3912 = ~w13184 & ~w7138;
assign w3913 = ~w13231 & pi0571;
assign w3914 = ~w9275 & ~w17997;
assign w3915 = ~w8705 & ~w14386;
assign w3916 = ~w153 & ~w4352;
assign w3917 = ~w11896 & ~w9802;
assign w3918 = ~w18371 & w11260;
assign w3919 = pi3514 & pi3515;
assign w3920 = w9440 & pi0170;
assign w3921 = w2725 & ~w9852;
assign w3922 = ~w14523 & ~w8290;
assign w3923 = ~pi2130 & w16041;
assign w3924 = (pi0544 & ~w13509) | (pi0544 & w8279) | (~w13509 & w8279);
assign w3925 = ~w5425 & ~w14655;
assign w3926 = ~w15808 & pi0756;
assign w3927 = ~w9724 & ~w5677;
assign w3928 = (pi1067 & ~w13509) | (pi1067 & w14907) | (~w13509 & w14907);
assign w3929 = ~w13231 & pi1095;
assign w3930 = w922 & w8259;
assign w3931 = (~w13564 & ~w9420) | (~w13564 & w8877) | (~w9420 & w8877);
assign w3932 = (pi1132 & ~w5437) | (pi1132 & w15617) | (~w5437 & w15617);
assign w3933 = w3375 & w4135;
assign w3934 = ~w1692 & ~w18247;
assign w3935 = ~pi3166 & w3805;
assign w3936 = ~pi3052 & w226;
assign w3937 = ~pi3050 & w3555;
assign w3938 = ~w389 & w7808;
assign w3939 = w934 & pi0423;
assign w3940 = (pi0733 & ~w13509) | (pi0733 & w7920) | (~w13509 & w7920);
assign w3941 = ~pi0735 & w17899;
assign w3942 = pi1992 & ~w9414;
assign w3943 = (pi0688 & ~w13509) | (pi0688 & w5237) | (~w13509 & w5237);
assign w3944 = w13509 & w11758;
assign w3945 = ~w15525 & ~w8443;
assign w3946 = ~pi0265 & w18262;
assign w3947 = w5292 & w5043;
assign w3948 = ~w10001 & ~w8727;
assign w3949 = pi1171 & pi3209;
assign w3950 = w13509 & w1060;
assign w3951 = ~w4233 & ~w14724;
assign w3952 = ~w16506 & pi1134;
assign w3953 = w16182 & w7741;
assign w3954 = ~w10739 & ~w14205;
assign w3955 = ~pi1103 & w17899;
assign w3956 = ~w16251 & ~w9575;
assign w3957 = pi1469 & ~w7090;
assign w3958 = ~w10267 & ~w12570;
assign w3959 = w13509 & w8531;
assign w3960 = w18111 & w2199;
assign w3961 = ~w13316 & ~w926;
assign w3962 = ~pi1694 & pi1695;
assign w3963 = ~pi2397 & w9340;
assign w3964 = w13509 & w927;
assign w3965 = ~pi2317 & w8617;
assign w3966 = ~w4030 & ~w897;
assign w3967 = w13509 & w4604;
assign w3968 = ~pi1132 & ~pi2938;
assign w3969 = pi1760 & pi3153;
assign w3970 = w4850 & w12633;
assign w3971 = w13509 & w9046;
assign w3972 = (~pi0513 & w17577) | (~pi0513 & w13662) | (w17577 & w13662);
assign w3973 = ~pi2744 & w13343;
assign w3974 = pi0257 & w5274;
assign w3975 = pi2896 & ~w3555;
assign w3976 = ~pi3166 & w17993;
assign w3977 = w13584 & w14800;
assign w3978 = w6352 & w882;
assign w3979 = w13509 & w13672;
assign w3980 = ~w15477 & w15272;
assign w3981 = pi1828 & w7858;
assign w3982 = ~w4020 & w15271;
assign w3983 = w12460 & w10405;
assign w3984 = ~w4512 & ~w16847;
assign w3985 = ~w1807 & ~w11039;
assign w3986 = ~pi3053 & w16815;
assign w3987 = pi3130 & w545;
assign w3988 = pi1167 & pi1176;
assign w3989 = ~w5975 & w11403;
assign w3990 = ~pi3054 & w15235;
assign w3991 = ~pi2273 & w12724;
assign w3992 = w11383 & w10386;
assign w3993 = w5865 & w14303;
assign w3994 = w7164 & w359;
assign w3995 = (~w13367 & w17577) | (~w13367 & w12879) | (w17577 & w12879);
assign w3996 = ~w17810 & ~w4098;
assign w3997 = ~pi3146 & w8515;
assign w3998 = pi1463 & w13753;
assign w3999 = ~pi3084 & w6463;
assign w4000 = ~w5855 & ~w18364;
assign w4001 = ~pi0290 & w2196;
assign w4002 = ~w732 & ~w8766;
assign w4003 = w12705 & w17040;
assign w4004 = ~pi2524 & w735;
assign w4005 = ~w18020 & ~w12285;
assign w4006 = w14560 & pi0356;
assign w4007 = ~pi3315 & w7090;
assign w4008 = pi3508 & w13367;
assign w4009 = pi1161 & w14352;
assign w4010 = ~w7918 & w13140;
assign w4011 = w13509 & w14694;
assign w4012 = pi2443 & ~w10299;
assign w4013 = ~w14100 & ~w10286;
assign w4014 = (pi1186 & ~w5437) | (pi1186 & w2147) | (~w5437 & w2147);
assign w4015 = w16939 & w8324;
assign w4016 = ~w968 & ~w1934;
assign w4017 = pi1551 & w13753;
assign w4018 = w13509 & w1553;
assign w4019 = w9366 & w6481;
assign w4020 = pi3027 & ~pi3201;
assign w4021 = ~w5855 & w4020;
assign w4022 = ~pi2134 & w12941;
assign w4023 = ~w14640 & ~w8162;
assign w4024 = ~pi3128 & w9504;
assign w4025 = ~w1140 & ~w5409;
assign w4026 = ~w5736 & ~w5222;
assign w4027 = ~pi0810 & w1147;
assign w4028 = ~w7019 & ~w2220;
assign w4029 = ~w17921 & ~w11643;
assign w4030 = (pi0751 & ~w13509) | (pi0751 & w694) | (~w13509 & w694);
assign w4031 = ~w440 & ~w8693;
assign w4032 = w1329 & ~w7760;
assign w4033 = pi1337 & pi0304;
assign w4034 = ~w7227 & ~w1746;
assign w4035 = ~w13373 & w1106;
assign w4036 = ~w15044 & ~w600;
assign w4037 = ~w17665 & ~w5539;
assign w4038 = w9720 & pi1710;
assign w4039 = ~w17874 & w13321;
assign w4040 = pi1715 & ~w619;
assign w4041 = ~w888 & ~w9106;
assign w4042 = ~w14187 & ~w7819;
assign w4043 = ~pi1289 & pi1345;
assign w4044 = w3203 & ~w1340;
assign w4045 = ~pi2120 & w12755;
assign w4046 = ~w17 & ~w7344;
assign w4047 = ~w11418 & ~w12086;
assign w4048 = ~pi3094 & w3555;
assign w4049 = w384 & w16609;
assign w4050 = w13509 & w11551;
assign w4051 = ~w2613 & pi1176;
assign w4052 = ~w17666 & ~w8381;
assign w4053 = ~w8968 & ~w15447;
assign w4054 = pi2288 & ~w18123;
assign w4055 = ~w1482 & ~w13923;
assign w4056 = ~w9544 & ~w3187;
assign w4057 = ~pi3171 & w13570;
assign w4058 = ~w325 & ~w17327;
assign w4059 = w2611 & w2026;
assign w4060 = ~pi1029 & w17899;
assign w4061 = pi2776 & ~w15235;
assign w4062 = w11345 & w18365;
assign w4063 = ~w6138 & ~w17324;
assign w4064 = w1962 & ~w4043;
assign w4065 = ~w14848 & ~w7349;
assign w4066 = pi1858 & w13691;
assign w4067 = w1766 & w6203;
assign w4068 = ~w590 & ~w16929;
assign w4069 = ~pi1695 & ~w11760;
assign w4070 = ~w1391 & pi0772;
assign w4071 = pi2323 & ~w4508;
assign w4072 = pi1480 & ~w9781;
assign w4073 = ~w17116 & ~w37;
assign w4074 = (pi1889 & w2014) | (pi1889 & w3361) | (w2014 & w3361);
assign w4075 = pi1426 & ~w13753;
assign w4076 = ~w10275 & ~w16380;
assign w4077 = (w15379 & w8931) | (w15379 & w16207) | (w8931 & w16207);
assign w4078 = ~w14228 & pi1005;
assign w4079 = ~w11700 & ~w5988;
assign w4080 = ~w12975 & w11937;
assign w4081 = ~w9560 & ~w529;
assign w4082 = ~w7077 & pi1043;
assign w4083 = ~w6248 & ~w4596;
assign w4084 = w17741 & w7839;
assign w4085 = ~pi2223 & w2151;
assign w4086 = pi1209 & pi1195;
assign w4087 = ~w16455 & ~w8777;
assign w4088 = w13509 & w9157;
assign w4089 = ~pi3336 & w7090;
assign w4090 = ~w15730 & ~w15437;
assign w4091 = ~pi0879 & w1126;
assign w4092 = pi2507 & ~w9504;
assign w4093 = w2725 & ~w12800;
assign w4094 = pi1512 & ~w16922;
assign w4095 = pi2923 & w6045;
assign w4096 = ~pi3018 & ~pi3160;
assign w4097 = w2742 & ~w12577;
assign w4098 = pi3160 & ~pi3497;
assign w4099 = ~w17665 & ~w1001;
assign w4100 = ~w1391 & pi1093;
assign w4101 = w3203 & ~w14597;
assign w4102 = pi1320 & w458;
assign w4103 = ~w15826 & ~w725;
assign w4104 = ~pi3159 & w17669;
assign w4105 = w14648 & ~pi2493;
assign w4106 = pi1910 & ~w14524;
assign w4107 = ~w16506 & pi1269;
assign w4108 = ~w9095 & ~w8057;
assign w4109 = pi2483 & ~w5274;
assign w4110 = pi0272 & w5113;
assign w4111 = ~pi2946 & w16815;
assign w4112 = w2341 & w15609;
assign w4113 = ~pi3158 & w17669;
assign w4114 = pi2591 & ~w5274;
assign w4115 = ~pi3147 & w14753;
assign w4116 = w15896 & w7113;
assign w4117 = ~pi3340 & w14918;
assign w4118 = pi1630 & ~w13753;
assign w4119 = w13509 & w17454;
assign w4120 = w5642 & w12281;
assign w4121 = ~pi3075 & pi3170;
assign w4122 = ~w15813 & ~w8552;
assign w4123 = ~w7629 & ~w10839;
assign w4124 = ~w15889 & w2008;
assign w4125 = pi0248 & w5113;
assign w4126 = ~w4060 & ~w11071;
assign w4127 = ~w7844 & pi0605;
assign w4128 = ~w1791 & w7655;
assign w4129 = w9158 & w7289;
assign w4130 = w2725 & ~w1236;
assign w4131 = ~pi2570 & pi2966;
assign w4132 = w384 & w11955;
assign w4133 = pi3139 & w10389;
assign w4134 = pi2919 & pi2925;
assign w4135 = w14298 & w15840;
assign w4136 = pi1969 & ~w7177;
assign w4137 = ~w7494 & ~w13844;
assign w4138 = ~pi3170 & w17669;
assign w4139 = ~pi1335 & ~w3987;
assign w4140 = w16893 & w5262;
assign w4141 = w709 & pi1873;
assign w4142 = (pi1782 & w7215) | (pi1782 & w11912) | (w7215 & w11912);
assign w4143 = ~w5721 & ~w10594;
assign w4144 = pi2686 & ~w15235;
assign w4145 = w384 & w7530;
assign w4146 = w4750 & w8947;
assign w4147 = ~pi0900 & w12825;
assign w4148 = ~w1391 & pi0775;
assign w4149 = ~w15719 & ~w1372;
assign w4150 = pi1535 & w13753;
assign w4151 = (pi1004 & ~w13509) | (pi1004 & w13950) | (~w13509 & w13950);
assign w4152 = w7703 & w3513;
assign w4153 = ~pi2423 & w13204;
assign w4154 = ~pi0873 & w1126;
assign w4155 = pi0041 & ~w14148;
assign w4156 = ~w7116 & w8661;
assign w4157 = ~w15608 & ~w6908;
assign w4158 = w13509 & w493;
assign w4159 = ~w6769 & ~w5552;
assign w4160 = ~w13575 & ~w17799;
assign w4161 = w10299 & w14078;
assign w4162 = w7158 & w10802;
assign w4163 = (pi1271 & ~w545) | (pi1271 & w3331) | (~w545 & w3331);
assign w4164 = pi3066 & ~pi3163;
assign w4165 = ~w12435 & ~w13325;
assign w4166 = ~w1391 & pi0759;
assign w4167 = ~w12667 & w6664;
assign w4168 = w16506 & ~w6647;
assign w4169 = ~pi3170 & w12427;
assign w4170 = ~w6303 & w5996;
assign w4171 = ~w7986 & ~w13037;
assign w4172 = (~pi0956 & ~w13509) | (~pi0956 & w3036) | (~w13509 & w3036);
assign w4173 = ~w3749 & ~w12015;
assign w4174 = ~pi3298 & w9781;
assign w4175 = ~pi2042 & w13204;
assign w4176 = ~w9632 & w10171;
assign w4177 = pi1865 & ~w15036;
assign w4178 = pi1793 & w8658;
assign w4179 = pi1321 & pi1345;
assign w4180 = ~w9805 & ~w11726;
assign w4181 = w9192 & w11328;
assign w4182 = pi0094 & w9284;
assign w4183 = ~pi3335 & w14918;
assign w4184 = ~w7512 & ~w16977;
assign w4185 = pi3145 & pi3207;
assign w4186 = ~w7266 & ~w8759;
assign w4187 = ~w14894 & ~w7675;
assign w4188 = pi1731 & ~w4058;
assign w4189 = ~w13027 & ~w7981;
assign w4190 = ~w6836 & ~w8769;
assign w4191 = ~w10753 & ~w18058;
assign w4192 = ~pi0259 & w5113;
assign w4193 = pi0260 & w5113;
assign w4194 = (pi1376 & ~w11505) | (pi1376 & w12169) | (~w11505 & w12169);
assign w4195 = pi0272 & w5274;
assign w4196 = ~pi3048 & w11406;
assign w4197 = ~w217 & ~w11115;
assign w4198 = ~w5560 & w3071;
assign w4199 = w13509 & w5960;
assign w4200 = w1421 & w17971;
assign w4201 = w13231 & w15609;
assign w4202 = w13509 & w5165;
assign w4203 = pi1872 & ~w15036;
assign w4204 = w14109 & pi0414;
assign w4205 = w1962 & ~w6680;
assign w4206 = w13509 & w5016;
assign w4207 = ~w12098 & ~w14492;
assign w4208 = (pi0921 & ~w13509) | (pi0921 & w1218) | (~w13509 & w1218);
assign w4209 = w7307 & w14545;
assign w4210 = w6857 & w10034;
assign w4211 = (~pi1182 & ~w11010) | (~pi1182 & w4988) | (~w11010 & w4988);
assign w4212 = ~w3619 & ~w11518;
assign w4213 = ~w15122 & ~pi2824;
assign w4214 = w10647 & ~w6213;
assign w4215 = w13509 & w2386;
assign w4216 = ~w3472 & ~w16192;
assign w4217 = ~pi3050 & w16815;
assign w4218 = (~pi0502 & ~w11345) | (~pi0502 & w14237) | (~w11345 & w14237);
assign w4219 = pi1265 & ~pi1332;
assign w4220 = pi1703 & ~w18497;
assign w4221 = ~w7398 & ~w3647;
assign w4222 = (~w13166 & ~w5517) | (~w13166 & w5868) | (~w5517 & w5868);
assign w4223 = ~pi3110 & ~w3987;
assign w4224 = (w7799 & w4287) | (w7799 & w11137) | (w4287 & w11137);
assign w4225 = w4420 & w614;
assign w4226 = ~w18421 & ~w10041;
assign w4227 = w15450 & pi1178;
assign w4228 = ~w17225 & ~w8908;
assign w4229 = ~w12965 & w2747;
assign w4230 = ~w12229 & ~w7263;
assign w4231 = pi1339 & ~w2848;
assign w4232 = (pi0307 & ~w325) | (pi0307 & w2160) | (~w325 & w2160);
assign w4233 = (pi0880 & ~w13509) | (pi0880 & w18337) | (~w13509 & w18337);
assign w4234 = ~pi0495 & ~pi1345;
assign w4235 = ~w5453 & ~pi1763;
assign w4236 = w10647 & ~w4877;
assign w4237 = ~w8879 & ~w9868;
assign w4238 = ~w17812 & ~w8643;
assign w4239 = pi1462 & ~w7090;
assign w4240 = w11800 & w447;
assign w4241 = (pi0729 & ~w13509) | (pi0729 & w7714) | (~w13509 & w7714);
assign w4242 = pi1412 & ~w13753;
assign w4243 = ~w15011 & w9445;
assign w4244 = ~w5077 & w14133;
assign w4245 = ~pi2366 & w8617;
assign w4246 = pi1530 & ~w14918;
assign w4247 = pi2804 & ~w11406;
assign w4248 = ~w1702 & ~w14457;
assign w4249 = ~w10099 & ~w10177;
assign w4250 = w10189 & pi0409;
assign w4251 = w9571 & w11963;
assign w4252 = ~w13369 & ~w18051;
assign w4253 = ~pi3138 & w17387;
assign w4254 = pi1828 & pi1984;
assign w4255 = pi1196 & ~w11010;
assign w4256 = w9653 & w876;
assign w4257 = ~w13086 & ~pi2920;
assign w4258 = w1516 & w726;
assign w4259 = ~pi1077 & w543;
assign w4260 = ~w13791 & ~w18598;
assign w4261 = ~pi2815 & w13343;
assign w4262 = ~w9029 & ~w17879;
assign w4263 = w2823 & w654;
assign w4264 = ~pi0554 & w11739;
assign w4265 = (~pi1774 & ~w7799) | (~pi1774 & w1948) | (~w7799 & w1948);
assign w4266 = ~w7681 & w15450;
assign w4267 = ~w12063 & ~w10283;
assign w4268 = pi1166 & pi3198;
assign w4269 = ~w3243 & pi0317;
assign w4270 = w8087 & ~pi0359;
assign w4271 = pi2429 & ~w17646;
assign w4272 = (w2460 & ~w384) | (w2460 & w1034) | (~w384 & w1034);
assign w4273 = w14374 & w5807;
assign w4274 = (pi0888 & ~w13509) | (pi0888 & w3911) | (~w13509 & w3911);
assign w4275 = ~w16353 & ~w1484;
assign w4276 = ~w14957 & ~w5023;
assign w4277 = w10189 & pi0398;
assign w4278 = ~pi3154 & w15839;
assign w4279 = ~w1343 & w6203;
assign w4280 = w10158 & w6320;
assign w4281 = ~w16154 & ~w7082;
assign w4282 = pi1241 & ~w11655;
assign w4283 = (pi0378 & w5560) | (pi0378 & w6643) | (w5560 & w6643);
assign w4284 = (pi0787 & ~w13509) | (pi0787 & w3412) | (~w13509 & w3412);
assign w4285 = pi1611 & w13753;
assign w4286 = pi1467 & ~w7090;
assign w4287 = pi1793 & pi1797;
assign w4288 = ~w8588 & w4420;
assign w4289 = ~w7691 & ~w9595;
assign w4290 = ~pi3160 & ~pi3170;
assign w4291 = ~pi3061 & w226;
assign w4292 = ~w4559 & ~w7206;
assign w4293 = ~pi0662 & w12197;
assign w4294 = pi1656 & ~w13753;
assign w4295 = (pi0337 & w3055) | (pi0337 & w7168) | (w3055 & w7168);
assign w4296 = ~w11452 & ~w12816;
assign w4297 = ~w18178 & ~w16762;
assign w4298 = ~w14648 & ~pi2158;
assign w4299 = ~w14235 & ~w7769;
assign w4300 = ~w5001 & ~w2070;
assign w4301 = ~pi3353 & w6448;
assign w4302 = ~w5453 & ~pi1802;
assign w4303 = w9720 & pi1715;
assign w4304 = w13569 & w15176;
assign w4305 = pi0256 & w5274;
assign w4306 = (pi1190 & ~w13509) | (pi1190 & w11131) | (~w13509 & w11131);
assign w4307 = ~w14456 & ~w5095;
assign w4308 = w1792 & ~w8789;
assign w4309 = ~w17135 & ~w7429;
assign w4310 = ~w4020 & w412;
assign w4311 = pi2315 & ~w15883;
assign w4312 = ~w10559 & ~w13898;
assign w4313 = pi1735 & ~w4058;
assign w4314 = pi3044 & ~w16502;
assign w4315 = (~w12581 & ~w9420) | (~w12581 & w13552) | (~w9420 & w13552);
assign w4316 = ~w2015 & ~w5119;
assign w4317 = (pi0341 & w6195) | (pi0341 & w893) | (w6195 & w893);
assign w4318 = w11209 & ~w14173;
assign w4319 = ~w18003 & ~w8582;
assign w4320 = w12466 & w11711;
assign w4321 = ~pi2445 & w5384;
assign w4322 = w14648 & ~pi2726;
assign w4323 = ~w10794 & ~w13042;
assign w4324 = w17413 & w876;
assign w4325 = ~w15943 & w11975;
assign w4326 = pi1783 & ~w8829;
assign w4327 = w17562 & pi2572;
assign w4328 = ~w5019 & w11312;
assign w4329 = ~pi3343 & w9781;
assign w4330 = pi2285 & ~w5274;
assign w4331 = ~w17688 & w12208;
assign w4332 = w15450 & pi1165;
assign w4333 = ~w458 & w13072;
assign w4334 = ~w9165 & ~w1900;
assign w4335 = pi3038 & w16502;
assign w4336 = ~pi2730 & w15122;
assign w4337 = ~pi1097 & w17490;
assign w4338 = ~w4574 & ~w1208;
assign w4339 = w2341 & ~w13028;
assign w4340 = ~w16535 & ~w3524;
assign w4341 = ~pi1314 & ~pi1302;
assign w4342 = w14043 & w11901;
assign w4343 = pi1907 & ~w10299;
assign w4344 = (pi0368 & w6195) | (pi0368 & w10464) | (w6195 & w10464);
assign w4345 = ~w6761 & ~w11861;
assign w4346 = w14782 & w936;
assign w4347 = ~w530 & ~w13408;
assign w4348 = w2363 & w7498;
assign w4349 = ~w3577 & ~w9724;
assign w4350 = pi1412 & ~w6072;
assign w4351 = pi2871 & w14148;
assign w4352 = ~pi3321 & w16922;
assign w4353 = (pi1087 & ~w13509) | (pi1087 & w17339) | (~w13509 & w17339);
assign w4354 = pi2668 & ~w6463;
assign w4355 = ~w10746 & ~w12927;
assign w4356 = ~pi3060 & w9504;
assign w4357 = pi2118 & ~w412;
assign w4358 = ~w16776 & ~w5731;
assign w4359 = ~pi0100 & w9284;
assign w4360 = pi0101 & w9284;
assign w4361 = w934 & pi0442;
assign w4362 = (pi0574 & ~w13509) | (pi0574 & w13033) | (~w13509 & w13033);
assign w4363 = ~w17819 & w11362;
assign w4364 = w5968 & ~pi1337;
assign w4365 = ~pi2450 & w5384;
assign w4366 = ~w16911 & ~w12047;
assign w4367 = ~pi3089 & w11406;
assign w4368 = ~w9456 & ~w1674;
assign w4369 = pi1164 & ~pi3222;
assign w4370 = pi0499 & pi0515;
assign w4371 = ~w15423 & ~w43;
assign w4372 = w10920 & w12549;
assign w4373 = w6697 & ~w14978;
assign w4374 = pi0258 & w11952;
assign w4375 = (w3078 & w17573) | (w3078 & w12540) | (w17573 & w12540);
assign w4376 = ~pi3139 & w4310;
assign w4377 = ~w10691 & ~w4119;
assign w4378 = pi0305 & w5274;
assign w4379 = pi3143 & w3987;
assign w4380 = w10647 & ~w5068;
assign w4381 = ~w9062 & ~w3439;
assign w4382 = w384 & w7993;
assign w4383 = w17248 & ~w4179;
assign w4384 = (pi1124 & ~w13509) | (pi1124 & w10638) | (~w13509 & w10638);
assign w4385 = ~pi1366 & ~pi2966;
assign w4386 = ~w8770 & ~w9328;
assign w4387 = pi2037 & ~w17646;
assign w4388 = ~pi3103 & w3555;
assign w4389 = ~pi2413 & w9340;
assign w4390 = ~w6387 & ~w4388;
assign w4391 = ~w12411 & ~w10463;
assign w4392 = ~w10552 & ~w5086;
assign w4393 = ~w1962 & pi0645;
assign w4394 = ~w15122 & ~pi2678;
assign w4395 = pi3150 & w10992;
assign w4396 = w11383 & w17190;
assign w4397 = (pi0812 & ~w13509) | (pi0812 & w6842) | (~w13509 & w6842);
assign w4398 = ~w12460 & w17067;
assign w4399 = pi1858 & ~pi0274;
assign w4400 = ~w816 & ~w9630;
assign w4401 = w12237 & w10527;
assign w4402 = ~pi2396 & w13204;
assign w4403 = w968 & ~pi0288;
assign w4404 = ~w16383 & ~w9871;
assign w4405 = pi2435 & ~w3223;
assign w4406 = ~w9331 & ~w9999;
assign w4407 = pi0031 & ~w14148;
assign w4408 = pi2821 & ~w226;
assign w4409 = ~pi0286 & w2196;
assign w4410 = (~pi2911 & w5607) | (~pi2911 & w14251) | (w5607 & w14251);
assign w4411 = ~w17740 & ~w17298;
assign w4412 = (~pi0510 & w17577) | (~pi0510 & w9483) | (w17577 & w9483);
assign w4413 = ~w16830 & w12922;
assign w4414 = pi0147 & w8912;
assign w4415 = ~w14688 & w8109;
assign w4416 = ~w6898 & ~w12896;
assign w4417 = w8437 & w6018;
assign w4418 = ~w13120 & ~w3561;
assign w4419 = pi2255 & ~w11671;
assign w4420 = w13090 & w14342;
assign w4421 = ~w16581 & ~w16901;
assign w4422 = ~pi0688 & w9110;
assign w4423 = ~w3203 & pi1080;
assign w4424 = ~w12906 & ~w5606;
assign w4425 = ~pi2380 & w12755;
assign w4426 = ~w2315 & ~w6107;
assign w4427 = w14560 & pi0374;
assign w4428 = ~w1962 & pi1010;
assign w4429 = ~w5838 & ~w8136;
assign w4430 = ~pi3157 & w14753;
assign w4431 = ~pi1056 & w1126;
assign w4432 = ~w7844 & pi0599;
assign w4433 = pi3379 & w13367;
assign w4434 = w14109 & pi0418;
assign w4435 = w16699 & w758;
assign w4436 = pi2501 & ~w5274;
assign w4437 = pi1906 & ~w15271;
assign w4438 = w6649 & ~w1589;
assign w4439 = ~pi1693 & w317;
assign w4440 = ~pi3166 & w13570;
assign w4441 = ~pi2475 & w16041;
assign w4442 = w7077 & ~w16498;
assign w4443 = ~w15569 & ~w768;
assign w4444 = ~w2558 & w11062;
assign w4445 = ~w9986 & ~w10889;
assign w4446 = ~w709 & pi1281;
assign w4447 = ~w15503 & ~w17593;
assign w4448 = w10074 & w5108;
assign w4449 = ~pi3347 & w14918;
assign w4450 = ~w6034 & ~w11183;
assign w4451 = pi1822 & ~w653;
assign w4452 = pi2403 & ~w412;
assign w4453 = ~w14854 & ~w11374;
assign w4454 = ~w15722 & ~w14861;
assign w4455 = ~pi0122 & w9284;
assign w4456 = w2341 & ~w6647;
assign w4457 = ~w8619 & ~w2217;
assign w4458 = ~pi0811 & w1147;
assign w4459 = w715 & w4560;
assign w4460 = w2725 & ~w7707;
assign w4461 = ~w14560 & pi0246;
assign w4462 = ~pi0908 & w543;
assign w4463 = pi1803 & ~w5457;
assign w4464 = pi1794 & ~w435;
assign w4465 = ~w11390 & ~w13760;
assign w4466 = ~pi2296 & w5075;
assign w4467 = ~w5888 & ~w7632;
assign w4468 = ~w2320 & ~w10630;
assign w4469 = pi0507 & w9084;
assign w4470 = ~w13620 & ~w458;
assign w4471 = ~w9648 & ~w4182;
assign w4472 = w13231 & ~w7020;
assign w4473 = ~pi3295 & w17935;
assign w4474 = ~w17119 & ~w40;
assign w4475 = w9475 & w16058;
assign w4476 = ~w15190 & ~w4939;
assign w4477 = pi1963 & ~w14833;
assign w4478 = w18163 & pi0489;
assign w4479 = ~w2933 & ~w10223;
assign w4480 = ~w14648 & ~pi2724;
assign w4481 = pi2337 & ~w17683;
assign w4482 = pi2781 & ~w16815;
assign w4483 = pi1884 & ~w11406;
assign w4484 = pi1305 & ~w14094;
assign w4485 = ~w16506 & pi1264;
assign w4486 = w2206 & ~w170;
assign w4487 = ~pi2216 & w11313;
assign w4488 = ~pi2176 & w5384;
assign w4489 = ~pi0694 & w9110;
assign w4490 = ~pi0961 & w12197;
assign w4491 = ~w9004 & ~w15849;
assign w4492 = pi2962 & w8003;
assign w4493 = w6649 & ~w13693;
assign w4494 = ~w3660 & ~w3465;
assign w4495 = w13509 & w14502;
assign w4496 = pi1320 & pi1345;
assign w4497 = pi1783 & ~w16995;
assign w4498 = ~w18095 & ~w10212;
assign w4499 = w10818 & ~w5645;
assign w4500 = pi1534 & w13753;
assign w4501 = ~w525 & ~w13367;
assign w4502 = (pi0822 & ~w13509) | (pi0822 & w4897) | (~w13509 & w4897);
assign w4503 = (~pi0262 & ~w325) | (~pi0262 & w11167) | (~w325 & w11167);
assign w4504 = ~w14648 & ~pi2825;
assign w4505 = ~w6486 & ~w15832;
assign w4506 = pi2247 & ~w18123;
assign w4507 = ~pi3054 & w11406;
assign w4508 = w14244 & w3167;
assign w4509 = w13509 & w17284;
assign w4510 = ~w3957 & ~w9749;
assign w4511 = ~pi0778 & w6200;
assign w4512 = ~pi0333 & w2196;
assign w4513 = (pi1072 & ~w13509) | (pi1072 & w11155) | (~w13509 & w11155);
assign w4514 = ~w4312 & w11879;
assign w4515 = w6857 & w9519;
assign w4516 = ~w3203 & pi0998;
assign w4517 = pi1367 & w5043;
assign w4518 = ~w14691 & w5477;
assign w4519 = ~pi0483 & pi3407;
assign w4520 = ~w17611 & ~w14987;
assign w4521 = ~w17132 & ~w10985;
assign w4522 = ~w9154 & w6760;
assign w4523 = ~w15122 & ~pi2513;
assign w4524 = ~w4258 & ~w5340;
assign w4525 = ~w16011 & ~w956;
assign w4526 = ~pi3172 & pi3207;
assign w4527 = pi1371 & ~pi2913;
assign w4528 = ~w14560 & pi0234;
assign w4529 = pi2291 & ~w4508;
assign w4530 = w13964 & w2004;
assign w4531 = ~w12099 & ~w7822;
assign w4532 = ~pi0831 & w93;
assign w4533 = ~w12853 & ~w1809;
assign w4534 = w15842 & pi1354;
assign w4535 = ~w8221 & w1179;
assign w4536 = ~w7917 & ~w12394;
assign w4537 = ~w6386 & ~w14708;
assign w4538 = ~w10361 & ~w9940;
assign w4539 = ~w6024 & ~w13955;
assign w4540 = pi2376 & ~w18123;
assign w4541 = pi0378 & w871;
assign w4542 = ~w16506 & pi1150;
assign w4543 = pi2640 & ~w3555;
assign w4544 = ~pi0202 & ~w9954;
assign w4545 = ~pi1838 & ~w3223;
assign w4546 = w9440 & pi0143;
assign w4547 = pi2705 & ~w5274;
assign w4548 = ~w885 & ~w15338;
assign w4549 = (pi1023 & ~w13509) | (pi1023 & w8284) | (~w13509 & w8284);
assign w4550 = pi0102 & w3748;
assign w4551 = ~w7846 & ~w8124;
assign w4552 = w9720 & pi1752;
assign w4553 = ~w2725 & pi0789;
assign w4554 = ~pi1271 & ~pi3024;
assign w4555 = ~w13231 & pi0993;
assign w4556 = ~pi3171 & w15048;
assign w4557 = ~pi2649 & w15122;
assign w4558 = (pi0346 & w6195) | (pi0346 & w10834) | (w6195 & w10834);
assign w4559 = (pi0377 & w5560) | (pi0377 & w5317) | (w5560 & w5317);
assign w4560 = w13720 & w10747;
assign w4561 = pi2864 & w14148;
assign w4562 = (pi0854 & ~w13509) | (pi0854 & w6113) | (~w13509 & w6113);
assign w4563 = w13509 & w1422;
assign w4564 = pi2539 & w14148;
assign w4565 = ~pi2857 & w15122;
assign w4566 = ~w12392 & ~w16008;
assign w4567 = ~w10279 & ~w9489;
assign w4568 = (~w9737 & ~w14073) | (~w9737 & w14759) | (~w14073 & w14759);
assign w4569 = ~w13333 & ~w15788;
assign w4570 = ~w16417 & ~w6823;
assign w4571 = w709 & pi1899;
assign w4572 = pi2141 & ~w15883;
assign w4573 = pi1435 & ~w13753;
assign w4574 = pi1704 & ~w18497;
assign w4575 = ~w8588 & w9414;
assign w4576 = ~w6902 & ~w17075;
assign w4577 = ~pi0629 & w14641;
assign w4578 = ~pi0264 & w4058;
assign w4579 = ~w4513 & ~w15086;
assign w4580 = pi2805 & ~w6463;
assign w4581 = ~w709 & ~w1638;
assign w4582 = ~pi3159 & w17387;
assign w4583 = ~w5453 & ~pi1804;
assign w4584 = ~w10601 & ~w11934;
assign w4585 = pi1216 & ~w17367;
assign w4586 = ~w240 & ~w3974;
assign w4587 = pi1723 & ~w8113;
assign w4588 = (pi1376 & ~w11505) | (pi1376 & w5760) | (~w11505 & w5760);
assign w4589 = pi0017 & ~w3748;
assign w4590 = ~w12919 & w2810;
assign w4591 = w13509 & w6368;
assign w4592 = ~pi3124 & ~w5855;
assign w4593 = ~w16285 & w14680;
assign w4594 = ~pi2288 & w16041;
assign w4595 = ~w10353 & ~w4898;
assign w4596 = pi1249 & w11655;
assign w4597 = ~pi0832 & w93;
assign w4598 = ~pi0506 & ~pi1149;
assign w4599 = pi1858 & ~w968;
assign w4600 = pi2466 & ~w14524;
assign w4601 = (pi0868 & ~w13509) | (pi0868 & w9343) | (~w13509 & w9343);
assign w4602 = w15808 & ~w9852;
assign w4603 = ~pi1975 & w15122;
assign w4604 = w15808 & ~w4179;
assign w4605 = pi1617 & ~w16922;
assign w4606 = ~w18386 & ~w6115;
assign w4607 = pi3030 & ~w16502;
assign w4608 = pi3160 & ~pi3474;
assign w4609 = ~w2341 & pi0843;
assign w4610 = ~w2925 & ~w1544;
assign w4611 = w9462 & w9771;
assign w4612 = pi1930 & ~w11735;
assign w4613 = w9720 & pi1720;
assign w4614 = ~w6892 & ~w6492;
assign w4615 = pi1882 & ~w6463;
assign w4616 = ~w16689 & ~w17651;
assign w4617 = pi0010 & ~w14148;
assign w4618 = w1962 & ~w7449;
assign w4619 = ~pi3166 & w17669;
assign w4620 = pi2638 & ~w9504;
assign w4621 = ~w10046 & ~w8962;
assign w4622 = ~w15491 & ~w4335;
assign w4623 = ~pi2201 & w9340;
assign w4624 = w5189 & ~w16498;
assign w4625 = ~w14228 & ~pi0982;
assign w4626 = ~w6990 & ~w14997;
assign w4627 = w14009 & w8768;
assign w4628 = pi1215 & pi3220;
assign w4629 = ~pi0329 & w4058;
assign w4630 = ~pi1760 & ~pi3153;
assign w4631 = w13509 & w1850;
assign w4632 = w15808 & ~w17513;
assign w4633 = ~w7627 & w3319;
assign w4634 = pi2317 & ~w4508;
assign w4635 = ~w14961 & ~w5053;
assign w4636 = ~pi0489 & ~pi1345;
assign w4637 = ~w12975 & w10129;
assign w4638 = w13840 & w17741;
assign w4639 = pi0027 & ~w14148;
assign w4640 = ~w13593 & ~w12901;
assign w4641 = pi1753 & ~pi3138;
assign w4642 = w17562 & pi2501;
assign w4643 = w6857 & w934;
assign w4644 = (pi0936 & ~w13509) | (pi0936 & w8667) | (~w13509 & w8667);
assign w4645 = ~w14206 & ~w5667;
assign w4646 = ~pi0830 & w93;
assign w4647 = w6360 & w283;
assign w4648 = (pi1033 & ~w13509) | (pi1033 & w5355) | (~w13509 & w5355);
assign w4649 = ~w12460 & w18030;
assign w4650 = (pi1066 & ~w13509) | (pi1066 & w1456) | (~w13509 & w1456);
assign w4651 = ~pi0518 & w15707;
assign w4652 = w14198 & w1992;
assign w4653 = w9161 & w11342;
assign w4654 = w16575 & w9204;
assign w4655 = ~w15874 & w1455;
assign w4656 = ~w14852 & ~w10763;
assign w4657 = w14109 & pi0422;
assign w4658 = ~pi3158 & ~pi3160;
assign w4659 = pi1343 & w9440;
assign w4660 = ~w4931 & ~w14652;
assign w4661 = ~pi3091 & w9504;
assign w4662 = ~w7385 & ~w7834;
assign w4663 = w6785 & ~w2587;
assign w4664 = pi2427 & ~w3223;
assign w4665 = ~pi3052 & w3555;
assign w4666 = ~w12224 & ~w7676;
assign w4667 = ~w17534 & ~w11743;
assign w4668 = pi0011 & ~w14148;
assign w4669 = (pi0565 & ~w13509) | (pi0565 & w8080) | (~w13509 & w8080);
assign w4670 = (pi1054 & ~w13509) | (pi1054 & w5004) | (~w13509 & w5004);
assign w4671 = (~w18096 & w8928) | (~w18096 & w2018) | (w8928 & w2018);
assign w4672 = pi0253 & w5274;
assign w4673 = ~w13156 & ~w3496;
assign w4674 = ~w14383 & w12772;
assign w4675 = (pi1102 & ~w13509) | (pi1102 & w9950) | (~w13509 & w9950);
assign w4676 = pi2692 & ~w6463;
assign w4677 = ~pi2975 & w11671;
assign w4678 = ~w376 & ~w15932;
assign w4679 = ~pi3349 & w17935;
assign w4680 = pi3005 & ~pi3165;
assign w4681 = ~w10563 & w17731;
assign w4682 = ~w16278 & pi0706;
assign w4683 = w17741 & w11060;
assign w4684 = pi1462 & w13753;
assign w4685 = ~pi3328 & w6448;
assign w4686 = w1494 & w11906;
assign w4687 = w13509 & w17531;
assign w4688 = w13509 & w17532;
assign w4689 = (pi1003 & ~w13509) | (pi1003 & w15900) | (~w13509 & w15900);
assign w4690 = w12040 & ~w3430;
assign w4691 = w7307 & w14940;
assign w4692 = ~w18487 & ~w5964;
assign w4693 = ~w4931 & ~w12329;
assign w4694 = ~pi2132 & w16041;
assign w4695 = ~pi0667 & w12197;
assign w4696 = ~w13187 & ~w2467;
assign w4697 = pi2544 & w14148;
assign w4698 = ~w12460 & w3755;
assign w4699 = ~w11381 & ~w13088;
assign w4700 = ~w2336 & ~w13701;
assign w4701 = ~pi1316 & ~w2325;
assign w4702 = ~w6195 & w5071;
assign w4703 = pi0263 & w7807;
assign w4704 = ~pi2490 & w17213;
assign w4705 = ~w14035 & ~w1238;
assign w4706 = ~w13771 & w5483;
assign w4707 = w7844 & ~w11978;
assign w4708 = (pi1888 & w2014) | (pi1888 & w15134) | (w2014 & w15134);
assign w4709 = pi0040 & ~w14148;
assign w4710 = ~w3000 & ~pi1882;
assign w4711 = ~w987 & w6252;
assign w4712 = pi3011 & ~w3987;
assign w4713 = w9440 & pi0175;
assign w4714 = w968 & ~pi0281;
assign w4715 = ~w6325 & ~w2500;
assign w4716 = ~pi2880 & w15122;
assign w4717 = ~w5208 & w14486;
assign w4718 = w13509 & w3070;
assign w4719 = pi0263 & w5113;
assign w4720 = pi2913 & ~w17729;
assign w4721 = pi2211 & ~w3223;
assign w4722 = ~pi0296 & w4058;
assign w4723 = ~pi2524 & w14148;
assign w4724 = ~pi3138 & w17669;
assign w4725 = (pi0947 & ~w13509) | (pi0947 & w5127) | (~w13509 & w5127);
assign w4726 = ~w11143 & ~w8384;
assign w4727 = ~w5829 & ~w17525;
assign w4728 = ~w3203 & pi0995;
assign w4729 = pi1582 & ~w14918;
assign w4730 = pi2246 & ~w9414;
assign w4731 = ~w13456 & ~w14270;
assign w4732 = ~pi3100 & w226;
assign w4733 = (pi0600 & ~w13509) | (pi0600 & w11979) | (~w13509 & w11979);
assign w4734 = (~pi0980 & ~w13509) | (~pi0980 & w3088) | (~w13509 & w3088);
assign w4735 = ~w16866 & ~w16229;
assign w4736 = ~w6785 & pi0865;
assign w4737 = ~pi3092 & w3555;
assign w4738 = ~w18509 & w12436;
assign w4739 = ~w14598 & ~w2468;
assign w4740 = (pi0370 & w6195) | (pi0370 & w4932) | (w6195 & w4932);
assign w4741 = ~pi3057 & w9243;
assign w4742 = ~w196 & ~w10511;
assign w4743 = pi1340 & w735;
assign w4744 = w384 & w14748;
assign w4745 = w17788 & w7924;
assign w4746 = w2584 & w4190;
assign w4747 = ~w5782 & w17359;
assign w4748 = ~w17151 & ~w3782;
assign w4749 = pi2357 & ~w412;
assign w4750 = w17747 & w12815;
assign w4751 = pi1244 & ~w11655;
assign w4752 = w13509 & w14007;
assign w4753 = ~pi3135 & w12427;
assign w4754 = ~w6883 & ~w17011;
assign w4755 = ~pi0784 & w543;
assign w4756 = ~w17534 & pi0137;
assign w4757 = ~pi3093 & w3555;
assign w4758 = ~w1930 & ~w11882;
assign w4759 = w14833 & w3515;
assign w4760 = ~pi2190 & w2151;
assign w4761 = ~w17234 & ~w18302;
assign w4762 = ~pi2786 & w15122;
assign w4763 = ~w15865 & ~w3752;
assign w4764 = ~pi3153 & ~pi3160;
assign w4765 = ~w9844 & w14911;
assign w4766 = w6277 & w6525;
assign w4767 = pi2942 & ~w6045;
assign w4768 = w1468 & w13224;
assign w4769 = (pi1139 & ~w5437) | (pi1139 & w2951) | (~w5437 & w2951);
assign w4770 = (pi1270 & ~w14158) | (pi1270 & w16457) | (~w14158 & w16457);
assign w4771 = pi2809 & ~w6463;
assign w4772 = ~pi0337 & ~pi0338;
assign w4773 = ~w296 & w9257;
assign w4774 = ~pi3096 & w261;
assign w4775 = w384 & w5134;
assign w4776 = (pi1311 & ~w14094) | (pi1311 & w9539) | (~w14094 & w9539);
assign w4777 = ~pi3103 & w16815;
assign w4778 = w15122 & ~pi2698;
assign w4779 = pi1683 & ~w7212;
assign w4780 = ~pi3084 & w11406;
assign w4781 = ~w17794 & ~w9801;
assign w4782 = pi2340 & ~w3223;
assign w4783 = ~w13252 & w6374;
assign w4784 = ~pi3335 & w16922;
assign w4785 = pi1455 & w13753;
assign w4786 = ~w12333 & ~w13310;
assign w4787 = pi0503 & pi0514;
assign w4788 = ~pi2424 & w13204;
assign w4789 = pi1795 & ~w9103;
assign w4790 = ~pi2094 & w12724;
assign w4791 = ~w6697 & pi0671;
assign w4792 = ~w9236 & ~w18014;
assign w4793 = ~w3797 & ~w16885;
assign w4794 = (pi0991 & ~w13509) | (pi0991 & w2394) | (~w13509 & w2394);
assign w4795 = pi3026 & ~pi3166;
assign w4796 = (~pi2913 & ~w1598) | (~pi2913 & w17158) | (~w1598 & w17158);
assign w4797 = w1962 & ~w14597;
assign w4798 = (pi0405 & w5560) | (pi0405 & w17254) | (w5560 & w17254);
assign w4799 = w7077 & ~w6922;
assign w4800 = w16634 & w8534;
assign w4801 = ~w6785 & pi0860;
assign w4802 = pi2386 & ~w18123;
assign w4803 = ~w15369 & ~w4131;
assign w4804 = w13509 & w1784;
assign w4805 = ~w4397 & ~w684;
assign w4806 = ~w6184 & ~w7925;
assign w4807 = ~w17222 & ~w13638;
assign w4808 = ~w16389 & ~w5597;
assign w4809 = ~w3844 & ~w12012;
assign w4810 = ~pi0912 & w12197;
assign w4811 = w5189 & ~w1340;
assign w4812 = pi0073 & ~w14148;
assign w4813 = ~w16131 & ~w2428;
assign w4814 = ~w5662 & ~w11109;
assign w4815 = ~pi3286 & w18259;
assign w4816 = pi2908 & ~pi3175;
assign w4817 = w902 & w15329;
assign w4818 = w5968 & w10038;
assign w4819 = (pi1892 & w2014) | (pi1892 & w7697) | (w2014 & w7697);
assign w4820 = ~pi2019 & w11688;
assign w4821 = ~pi3139 & w17993;
assign w4822 = pi2517 & ~w9504;
assign w4823 = pi1395 & ~w6853;
assign w4824 = pi2305 & ~w15883;
assign w4825 = w16278 & ~w15296;
assign w4826 = ~pi2387 & w12755;
assign w4827 = pi1432 & ~w6448;
assign w4828 = ~w2738 & w9061;
assign w4829 = w17562 & pi2561;
assign w4830 = ~w1573 & ~w12157;
assign w4831 = (pi0794 & ~w13509) | (pi0794 & w1134) | (~w13509 & w1134);
assign w4832 = (~w14698 & ~w14073) | (~w14698 & w2931) | (~w14073 & w2931);
assign w4833 = pi0056 & pi0055;
assign w4834 = ~pi3328 & w16922;
assign w4835 = w12284 & w4263;
assign w4836 = w17782 & w10519;
assign w4837 = ~w1861 & ~w1928;
assign w4838 = ~pi2945 & pi3199;
assign w4839 = (pi0914 & ~w13509) | (pi0914 & w18458) | (~w13509 & w18458);
assign w4840 = w604 & w2549;
assign w4841 = ~pi1828 & w9165;
assign w4842 = w2725 & ~w3430;
assign w4843 = w9864 & w14304;
assign w4844 = ~w17483 & ~w14239;
assign w4845 = ~w3562 & ~w4530;
assign w4846 = ~w7752 & ~w16509;
assign w4847 = w11209 & ~w8316;
assign w4848 = ~w13857 & ~w13126;
assign w4849 = pi2088 & ~w4420;
assign w4850 = (w5855 & w1295) | (w5855 & w7371) | (w1295 & w7371);
assign w4851 = pi2592 & ~w5274;
assign w4852 = ~w5634 & ~w2032;
assign w4853 = ~w18048 & w16653;
assign w4854 = w16047 & w11784;
assign w4855 = ~pi0567 & w11739;
assign w4856 = ~pi0952 & w11739;
assign w4857 = ~w8171 & pi1204;
assign w4858 = ~pi2022 & w7455;
assign w4859 = ~pi3311 & w18259;
assign w4860 = ~pi0768 & w6200;
assign w4861 = w7077 & ~w10947;
assign w4862 = ~pi0145 & ~pi0195;
assign w4863 = ~w17880 & ~w14394;
assign w4864 = ~w17239 & ~w2792;
assign w4865 = ~w15471 & ~w3950;
assign w4866 = pi2900 & ~w226;
assign w4867 = pi1167 & w13509;
assign w4868 = ~w4592 & ~w5842;
assign w4869 = ~w8142 & ~w6533;
assign w4870 = ~w16806 & ~w10141;
assign w4871 = pi2531 & w15191;
assign w4872 = (pi0746 & ~w13509) | (pi0746 & w5479) | (~w13509 & w5479);
assign w4873 = ~pi3354 & w7090;
assign w4874 = w934 & pi0437;
assign w4875 = pi1616 & w13753;
assign w4876 = w5189 & ~w12800;
assign w4877 = pi1487 & w13753;
assign w4878 = w16278 & ~w2587;
assign w4879 = ~w7089 & ~w11373;
assign w4880 = ~pi1218 & pi2486;
assign w4881 = ~w15282 & ~w755;
assign w4882 = ~w12040 & pi0681;
assign w4883 = ~pi2221 & w11313;
assign w4884 = w1391 & ~w14465;
assign w4885 = pi0110 & w9284;
assign w4886 = w7121 & w6165;
assign w4887 = pi1870 & ~w458;
assign w4888 = ~w16575 & w4250;
assign w4889 = ~w1937 & ~w4217;
assign w4890 = ~pi3154 & w11132;
assign w4891 = ~pi0595 & w12825;
assign w4892 = ~pi2969 & w3479;
assign w4893 = (pi0604 & ~w13509) | (pi0604 & w15283) | (~w13509 & w15283);
assign w4894 = ~w12460 & w9523;
assign w4895 = ~pi0497 & ~pi1345;
assign w4896 = w12460 & w5168;
assign w4897 = ~w7077 & pi0822;
assign w4898 = pi3162 & w3987;
assign w4899 = pi3191 & w8042;
assign w4900 = ~w7884 & ~w10197;
assign w4901 = ~w15916 & w703;
assign w4902 = ~w16838 & ~w1230;
assign w4903 = ~w10633 & ~w11916;
assign w4904 = pi1256 & w11655;
assign w4905 = ~w1225 & w3125;
assign w4906 = ~pi1255 & w11655;
assign w4907 = w7703 & w3063;
assign w4908 = (pi0899 & ~w13509) | (pi0899 & w9120) | (~w13509 & w9120);
assign w4909 = ~pi2323 & w8617;
assign w4910 = ~w17218 & ~w8289;
assign w4911 = (~w14403 & ~w7692) | (~w14403 & w9013) | (~w7692 & w9013);
assign w4912 = ~w9991 & w13670;
assign w4913 = ~w4192 & ~w16813;
assign w4914 = w1368 & pi0395;
assign w4915 = ~pi3084 & w3555;
assign w4916 = pi1521 & ~w14918;
assign w4917 = ~w17677 & ~w10400;
assign w4918 = ~w14428 & ~w4495;
assign w4919 = w12460 & w9305;
assign w4920 = ~pi1355 & w15842;
assign w4921 = pi1369 & ~pi2913;
assign w4922 = ~w6263 & w1326;
assign w4923 = ~w4178 & ~w9268;
assign w4924 = ~pi3328 & w6072;
assign w4925 = ~w8125 & w16822;
assign w4926 = w539 & ~w728;
assign w4927 = w12188 & w4731;
assign w4928 = pi2945 & ~pi3199;
assign w4929 = pi0030 & ~w14148;
assign w4930 = ~w14259 & ~w14711;
assign w4931 = w5968 & pi1858;
assign w4932 = w14560 & pi0370;
assign w4933 = ~w17326 & ~w13367;
assign w4934 = pi1140 & pi2941;
assign w4935 = ~w16506 & pi1192;
assign w4936 = w9476 & w15081;
assign w4937 = pi0019 & ~w3748;
assign w4938 = pi1327 & pi1345;
assign w4939 = ~pi0704 & w3106;
assign w4940 = pi1337 & pi0260;
assign w4941 = ~w4667 & ~w13394;
assign w4942 = pi2031 & ~w17646;
assign w4943 = ~w17346 & w18185;
assign w4944 = w11345 & w15021;
assign w4945 = ~pi3153 & w1843;
assign w4946 = ~w11673 & ~w16940;
assign w4947 = ~pi0066 & w922;
assign w4948 = pi2165 & ~w9414;
assign w4949 = pi3082 & w3555;
assign w4950 = pi1722 & ~pi3133;
assign w4951 = w9440 & pi0163;
assign w4952 = ~w10308 & w15675;
assign w4953 = ~w12946 & w17097;
assign w4954 = pi0045 & ~pi0048;
assign w4955 = pi1653 & ~w13753;
assign w4956 = ~pi1212 & pi1221;
assign w4957 = w4786 & w970;
assign w4958 = ~pi1833 & w2151;
assign w4959 = ~w11509 & ~w15059;
assign w4960 = ~pi0281 & w2196;
assign w4961 = ~w13746 & ~w3532;
assign w4962 = pi0037 & ~w3748;
assign w4963 = w6857 & w14816;
assign w4964 = w14158 & w485;
assign w4965 = ~w5517 & w8757;
assign w4966 = w10189 & pi0382;
assign w4967 = pi2298 & ~w15883;
assign w4968 = w8337 & pi3358;
assign w4969 = ~w14842 & w7323;
assign w4970 = ~w818 & ~w10073;
assign w4971 = ~w15795 & ~w4199;
assign w4972 = pi0130 & ~pi0153;
assign w4973 = w17562 & pi1817;
assign w4974 = ~w5025 & ~w18427;
assign w4975 = pi2324 & ~w4508;
assign w4976 = ~w17684 & ~w1281;
assign w4977 = ~w1791 & w12687;
assign w4978 = w2609 & w4763;
assign w4979 = (pi0403 & w5560) | (pi0403 & w14649) | (w5560 & w14649);
assign w4980 = pi1563 & ~w13753;
assign w4981 = w4364 & ~pi0435;
assign w4982 = pi1373 & w657;
assign w4983 = ~w5232 & ~w16396;
assign w4984 = ~w16611 & w11591;
assign w4985 = pi2545 & w605;
assign w4986 = w13509 & w2831;
assign w4987 = ~pi3321 & w9781;
assign w4988 = pi1209 & ~pi1182;
assign w4989 = ~w15504 & ~w14294;
assign w4990 = pi1599 & w13753;
assign w4991 = w7703 & w12473;
assign w4992 = w6785 & ~w6922;
assign w4993 = ~w17705 & ~w7153;
assign w4994 = ~w11361 & ~w7421;
assign w4995 = ~w6604 & ~w9032;
assign w4996 = ~w517 & ~w17098;
assign w4997 = pi2594 & ~w8304;
assign w4998 = pi1807 & ~w8097;
assign w4999 = ~w2095 & w18561;
assign w5000 = ~w3054 & w14969;
assign w5001 = (pi0662 & ~w13509) | (pi0662 & w14531) | (~w13509 & w14531);
assign w5002 = pi1575 & ~w16922;
assign w5003 = ~pi0826 & w93;
assign w5004 = ~w17248 & pi1054;
assign w5005 = ~pi2142 & w12941;
assign w5006 = ~pi2035 & w7455;
assign w5007 = ~w13583 & ~w8707;
assign w5008 = pi3039 & w16502;
assign w5009 = ~w12040 & pi0696;
assign w5010 = (~w1542 & ~w5517) | (~w1542 & w6703) | (~w5517 & w6703);
assign w5011 = w6785 & ~w15296;
assign w5012 = ~w5855 & w3442;
assign w5013 = ~w6953 & ~w11246;
assign w5014 = w3674 & w11142;
assign w5015 = w3333 & pi0506;
assign w5016 = w17248 & w11302;
assign w5017 = ~w7538 & w5225;
assign w5018 = (pi1783 & w7215) | (pi1783 & w12953) | (w7215 & w12953);
assign w5019 = pi3369 & w15974;
assign w5020 = ~pi2005 & w3019;
assign w5021 = ~pi0178 & pi0190;
assign w5022 = w7307 & w10517;
assign w5023 = w539 & ~w13386;
assign w5024 = ~pi2063 & w8617;
assign w5025 = ~pi2266 & w13065;
assign w5026 = ~w18028 & ~w13493;
assign w5027 = pi1486 & w13753;
assign w5028 = w539 & ~w7640;
assign w5029 = (pi1019 & ~w13509) | (pi1019 & w8800) | (~w13509 & w8800);
assign w5030 = w13509 & w12141;
assign w5031 = pi1238 & pi1257;
assign w5032 = ~w10320 & ~w13216;
assign w5033 = ~w5453 & ~pi1799;
assign w5034 = (pi0768 & ~w13509) | (pi0768 & w2045) | (~w13509 & w2045);
assign w5035 = ~w3243 & pi0315;
assign w5036 = pi1719 & ~w8113;
assign w5037 = pi1509 & ~w13753;
assign w5038 = ~pi3314 & w14918;
assign w5039 = ~pi3313 & w9781;
assign w5040 = w7844 & ~w305;
assign w5041 = w11383 & w15820;
assign w5042 = ~w10056 & w12531;
assign w5043 = pi2968 & ~w15476;
assign w5044 = pi1504 & ~w13753;
assign w5045 = (pi0785 & ~w13509) | (pi0785 & w2303) | (~w13509 & w2303);
assign w5046 = ~w7213 & ~w2133;
assign w5047 = ~w1982 & w5220;
assign w5048 = ~w5453 & ~w2024;
assign w5049 = ~pi0560 & w11739;
assign w5050 = pi1954 & ~w14833;
assign w5051 = w17562 & pi1853;
assign w5052 = (pi0776 & ~w13509) | (pi0776 & w6164) | (~w13509 & w6164);
assign w5053 = ~pi3042 & w18559;
assign w5054 = ~w14228 & pi0620;
assign w5055 = ~pi1223 & w5566;
assign w5056 = pi1457 & w13753;
assign w5057 = ~w15122 & ~pi2833;
assign w5058 = ~w10703 & ~w3309;
assign w5059 = pi3163 & w11272;
assign w5060 = ~w13231 & pi0913;
assign w5061 = pi2872 & w15191;
assign w5062 = ~pi3097 & w226;
assign w5063 = ~w456 & ~w8081;
assign w5064 = ~pi0559 & w11739;
assign w5065 = w2971 & w4534;
assign w5066 = ~w11984 & ~w3053;
assign w5067 = w10189 & ~pi0471;
assign w5068 = pi1491 & w13753;
assign w5069 = ~pi3293 & w17935;
assign w5070 = ~w5453 & ~pi1760;
assign w5071 = ~w14560 & pi0210;
assign w5072 = ~w13920 & ~w10021;
assign w5073 = ~w14164 & ~w12092;
assign w5074 = ~w9598 & ~w6347;
assign w5075 = w14138 & w5410;
assign w5076 = ~pi3436 & w15036;
assign w5077 = w7703 & w841;
assign w5078 = pi3083 & pi3129;
assign w5079 = w6857 & w4361;
assign w5080 = (pi1013 & ~w13509) | (pi1013 & w11970) | (~w13509 & w11970);
assign w5081 = (pi0361 & w6195) | (pi0361 & w14091) | (w6195 & w14091);
assign w5082 = w11952 & w2892;
assign w5083 = w11383 & w5752;
assign w5084 = ~w5164 & ~w1903;
assign w5085 = ~w10336 & ~w1593;
assign w5086 = pi2486 & ~w7212;
assign w5087 = pi1898 & ~w15036;
assign w5088 = ~w5993 & w18358;
assign w5089 = w16506 & ~w2776;
assign w5090 = ~w10798 & ~w9585;
assign w5091 = ~pi2967 & pi3029;
assign w5092 = ~w8418 & w16789;
assign w5093 = pi1337 & w6659;
assign w5094 = ~pi1685 & pi3246;
assign w5095 = ~pi2990 & w6225;
assign w5096 = ~w2301 & ~w14685;
assign w5097 = pi2525 & ~w13236;
assign w5098 = w12460 & w2153;
assign w5099 = ~w7212 & ~w11037;
assign w5100 = ~pi2444 & w9340;
assign w5101 = ~w10669 & ~w3630;
assign w5102 = ~w2123 & ~w12246;
assign w5103 = w13509 & w7818;
assign w5104 = ~w8314 & ~w4795;
assign w5105 = w5189 & ~w6922;
assign w5106 = (pi0997 & ~w13509) | (pi0997 & w1881) | (~w13509 & w1881);
assign w5107 = ~pi1842 & w12755;
assign w5108 = ~w5020 & ~w15910;
assign w5109 = ~pi0582 & w795;
assign w5110 = ~w9708 & ~w8694;
assign w5111 = ~w2417 & ~w11244;
assign w5112 = ~w13231 & pi1096;
assign w5113 = (w18583 & ~w12460) | (w18583 & w15548) | (~w12460 & w15548);
assign w5114 = ~w18554 & ~w9048;
assign w5115 = ~w15129 & ~w15884;
assign w5116 = w4655 & w2969;
assign w5117 = ~pi1106 & w3106;
assign w5118 = pi1650 & ~w13753;
assign w5119 = w13509 & w18529;
assign w5120 = w17248 & ~w17513;
assign w5121 = ~w9245 & ~w8333;
assign w5122 = ~w9021 & w6561;
assign w5123 = ~w3273 & ~w3959;
assign w5124 = ~w13834 & w5468;
assign w5125 = ~pi3150 & w1843;
assign w5126 = pi1542 & w13753;
assign w5127 = ~w17248 & pi0947;
assign w5128 = pi2625 & ~w16815;
assign w5129 = w16878 & w18162;
assign w5130 = w13509 & w14049;
assign w5131 = ~pi0754 & w17490;
assign w5132 = ~pi3142 & w14753;
assign w5133 = w4717 & w10686;
assign w5134 = w5453 & pi2856;
assign w5135 = ~pi2446 & w5384;
assign w5136 = ~pi3153 & w4310;
assign w5137 = ~w3777 & ~w16424;
assign w5138 = ~w17665 & ~w11053;
assign w5139 = ~pi3094 & w9504;
assign w5140 = ~pi2328 & w12941;
assign w5141 = w9514 & w9873;
assign w5142 = pi1727 & w1924;
assign w5143 = pi0247 & w5274;
assign w5144 = pi1405 & ~pi1966;
assign w5145 = ~pi1841 & w3019;
assign w5146 = w13509 & w1852;
assign w5147 = pi2633 & ~w9504;
assign w5148 = ~w11438 & ~w16608;
assign w5149 = ~w9886 & ~w1759;
assign w5150 = ~w9574 & ~w646;
assign w5151 = w6785 & ~w2776;
assign w5152 = pi0250 & w1516;
assign w5153 = pi1527 & ~w14918;
assign w5154 = ~w2014 & w14240;
assign w5155 = ~w17735 & ~w8202;
assign w5156 = w8383 & ~w13818;
assign w5157 = ~w1739 & ~w8156;
assign w5158 = ~w2980 & w2278;
assign w5159 = (~pi0277 & ~w6857) | (~pi0277 & w16126) | (~w6857 & w16126);
assign w5160 = w13509 & w14228;
assign w5161 = w16420 & w1092;
assign w5162 = (pi1089 & ~w13509) | (pi1089 & w8583) | (~w13509 & w8583);
assign w5163 = ~w14454 & w14981;
assign w5164 = (pi0647 & ~w13509) | (pi0647 & w12195) | (~w13509 & w12195);
assign w5165 = w2341 & ~w2741;
assign w5166 = pi1132 & ~w17391;
assign w5167 = pi1654 & ~w6072;
assign w5168 = w9440 & pi0131;
assign w5169 = w8789 & pi0406;
assign w5170 = ~w8204 & w2460;
assign w5171 = pi1537 & ~w17935;
assign w5172 = ~w9580 & ~w1349;
assign w5173 = w384 & w623;
assign w5174 = (pi0343 & w6195) | (pi0343 & w13927) | (w6195 & w13927);
assign w5175 = (pi0684 & ~w13509) | (pi0684 & w10392) | (~w13509 & w10392);
assign w5176 = ~w5533 & w3987;
assign w5177 = (pi0360 & w5560) | (pi0360 & w15581) | (w5560 & w15581);
assign w5178 = w3203 & ~w12800;
assign w5179 = ~w1962 & pi0650;
assign w5180 = (pi0598 & ~w13509) | (pi0598 & w15601) | (~w13509 & w15601);
assign w5181 = ~w16506 & pi1218;
assign w5182 = ~pi1154 & w13509;
assign w5183 = pi0069 & ~w14148;
assign w5184 = ~w7377 & ~w7442;
assign w5185 = ~pi3347 & w18259;
assign w5186 = pi1850 & ~w12558;
assign w5187 = ~w11907 & ~w8841;
assign w5188 = w3243 & pi0083;
assign w5189 = w15907 & w6676;
assign w5190 = ~pi2967 & w14446;
assign w5191 = w15842 & pi2555;
assign w5192 = w5466 & w17093;
assign w5193 = ~pi1252 & pi3228;
assign w5194 = pi3112 & ~w16502;
assign w5195 = ~pi0639 & w3791;
assign w5196 = ~w2238 & w15217;
assign w5197 = w291 & ~w11806;
assign w5198 = ~w4080 & w6522;
assign w5199 = (pi0778 & ~w13509) | (pi0778 & w12434) | (~w13509 & w12434);
assign w5200 = ~w2341 & pi0842;
assign w5201 = w3243 & pi0338;
assign w5202 = w13509 & w11278;
assign w5203 = ~w11913 & ~w4529;
assign w5204 = w1391 & ~w6033;
assign w5205 = pi2547 & w605;
assign w5206 = pi1337 & ~pi0298;
assign w5207 = ~pi3117 & pi3207;
assign w5208 = w7307 & w10905;
assign w5209 = ~w7291 & ~w8835;
assign w5210 = pi3133 & w3987;
assign w5211 = w14560 & pi0348;
assign w5212 = ~w2319 & ~w1609;
assign w5213 = w13509 & w699;
assign w5214 = w4846 & w15736;
assign w5215 = ~pi2112 & w12755;
assign w5216 = ~pi1054 & w1126;
assign w5217 = ~pi1161 & w678;
assign w5218 = w735 & pi3177;
assign w5219 = ~w1368 & ~pi0471;
assign w5220 = (~w10678 & ~w5517) | (~w10678 & w10525) | (~w5517 & w10525);
assign w5221 = ~w1213 & ~w1243;
assign w5222 = ~w2701 & w11135;
assign w5223 = w553 & ~pi1303;
assign w5224 = pi2904 & ~w5274;
assign w5225 = ~w9704 & ~w9360;
assign w5226 = ~pi2283 & w5075;
assign w5227 = ~pi1120 & w1126;
assign w5228 = ~w14388 & ~w4110;
assign w5229 = ~w709 & pi1277;
assign w5230 = ~w10779 & ~w2898;
assign w5231 = ~w7180 & ~w13444;
assign w5232 = (pi0318 & w3055) | (pi0318 & w9111) | (w3055 & w9111);
assign w5233 = ~pi0774 & w6200;
assign w5234 = w13509 & w8748;
assign w5235 = ~w6487 & w18049;
assign w5236 = ~w15137 & ~w9967;
assign w5237 = ~w12040 & pi0688;
assign w5238 = ~w10748 & ~w11101;
assign w5239 = ~w4020 & ~w3671;
assign w5240 = ~pi3169 & w17387;
assign w5241 = ~w16086 & ~w16557;
assign w5242 = ~pi3087 & w6463;
assign w5243 = ~w5000 & w8320;
assign w5244 = ~w13367 & ~w1648;
assign w5245 = pi1880 & ~w261;
assign w5246 = pi3143 & ~pi3157;
assign w5247 = ~pi1076 & w795;
assign w5248 = ~w7844 & pi0900;
assign w5249 = (pi1189 & ~w13509) | (pi1189 & w12592) | (~w13509 & w12592);
assign w5250 = pi1637 & ~w18259;
assign w5251 = ~w4934 & ~w16676;
assign w5252 = w7844 & ~w12800;
assign w5253 = ~pi3138 & w15839;
assign w5254 = pi2077 & ~w17683;
assign w5255 = pi2187 & ~w11735;
assign w5256 = ~pi2846 & w14148;
assign w5257 = pi2847 & w14148;
assign w5258 = w5491 & w11006;
assign w5259 = ~w6697 & pi0668;
assign w5260 = w13509 & w3052;
assign w5261 = (w2460 & ~w384) | (w2460 & w15192) | (~w384 & w15192);
assign w5262 = w5383 & w735;
assign w5263 = ~w5560 & w2620;
assign w5264 = ~w17620 & ~w14958;
assign w5265 = w1912 & w7610;
assign w5266 = pi1578 & ~w14918;
assign w5267 = pi0171 & ~pi0177;
assign w5268 = ~w14213 & w12959;
assign w5269 = ~pi3133 & w14753;
assign w5270 = ~w8997 & ~w5781;
assign w5271 = pi2861 & w15191;
assign w5272 = w7844 & ~w2741;
assign w5273 = w9720 & pi1668;
assign w5274 = pi1858 & ~w6523;
assign w5275 = ~w16918 & ~w6914;
assign w5276 = ~w18007 & ~w14862;
assign w5277 = w16506 & ~w17210;
assign w5278 = ~pi3101 & w16815;
assign w5279 = ~pi1832 & ~w14524;
assign w5280 = ~pi3164 & w3982;
assign w5281 = (pi0829 & ~w13509) | (pi0829 & w11327) | (~w13509 & w11327);
assign w5282 = ~w1186 & ~w11426;
assign w5283 = ~w5453 & ~pi1801;
assign w5284 = w17768 & w15114;
assign w5285 = ~pi3162 & w15839;
assign w5286 = ~w15654 & ~w3904;
assign w5287 = ~w4803 & pi2920;
assign w5288 = (pi0615 & ~w13509) | (pi0615 & w12997) | (~w13509 & w12997);
assign w5289 = (pi0656 & ~w13509) | (pi0656 & w9945) | (~w13509 & w9945);
assign w5290 = w16506 & pi2955;
assign w5291 = (pi0884 & ~w13509) | (pi0884 & w1781) | (~w13509 & w1781);
assign w5292 = ~w1598 & ~w3400;
assign w5293 = ~w13812 & pi1337;
assign w5294 = ~pi3017 & ~pi3207;
assign w5295 = w5453 & pi2901;
assign w5296 = ~pi1907 & w9340;
assign w5297 = ~w2860 & ~w16096;
assign w5298 = w7703 & w10151;
assign w5299 = ~w10718 & w11186;
assign w5300 = w13509 & w2274;
assign w5301 = w13509 & w13129;
assign w5302 = ~w6286 & ~w742;
assign w5303 = ~pi3413 & w15036;
assign w5304 = ~w18429 & ~w128;
assign w5305 = ~w3058 & ~w8260;
assign w5306 = w11383 & w2888;
assign w5307 = pi2222 & ~w11735;
assign w5308 = w6359 & w14026;
assign w5309 = pi2325 & ~w18123;
assign w5310 = ~pi0067 & w922;
assign w5311 = ~w18444 & ~w6704;
assign w5312 = ~w5901 & w10588;
assign w5313 = ~pi0869 & w15707;
assign w5314 = ~w13392 & ~w7937;
assign w5315 = w2341 & ~w16498;
assign w5316 = pi2347 & ~w15883;
assign w5317 = w1368 & pi0377;
assign w5318 = ~w3055 & w5201;
assign w5319 = w14648 & ~pi2609;
assign w5320 = ~w11799 & ~w15457;
assign w5321 = w2341 & ~w4043;
assign w5322 = pi3170 & w10389;
assign w5323 = w14679 & w15158;
assign w5324 = ~pi3087 & w9504;
assign w5325 = pi0094 & w3748;
assign w5326 = ~pi2256 & w13065;
assign w5327 = pi1518 & w13753;
assign w5328 = ~w3391 & ~w3692;
assign w5329 = ~w9666 & w12382;
assign w5330 = w13509 & w15004;
assign w5331 = ~w13460 & ~w13490;
assign w5332 = ~w8417 & w3241;
assign w5333 = ~w13231 & pi0561;
assign w5334 = ~w7300 & ~w12928;
assign w5335 = w13509 & w2222;
assign w5336 = ~w16278 & pi0716;
assign w5337 = w13509 & w15006;
assign w5338 = w13539 & w5251;
assign w5339 = w9748 & w11754;
assign w5340 = ~w9746 & w11755;
assign w5341 = w3596 & w15072;
assign w5342 = ~w7155 & ~w17923;
assign w5343 = ~w17891 & ~w13219;
assign w5344 = ~w18238 & w8208;
assign w5345 = ~w17136 & ~w15422;
assign w5346 = ~w12375 & ~w1347;
assign w5347 = ~w13367 & ~w3311;
assign w5348 = ~w5562 & ~w15643;
assign w5349 = ~w13669 & ~w12605;
assign w5350 = ~pi2150 & w13065;
assign w5351 = ~pi3098 & w11406;
assign w5352 = (~w10463 & ~w5517) | (~w10463 & w4391) | (~w5517 & w4391);
assign w5353 = ~w709 & ~pi1290;
assign w5354 = pi3141 & w10389;
assign w5355 = ~w15808 & pi1033;
assign w5356 = ~w11478 & ~w2347;
assign w5357 = w13840 & pi1699;
assign w5358 = ~pi3340 & w6448;
assign w5359 = w10772 & w17455;
assign w5360 = ~w13011 & ~w16397;
assign w5361 = ~w8588 & w15883;
assign w5362 = ~w14228 & pi0625;
assign w5363 = pi1562 & ~w18259;
assign w5364 = pi2995 & ~w3987;
assign w5365 = ~w4798 & ~w5878;
assign w5366 = ~w5855 & w5968;
assign w5367 = w968 & ~pi0329;
assign w5368 = w10811 & w2565;
assign w5369 = (~pi1777 & ~w7799) | (~pi1777 & w1168) | (~w7799 & w1168);
assign w5370 = ~pi1008 & w3791;
assign w5371 = pi1557 & ~w18259;
assign w5372 = ~w5363 & ~w2914;
assign w5373 = pi2959 & ~w458;
assign w5374 = pi1801 & ~w14951;
assign w5375 = ~pi3142 & w17669;
assign w5376 = pi3077 & ~w3987;
assign w5377 = (pi1078 & ~w13509) | (pi1078 & w8196) | (~w13509 & w8196);
assign w5378 = w13509 & w6070;
assign w5379 = ~w8712 & ~w16073;
assign w5380 = ~w7444 & ~w13479;
assign w5381 = w13509 & w9370;
assign w5382 = w3111 & ~pi3369;
assign w5383 = pi2981 & pi2982;
assign w5384 = w3556 & w5767;
assign w5385 = pi1955 & ~w14833;
assign w5386 = w735 & w3411;
assign w5387 = (pi0876 & ~w13509) | (pi0876 & w16151) | (~w13509 & w16151);
assign w5388 = (pi1049 & ~w13509) | (pi1049 & w13795) | (~w13509 & w13795);
assign w5389 = w5189 & ~w15173;
assign w5390 = ~pi2599 & w1333;
assign w5391 = ~pi2844 & w13343;
assign w5392 = pi2242 & ~w15883;
assign w5393 = w10647 & ~w6163;
assign w5394 = pi2057 & ~w10158;
assign w5395 = ~pi3326 & w7090;
assign w5396 = w13318 & w13176;
assign w5397 = w11209 & ~w10322;
assign w5398 = w10647 & ~w15198;
assign w5399 = pi1355 & w11685;
assign w5400 = ~w3899 & ~w14924;
assign w5401 = ~pi2078 & w17439;
assign w5402 = w11209 & ~w18264;
assign w5403 = ~w12890 & w3723;
assign w5404 = pi1305 & pi1266;
assign w5405 = pi2961 & w8789;
assign w5406 = w11383 & w17994;
assign w5407 = w934 & pi0432;
assign w5408 = ~w8273 & ~w6208;
assign w5409 = w7307 & w6517;
assign w5410 = ~w16650 & w1929;
assign w5411 = w2206 & ~w10296;
assign w5412 = ~w123 & ~w11094;
assign w5413 = pi2759 & ~w6463;
assign w5414 = ~w14648 & ~pi2697;
assign w5415 = pi2536 & w15191;
assign w5416 = w17562 & pi2518;
assign w5417 = w13509 & w7450;
assign w5418 = ~w12201 & ~w5279;
assign w5419 = ~pi0495 & pi1142;
assign w5420 = ~w15446 & ~w102;
assign w5421 = ~pi0083 & pi0084;
assign w5422 = w384 & w11392;
assign w5423 = ~w17442 & ~w2940;
assign w5424 = ~pi0120 & pi1220;
assign w5425 = w12460 & w7315;
assign w5426 = ~w18345 & ~w6499;
assign w5427 = ~w14423 & ~w1499;
assign w5428 = pi1779 & ~w18343;
assign w5429 = ~w541 & w3180;
assign w5430 = (pi0561 & ~w13509) | (pi0561 & w5333) | (~w13509 & w5333);
assign w5431 = ~w6498 & ~w15821;
assign w5432 = ~pi3079 & ~pi3207;
assign w5433 = ~w10899 & ~w12313;
assign w5434 = ~w3809 & ~w17515;
assign w5435 = ~w11646 & ~w8863;
assign w5436 = ~w9122 & ~w1476;
assign w5437 = ~w7033 & w18454;
assign w5438 = ~w15573 & ~w8986;
assign w5439 = ~w4369 & ~w17163;
assign w5440 = ~pi0823 & w1147;
assign w5441 = w13509 & w6027;
assign w5442 = ~pi3293 & w14918;
assign w5443 = ~w13367 & ~w1030;
assign w5444 = w10818 & ~w9197;
assign w5445 = pi1399 & ~w13786;
assign w5446 = ~pi0308 & ~w291;
assign w5447 = ~pi0898 & w93;
assign w5448 = ~pi2255 & w13065;
assign w5449 = ~w6459 & ~w4561;
assign w5450 = pi1593 & ~w13753;
assign w5451 = ~w12239 & ~w9379;
assign w5452 = w3960 & w8595;
assign w5453 = ~pi2920 & pi2966;
assign w5454 = ~pi0668 & w12197;
assign w5455 = ~w16278 & pi1105;
assign w5456 = ~pi3020 & pi3207;
assign w5457 = w9227 & w8658;
assign w5458 = pi2238 & ~w11735;
assign w5459 = ~w14185 & w13993;
assign w5460 = ~w514 & ~w8914;
assign w5461 = ~w11960 & ~w14260;
assign w5462 = w5453 & pi2591;
assign w5463 = pi1436 & ~w6448;
assign w5464 = ~w5375 & ~w1335;
assign w5465 = ~w3054 & w9817;
assign w5466 = w14296 & w15837;
assign w5467 = w13509 & w10615;
assign w5468 = w62 & ~w4770;
assign w5469 = ~w5050 & ~w9339;
assign w5470 = ~w16506 & pi1145;
assign w5471 = w1962 & ~w13195;
assign w5472 = pi3155 & w15767;
assign w5473 = pi2787 & ~w5274;
assign w5474 = w13509 & w18228;
assign w5475 = ~pi3150 & w15048;
assign w5476 = ~w213 & ~w17647;
assign w5477 = ~pi1858 & w12329;
assign w5478 = ~w14696 & ~w8075;
assign w5479 = ~w15808 & pi0746;
assign w5480 = pi1631 & ~w6448;
assign w5481 = ~w16278 & pi0701;
assign w5482 = w9440 & pi0180;
assign w5483 = ~w398 & w13217;
assign w5484 = pi2301 & ~w18123;
assign w5485 = w7703 & w6019;
assign w5486 = ~w8718 & ~w3765;
assign w5487 = ~pi3347 & w17935;
assign w5488 = w17562 & pi2575;
assign w5489 = ~pi1019 & w9110;
assign w5490 = pi1625 & ~w13753;
assign w5491 = ~w14356 & ~w6510;
assign w5492 = (~w13367 & w17577) | (~w13367 & w8451) | (w17577 & w8451);
assign w5493 = ~w4014 & ~w13937;
assign w5494 = ~w16404 & w15238;
assign w5495 = ~w594 & ~w7511;
assign w5496 = ~pi2943 & ~w13070;
assign w5497 = w15122 & ~pi1689;
assign w5498 = w7077 & ~w13195;
assign w5499 = ~pi3343 & w6448;
assign w5500 = pi1663 & ~w4058;
assign w5501 = w13509 & w10303;
assign w5502 = ~w8920 & w6896;
assign w5503 = pi1620 & w13753;
assign w5504 = w5190 & pi3115;
assign w5505 = ~w2293 & ~w18118;
assign w5506 = ~w14276 & ~w18413;
assign w5507 = pi0012 & ~w14148;
assign w5508 = ~w2316 & w7593;
assign w5509 = ~w7844 & pi1200;
assign w5510 = ~pi0503 & ~pi1155;
assign w5511 = ~w10448 & w2998;
assign w5512 = pi1495 & ~w13753;
assign w5513 = ~w10202 & ~w1247;
assign w5514 = w4348 & ~w322;
assign w5515 = ~w13039 & ~w16894;
assign w5516 = pi1455 & ~w7090;
assign w5517 = w12239 & w3228;
assign w5518 = ~w6418 & ~w16014;
assign w5519 = w13509 & w11705;
assign w5520 = ~pi3088 & w16815;
assign w5521 = (w3770 & ~w11247) | (w3770 & w17658) | (~w11247 & w17658);
assign w5522 = (~w13367 & w17577) | (~w13367 & w4933) | (w17577 & w4933);
assign w5523 = ~w2093 & ~w15507;
assign w5524 = ~pi2247 & w16041;
assign w5525 = ~w16278 & pi0927;
assign w5526 = pi1594 & ~w16922;
assign w5527 = ~w16790 & w15277;
assign w5528 = (w15056 & ~w32) | (w15056 & w16477) | (~w32 & w16477);
assign w5529 = ~w6405 & ~w3536;
assign w5530 = w13509 & w2932;
assign w5531 = ~w12329 & ~w6838;
assign w5532 = ~pi3162 & w1843;
assign w5533 = w2204 & w15996;
assign w5534 = ~w8844 & ~w2755;
assign w5535 = w384 & w1502;
assign w5536 = ~w11476 & w12665;
assign w5537 = ~w18175 & ~w8222;
assign w5538 = w7307 & w7659;
assign w5539 = ~w12460 & w8288;
assign w5540 = pi0009 & ~w3748;
assign w5541 = w6785 & ~w17210;
assign w5542 = (pi1122 & ~w13509) | (pi1122 & w6181) | (~w13509 & w6181);
assign w5543 = ~w13231 & pi1197;
assign w5544 = ~pi2537 & w15842;
assign w5545 = w17562 & pi1825;
assign w5546 = ~pi0605 & w12825;
assign w5547 = w485 & ~pi1299;
assign w5548 = ~pi3155 & w1843;
assign w5549 = pi3147 & w3987;
assign w5550 = ~w16467 & ~w13133;
assign w5551 = (pi1303 & ~w17477) | (pi1303 & w9362) | (~w17477 & w9362);
assign w5552 = ~pi3096 & w6463;
assign w5553 = ~w2381 & ~w6629;
assign w5554 = ~w14343 & ~w391;
assign w5555 = pi2098 & ~w4420;
assign w5556 = w14228 & ~w10947;
assign w5557 = (~w8011 & ~w9420) | (~w8011 & w13628) | (~w9420 & w13628);
assign w5558 = pi1485 & w13753;
assign w5559 = pi1222 & pi3204;
assign w5560 = ~w14420 & w13690;
assign w5561 = pi1896 & ~w15036;
assign w5562 = ~w11147 & w9006;
assign w5563 = ~w1791 & w16997;
assign w5564 = ~pi3172 & w3982;
assign w5565 = w12185 & w11598;
assign w5566 = (pi2913 & w5560) | (pi2913 & w1629) | (w5560 & w1629);
assign w5567 = ~w14865 & ~w15280;
assign w5568 = pi1985 & ~w4254;
assign w5569 = ~pi2967 & ~pi3114;
assign w5570 = w13509 & w6076;
assign w5571 = pi3136 & pi3207;
assign w5572 = ~pi3135 & pi3207;
assign w5573 = pi1891 & ~w15036;
assign w5574 = ~w10224 & ~w8746;
assign w5575 = ~w12945 & ~w14272;
assign w5576 = ~pi3138 & w3982;
assign w5577 = pi0301 & pi0260;
assign w5578 = ~w3203 & pi0578;
assign w5579 = ~w17806 & ~w17680;
assign w5580 = ~w3448 & w7817;
assign w5581 = ~pi2241 & w12724;
assign w5582 = pi2981 & ~w3987;
assign w5583 = pi0058 & ~w14148;
assign w5584 = ~w10304 & ~w16758;
assign w5585 = ~pi2509 & w17213;
assign w5586 = w16278 & ~w17210;
assign w5587 = w11266 & w13161;
assign w5588 = ~w11274 & ~w8980;
assign w5589 = (w5855 & w18597) | (w5855 & w16174) | (w18597 & w16174);
assign w5590 = ~pi0892 & w1126;
assign w5591 = ~w17503 & w18128;
assign w5592 = w934 & pi0412;
assign w5593 = w8432 & w14016;
assign w5594 = pi0146 & w5274;
assign w5595 = pi1767 & pi3154;
assign w5596 = w4809 & w7130;
assign w5597 = ~pi3097 & w16815;
assign w5598 = ~pi3434 & w15036;
assign w5599 = ~w7902 & ~w13414;
assign w5600 = pi0248 & w5274;
assign w5601 = w6785 & ~w14978;
assign w5602 = ~w2725 & pi1083;
assign w5603 = ~pi3170 & w8515;
assign w5604 = ~w5688 & ~w6965;
assign w5605 = ~w18106 & ~w13044;
assign w5606 = ~pi0075 & w922;
assign w5607 = pi1218 & ~pi2519;
assign w5608 = pi2412 & ~w10158;
assign w5609 = ~pi2310 & w3019;
assign w5610 = w2341 & ~w7020;
assign w5611 = ~w3728 & ~w17883;
assign w5612 = pi1153 & w13509;
assign w5613 = ~w16094 & ~w16780;
assign w5614 = ~w10771 & w4375;
assign w5615 = w6697 & ~w13028;
assign w5616 = pi2406 & ~w3223;
assign w5617 = (pi1034 & ~w13509) | (pi1034 & w2643) | (~w13509 & w2643);
assign w5618 = ~pi3163 & w3982;
assign w5619 = ~w1601 & ~w9977;
assign w5620 = ~w6450 & w1332;
assign w5621 = ~w1368 & ~pi0474;
assign w5622 = ~pi3145 & w11701;
assign w5623 = ~w15697 & ~w7869;
assign w5624 = w1127 & ~w5126;
assign w5625 = ~w10330 & ~w11201;
assign w5626 = ~w1962 & pi1116;
assign w5627 = pi1424 & ~w6072;
assign w5628 = (pi1020 & ~w13509) | (pi1020 & w17236) | (~w13509 & w17236);
assign w5629 = pi0114 & w3748;
assign w5630 = ~w3145 & ~w1299;
assign w5631 = pi1513 & ~w14918;
assign w5632 = ~w12686 & ~w3871;
assign w5633 = ~pi0726 & w17899;
assign w5634 = pi1814 & ~w2732;
assign w5635 = ~pi1066 & w93;
assign w5636 = pi2817 & ~w15235;
assign w5637 = ~w13056 & ~w17068;
assign w5638 = w8337 & pi3276;
assign w5639 = ~w9570 & ~w14443;
assign w5640 = pi1426 & ~w6072;
assign w5641 = ~w12460 & w6317;
assign w5642 = w17103 & w3266;
assign w5643 = pi1672 & ~w4058;
assign w5644 = pi3210 & pi3351;
assign w5645 = pi1583 & w13753;
assign w5646 = pi1948 & ~w14833;
assign w5647 = ~w6349 & ~w18570;
assign w5648 = ~pi2066 & w8617;
assign w5649 = w6649 & ~w5846;
assign w5650 = ~pi1129 & ~pi1177;
assign w5651 = pi1574 & ~w13753;
assign w5652 = w6111 & w2380;
assign w5653 = ~pi1034 & w17490;
assign w5654 = ~pi3298 & w7090;
assign w5655 = pi2546 & w14148;
assign w5656 = ~w3672 & ~w7453;
assign w5657 = pi1162 & ~w14073;
assign w5658 = ~pi2246 & w3019;
assign w5659 = pi2916 & ~pi3205;
assign w5660 = w6697 & ~w13195;
assign w5661 = ~w8799 & w6202;
assign w5662 = (pi1146 & ~w5437) | (pi1146 & w9030) | (~w5437 & w9030);
assign w5663 = w10158 & w614;
assign w5664 = ~w6056 & w5421;
assign w5665 = (pi1204 & w4470) | (pi1204 & w4857) | (w4470 & w4857);
assign w5666 = pi1629 & ~w13753;
assign w5667 = (~pi0978 & ~w13509) | (~pi0978 & w7584) | (~w13509 & w7584);
assign w5668 = pi1773 & ~w10389;
assign w5669 = ~pi2335 & w8617;
assign w5670 = w13509 & w5105;
assign w5671 = ~w6195 & w11773;
assign w5672 = (pi1091 & ~w13509) | (pi1091 & w7704) | (~w13509 & w7704);
assign w5673 = w13840 & w15842;
assign w5674 = ~pi2210 & w5075;
assign w5675 = pi2923 & w2276;
assign w5676 = ~w6373 & ~w9799;
assign w5677 = w12460 & w7573;
assign w5678 = w11345 & w1112;
assign w5679 = ~w9944 & ~w12380;
assign w5680 = (pi1786 & w7215) | (pi1786 & w16134) | (w7215 & w16134);
assign w5681 = w14109 & pi0433;
assign w5682 = w17646 & w3515;
assign w5683 = pi1862 & ~w458;
assign w5684 = ~pi2033 & w7455;
assign w5685 = w11122 & w4289;
assign w5686 = pi3030 & ~pi3138;
assign w5687 = w16575 & w2168;
assign w5688 = ~pi0918 & w17490;
assign w5689 = ~pi3098 & w261;
assign w5690 = ~w2706 & ~w3873;
assign w5691 = pi0305 & w18583;
assign w5692 = ~w17827 & w14265;
assign w5693 = w6649 & ~w9796;
assign w5694 = w4957 & w13796;
assign w5695 = ~w10269 & w11292;
assign w5696 = pi3037 & ~w16502;
assign w5697 = ~w6682 & w17350;
assign w5698 = ~pi0872 & w15707;
assign w5699 = ~w16506 & pi1187;
assign w5700 = w13509 & w11569;
assign w5701 = ~w7276 & ~w6408;
assign w5702 = pi1298 & ~w14158;
assign w5703 = ~w11783 & ~w5447;
assign w5704 = pi1295 & pi1345;
assign w5705 = ~w17248 & pi0874;
assign w5706 = w13509 & w4201;
assign w5707 = pi2106 & ~w4420;
assign w5708 = w9440 & pi0168;
assign w5709 = ~w6324 & ~w7415;
assign w5710 = ~pi3139 & pi3207;
assign w5711 = ~w6472 & ~w4193;
assign w5712 = ~w3373 & ~w5448;
assign w5713 = ~w5646 & ~w1460;
assign w5714 = ~pi3062 & w6463;
assign w5715 = w15122 & ~pi2629;
assign w5716 = pi0195 & w5274;
assign w5717 = pi2561 & ~w5274;
assign w5718 = ~w18548 & ~w8924;
assign w5719 = pi1711 & ~pi3132;
assign w5720 = w13509 & w4992;
assign w5721 = pi1980 & ~w11406;
assign w5722 = (pi0743 & ~w13509) | (pi0743 & w14744) | (~w13509 & w14744);
assign w5723 = ~w16278 & pi1025;
assign w5724 = ~pi1750 & ~w3633;
assign w5725 = w11383 & w5950;
assign w5726 = w7703 & w7889;
assign w5727 = ~w5189 & pi0922;
assign w5728 = w10647 & ~w6591;
assign w5729 = ~w3203 & pi0588;
assign w5730 = ~w7077 & pi0820;
assign w5731 = ~pi3295 & w16922;
assign w5732 = ~pi3123 & ~w6801;
assign w5733 = ~w674 & ~w11841;
assign w5734 = pi0483 & pi0501;
assign w5735 = pi3160 & ~pi3503;
assign w5736 = ~w18082 & w11096;
assign w5737 = w8211 & w16318;
assign w5738 = ~w2216 & ~w16355;
assign w5739 = ~w8588 & w11671;
assign w5740 = pi0203 & w5274;
assign w5741 = (pi0990 & ~w13509) | (pi0990 & w9431) | (~w13509 & w9431);
assign w5742 = ~pi1337 & ~w3655;
assign w5743 = w17279 & w17266;
assign w5744 = w13509 & w16932;
assign w5745 = ~w7814 & w1895;
assign w5746 = w10887 & w3182;
assign w5747 = ~w10701 & ~w3901;
assign w5748 = ~w7224 & ~w8;
assign w5749 = w13509 & w11959;
assign w5750 = ~w14134 & w6776;
assign w5751 = ~pi1127 & w14641;
assign w5752 = ~w14648 & ~pi2284;
assign w5753 = ~pi2851 & w735;
assign w5754 = ~w625 & ~pi0496;
assign w5755 = ~w7844 & pi1065;
assign w5756 = ~pi1778 & w10335;
assign w5757 = (pi0369 & w6195) | (pi0369 & w12956) | (w6195 & w12956);
assign w5758 = ~pi2036 & w7455;
assign w5759 = ~w2115 & ~w11382;
assign w5760 = ~w5031 & pi1376;
assign w5761 = ~pi3091 & w11406;
assign w5762 = w8211 & w876;
assign w5763 = w5944 & pi0078;
assign w5764 = w11383 & w11845;
assign w5765 = w6785 & ~w14143;
assign w5766 = w11209 & ~w1853;
assign w5767 = w7681 & w8067;
assign w5768 = ~pi1409 & ~pi2913;
assign w5769 = pi1410 & ~pi2913;
assign w5770 = pi2984 & ~w3987;
assign w5771 = pi2465 & ~w603;
assign w5772 = ~w2462 & ~w3713;
assign w5773 = w1391 & ~w4043;
assign w5774 = ~pi1261 & ~w3987;
assign w5775 = pi1929 & ~w10299;
assign w5776 = ~pi2789 & w13343;
assign w5777 = w9440 & pi0136;
assign w5778 = ~pi0500 & pi0508;
assign w5779 = w13509 & w1270;
assign w5780 = ~w15319 & ~w16926;
assign w5781 = w13509 & w10668;
assign w5782 = w11383 & w3559;
assign w5783 = w11383 & w3560;
assign w5784 = w15946 & w17820;
assign w5785 = ~pi1110 & w12197;
assign w5786 = ~w10160 & ~w3688;
assign w5787 = ~w14132 & ~w831;
assign w5788 = pi1638 & ~w6448;
assign w5789 = ~w16876 & ~w4572;
assign w5790 = (~pi1221 & w5560) | (~pi1221 & w15058) | (w5560 & w15058);
assign w5791 = w1962 & ~w3374;
assign w5792 = ~w1547 & ~w8659;
assign w5793 = ~w2725 & pi0780;
assign w5794 = ~w9381 & ~w11914;
assign w5795 = ~w9996 & ~w6685;
assign w5796 = pi3160 & ~pi3499;
assign w5797 = ~pi3171 & w3982;
assign w5798 = ~w12938 & ~w6017;
assign w5799 = ~pi2358 & ~w7858;
assign w5800 = ~pi3060 & w261;
assign w5801 = ~w15605 & ~w9460;
assign w5802 = ~w1487 & ~w1683;
assign w5803 = w4035 & w12738;
assign w5804 = ~w2657 & ~w18350;
assign w5805 = ~pi3134 & ~pi3160;
assign w5806 = ~pi2463 & ~pi2526;
assign w5807 = w14814 & w6913;
assign w5808 = (pi0925 & ~w13509) | (pi0925 & w1304) | (~w13509 & w1304);
assign w5809 = ~w16413 & ~w3327;
assign w5810 = w16965 & ~pi3016;
assign w5811 = ~w2392 & ~w14555;
assign w5812 = pi0059 & w17103;
assign w5813 = (pi0834 & ~w13509) | (pi0834 & w30) | (~w13509 & w30);
assign w5814 = w10647 & ~w81;
assign w5815 = ~w12040 & pi0543;
assign w5816 = ~w6697 & pi0665;
assign w5817 = ~w16665 & ~w13021;
assign w5818 = w5968 & pi0444;
assign w5819 = w1962 & ~w16498;
assign w5820 = pi2576 & ~w5274;
assign w5821 = w13231 & ~w10947;
assign w5822 = pi1336 & w13250;
assign w5823 = pi2417 & ~w3223;
assign w5824 = pi2810 & ~w226;
assign w5825 = w6785 & ~w15173;
assign w5826 = w14228 & ~w17210;
assign w5827 = ~w18047 & ~w4084;
assign w5828 = w3298 & w13586;
assign w5829 = ~pi1908 & w5075;
assign w5830 = w11209 & ~w6480;
assign w5831 = ~w16939 & pi0004;
assign w5832 = w17562 & pi2733;
assign w5833 = ~w7052 & ~w11965;
assign w5834 = ~pi3003 & ~pi3207;
assign w5835 = ~w14885 & ~w10876;
assign w5836 = ~w15934 & w13139;
assign w5837 = ~w5823 & ~w3051;
assign w5838 = pi3158 & w14980;
assign w5839 = ~w2444 & ~pi0485;
assign w5840 = w13509 & w2389;
assign w5841 = pi0076 & ~pi3366;
assign w5842 = pi2924 & w11760;
assign w5843 = ~pi0174 & ~pi0175;
assign w5844 = ~w12669 & ~w4115;
assign w5845 = ~pi2967 & pi3078;
assign w5846 = pi1459 & w13753;
assign w5847 = pi1428 & ~w13753;
assign w5848 = pi2844 & ~w11406;
assign w5849 = w7844 & ~w6680;
assign w5850 = ~w16278 & pi0932;
assign w5851 = ~w14201 & ~w12364;
assign w5852 = ~w13137 & ~w18398;
assign w5853 = ~pi3163 & w15839;
assign w5854 = w7307 & w9036;
assign w5855 = ~w11743 & ~w11760;
assign w5856 = ~w17694 & ~w15993;
assign w5857 = w11383 & w949;
assign w5858 = pi0311 & ~pi0312;
assign w5859 = w13509 & w1464;
assign w5860 = ~w3243 & pi0313;
assign w5861 = pi3158 & w3358;
assign w5862 = ~w5560 & w10456;
assign w5863 = w539 & ~w9254;
assign w5864 = w16970 & w10960;
assign w5865 = ~w13260 & ~w568;
assign w5866 = ~pi2138 & w12941;
assign w5867 = w18514 & w142;
assign w5868 = ~w6306 & ~w13166;
assign w5869 = ~w17039 & ~w10993;
assign w5870 = ~pi0852 & w15707;
assign w5871 = ~w8369 & ~w6342;
assign w5872 = ~w7047 & ~w9671;
assign w5873 = pi1745 & ~w4058;
assign w5874 = w17378 & w1250;
assign w5875 = w13509 & w16300;
assign w5876 = ~w12914 & ~w15498;
assign w5877 = pi0065 & ~w14148;
assign w5878 = ~w5560 & w599;
assign w5879 = ~w15122 & ~pi2677;
assign w5880 = ~pi2013 & w11688;
assign w5881 = ~w17248 & pi0883;
assign w5882 = w11209 & ~w13426;
assign w5883 = ~w15944 & ~w14257;
assign w5884 = ~w15541 & ~w12351;
assign w5885 = ~w5034 & ~w1296;
assign w5886 = ~w16362 & ~w16105;
assign w5887 = ~w14843 & w7716;
assign w5888 = (pi0587 & ~w13509) | (pi0587 & w3486) | (~w13509 & w3486);
assign w5889 = pi2248 & ~w15883;
assign w5890 = ~w2341 & pi0841;
assign w5891 = pi1847 & ~w12558;
assign w5892 = pi1998 & ~w9414;
assign w5893 = ~w6939 & ~w18442;
assign w5894 = pi0116 & w3748;
assign w5895 = ~pi0775 & w6200;
assign w5896 = pi1694 & ~w15379;
assign w5897 = (~pi0951 & ~w13509) | (~pi0951 & w7085) | (~w13509 & w7085);
assign w5898 = pi2079 & ~w17683;
assign w5899 = pi3160 & ~pi3505;
assign w5900 = ~w18115 & w544;
assign w5901 = w6111 & ~w4156;
assign w5902 = ~pi3055 & w9504;
assign w5903 = (pi0715 & ~w13509) | (pi0715 & w16322) | (~w13509 & w16322);
assign w5904 = (pi0591 & ~w13509) | (pi0591 & w14784) | (~w13509 & w14784);
assign w5905 = w13509 & w2091;
assign w5906 = ~w6380 & ~w6278;
assign w5907 = ~pi3330 & w6448;
assign w5908 = ~pi0483 & pi3383;
assign w5909 = ~w3557 & ~w353;
assign w5910 = ~w11339 & ~w6936;
assign w5911 = w384 & w1841;
assign w5912 = w16575 & w9912;
assign w5913 = w4103 & w13711;
assign w5914 = ~pi1724 & w18503;
assign w5915 = ~w4872 & ~w16673;
assign w5916 = ~w3405 & ~w1252;
assign w5917 = ~w17204 & ~w5370;
assign w5918 = ~w9867 & ~w12121;
assign w5919 = ~w8293 & ~w3263;
assign w5920 = w14648 & ~pi1880;
assign w5921 = ~w17665 & ~w9409;
assign w5922 = ~w5560 & w15415;
assign w5923 = ~w11367 & w16868;
assign w5924 = ~w14067 & w6983;
assign w5925 = ~w7556 & ~w2328;
assign w5926 = ~pi3142 & w17387;
assign w5927 = ~pi3155 & w14753;
assign w5928 = pi1486 & ~w9781;
assign w5929 = ~w13692 & ~w7156;
assign w5930 = ~pi2812 & w17213;
assign w5931 = ~pi3287 & w7090;
assign w5932 = ~w1038 & ~w656;
assign w5933 = w17683 & w3515;
assign w5934 = pi1858 & w4021;
assign w5935 = pi3160 & ~pi3476;
assign w5936 = pi1754 & ~w619;
assign w5937 = pi2952 & ~w13367;
assign w5938 = ~w5516 & ~w2743;
assign w5939 = w11383 & w1955;
assign w5940 = w13509 & w15987;
assign w5941 = pi2452 & ~w10299;
assign w5942 = w13509 & w3458;
assign w5943 = pi3065 & ~w3987;
assign w5944 = (pi1318 & ~w8087) | (pi1318 & w18527) | (~w8087 & w18527);
assign w5945 = pi1576 & ~w14918;
assign w5946 = ~w661 & ~w7128;
assign w5947 = pi1251 & ~w11655;
assign w5948 = ~w7677 & ~w7373;
assign w5949 = pi0044 & pi0057;
assign w5950 = ~w14648 & ~pi2623;
assign w5951 = ~pi0675 & w12197;
assign w5952 = pi2023 & ~w17646;
assign w5953 = ~pi3024 & ~pi3207;
assign w5954 = ~pi2778 & w15122;
assign w5955 = pi0059 & ~w14148;
assign w5956 = w15122 & ~pi2517;
assign w5957 = w6649 & ~w2433;
assign w5958 = pi3023 & w16502;
assign w5959 = ~w11678 & w10665;
assign w5960 = w14228 & ~w6033;
assign w5961 = pi1518 & ~w14918;
assign w5962 = pi1460 & ~w7090;
assign w5963 = ~w6354 & ~w3282;
assign w5964 = ~pi2080 & w17439;
assign w5965 = w6697 & ~w17210;
assign w5966 = pi1561 & ~w18259;
assign w5967 = pi0093 & w9284;
assign w5968 = ~pi3042 & ~pi3118;
assign w5969 = ~w6690 & ~w2721;
assign w5970 = ~w7308 & ~w8666;
assign w5971 = ~pi3146 & w12427;
assign w5972 = w2037 & w12913;
assign w5973 = w968 & ~pi0286;
assign w5974 = w12460 & w12782;
assign w5975 = (w8645 & ~w1516) | (w8645 & w11007) | (~w1516 & w11007);
assign w5976 = ~w11519 & ~w1439;
assign w5977 = w14109 & pi0437;
assign w5978 = pi1634 & ~w13753;
assign w5979 = w2528 & w8145;
assign w5980 = ~w17569 & ~w6449;
assign w5981 = pi3018 & ~w858;
assign w5982 = (pi0622 & ~w13509) | (pi0622 & w1098) | (~w13509 & w1098);
assign w5983 = w18274 & w13035;
assign w5984 = ~w17128 & w3876;
assign w5985 = ~w15003 & w12430;
assign w5986 = ~w33 & ~w17056;
assign w5987 = ~w17645 & ~w14532;
assign w5988 = ~pi3090 & w3555;
assign w5989 = ~w11018 & ~w569;
assign w5990 = ~w11059 & ~w10608;
assign w5991 = ~w4856 & ~w8756;
assign w5992 = ~pi3293 & w7090;
assign w5993 = pi1622 & ~w13753;
assign w5994 = pi2802 & ~w6463;
assign w5995 = w10232 & w17955;
assign w5996 = w1127 & ~w17060;
assign w5997 = pi0143 & ~pi0198;
assign w5998 = pi2244 & ~w17683;
assign w5999 = ~w1108 & ~w825;
assign w6000 = ~w345 & ~w6183;
assign w6001 = pi1337 & ~w13236;
assign w6002 = ~pi1813 & pi3034;
assign w6003 = ~w6785 & pi0859;
assign w6004 = w4647 & w9123;
assign w6005 = pi3010 & w16502;
assign w6006 = ~w18177 & ~w1461;
assign w6007 = ~w959 & ~w9198;
assign w6008 = ~w12884 & ~w2121;
assign w6009 = ~w8703 & ~w12076;
assign w6010 = w606 & w10288;
assign w6011 = ~w7973 & ~w17761;
assign w6012 = pi1549 & w13753;
assign w6013 = pi1556 & ~w13753;
assign w6014 = pi1540 & w13753;
assign w6015 = w5437 & w12253;
assign w6016 = w17581 & ~w7882;
assign w6017 = ~pi3336 & w17935;
assign w6018 = ~w1906 & ~w1002;
assign w6019 = ~w15122 & ~pi2883;
assign w6020 = (pi0752 & ~w13509) | (pi0752 & w16248) | (~w13509 & w16248);
assign w6021 = ~pi0490 & ~pi1345;
assign w6022 = pi1505 & ~w13753;
assign w6023 = ~w6697 & pi0942;
assign w6024 = ~pi1367 & w11747;
assign w6025 = ~w10932 & ~w2659;
assign w6026 = w13509 & w17459;
assign w6027 = w1962 & ~w1236;
assign w6028 = pi2469 & ~w14524;
assign w6029 = w11209 & ~w281;
assign w6030 = ~pi0670 & w12197;
assign w6031 = ~w2563 & ~w3564;
assign w6032 = ~w13231 & pi0562;
assign w6033 = ~w1518 & ~w4636;
assign w6034 = ~pi2290 & w3019;
assign w6035 = w18412 & w6295;
assign w6036 = ~w9413 & w221;
assign w6037 = ~w375 & ~w12115;
assign w6038 = pi1181 & w14073;
assign w6039 = w8337 & pi3281;
assign w6040 = pi3151 & w8113;
assign w6041 = ~w919 & ~w1008;
assign w6042 = pi1609 & w13753;
assign w6043 = ~w7077 & pi1071;
assign w6044 = ~w15320 & ~w8735;
assign w6045 = pi1306 & ~w9704;
assign w6046 = ~pi1049 & w15707;
assign w6047 = ~pi0581 & w795;
assign w6048 = w7077 & ~w15296;
assign w6049 = pi2526 & ~w13394;
assign w6050 = pi0174 & w5274;
assign w6051 = ~pi2002 & w3019;
assign w6052 = pi1644 & ~w13753;
assign w6053 = ~w11087 & ~w5740;
assign w6054 = pi1210 & pi3362;
assign w6055 = ~pi1980 & w13343;
assign w6056 = ~w18010 & ~w14012;
assign w6057 = pi0129 & ~pi0223;
assign w6058 = w13509 & w12324;
assign w6059 = pi3146 & pi3207;
assign w6060 = w12460 & w10037;
assign w6061 = w384 & w17417;
assign w6062 = (pi0937 & ~w13509) | (pi0937 & w1415) | (~w13509 & w1415);
assign w6063 = ~w9745 & ~w13419;
assign w6064 = ~w4492 & w1326;
assign w6065 = ~w1962 & pi0655;
assign w6066 = pi2740 & ~w6463;
assign w6067 = w13509 & w18474;
assign w6068 = ~w309 & ~w10123;
assign w6069 = w1697 & w4034;
assign w6070 = w6697 & ~w17513;
assign w6071 = (pi0305 & w15203) | (pi0305 & w18276) | (w15203 & w18276);
assign w6072 = ~pi1371 & w6024;
assign w6073 = w10189 & pi0407;
assign w6074 = ~w17529 & ~w12526;
assign w6075 = ~pi0766 & w6200;
assign w6076 = w17248 & ~w10235;
assign w6077 = (w15450 & w14073) | (w15450 & w8973) | (w14073 & w8973);
assign w6078 = ~w14742 & w1326;
assign w6079 = pi1565 & ~w13753;
assign w6080 = ~w13984 & w17910;
assign w6081 = ~w14120 & ~w3272;
assign w6082 = ~pi3346 & w6072;
assign w6083 = w13509 & w14631;
assign w6084 = ~w11883 & ~w14621;
assign w6085 = w17562 & pi1850;
assign w6086 = ~w523 & ~w14575;
assign w6087 = ~pi3435 & w15036;
assign w6088 = ~pi2169 & w11313;
assign w6089 = w13509 & w1680;
assign w6090 = ~w5855 & w4364;
assign w6091 = pi1447 & ~w6448;
assign w6092 = (~pi0508 & w17577) | (~pi0508 & w14860) | (w17577 & w14860);
assign w6093 = w9627 & w1745;
assign w6094 = ~pi1589 & ~pi1712;
assign w6095 = w16620 & pi0504;
assign w6096 = ~w11530 & ~w14754;
assign w6097 = ~pi1371 & w5043;
assign w6098 = pi0012 & ~w3748;
assign w6099 = ~w4109 & ~w3176;
assign w6100 = ~w1962 & ~pi0959;
assign w6101 = ~w16770 & ~w2240;
assign w6102 = ~pi1070 & w1147;
assign w6103 = ~pi3056 & w9504;
assign w6104 = (~pi0312 & ~w13184) | (~pi0312 & w5858) | (~w13184 & w5858);
assign w6105 = ~w15150 & ~w6110;
assign w6106 = ~pi2829 & w15122;
assign w6107 = w13509 & w4825;
assign w6108 = ~w17248 & pi0892;
assign w6109 = w15292 & pi1240;
assign w6110 = w13509 & w14413;
assign w6111 = ~pi3366 & w15561;
assign w6112 = pi3132 & pi3146;
assign w6113 = ~w6785 & pi0854;
assign w6114 = ~w10344 & ~w15768;
assign w6115 = ~pi3045 & w15235;
assign w6116 = ~pi0643 & w3791;
assign w6117 = w1927 & w5141;
assign w6118 = pi2221 & ~w15271;
assign w6119 = ~pi3153 & w17387;
assign w6120 = ~pi1801 & ~pi3165;
assign w6121 = ~w11176 & ~w1931;
assign w6122 = ~w4802 & ~w5132;
assign w6123 = ~pi1123 & w17899;
assign w6124 = ~w13231 & pi1090;
assign w6125 = (pi0616 & ~w13509) | (pi0616 & w10987) | (~w13509 & w10987);
assign w6126 = ~w9846 & ~w3012;
assign w6127 = w17562 & pi1814;
assign w6128 = ~w1258 & ~w7885;
assign w6129 = ~w15688 & ~w7176;
assign w6130 = pi1524 & w13753;
assign w6131 = ~pi3353 & w18259;
assign w6132 = ~w1559 & ~w9235;
assign w6133 = ~w17665 & ~w531;
assign w6134 = ~w3162 & ~w2965;
assign w6135 = ~pi1345 & ~pi1762;
assign w6136 = ~pi3299 & w9781;
assign w6137 = w10189 & pi0396;
assign w6138 = (pi1069 & ~w13509) | (pi1069 & w10954) | (~w13509 & w10954);
assign w6139 = ~pi3158 & w11701;
assign w6140 = pi2799 & ~w6463;
assign w6141 = ~pi2098 & w12724;
assign w6142 = pi2972 & ~w3651;
assign w6143 = ~w1846 & w8823;
assign w6144 = ~pi0815 & w1147;
assign w6145 = ~w5227 & ~w5751;
assign w6146 = pi1762 & ~w7177;
assign w6147 = pi2986 & w3067;
assign w6148 = pi1470 & ~w7090;
assign w6149 = pi3160 & ~pi3496;
assign w6150 = w13509 & w17926;
assign w6151 = pi2032 & ~w17646;
assign w6152 = ~w4764 & ~w14017;
assign w6153 = pi1517 & w13753;
assign w6154 = ~pi3313 & w7090;
assign w6155 = ~pi2468 & w7455;
assign w6156 = ~w492 & ~w4944;
assign w6157 = w6785 & ~w305;
assign w6158 = ~pi0772 & w6200;
assign w6159 = ~w10847 & ~w8921;
assign w6160 = (w6203 & ~w8324) | (w6203 & w4279) | (~w8324 & w4279);
assign w6161 = ~w5453 & ~w11421;
assign w6162 = ~w8165 & ~w8016;
assign w6163 = pi1588 & w13753;
assign w6164 = ~w1391 & pi0776;
assign w6165 = ~w18189 & ~w5524;
assign w6166 = ~pi1947 & w7455;
assign w6167 = ~pi3061 & w9504;
assign w6168 = pi2279 & ~w15883;
assign w6169 = ~w1469 & ~w18254;
assign w6170 = ~w1391 & pi0760;
assign w6171 = ~pi2967 & ~pi3013;
assign w6172 = (pi1093 & ~w13509) | (pi1093 & w4100) | (~w13509 & w4100);
assign w6173 = pi2014 & ~w14833;
assign w6174 = ~w9740 & ~w56;
assign w6175 = pi1389 & ~w17935;
assign w6176 = ~w15122 & ~pi2893;
assign w6177 = w7307 & w16171;
assign w6178 = ~w9901 & ~w13478;
assign w6179 = ~w17377 & w13385;
assign w6180 = ~w4327 & w2460;
assign w6181 = ~w14228 & pi1122;
assign w6182 = w13231 & ~w7449;
assign w6183 = ~pi3293 & w16922;
assign w6184 = w6857 & w313;
assign w6185 = w14830 & w1101;
assign w6186 = ~pi3164 & w17669;
assign w6187 = ~w8393 & ~w4741;
assign w6188 = ~pi1696 & ~pi1697;
assign w6189 = ~pi3147 & w17387;
assign w6190 = ~w709 & pi1287;
assign w6191 = ~w10095 & ~w10355;
assign w6192 = ~w13163 & w2811;
assign w6193 = w12551 & ~w10593;
assign w6194 = ~w10720 & ~w15696;
assign w6195 = (~pi0359 & w860) | (~pi0359 & w4270) | (w860 & w4270);
assign w6196 = pi2138 & ~w15883;
assign w6197 = ~w11846 & ~w3456;
assign w6198 = w1127 & ~w6014;
assign w6199 = w5437 & w367;
assign w6200 = w134 & w9110;
assign w6201 = ~w10287 & ~w4665;
assign w6202 = w1127 & ~w14551;
assign w6203 = ~w14783 & w3886;
assign w6204 = w13509 & w17886;
assign w6205 = ~w1391 & pi0763;
assign w6206 = pi1703 & w4667;
assign w6207 = ~pi1702 & w4667;
assign w6208 = ~pi0813 & w1147;
assign w6209 = ~w6242 & ~w9839;
assign w6210 = pi0442 & w17173;
assign w6211 = ~pi0441 & w17173;
assign w6212 = ~w12403 & w12369;
assign w6213 = pi1489 & w13753;
assign w6214 = ~pi1681 & w7199;
assign w6215 = pi0023 & ~w3748;
assign w6216 = ~pi0987 & w15707;
assign w6217 = ~w16620 & ~pi0504;
assign w6218 = ~w10357 & ~w11961;
assign w6219 = w3243 & ~pi0315;
assign w6220 = w3243 & pi0316;
assign w6221 = ~pi1020 & w9110;
assign w6222 = ~pi3321 & w6448;
assign w6223 = ~w3581 & ~w803;
assign w6224 = w5593 & w7409;
assign w6225 = ~pi3025 & w5953;
assign w6226 = w16684 & w7376;
assign w6227 = ~w4821 & ~w18533;
assign w6228 = ~pi2984 & ~w7322;
assign w6229 = w1368 & pi0396;
assign w6230 = ~pi3163 & w17993;
assign w6231 = pi1276 & pi1345;
assign w6232 = pi3160 & ~pi3502;
assign w6233 = ~w3146 & ~w454;
assign w6234 = ~w3690 & ~w11080;
assign w6235 = (pi0394 & w5560) | (pi0394 & w3662) | (w5560 & w3662);
assign w6236 = ~w930 & ~w4735;
assign w6237 = ~pi3166 & w15839;
assign w6238 = ~w15671 & ~w898;
assign w6239 = ~w127 & ~w15762;
assign w6240 = pi3165 & w653;
assign w6241 = ~w13485 & ~w18389;
assign w6242 = (pi0638 & ~w13509) | (pi0638 & w14480) | (~w13509 & w14480);
assign w6243 = ~pi3103 & w11406;
assign w6244 = ~pi3154 & w4310;
assign w6245 = pi2969 & ~pi0484;
assign w6246 = pi3138 & w3987;
assign w6247 = ~w13883 & ~w15742;
assign w6248 = pi1246 & ~w11655;
assign w6249 = ~w15808 & pi1207;
assign w6250 = w3987 & w563;
assign w6251 = (pi0557 & ~w13509) | (pi0557 & w10927) | (~w13509 & w10927);
assign w6252 = ~w17665 & ~w18493;
assign w6253 = ~pi2224 & w2151;
assign w6254 = pi2178 & ~w14524;
assign w6255 = ~w15229 & ~w13182;
assign w6256 = ~pi3166 & w11132;
assign w6257 = ~w4980 & w8786;
assign w6258 = ~pi3163 & w14753;
assign w6259 = ~pi3026 & pi3166;
assign w6260 = pi1262 & ~pi2955;
assign w6261 = pi1267 & w11655;
assign w6262 = ~w991 & ~w16150;
assign w6263 = pi2979 & w6147;
assign w6264 = ~pi0804 & w1147;
assign w6265 = ~w12288 & w13595;
assign w6266 = ~w14228 & pi1061;
assign w6267 = w4420 & w6320;
assign w6268 = w12460 & w5708;
assign w6269 = w5129 & w3767;
assign w6270 = pi1904 & ~w15235;
assign w6271 = ~pi3106 & ~pi3207;
assign w6272 = ~w11506 & ~w11707;
assign w6273 = ~w2668 & ~w16354;
assign w6274 = ~w17717 & w14612;
assign w6275 = ~w7062 & ~w5585;
assign w6276 = ~w3000 & ~pi2740;
assign w6277 = ~w1612 & w903;
assign w6278 = ~pi3045 & w9504;
assign w6279 = w8462 & w17789;
assign w6280 = (pi0254 & ~w325) | (pi0254 & w937) | (~w325 & w937);
assign w6281 = w5189 & w15609;
assign w6282 = ~pi3247 & w9250;
assign w6283 = pi2766 & w14148;
assign w6284 = ~w1192 & ~w946;
assign w6285 = ~w11664 & ~w11179;
assign w6286 = ~pi0658 & w12197;
assign w6287 = ~w1630 & w1866;
assign w6288 = w5642 & w13029;
assign w6289 = ~w8502 & ~w10440;
assign w6290 = w13509 & w1600;
assign w6291 = pi2716 & ~w15235;
assign w6292 = w11383 & w1943;
assign w6293 = w8789 & pi0469;
assign w6294 = w8789 & ~pi0468;
assign w6295 = ~w4431 & ~w13770;
assign w6296 = ~w16468 & ~w5394;
assign w6297 = w7177 & w11685;
assign w6298 = pi2250 & ~w9414;
assign w6299 = ~pi3172 & w8515;
assign w6300 = pi2665 & ~w6463;
assign w6301 = ~pi2193 & w9340;
assign w6302 = w1391 & ~w6922;
assign w6303 = pi1500 & ~w13753;
assign w6304 = ~pi0513 & ~pi1144;
assign w6305 = w5338 & w10273;
assign w6306 = ~pi2967 & pi3067;
assign w6307 = ~w5099 & w2088;
assign w6308 = pi0152 & pi0203;
assign w6309 = pi1393 & w13753;
assign w6310 = pi1927 & ~w10299;
assign w6311 = ~pi3128 & w6463;
assign w6312 = pi0498 & ~pi1145;
assign w6313 = ~w10301 & ~w9906;
assign w6314 = pi1147 & w9420;
assign w6315 = pi2500 & ~w9504;
assign w6316 = pi2627 & ~w9504;
assign w6317 = w14109 & pi0441;
assign w6318 = w7077 & ~w14143;
assign w6319 = w10189 & pi0385;
assign w6320 = ~pi3134 & ~w4020;
assign w6321 = ~w17760 & ~w17596;
assign w6322 = pi2391 & ~w18123;
assign w6323 = pi2813 & ~w11406;
assign w6324 = ~pi3146 & w13730;
assign w6325 = pi1538 & ~w17935;
assign w6326 = ~pi3165 & w8515;
assign w6327 = ~pi3169 & w8515;
assign w6328 = w8789 & ~pi0381;
assign w6329 = ~w2756 & ~w6168;
assign w6330 = pi2768 & ~w226;
assign w6331 = ~w6054 & ~w9422;
assign w6332 = ~w10249 & ~w11480;
assign w6333 = ~w6954 & ~w12035;
assign w6334 = w14648 & ~pi2619;
assign w6335 = ~w2309 & ~w9118;
assign w6336 = w11383 & w12716;
assign w6337 = pi0197 & w9653;
assign w6338 = ~w16904 & ~w14313;
assign w6339 = ~w8790 & w2651;
assign w6340 = ~w15156 & w10606;
assign w6341 = ~pi2185 & w2151;
assign w6342 = w13509 & w1954;
assign w6343 = ~pi2934 & pi3208;
assign w6344 = ~w15712 & w1131;
assign w6345 = ~w740 & w13659;
assign w6346 = ~w10257 & ~w1043;
assign w6347 = (~pi1242 & w11655) | (~pi1242 & w8860) | (w11655 & w8860);
assign w6348 = ~pi2394 & w5075;
assign w6349 = ~pi1079 & w1147;
assign w6350 = ~pi1829 & ~w14833;
assign w6351 = (pi1021 & ~w13509) | (pi1021 & w6938) | (~w13509 & w6938);
assign w6352 = ~w17205 & ~w17983;
assign w6353 = ~w15248 & ~w7977;
assign w6354 = ~pi3063 & ~pi3207;
assign w6355 = pi3164 & w619;
assign w6356 = ~pi0949 & w1126;
assign w6357 = w11077 & ~w4554;
assign w6358 = ~w12937 & w8092;
assign w6359 = w11743 & w11921;
assign w6360 = w208 & w16648;
assign w6361 = ~w1791 & w14371;
assign w6362 = ~w11831 & ~w11988;
assign w6363 = ~w15546 & ~w9808;
assign w6364 = ~w15828 & w12318;
assign w6365 = w7498 & w7820;
assign w6366 = ~w15807 & ~w18489;
assign w6367 = pi1642 & ~w18259;
assign w6368 = w1962 & ~w17210;
assign w6369 = pi1496 & ~w16922;
assign w6370 = pi2481 & ~w15235;
assign w6371 = w17038 & w2836;
assign w6372 = w13509 & w16364;
assign w6373 = ~w16987 & w10557;
assign w6374 = w1127 & ~w318;
assign w6375 = pi1667 & ~w4058;
assign w6376 = pi1934 & ~w4420;
assign w6377 = w11383 & w5414;
assign w6378 = w6857 & w13866;
assign w6379 = ~w17825 & ~w9635;
assign w6380 = pi2695 & ~w9504;
assign w6381 = w13683 & ~w9485;
assign w6382 = (~w12368 & ~w9420) | (~w12368 & w6847) | (~w9420 & w6847);
assign w6383 = pi2366 & ~w4508;
assign w6384 = ~w17023 & ~w16373;
assign w6385 = ~w16257 & ~w9957;
assign w6386 = ~w1791 & w4336;
assign w6387 = pi2857 & ~w3555;
assign w6388 = (pi1123 & ~w13509) | (pi1123 & w7361) | (~w13509 & w7361);
assign w6389 = pi0074 & ~w14148;
assign w6390 = w7307 & w9956;
assign w6391 = ~w11215 & ~w7745;
assign w6392 = ~w17219 & ~w10175;
assign w6393 = pi0051 & pi0052;
assign w6394 = ~w13611 & ~w13572;
assign w6395 = w9414 & w14078;
assign w6396 = ~w2422 & w1966;
assign w6397 = w16062 & w395;
assign w6398 = ~pi0310 & pi3218;
assign w6399 = ~w17925 & w4236;
assign w6400 = w13509 & w1489;
assign w6401 = ~w16803 & ~w1932;
assign w6402 = ~w14553 & w5398;
assign w6403 = w1391 & ~w3374;
assign w6404 = w709 & pi1893;
assign w6405 = pi0034 & ~w14148;
assign w6406 = (~pi0298 & ~w325) | (~pi0298 & w5206) | (~w325 & w5206);
assign w6407 = ~w17594 & ~w9754;
assign w6408 = w13867 & w13344;
assign w6409 = ~w18467 & ~w7370;
assign w6410 = pi1825 & ~w2732;
assign w6411 = ~w12699 & ~w16586;
assign w6412 = ~w3847 & ~w12345;
assign w6413 = ~w11396 & ~w3558;
assign w6414 = pi1638 & ~w13753;
assign w6415 = ~pi3414 & w15036;
assign w6416 = ~w12700 & ~w11378;
assign w6417 = ~pi2654 & w17213;
assign w6418 = ~pi2790 & w13343;
assign w6419 = w9440 & pi0141;
assign w6420 = ~w12004 & ~w7439;
assign w6421 = pi1555 & ~w18259;
assign w6422 = w12915 & w16388;
assign w6423 = w3120 & w4961;
assign w6424 = ~w5747 & w17697;
assign w6425 = ~pi0114 & w9284;
assign w6426 = pi0115 & w9284;
assign w6427 = ~w1368 & ~pi0456;
assign w6428 = ~w7838 & ~w6606;
assign w6429 = ~w3225 & ~w7404;
assign w6430 = w13509 & w4460;
assign w6431 = ~w16908 & w4497;
assign w6432 = ~w1417 & ~w9900;
assign w6433 = (pi0603 & ~w13509) | (pi0603 & w7749) | (~w13509 & w7749);
assign w6434 = ~w11926 & w12648;
assign w6435 = pi0092 & w3748;
assign w6436 = ~pi2741 & w17213;
assign w6437 = ~w15871 & ~w13457;
assign w6438 = ~w5643 & ~w4629;
assign w6439 = pi2672 & ~w6463;
assign w6440 = ~w11676 & ~w6341;
assign w6441 = ~w6670 & w6511;
assign w6442 = w7643 & w18366;
assign w6443 = ~w1160 & ~w13254;
assign w6444 = pi1400 & ~w7946;
assign w6445 = ~w18299 & ~w162;
assign w6446 = pi1578 & w13753;
assign w6447 = w15842 & w13584;
assign w6448 = pi1371 & w6024;
assign w6449 = pi2473 & ~w10299;
assign w6450 = w7703 & w2239;
assign w6451 = ~w5766 & ~w2282;
assign w6452 = ~w8549 & ~w10203;
assign w6453 = pi2820 & ~w15235;
assign w6454 = ~w12643 & ~w6728;
assign w6455 = ~pi2258 & w13065;
assign w6456 = w2341 & ~w6680;
assign w6457 = w6788 & w13274;
assign w6458 = ~pi1985 & ~w7140;
assign w6459 = pi0070 & ~w14148;
assign w6460 = ~pi3138 & pi0002;
assign w6461 = w1063 & w15038;
assign w6462 = w11232 & w10801;
assign w6463 = ~pi2949 & w7912;
assign w6464 = ~w3054 & w2226;
assign w6465 = pi2166 & ~w15271;
assign w6466 = pi0008 & ~w14148;
assign w6467 = ~w16440 & ~w11756;
assign w6468 = w8214 & w18109;
assign w6469 = ~w5391 & ~w14682;
assign w6470 = ~pi3095 & w6463;
assign w6471 = ~w5595 & w193;
assign w6472 = ~pi0294 & w2196;
assign w6473 = ~w1688 & w9158;
assign w6474 = ~pi2282 & w13065;
assign w6475 = w6697 & ~w2587;
assign w6476 = ~w3243 & ~w3351;
assign w6477 = (w7693 & ~w10247) | (w7693 & w11645) | (~w10247 & w11645);
assign w6478 = ~pi3055 & w3555;
assign w6479 = ~w14560 & pi0235;
assign w6480 = w3948 & w10888;
assign w6481 = ~w8496 & ~w12322;
assign w6482 = ~w14746 & ~w3207;
assign w6483 = pi2872 & w14148;
assign w6484 = w7077 & ~w3374;
assign w6485 = w14228 & ~w3430;
assign w6486 = ~w12760 & w108;
assign w6487 = ~pi1304 & ~w17477;
assign w6488 = ~w965 & ~w11868;
assign w6489 = ~pi2199 & w9340;
assign w6490 = pi1646 & ~w13753;
assign w6491 = ~pi2012 & w11688;
assign w6492 = w13509 & w7832;
assign w6493 = w384 & w6694;
assign w6494 = ~w5309 & ~w8300;
assign w6495 = w13262 & w6683;
assign w6496 = ~pi1002 & w12825;
assign w6497 = ~w9707 & ~w12834;
assign w6498 = pi1922 & ~w10299;
assign w6499 = pi1762 & pi2465;
assign w6500 = ~w16506 & pi1140;
assign w6501 = pi1411 & ~w6072;
assign w6502 = ~w18096 & ~w8063;
assign w6503 = ~w11095 & w15097;
assign w6504 = ~w8436 & ~w18143;
assign w6505 = w13509 & w11808;
assign w6506 = ~w12332 & ~w6146;
assign w6507 = ~pi3131 & w1843;
assign w6508 = w17741 & w5357;
assign w6509 = w14560 & pi0357;
assign w6510 = ~pi0711 & w3106;
assign w6511 = w10647 & ~w7602;
assign w6512 = ~w2592 & ~w2941;
assign w6513 = ~w11317 & ~w14910;
assign w6514 = ~w16278 & pi0983;
assign w6515 = w9440 & pi0173;
assign w6516 = w13509 & w18193;
assign w6517 = ~w3000 & ~pi2798;
assign w6518 = w13509 & w8854;
assign w6519 = w7307 & w15340;
assign w6520 = w13509 & w4112;
assign w6521 = ~pi3145 & w13570;
assign w6522 = pi0307 & ~w4667;
assign w6523 = ~w4021 & ~w3408;
assign w6524 = w1846 & ~w8823;
assign w6525 = ~w11990 & ~w4323;
assign w6526 = pi2155 & ~w11671;
assign w6527 = ~w12217 & w8994;
assign w6528 = ~pi3146 & w17387;
assign w6529 = (pi0819 & ~w13509) | (pi0819 & w1000) | (~w13509 & w1000);
assign w6530 = ~w8242 & ~w8439;
assign w6531 = ~w3248 & ~w4697;
assign w6532 = ~w6056 & ~pi0085;
assign w6533 = ~pi3287 & w6448;
assign w6534 = pi2063 & ~w4508;
assign w6535 = pi2370 & ~w18123;
assign w6536 = pi1265 & pi2960;
assign w6537 = ~w3753 & ~w1369;
assign w6538 = ~pi3155 & w13730;
assign w6539 = w11812 & w16042;
assign w6540 = w13509 & w8977;
assign w6541 = ~pi3088 & w15235;
assign w6542 = ~w1197 & ~w9670;
assign w6543 = ~pi3092 & w226;
assign w6544 = ~w9000 & ~w14644;
assign w6545 = pi2283 & ~w3223;
assign w6546 = ~w1953 & w16594;
assign w6547 = ~w2341 & pi0840;
assign w6548 = ~w962 & ~w16440;
assign w6549 = w16506 & ~w14978;
assign w6550 = ~pi0776 & w6200;
assign w6551 = ~w8848 & ~w3115;
assign w6552 = ~w18565 & ~w2963;
assign w6553 = ~w18559 & ~w2929;
assign w6554 = w934 & pi0446;
assign w6555 = ~w2650 & w120;
assign w6556 = (pi0619 & ~w13509) | (pi0619 & w15339) | (~w13509 & w15339);
assign w6557 = ~w3325 & ~w16302;
assign w6558 = ~w7538 & ~w18139;
assign w6559 = pi3158 & w3987;
assign w6560 = (w5517 & w17230) | (w5517 & w11116) | (w17230 & w11116);
assign w6561 = pi1858 & ~pi0273;
assign w6562 = w16575 & w18216;
assign w6563 = ~w11193 & ~w14925;
assign w6564 = (pi1158 & ~w5437) | (pi1158 & w14274) | (~w5437 & w14274);
assign w6565 = ~w790 & ~w7467;
assign w6566 = ~w7264 & ~w812;
assign w6567 = w14782 & w2920;
assign w6568 = (pi0357 & w6195) | (pi0357 & w6509) | (w6195 & w6509);
assign w6569 = pi0054 & pi0066;
assign w6570 = pi0512 & pi1150;
assign w6571 = pi3188 & pi3243;
assign w6572 = ~w11529 & ~w4356;
assign w6573 = ~pi0309 & pi0265;
assign w6574 = ~w759 & w11672;
assign w6575 = ~w8504 & ~w18142;
assign w6576 = ~pi0687 & w9110;
assign w6577 = ~w3223 & ~w7829;
assign w6578 = ~w15122 & ~pi2504;
assign w6579 = ~w8725 & ~w15482;
assign w6580 = ~pi0609 & w12825;
assign w6581 = pi1319 & w458;
assign w6582 = w15808 & ~w12800;
assign w6583 = pi1473 & ~w9781;
assign w6584 = w7698 & w14647;
assign w6585 = w15808 & ~w7449;
assign w6586 = ~w15206 & ~w16473;
assign w6587 = ~w17940 & w12557;
assign w6588 = pi0093 & w3748;
assign w6589 = pi0101 & w3748;
assign w6590 = ~w5180 & ~w8937;
assign w6591 = pi1493 & w13753;
assign w6592 = ~w1980 & ~w10106;
assign w6593 = w16771 & ~w11102;
assign w6594 = ~w7077 & pi0818;
assign w6595 = (pi0826 & ~w13509) | (pi0826 & w13263) | (~w13509 & w13263);
assign w6596 = ~w16497 & ~w7661;
assign w6597 = ~w5631 & ~w10090;
assign w6598 = ~w9962 & ~w18154;
assign w6599 = ~w9536 & ~w7244;
assign w6600 = ~w7018 & ~w11571;
assign w6601 = ~w15220 & ~w16098;
assign w6602 = w4364 & ~pi0436;
assign w6603 = w709 & pi2958;
assign w6604 = ~pi0584 & w795;
assign w6605 = ~w9750 & ~w17650;
assign w6606 = ~pi1194 & ~w11010;
assign w6607 = w17857 & w13568;
assign w6608 = ~w4439 & w6223;
assign w6609 = ~w16278 & pi0710;
assign w6610 = pi2116 & ~w412;
assign w6611 = w11876 & w11552;
assign w6612 = ~w16575 & w7893;
assign w6613 = pi2936 & w6045;
assign w6614 = ~w4562 & ~w16627;
assign w6615 = pi1660 & ~w13753;
assign w6616 = (~pi1199 & ~w13509) | (~pi1199 & w16741) | (~w13509 & w16741);
assign w6617 = pi3117 & ~pi3120;
assign w6618 = ~w17847 & ~w16437;
assign w6619 = ~pi2988 & w15235;
assign w6620 = ~pi1071 & w1147;
assign w6621 = ~w4733 & ~w183;
assign w6622 = ~w14976 & ~w11611;
assign w6623 = (pi0583 & ~w13509) | (pi0583 & w10926) | (~w13509 & w10926);
assign w6624 = pi1397 & w12817;
assign w6625 = ~w4211 & ~w15396;
assign w6626 = w10676 & w15213;
assign w6627 = w6045 & w2004;
assign w6628 = ~w6785 & ~pi0950;
assign w6629 = w13509 & w11604;
assign w6630 = pi1947 & ~w17646;
assign w6631 = ~pi3059 & w226;
assign w6632 = ~pi3164 & pi3207;
assign w6633 = ~pi0932 & w3106;
assign w6634 = ~w6785 & pi1048;
assign w6635 = pi2898 & ~w3555;
assign w6636 = ~w7537 & ~w8613;
assign w6637 = ~pi3139 & w13570;
assign w6638 = ~pi2822 & w13343;
assign w6639 = ~w11341 & ~w5006;
assign w6640 = pi1392 & ~w17935;
assign w6641 = ~pi2922 & w4095;
assign w6642 = ~pi3133 & pi3165;
assign w6643 = w1368 & pi0378;
assign w6644 = ~pi0645 & w3791;
assign w6645 = w12708 & w7154;
assign w6646 = (~pi1313 & ~w11356) | (~pi1313 & w7389) | (~w11356 & w7389);
assign w6647 = ~w6231 & ~w823;
assign w6648 = ~pi2351 & w12755;
assign w6649 = w8430 & w16095;
assign w6650 = pi2459 & ~w11671;
assign w6651 = ~pi1094 & w17490;
assign w6652 = ~w6441 & ~w10459;
assign w6653 = ~pi0751 & w17490;
assign w6654 = w13509 & w15091;
assign w6655 = w12460 & w338;
assign w6656 = pi1606 & ~w7090;
assign w6657 = ~w12128 & w16801;
assign w6658 = ~w4620 & ~w12843;
assign w6659 = w13691 & ~w16459;
assign w6660 = ~w9806 & ~w1968;
assign w6661 = w9151 & w6394;
assign w6662 = ~w6785 & pi0518;
assign w6663 = pi3015 & ~w3987;
assign w6664 = (pi2920 & ~w384) | (pi2920 & w12754) | (~w384 & w12754);
assign w6665 = ~w2727 & ~w12240;
assign w6666 = ~w2211 & ~w9359;
assign w6667 = (pi0391 & w5560) | (pi0391 & w10306) | (w5560 & w10306);
assign w6668 = w13509 & w1399;
assign w6669 = pi2142 & ~w15883;
assign w6670 = pi1641 & ~w13753;
assign w6671 = (pi1096 & ~w13509) | (pi1096 & w5112) | (~w13509 & w5112);
assign w6672 = w7844 & ~w10235;
assign w6673 = ~pi2922 & ~w6045;
assign w6674 = ~pi3010 & ~pi3207;
assign w6675 = ~w1005 & ~w15066;
assign w6676 = pi1152 & ~pi1154;
assign w6677 = ~pi1011 & w3791;
assign w6678 = ~w12654 & ~w1624;
assign w6679 = pi2738 & ~w5274;
assign w6680 = ~w3853 & ~w11973;
assign w6681 = ~pi3164 & w11132;
assign w6682 = w9884 & w7700;
assign w6683 = ~w3923 & ~w7840;
assign w6684 = pi2163 & ~w9504;
assign w6685 = w14833 & w9407;
assign w6686 = pi2843 & w14148;
assign w6687 = w12193 & w8275;
assign w6688 = w3402 & ~w18501;
assign w6689 = ~w14330 & ~w9731;
assign w6690 = ~pi1207 & w17490;
assign w6691 = w17562 & pi1822;
assign w6692 = ~w9842 & ~w9803;
assign w6693 = ~w8135 & ~w12106;
assign w6694 = w15842 & pi2482;
assign w6695 = ~w15392 & w7696;
assign w6696 = w11383 & w2981;
assign w6697 = w28 & w13679;
assign w6698 = pi1265 & w10552;
assign w6699 = pi0043 & w15064;
assign w6700 = w13231 & ~w14143;
assign w6701 = ~pi2716 & w17213;
assign w6702 = pi1445 & ~w13753;
assign w6703 = ~w1104 & ~w1542;
assign w6704 = w17646 & w9407;
assign w6705 = ~w7007 & ~w15611;
assign w6706 = w10189 & ~pi0474;
assign w6707 = ~w4376 & ~w2628;
assign w6708 = ~w1077 & ~w18319;
assign w6709 = pi0113 & ~w17632;
assign w6710 = ~w13613 & ~w16804;
assign w6711 = pi2621 & ~w16815;
assign w6712 = ~w4650 & ~w1874;
assign w6713 = pi2833 & ~w226;
assign w6714 = ~w1623 & ~w11636;
assign w6715 = w9440 & pi0200;
assign w6716 = ~pi2180 & w5384;
assign w6717 = ~w1302 & ~w9314;
assign w6718 = pi1676 & ~w17062;
assign w6719 = ~pi2655 & w17213;
assign w6720 = pi2931 & ~w16815;
assign w6721 = ~w5081 & ~w3242;
assign w6722 = pi1403 & w4683;
assign w6723 = pi1452 & w13753;
assign w6724 = pi2351 & ~w412;
assign w6725 = w1962 & ~w14465;
assign w6726 = w14275 & ~w15689;
assign w6727 = w5437 & w8684;
assign w6728 = ~pi1833 & ~w11735;
assign w6729 = w15758 & w7022;
assign w6730 = ~w18585 & ~w7202;
assign w6731 = pi1581 & ~w14918;
assign w6732 = ~pi3050 & w11406;
assign w6733 = (pi0382 & w5560) | (pi0382 & w1272) | (w5560 & w1272);
assign w6734 = w13231 & ~w6680;
assign w6735 = ~w13096 & ~w13462;
assign w6736 = pi2287 & ~w4508;
assign w6737 = w16575 & w7570;
assign w6738 = ~pi2189 & w2151;
assign w6739 = ~w5560 & w14585;
assign w6740 = pi0452 & pi3364;
assign w6741 = ~w12909 & ~w10707;
assign w6742 = ~w17558 & ~w13610;
assign w6743 = ~w13231 & pi0563;
assign w6744 = ~w1962 & pi0636;
assign w6745 = (pi0699 & ~w13509) | (pi0699 & w8675) | (~w13509 & w8675);
assign w6746 = ~w8569 & w1326;
assign w6747 = ~pi3030 & pi3138;
assign w6748 = ~w7656 & pi1212;
assign w6749 = pi1341 & ~w5762;
assign w6750 = pi2850 & w14148;
assign w6751 = w17248 & ~w3374;
assign w6752 = ~w5952 & ~w12876;
assign w6753 = w6649 & ~w7297;
assign w6754 = ~w10391 & w5010;
assign w6755 = w18127 & w194;
assign w6756 = (~w10679 & ~w5517) | (~w10679 & w11019) | (~w5517 & w11019);
assign w6757 = w13509 & w8942;
assign w6758 = pi0302 & w5274;
assign w6759 = pi1709 & ~w7946;
assign w6760 = ~pi1811 & w8230;
assign w6761 = ~pi1204 & w795;
assign w6762 = ~pi3056 & w261;
assign w6763 = w14293 & w5809;
assign w6764 = ~pi0705 & w3106;
assign w6765 = pi1422 & ~w6072;
assign w6766 = ~pi3045 & w11406;
assign w6767 = pi0008 & ~w3748;
assign w6768 = (pi1187 & ~w5437) | (pi1187 & w5699) | (~w5437 & w5699);
assign w6769 = pi2751 & ~w6463;
assign w6770 = w15808 & ~w2776;
assign w6771 = w13509 & w17736;
assign w6772 = ~w3750 & ~w9972;
assign w6773 = ~w4675 & ~w7823;
assign w6774 = ~w4243 & ~w2243;
assign w6775 = pi3151 & pi3158;
assign w6776 = ~w16482 & ~w8782;
assign w6777 = ~pi3142 & w1843;
assign w6778 = ~pi2899 & w17213;
assign w6779 = w12040 & ~w13195;
assign w6780 = ~pi3166 & w13730;
assign w6781 = ~pi1169 & ~pi3198;
assign w6782 = ~pi1095 & w11739;
assign w6783 = ~w17248 & pi1125;
assign w6784 = ~pi2064 & w8617;
assign w6785 = w2613 & w3988;
assign w6786 = (pi0945 & ~w13509) | (pi0945 & w17759) | (~w13509 & w17759);
assign w6787 = ~pi2909 & ~pi2919;
assign w6788 = w14880 & w2919;
assign w6789 = ~w11281 & w11544;
assign w6790 = ~w5250 & ~w5185;
assign w6791 = w11671 & w17115;
assign w6792 = w7519 & w11982;
assign w6793 = ~w15808 & pi0749;
assign w6794 = ~pi3154 & w15048;
assign w6795 = ~pi0897 & w12825;
assign w6796 = ~w9512 & ~w10187;
assign w6797 = ~w132 & ~w2674;
assign w6798 = ~pi3299 & w16922;
assign w6799 = ~pi0515 & ~w13367;
assign w6800 = ~w2822 & ~w7680;
assign w6801 = pi1344 & ~pi3120;
assign w6802 = (~pi0950 & ~w13509) | (~pi0950 & w6628) | (~w13509 & w6628);
assign w6803 = w13509 & w8217;
assign w6804 = w13175 & ~w5614;
assign w6805 = ~pi0483 & pi3406;
assign w6806 = ~w2740 & ~w12566;
assign w6807 = ~w12500 & ~w17492;
assign w6808 = w15808 & ~w305;
assign w6809 = ~pi2020 & w11688;
assign w6810 = ~w15122 & ~pi2764;
assign w6811 = ~w17320 & w998;
assign w6812 = ~pi1263 & w4880;
assign w6813 = w1391 & ~w7707;
assign w6814 = ~w17889 & w6571;
assign w6815 = (pi1871 & w2014) | (pi1871 & w17291) | (w2014 & w17291);
assign w6816 = ~pi2915 & pi2917;
assign w6817 = w1391 & ~w1340;
assign w6818 = ~pi3286 & w6072;
assign w6819 = w8337 & pi3356;
assign w6820 = ~w11580 & ~w3895;
assign w6821 = w13509 & w10648;
assign w6822 = ~w16759 & w15922;
assign w6823 = ~pi3095 & w226;
assign w6824 = w13801 & w13949;
assign w6825 = w14109 & pi0413;
assign w6826 = ~pi1686 & ~w4899;
assign w6827 = w5383 & pi2966;
assign w6828 = pi1532 & w13753;
assign w6829 = (pi0911 & ~w13509) | (pi0911 & w9669) | (~w13509 & w9669);
assign w6830 = ~pi3354 & w6448;
assign w6831 = ~pi3138 & w14753;
assign w6832 = w13509 & w8711;
assign w6833 = ~w17185 & ~w12102;
assign w6834 = w9440 & pi0161;
assign w6835 = pi2112 & ~w412;
assign w6836 = ~pi1057 & w1126;
assign w6837 = ~w10236 & w16819;
assign w6838 = ~w7212 & w13430;
assign w6839 = ~pi1840 & ~w11671;
assign w6840 = pi0309 & ~w18262;
assign w6841 = ~w16644 & ~w11112;
assign w6842 = ~w7077 & pi0812;
assign w6843 = w11345 & w8261;
assign w6844 = w11345 & w8262;
assign w6845 = ~w11284 & ~w8771;
assign w6846 = pi1501 & ~w13753;
assign w6847 = pi1183 & ~w12368;
assign w6848 = ~pi2993 & ~pi3207;
assign w6849 = pi1717 & ~pi3153;
assign w6850 = w7844 & ~w4043;
assign w6851 = ~w14535 & ~w7217;
assign w6852 = ~w3243 & pi0324;
assign w6853 = w12817 & w876;
assign w6854 = ~w8606 & ~w1200;
assign w6855 = ~w7844 & pi0610;
assign w6856 = ~w2129 & ~w5213;
assign w6857 = ~w325 & ~w16897;
assign w6858 = ~w13301 & ~w5930;
assign w6859 = ~w8033 & ~w15490;
assign w6860 = ~w13159 & ~w3074;
assign w6861 = ~w12519 & ~w1616;
assign w6862 = ~w2 & ~w15128;
assign w6863 = ~pi3169 & pi3171;
assign w6864 = pi1514 & w13753;
assign w6865 = pi2966 & pi2584;
assign w6866 = ~w14228 & pi0549;
assign w6867 = ~w18349 & ~w13105;
assign w6868 = (~pi0335 & w3055) | (~pi0335 & w12746) | (w3055 & w12746);
assign w6869 = w8596 & w6423;
assign w6870 = ~pi0492 & w4501;
assign w6871 = ~w11057 & ~w6719;
assign w6872 = ~pi1307 & ~pi3213;
assign w6873 = w16703 & pi0066;
assign w6874 = w384 & w9215;
assign w6875 = w417 & w10695;
assign w6876 = pi3147 & w12558;
assign w6877 = w13193 & ~w18088;
assign w6878 = ~w12550 & ~w13475;
assign w6879 = pi2995 & w2460;
assign w6880 = pi3018 & w3987;
assign w6881 = ~w5402 & ~w2869;
assign w6882 = w13509 & w9057;
assign w6883 = pi1491 & ~w9781;
assign w6884 = pi2308 & ~w15883;
assign w6885 = pi2478 & ~w14524;
assign w6886 = ~pi0496 & ~pi1345;
assign w6887 = ~w1368 & ~pi0465;
assign w6888 = ~pi3094 & w226;
assign w6889 = ~w2593 & ~w14041;
assign w6890 = ~w1989 & ~w9042;
assign w6891 = ~pi0985 & w15707;
assign w6892 = (pi1097 & ~w13509) | (pi1097 & w14318) | (~w13509 & w14318);
assign w6893 = pi1342 & ~w18281;
assign w6894 = w12040 & ~w11978;
assign w6895 = pi2527 & w15191;
assign w6896 = w17955 & ~w11129;
assign w6897 = ~w1095 & ~w15737;
assign w6898 = (pi0702 & ~w13509) | (pi0702 & w2818) | (~w13509 & w2818);
assign w6899 = ~w1090 & ~w14872;
assign w6900 = ~pi2030 & w7455;
assign w6901 = pi1546 & ~w17935;
assign w6902 = ~pi1884 & w13343;
assign w6903 = ~w12460 & w1584;
assign w6904 = ~w6521 & ~w12731;
assign w6905 = ~w13964 & ~w10143;
assign w6906 = ~w14670 & pi1198;
assign w6907 = ~w14766 & ~w10696;
assign w6908 = ~pi0798 & w543;
assign w6909 = ~w2154 & ~w11001;
assign w6910 = ~w16693 & ~w10033;
assign w6911 = ~w3682 & ~w17496;
assign w6912 = w10818 & ~w14476;
assign w6913 = pi0249 & pi0263;
assign w6914 = ~pi2376 & w16041;
assign w6915 = ~pi3157 & w13730;
assign w6916 = pi0120 & pi3207;
assign w6917 = (~pi1302 & ~w11356) | (~pi1302 & w4341) | (~w11356 & w4341);
assign w6918 = ~w337 & ~w775;
assign w6919 = pi1713 & ~w619;
assign w6920 = w7799 & w17562;
assign w6921 = ~w2903 & w9249;
assign w6922 = ~w9194 & ~w14131;
assign w6923 = w968 & ~pi0327;
assign w6924 = w14648 & ~pi2718;
assign w6925 = w412 & w17115;
assign w6926 = w772 & w8187;
assign w6927 = ~pi2304 & w8617;
assign w6928 = (~w1698 & ~w1206) | (~w1698 & w12422) | (~w1206 & w12422);
assign w6929 = ~pi2395 & w16041;
assign w6930 = ~w12054 & ~w7392;
assign w6931 = (pi1117 & ~w13509) | (pi1117 & w9982) | (~w13509 & w9982);
assign w6932 = ~pi0982 & w14641;
assign w6933 = pi2696 & ~w9504;
assign w6934 = w14560 & pi0375;
assign w6935 = ~pi0511 & ~pi1345;
assign w6936 = ~pi3058 & w3555;
assign w6937 = ~w2725 & pi0797;
assign w6938 = ~w12040 & pi1021;
assign w6939 = pi2217 & ~w11735;
assign w6940 = ~w12385 & ~w10430;
assign w6941 = ~w16064 & ~w8926;
assign w6942 = ~w13658 & ~w14050;
assign w6943 = pi2401 & ~w14524;
assign w6944 = ~pi3096 & w226;
assign w6945 = pi3139 & ~pi3141;
assign w6946 = w12460 & w12934;
assign w6947 = ~w15495 & ~w4102;
assign w6948 = ~w18534 & ~w3368;
assign w6949 = ~w1430 & ~w17922;
assign w6950 = (pi0492 & ~w11345) | (pi0492 & w10166) | (~w11345 & w10166);
assign w6951 = w7844 & ~w15296;
assign w6952 = ~w2725 & pi0782;
assign w6953 = (pi0926 & ~w13509) | (pi0926 & w13851) | (~w13509 & w13851);
assign w6954 = ~pi3014 & ~pi3207;
assign w6955 = ~w7897 & ~w10397;
assign w6956 = ~w7212 & ~w11288;
assign w6957 = (~pi0328 & ~w6857) | (~pi0328 & w11398) | (~w6857 & w11398);
assign w6958 = pi0133 & w9653;
assign w6959 = w1127 & ~w14183;
assign w6960 = w16759 & w16235;
assign w6961 = ~pi1083 & w543;
assign w6962 = pi3041 & w16502;
assign w6963 = (pi0713 & ~w13509) | (pi0713 & w809) | (~w13509 & w809);
assign w6964 = ~w9661 & ~w8112;
assign w6965 = ~pi0644 & w3791;
assign w6966 = w10904 & w11126;
assign w6967 = ~w7836 & ~w15168;
assign w6968 = (pi0860 & ~w13509) | (pi0860 & w4801) | (~w13509 & w4801);
assign w6969 = w6785 & ~w14465;
assign w6970 = ~w11889 & ~w12066;
assign w6971 = ~w15115 & ~w8688;
assign w6972 = pi1380 & ~w9781;
assign w6973 = w13509 & w12065;
assign w6974 = ~pi0598 & w12825;
assign w6975 = ~w5926 & ~w12936;
assign w6976 = ~w18546 & ~w9465;
assign w6977 = ~w7195 & ~w7580;
assign w6978 = ~w2060 & ~w15367;
assign w6979 = pi2671 & ~w6463;
assign w6980 = ~w9071 & ~w6483;
assign w6981 = pi3366 & w7536;
assign w6982 = ~w12492 & ~w4623;
assign w6983 = ~w8229 & w1326;
assign w6984 = pi0049 & w4954;
assign w6985 = pi1729 & ~w4058;
assign w6986 = ~w9964 & ~w10914;
assign w6987 = pi1380 & w13753;
assign w6988 = ~w17982 & ~w14032;
assign w6989 = ~w1661 & ~w8058;
assign w6990 = ~pi2803 & w13343;
assign w6991 = ~w1552 & ~w4311;
assign w6992 = pi2715 & ~w9504;
assign w6993 = ~pi1112 & w14641;
assign w6994 = w16278 & ~w4179;
assign w6995 = ~pi3343 & w17935;
assign w6996 = ~pi3084 & w226;
assign w6997 = ~w1835 & ~w13017;
assign w6998 = ~pi0969 & w17899;
assign w6999 = ~w14699 & ~w11357;
assign w7000 = ~w8958 & ~w16309;
assign w7001 = ~pi0483 & pi3396;
assign w7002 = w17248 & ~w13028;
assign w7003 = ~w2099 & w12955;
assign w7004 = ~w6071 & ~w5446;
assign w7005 = pi2815 & ~w11406;
assign w7006 = pi1764 & pi3171;
assign w7007 = pi2393 & ~w14524;
assign w7008 = ~pi0744 & w17490;
assign w7009 = (pi0802 & ~w13509) | (pi0802 & w13947) | (~w13509 & w13947);
assign w7010 = w3196 & w754;
assign w7011 = pi2562 & ~w5274;
assign w7012 = ~pi1797 & ~pi3158;
assign w7013 = w14109 & pi0417;
assign w7014 = ~w14920 & ~w12238;
assign w7015 = ~pi0507 & ~w13843;
assign w7016 = w16965 & ~pi3070;
assign w7017 = pi2906 & w8304;
assign w7018 = w16575 & w8634;
assign w7019 = pi3145 & w3987;
assign w7020 = ~pi1290 & pi1345;
assign w7021 = pi1291 & pi1345;
assign w7022 = ~w15650 & ~w11255;
assign w7023 = w13509 & w18172;
assign w7024 = ~w10587 & ~w8038;
assign w7025 = (w10417 & ~w13878) | (w10417 & w10590) | (~w13878 & w10590);
assign w7026 = ~w15808 & pi0755;
assign w7027 = ~pi2007 & w11688;
assign w7028 = pi3160 & ~pi3479;
assign w7029 = ~pi2471 & w5384;
assign w7030 = ~w642 & ~w9082;
assign w7031 = ~pi0515 & ~pi0503;
assign w7032 = ~w16555 & ~w6199;
assign w7033 = w14705 & ~w1225;
assign w7034 = (pi0940 & ~w13509) | (pi0940 & w7650) | (~w13509 & w7650);
assign w7035 = ~w14560 & pi0211;
assign w7036 = ~w1673 & ~w7207;
assign w7037 = ~w3000 & ~pi2742;
assign w7038 = w934 & pi0421;
assign w7039 = w6857 & w14357;
assign w7040 = pi1337 & ~pi0256;
assign w7041 = pi1337 & pi0257;
assign w7042 = pi2133 & ~w15883;
assign w7043 = ~pi2126 & w16041;
assign w7044 = ~w7572 & ~w7985;
assign w7045 = pi0266 & ~pi3217;
assign w7046 = ~pi1841 & ~w9414;
assign w7047 = ~pi1331 & ~w3987;
assign w7048 = ~w15131 & ~w9678;
assign w7049 = pi1488 & ~w9781;
assign w7050 = pi2529 & w15191;
assign w7051 = pi1484 & w13753;
assign w7052 = pi2902 & ~w226;
assign w7053 = ~w17203 & ~w17951;
assign w7054 = (pi0625 & ~w13509) | (pi0625 & w5362) | (~w13509 & w5362);
assign w7055 = w934 & pi0441;
assign w7056 = w10313 & w10412;
assign w7057 = w11345 & w2283;
assign w7058 = pi1866 & ~w458;
assign w7059 = ~pi3341 & w6448;
assign w7060 = w14269 & ~w1225;
assign w7061 = ~pi3350 & w14918;
assign w7062 = ~w1791 & w15901;
assign w7063 = ~pi3298 & w18259;
assign w7064 = ~w2944 & ~w16538;
assign w7065 = pi2262 & ~w11671;
assign w7066 = w14986 & w13477;
assign w7067 = ~w15042 & ~w14837;
assign w7068 = pi2453 & ~w14524;
assign w7069 = ~w7194 & ~w2362;
assign w7070 = ~pi3155 & w3982;
assign w7071 = ~w8201 & ~w8170;
assign w7072 = pi2089 & ~w4420;
assign w7073 = ~pi1092 & w11739;
assign w7074 = w11383 & w1868;
assign w7075 = ~w12225 & ~w2515;
assign w7076 = ~w11750 & ~w11996;
assign w7077 = w28 & w3988;
assign w7078 = pi1495 & ~w16922;
assign w7079 = w12460 & w6715;
assign w7080 = w13509 & w3076;
assign w7081 = ~w179 & ~w2017;
assign w7082 = ~pi2278 & w5384;
assign w7083 = pi3160 & ~w489;
assign w7084 = w12460 & w11086;
assign w7085 = ~w13231 & ~pi0951;
assign w7086 = ~w4306 & ~w15850;
assign w7087 = pi2477 & ~w14524;
assign w7088 = ~w1886 & w9337;
assign w7089 = (pi1125 & ~w13509) | (pi1125 & w6783) | (~w13509 & w6783);
assign w7090 = w667 & w4517;
assign w7091 = ~pi3353 & w6072;
assign w7092 = w8337 & pi3344;
assign w7093 = pi0335 & ~pi0338;
assign w7094 = ~pi1314 & ~w11356;
assign w7095 = w11722 & w5925;
assign w7096 = pi2273 & ~w4420;
assign w7097 = ~pi3131 & ~pi3160;
assign w7098 = pi0489 & pi0490;
assign w7099 = ~w3203 & pi0575;
assign w7100 = ~w14647 & ~w5953;
assign w7101 = w6432 & w4450;
assign w7102 = pi2300 & ~w18123;
assign w7103 = pi2538 & w14148;
assign w7104 = ~pi2378 & w12755;
assign w7105 = ~w5413 & ~w2934;
assign w7106 = ~w7077 & pi1079;
assign w7107 = w13509 & w13833;
assign w7108 = ~w1520 & ~w13314;
assign w7109 = pi0298 & w5113;
assign w7110 = (pi0518 & ~w13509) | (pi0518 & w6662) | (~w13509 & w6662);
assign w7111 = w13509 & w5660;
assign w7112 = ~w9541 & ~w3147;
assign w7113 = w5339 & w8379;
assign w7114 = ~w14756 & ~w4007;
assign w7115 = ~w16359 & ~w17340;
assign w7116 = ~pi3007 & ~pi3102;
assign w7117 = w14560 & pi0353;
assign w7118 = w15122 & ~pi2292;
assign w7119 = ~w3839 & ~w3178;
assign w7120 = ~pi1369 & w5043;
assign w7121 = ~w5880 & ~w11875;
assign w7122 = ~pi0141 & pi0189;
assign w7123 = ~w3482 & ~w14169;
assign w7124 = w16575 & w16425;
assign w7125 = w17562 & pi1847;
assign w7126 = ~w6389 & ~w8532;
assign w7127 = w12058 & w1722;
assign w7128 = ~pi0073 & w922;
assign w7129 = pi1472 & w13753;
assign w7130 = ~w5648 & ~w7690;
assign w7131 = pi2111 & ~w412;
assign w7132 = ~w2597 & ~w14369;
assign w7133 = pi2537 & w14148;
assign w7134 = ~w1537 & w542;
assign w7135 = ~w15568 & ~w17604;
assign w7136 = w14903 & w18336;
assign w7137 = pi2783 & ~w11406;
assign w7138 = (pi0267 & w3055) | (pi0267 & w14614) | (w3055 & w14614);
assign w7139 = ~w17730 & ~w13363;
assign w7140 = pi1984 & w3981;
assign w7141 = ~pi3058 & w11406;
assign w7142 = ~pi3146 & w4310;
assign w7143 = ~pi2972 & w13207;
assign w7144 = ~w13663 & ~w3506;
assign w7145 = ~w18472 & ~w8138;
assign w7146 = w1391 & ~w10235;
assign w7147 = ~w14648 & ~pi2720;
assign w7148 = ~w6534 & ~w8248;
assign w7149 = pi2225 & ~w15271;
assign w7150 = pi2887 & ~w226;
assign w7151 = w384 & w15698;
assign w7152 = pi1385 & ~w17935;
assign w7153 = w17646 & w17115;
assign w7154 = ~w4695 & ~w9251;
assign w7155 = pi2708 & ~w3555;
assign w7156 = ~pi3049 & w226;
assign w7157 = ~w15473 & ~w10667;
assign w7158 = w4281 & w13813;
assign w7159 = ~w18424 & ~w4975;
assign w7160 = ~w10131 & ~w13054;
assign w7161 = ~pi2969 & w131;
assign w7162 = ~w3054 & w1919;
assign w7163 = ~w6702 & w4214;
assign w7164 = w15253 & w10468;
assign w7165 = ~w6697 & pi0920;
assign w7166 = pi1376 & ~w945;
assign w7167 = ~w368 & w9117;
assign w7168 = ~w3243 & pi0337;
assign w7169 = w1962 & ~w2776;
assign w7170 = pi2718 & ~w261;
assign w7171 = pi2611 & ~w261;
assign w7172 = ~pi2046 & w13204;
assign w7173 = w13509 & w15523;
assign w7174 = ~pi3139 & pi3141;
assign w7175 = pi2953 & w6045;
assign w7176 = pi3160 & ~pi3504;
assign w7177 = (w3003 & ~w14705) | (w3003 & w12703) | (~w14705 & w12703);
assign w7178 = (pi0998 & ~w13509) | (pi0998 & w4516) | (~w13509 & w4516);
assign w7179 = ~w9160 & ~w5663;
assign w7180 = pi2430 & ~w3223;
assign w7181 = pi2577 & ~w5274;
assign w7182 = w3203 & ~w2587;
assign w7183 = ~w6620 & ~w11781;
assign w7184 = pi1172 & pi3192;
assign w7185 = ~w2503 & ~w5720;
assign w7186 = ~pi0627 & w14641;
assign w7187 = (pi0673 & ~w13509) | (pi0673 & w1771) | (~w13509 & w1771);
assign w7188 = ~pi2975 & w10158;
assign w7189 = ~w14245 & ~w12298;
assign w7190 = ~w2341 & pi0839;
assign w7191 = pi0253 & w5113;
assign w7192 = ~w5097 & w3274;
assign w7193 = w539 & ~w9496;
assign w7194 = ~w16575 & w9252;
assign w7195 = pi0301 & w9853;
assign w7196 = ~w2138 & ~w12407;
assign w7197 = ~w8220 & ~w17752;
assign w7198 = ~w16506 & pi1156;
assign w7199 = ~pi1680 & pi2465;
assign w7200 = ~w17153 & w2610;
assign w7201 = w11578 & w8983;
assign w7202 = pi1369 & ~pi3233;
assign w7203 = ~w8880 & ~w7063;
assign w7204 = ~w839 & ~w3766;
assign w7205 = ~w10375 & ~w14554;
assign w7206 = ~w5560 & w16307;
assign w7207 = w13509 & w17961;
assign w7208 = pi2854 & w14148;
assign w7209 = ~pi0322 & ~pi3229;
assign w7210 = pi3051 & ~pi3158;
assign w7211 = (pi1044 & ~w13509) | (pi1044 & w9127) | (~w13509 & w9127);
assign w7212 = ~pi1337 & w325;
assign w7213 = ~w14401 & w10101;
assign w7214 = w11383 & w9649;
assign w7215 = w7799 & w5453;
assign w7216 = w13509 & w17072;
assign w7217 = w12460 & w4951;
assign w7218 = ~pi3155 & w12427;
assign w7219 = w16511 & w4913;
assign w7220 = w384 & w12576;
assign w7221 = pi2503 & ~w5274;
assign w7222 = ~pi1768 & pi3151;
assign w7223 = pi1552 & w13753;
assign w7224 = (pi0917 & ~w13509) | (pi0917 & w2327) | (~w13509 & w2327);
assign w7225 = ~w3203 & pi0585;
assign w7226 = ~w18297 & ~w12652;
assign w7227 = ~pi3066 & pi3163;
assign w7228 = ~w12370 & w10623;
assign w7229 = ~w13367 & ~w1007;
assign w7230 = pi2015 & ~w14833;
assign w7231 = ~w12059 & ~w6243;
assign w7232 = ~w17911 & ~w16465;
assign w7233 = (w15842 & ~w2971) | (w15842 & w4920) | (~w2971 & w4920);
assign w7234 = (pi1860 & w2014) | (pi1860 & w17663) | (w2014 & w17663);
assign w7235 = ~w6713 & ~w4291;
assign w7236 = w384 & w688;
assign w7237 = w17436 & w5625;
assign w7238 = w10818 & ~w1441;
assign w7239 = ~w10292 & ~w4867;
assign w7240 = w17043 & w4122;
assign w7241 = ~pi2340 & w5075;
assign w7242 = pi1730 & w1924;
assign w7243 = ~w13702 & ~w3902;
assign w7244 = ~pi2792 & w13343;
assign w7245 = ~pi1305 & w6352;
assign w7246 = ~w17373 & ~w5303;
assign w7247 = ~pi3088 & w261;
assign w7248 = w14738 & pi0325;
assign w7249 = w13509 & w16475;
assign w7250 = w8679 & pi1313;
assign w7251 = ~pi1062 & w12825;
assign w7252 = ~w5450 & w12448;
assign w7253 = w12359 & w8029;
assign w7254 = ~pi1152 & ~pi1154;
assign w7255 = ~w14795 & ~w7770;
assign w7256 = ~w11915 & w75;
assign w7257 = w15808 & ~w2587;
assign w7258 = pi1639 & ~w18259;
assign w7259 = pi2203 & ~w4420;
assign w7260 = (~pi0293 & ~w6857) | (~pi0293 & w16221) | (~w6857 & w16221);
assign w7261 = ~w5199 & ~w11873;
assign w7262 = ~pi3170 & w13570;
assign w7263 = ~w16575 & w13830;
assign w7264 = pi2602 & ~w16815;
assign w7265 = w16212 & w15180;
assign w7266 = ~pi0672 & w12197;
assign w7267 = ~w14151 & ~w2478;
assign w7268 = w10647 & ~w17088;
assign w7269 = ~w15784 & ~w17050;
assign w7270 = w16278 & ~w3430;
assign w7271 = (pi1055 & ~w13509) | (pi1055 & w1137) | (~w13509 & w1137);
assign w7272 = w12589 & w14669;
assign w7273 = ~pi3058 & w6463;
assign w7274 = (~w10377 & w9490) | (~w10377 & w13127) | (w9490 & w13127);
assign w7275 = ~w6433 & ~w7960;
assign w7276 = (pi1207 & ~w13509) | (pi1207 & w6249) | (~w13509 & w6249);
assign w7277 = w1225 & w14767;
assign w7278 = w3987 & w15106;
assign w7279 = ~w14136 & ~w1481;
assign w7280 = ~w3018 & ~w5441;
assign w7281 = pi2461 & ~w7399;
assign w7282 = ~w4317 & ~w5671;
assign w7283 = ~w393 & w3995;
assign w7284 = ~w3648 & ~w14232;
assign w7285 = (pi1147 & ~w5437) | (pi1147 & w12575) | (~w5437 & w12575);
assign w7286 = pi1597 & ~w16922;
assign w7287 = ~w13979 & ~w3740;
assign w7288 = ~pi0789 & w543;
assign w7289 = ~pi0484 & ~pi3117;
assign w7290 = (w17562 & ~w8098) | (w17562 & w15350) | (~w8098 & w15350);
assign w7291 = ~pi1199 & w17899;
assign w7292 = ~pi2133 & w12941;
assign w7293 = ~w7459 & ~w3589;
assign w7294 = ~w16274 & ~w6486;
assign w7295 = ~pi2976 & w11406;
assign w7296 = pi3156 & pi3249;
assign w7297 = pi1453 & w13753;
assign w7298 = ~w2588 & ~w16152;
assign w7299 = w9499 & w11332;
assign w7300 = pi1686 & pi2912;
assign w7301 = w7703 & w6176;
assign w7302 = ~w7656 & pi1180;
assign w7303 = pi2422 & ~w3223;
assign w7304 = ~w16575 & w17159;
assign w7305 = (pi1790 & w5453) | (pi1790 & w8322) | (w5453 & w8322);
assign w7306 = w17103 & w3335;
assign w7307 = ~w14648 & ~w15122;
assign w7308 = (pi0607 & ~w13509) | (pi0607 & w11065) | (~w13509 & w11065);
assign w7309 = ~w12745 & ~w13879;
assign w7310 = ~pi2281 & w13065;
assign w7311 = w5747 & ~w17697;
assign w7312 = ~w15224 & ~w4514;
assign w7313 = ~w4984 & ~w7558;
assign w7314 = ~pi1078 & w11739;
assign w7315 = w9440 & pi0178;
assign w7316 = ~w16865 & ~w15266;
assign w7317 = w968 & ~pi0291;
assign w7318 = ~w13279 & ~w16427;
assign w7319 = pi3023 & ~w3987;
assign w7320 = ~pi1013 & w12197;
assign w7321 = ~w8034 & ~w2629;
assign w7322 = pi1331 & pi2969;
assign w7323 = ~pi0040 & w922;
assign w7324 = w3398 & w17085;
assign w7325 = ~w1454 & ~w13082;
assign w7326 = w5437 & w17034;
assign w7327 = pi1338 & w7799;
assign w7328 = (w6406 & ~w7807) | (w6406 & w1530) | (~w7807 & w1530);
assign w7329 = pi2052 & ~w10158;
assign w7330 = ~pi0483 & pi3386;
assign w7331 = pi3033 & pi3155;
assign w7332 = pi2597 & ~w9504;
assign w7333 = w13509 & w18494;
assign w7334 = w6857 & w5592;
assign w7335 = w6857 & w17430;
assign w7336 = ~w4054 & ~w13496;
assign w7337 = pi2145 & ~w11671;
assign w7338 = ~w9440 & w10959;
assign w7339 = w7844 & ~w6922;
assign w7340 = w6785 & ~w2741;
assign w7341 = pi1676 & ~w9302;
assign w7342 = ~pi2068 & w8617;
assign w7343 = ~w4422 & ~w9925;
assign w7344 = ~pi3423 & w15036;
assign w7345 = ~pi1766 & pi3162;
assign w7346 = w14856 & w17618;
assign w7347 = ~pi1989 & w3019;
assign w7348 = w2482 & w4976;
assign w7349 = ~pi2369 & w17439;
assign w7350 = ~pi3169 & w17993;
assign w7351 = ~w13465 & ~w13660;
assign w7352 = ~w6785 & pi0853;
assign w7353 = ~w4972 & ~w16728;
assign w7354 = ~w3851 & ~w17091;
assign w7355 = w11383 & w14568;
assign w7356 = w1127 & ~w1109;
assign w7357 = ~w3109 & ~w3224;
assign w7358 = ~w1791 & w4557;
assign w7359 = w4667 & pi1232;
assign w7360 = ~pi3314 & w16922;
assign w7361 = ~w5189 & pi1123;
assign w7362 = ~w18037 & ~w1666;
assign w7363 = w4140 & w876;
assign w7364 = ~pi3133 & w13570;
assign w7365 = (~w13367 & w17577) | (~w13367 & w14110) | (w17577 & w14110);
assign w7366 = ~w14228 & pi0517;
assign w7367 = pi1651 & ~w13753;
assign w7368 = ~pi2170 & w11313;
assign w7369 = ~w8932 & ~w18547;
assign w7370 = pi3136 & w13786;
assign w7371 = pi0273 & w14001;
assign w7372 = pi2251 & ~w9414;
assign w7373 = pi2208 & ~w3223;
assign w7374 = pi1633 & ~w13753;
assign w7375 = ~pi3086 & w11406;
assign w7376 = w13147 & w974;
assign w7377 = pi1627 & ~w18259;
assign w7378 = ~pi3169 & w13730;
assign w7379 = ~w8302 & ~w1385;
assign w7380 = ~w2341 & ~pi0976;
assign w7381 = ~w15122 & ~pi2676;
assign w7382 = w1913 & w8789;
assign w7383 = ~pi1949 & w7455;
assign w7384 = w13509 & w17848;
assign w7385 = ~pi2438 & w9340;
assign w7386 = w13509 & w9978;
assign w7387 = ~w14427 & ~w7581;
assign w7388 = ~w17534 & ~w15084;
assign w7389 = ~w8679 & ~pi1313;
assign w7390 = w13509 & w5825;
assign w7391 = (~w11450 & ~w9420) | (~w11450 & w222) | (~w9420 & w222);
assign w7392 = w13509 & w12300;
assign w7393 = ~w8938 & w6916;
assign w7394 = ~w9592 & ~w11641;
assign w7395 = ~pi3139 & w17387;
assign w7396 = ~w7645 & w18057;
assign w7397 = ~w3000 & ~pi2800;
assign w7398 = pi0050 & ~w14148;
assign w7399 = ~pi2294 & w3229;
assign w7400 = w13509 & w10142;
assign w7401 = ~pi1909 & w5384;
assign w7402 = ~w5571 & ~w9149;
assign w7403 = pi2871 & w15191;
assign w7404 = ~pi0604 & w12825;
assign w7405 = ~pi0929 & w3106;
assign w7406 = ~w12585 & ~w14695;
assign w7407 = w3203 & ~w7707;
assign w7408 = pi2903 & ~w3555;
assign w7409 = w13870 & w7789;
assign w7410 = w2725 & w1217;
assign w7411 = ~pi3095 & w261;
assign w7412 = w15122 & ~pi2628;
assign w7413 = ~w6737 & ~w1849;
assign w7414 = ~w14801 & ~w7360;
assign w7415 = pi2156 & ~w11671;
assign w7416 = (pi0767 & ~w13509) | (pi0767 & w8274) | (~w13509 & w8274);
assign w7417 = ~pi3341 & w16922;
assign w7418 = pi1988 & ~w9414;
assign w7419 = w7307 & w15572;
assign w7420 = w15421 & ~w13967;
assign w7421 = ~pi0422 & w17173;
assign w7422 = pi0423 & w17173;
assign w7423 = (pi0397 & w5560) | (pi0397 & w7548) | (w5560 & w7548);
assign w7424 = ~w15052 & ~w8831;
assign w7425 = ~w2109 & ~w3759;
assign w7426 = w5437 & w16319;
assign w7427 = ~w13231 & pi0564;
assign w7428 = (pi0300 & ~w325) | (pi0300 & w10861) | (~w325 & w10861);
assign w7429 = w5437 & w10470;
assign w7430 = pi0152 & w5274;
assign w7431 = (pi0668 & ~w13509) | (pi0668 & w5259) | (~w13509 & w5259);
assign w7432 = ~w11050 & ~w7898;
assign w7433 = ~w3203 & pi0996;
assign w7434 = ~w3973 & w15310;
assign w7435 = ~w3055 & w12305;
assign w7436 = ~pi1126 & w14641;
assign w7437 = w13509 & w14305;
assign w7438 = ~w3434 & ~w17355;
assign w7439 = ~pi3053 & w15235;
assign w7440 = ~w16278 & pi0705;
assign w7441 = ~pi3347 & w9781;
assign w7442 = ~pi2994 & w18259;
assign w7443 = ~pi0992 & w11739;
assign w7444 = ~pi3020 & ~pi3160;
assign w7445 = ~pi1027 & w3106;
assign w7446 = ~pi3316 & w14918;
assign w7447 = ~w1196 & w9138;
assign w7448 = pi2866 & w15191;
assign w7449 = ~w12196 & ~w14879;
assign w7450 = w12040 & ~w7707;
assign w7451 = ~pi1751 & pi3158;
assign w7452 = pi0081 & ~w6536;
assign w7453 = w11345 & w6805;
assign w7454 = ~pi3162 & w3805;
assign w7455 = w13807 & w5767;
assign w7456 = w11671 & w9407;
assign w7457 = pi3171 & w14951;
assign w7458 = ~w12149 & ~w13627;
assign w7459 = ~pi1723 & pi3150;
assign w7460 = w10818 & ~w7717;
assign w7461 = ~w15579 & ~w3184;
assign w7462 = ~pi0907 & w795;
assign w7463 = w13509 & w5151;
assign w7464 = w13509 & w1944;
assign w7465 = w13509 & w1945;
assign w7466 = ~w2581 & ~w197;
assign w7467 = w5437 & w9601;
assign w7468 = pi3163 & w7946;
assign w7469 = ~w10900 & ~w2161;
assign w7470 = pi1477 & w13753;
assign w7471 = ~w11737 & ~w2132;
assign w7472 = ~w8696 & ~w14302;
assign w7473 = ~w6022 & w2633;
assign w7474 = w13509 & w13778;
assign w7475 = w9414 & w9407;
assign w7476 = w10534 & w6279;
assign w7477 = pi3185 & pi3250;
assign w7478 = pi2130 & ~w18123;
assign w7479 = ~pi2534 & pi2920;
assign w7480 = ~w14228 & pi0624;
assign w7481 = ~w12093 & ~w15515;
assign w7482 = pi1464 & ~w7090;
assign w7483 = ~w3055 & w16851;
assign w7484 = ~pi0147 & ~w8912;
assign w7485 = w2725 & ~w17513;
assign w7486 = pi0250 & w5113;
assign w7487 = w14560 & pi0371;
assign w7488 = ~pi0498 & pi1145;
assign w7489 = w4097 & w7232;
assign w7490 = (pi0852 & ~w13509) | (pi0852 & w433) | (~w13509 & w433);
assign w7491 = pi1881 & ~w15235;
assign w7492 = ~pi2171 & w11313;
assign w7493 = ~pi1363 & ~pi2920;
assign w7494 = ~pi1937 & w16041;
assign w7495 = pi2771 & ~w11406;
assign w7496 = w13509 & w18491;
assign w7497 = ~w3017 & w14419;
assign w7498 = w9474 & w12840;
assign w7499 = ~w9828 & ~w4488;
assign w7500 = pi1371 & ~w5043;
assign w7501 = ~w13779 & ~w5395;
assign w7502 = ~w7844 & pi0609;
assign w7503 = ~w7755 & ~w7400;
assign w7504 = ~w5997 & ~w18137;
assign w7505 = (~pi0264 & ~w6857) | (~pi0264 & w486) | (~w6857 & w486);
assign w7506 = ~w12346 & ~w4437;
assign w7507 = pi1724 & w1027;
assign w7508 = w432 & w14956;
assign w7509 = ~w6446 & w10818;
assign w7510 = ~w18499 & ~w7333;
assign w7511 = ~pi0496 & ~pi1143;
assign w7512 = ~pi3147 & w13730;
assign w7513 = (pi0503 & ~w7031) | (pi0503 & ~w17577) | (~w7031 & ~w17577);
assign w7514 = w10189 & pi0399;
assign w7515 = w1127 & ~w7223;
assign w7516 = ~w13189 & ~w8806;
assign w7517 = w13509 & w3144;
assign w7518 = w9720 & pi1753;
assign w7519 = w13265 & w4448;
assign w7520 = ~pi0502 & pi1148;
assign w7521 = w4692 & w16988;
assign w7522 = ~w15298 & ~w10806;
assign w7523 = pi1619 & ~w16922;
assign w7524 = ~w12040 & pi0679;
assign w7525 = w16506 & ~w13028;
assign w7526 = pi2628 & ~w9504;
assign w7527 = w17248 & ~w1340;
assign w7528 = w16429 & w6074;
assign w7529 = (pi1099 & ~w13509) | (pi1099 & w13978) | (~w13509 & w13978);
assign w7530 = w5453 & pi2581;
assign w7531 = w13509 & w4618;
assign w7532 = w7807 & w17376;
assign w7533 = w15540 & w3552;
assign w7534 = w6857 & w10264;
assign w7535 = ~pi3128 & w16815;
assign w7536 = ~pi3364 & ~pi3365;
assign w7537 = pi1868 & ~w15036;
assign w7538 = w11511 & w16521;
assign w7539 = ~w12636 & ~w14468;
assign w7540 = ~w5294 & ~w15635;
assign w7541 = w9474 & ~w17809;
assign w7542 = ~w16506 & pi1135;
assign w7543 = ~w16575 & w16198;
assign w7544 = ~w1962 & pi0641;
assign w7545 = ~pi3133 & w17993;
assign w7546 = ~w13829 & ~w15262;
assign w7547 = (w12732 & ~w4413) | (w12732 & w13155) | (~w4413 & w13155);
assign w7548 = w1368 & pi0397;
assign w7549 = w16278 & ~w17513;
assign w7550 = ~pi3056 & w3555;
assign w7551 = pi2192 & ~w11735;
assign w7552 = pi0037 & ~w14148;
assign w7553 = w9720 & pi1721;
assign w7554 = w18123 & w17115;
assign w7555 = ~w14478 & ~w6631;
assign w7556 = pi3147 & ~pi3168;
assign w7557 = pi1760 & ~w10389;
assign w7558 = pi1705 & w4667;
assign w7559 = ~w6195 & w1797;
assign w7560 = ~pi0301 & ~w1206;
assign w7561 = ~w12706 & ~w10433;
assign w7562 = ~pi1835 & ~w4508;
assign w7563 = ~w17913 & ~w5139;
assign w7564 = w17021 & w4576;
assign w7565 = (~w13367 & w17577) | (~w13367 & w13382) | (w17577 & w13382);
assign w7566 = ~w7258 & ~w14157;
assign w7567 = ~w17248 & pi1120;
assign w7568 = ~pi1917 & w11313;
assign w7569 = ~w5189 & ~pi0970;
assign w7570 = w10189 & ~pi0466;
assign w7571 = (pi0594 & ~w13509) | (pi0594 & w12269) | (~w13509 & w12269);
assign w7572 = pi1615 & ~w7090;
assign w7573 = w9440 & pi0166;
assign w7574 = ~pi0335 & pi0337;
assign w7575 = (pi0302 & ~w325) | (pi0302 & w3353) | (~w325 & w3353);
assign w7576 = ~w3455 & ~w11083;
assign w7577 = ~w10908 & ~w13466;
assign w7578 = ~pi2967 & ~pi3044;
assign w7579 = ~pi3053 & w3555;
assign w7580 = (pi0261 & ~w325) | (pi0261 & w177) | (~w325 & w177);
assign w7581 = ~pi0276 & w4058;
assign w7582 = ~w1705 & w408;
assign w7583 = ~w7015 & w7565;
assign w7584 = ~w2725 & ~pi0978;
assign w7585 = pi1806 & ~w7177;
assign w7586 = ~w10143 & ~w15886;
assign w7587 = ~w15172 & ~w15481;
assign w7588 = ~w16999 & ~w13459;
assign w7589 = w12040 & ~w16498;
assign w7590 = ~w12165 & ~w14584;
assign w7591 = ~w6195 & w438;
assign w7592 = w7799 & w6127;
assign w7593 = (~w13063 & ~w14073) | (~w13063 & w15653) | (~w14073 & w15653);
assign w7594 = ~pi3287 & w18259;
assign w7595 = ~w15246 & ~w14409;
assign w7596 = pi1561 & ~w13753;
assign w7597 = ~w5560 & w1915;
assign w7598 = ~pi3050 & w9504;
assign w7599 = w1326 & w1291;
assign w7600 = w539 & ~w1345;
assign w7601 = ~w6722 & w16719;
assign w7602 = pi1604 & w13753;
assign w7603 = w2341 & ~w15296;
assign w7604 = w5437 & w17500;
assign w7605 = w7077 & ~w17210;
assign w7606 = pi1864 & ~w458;
assign w7607 = w12460 & w16604;
assign w7608 = w8992 & w3494;
assign w7609 = ~w13562 & ~w13951;
assign w7610 = ~w3980 & ~w12137;
assign w7611 = ~pi2261 & w13065;
assign w7612 = pi2100 & ~w4420;
assign w7613 = w2341 & w11302;
assign w7614 = pi1675 & w1924;
assign w7615 = ~w7416 & ~w8210;
assign w7616 = w7307 & w6276;
assign w7617 = ~pi2988 & w11406;
assign w7618 = w968 & ~pi0284;
assign w7619 = ~w12040 & pi0694;
assign w7620 = ~pi1403 & ~pi1404;
assign w7621 = ~w11605 & ~w8366;
assign w7622 = pi1705 & ~w18497;
assign w7623 = ~pi2156 & w13065;
assign w7624 = ~pi3316 & w7090;
assign w7625 = ~w2176 & w1521;
assign w7626 = ~w14560 & pi0218;
assign w7627 = ~w9746 & ~w9300;
assign w7628 = w8789 & w9684;
assign w7629 = pi3070 & ~w16502;
assign w7630 = w17597 & w14189;
assign w7631 = w13476 & w18207;
assign w7632 = w13509 & w7182;
assign w7633 = ~pi1206 & w14641;
assign w7634 = w13509 & w16610;
assign w7635 = w6697 & w11302;
assign w7636 = ~w5361 & ~w15824;
assign w7637 = w8337 & pi3274;
assign w7638 = ~w17656 & w73;
assign w7639 = w10189 & pi0388;
assign w7640 = w7343 & w5276;
assign w7641 = ~w12793 & ~w6505;
assign w7642 = ~w7490 & ~w12289;
assign w7643 = w12684 & w4727;
assign w7644 = ~pi1951 & w7455;
assign w7645 = w11383 & w8952;
assign w7646 = pi3171 & w619;
assign w7647 = ~w14648 & ~pi1879;
assign w7648 = (pi1206 & w4470) | (pi1206 & w7955) | (w4470 & w7955);
assign w7649 = pi2613 & ~w261;
assign w7650 = ~w12040 & pi0940;
assign w7651 = ~w13649 & ~w13685;
assign w7652 = ~w5855 & w5818;
assign w7653 = pi0507 & pi1151;
assign w7654 = w17683 & w9407;
assign w7655 = ~pi2896 & w15122;
assign w7656 = ~w1368 & ~w13762;
assign w7657 = pi0411 & ~pi3376;
assign w7658 = pi0060 & pi0061;
assign w7659 = ~w3000 & ~pi1977;
assign w7660 = w13509 & w14995;
assign w7661 = w13509 & w15857;
assign w7662 = ~w17444 & ~w9146;
assign w7663 = ~pi3336 & w18259;
assign w7664 = ~pi1298 & w14158;
assign w7665 = pi1773 & ~pi3139;
assign w7666 = w1962 & ~w7707;
assign w7667 = ~w8324 & ~w4912;
assign w7668 = (pi2952 & w2014) | (pi2952 & w10185) | (w2014 & w10185);
assign w7669 = w934 & pi0416;
assign w7670 = ~w6195 & w18576;
assign w7671 = ~w7077 & pi0810;
assign w7672 = w6857 & w7038;
assign w7673 = w13509 & w13313;
assign w7674 = ~w12349 & ~w9045;
assign w7675 = w13509 & w10977;
assign w7676 = ~pi2352 & w12724;
assign w7677 = ~pi3154 & w1843;
assign w7678 = ~pi0800 & w543;
assign w7679 = ~w3808 & ~w16831;
assign w7680 = pi2115 & ~w412;
assign w7681 = ~w15427 & ~w6038;
assign w7682 = ~w11455 & w14254;
assign w7683 = ~w15122 & ~pi2902;
assign w7684 = pi2933 & ~w261;
assign w7685 = ~pi1721 & pi3135;
assign w7686 = pi0262 & w5113;
assign w7687 = ~w12274 & ~w12133;
assign w7688 = w6188 & w3962;
assign w7689 = ~pi2354 & w12724;
assign w7690 = ~pi2383 & w5384;
assign w7691 = w11209 & ~w13854;
assign w7692 = ~w2238 & w13284;
assign w7693 = ~w228 & ~w10408;
assign w7694 = (pi1046 & ~w13509) | (pi1046 & w15793) | (~w13509 & w15793);
assign w7695 = w3166 & w17528;
assign w7696 = ~pi0081 & ~w7296;
assign w7697 = w709 & pi1892;
assign w7698 = ~pi3120 & ~pi3129;
assign w7699 = ~w10226 & w12905;
assign w7700 = ~w16481 & w5243;
assign w7701 = ~w2163 & ~w11540;
assign w7702 = ~pi3040 & ~pi3207;
assign w7703 = w14648 & w3000;
assign w7704 = ~w1391 & pi1091;
assign w7705 = w4348 & w3138;
assign w7706 = ~w3946 & ~w12672;
assign w7707 = ~w16269 & ~w15051;
assign w7708 = pi2431 & ~w17646;
assign w7709 = ~w14648 & ~pi2516;
assign w7710 = ~w709 & pi1278;
assign w7711 = ~w15237 & ~w1195;
assign w7712 = ~pi2017 & w11688;
assign w7713 = ~pi0894 & w1126;
assign w7714 = ~w5189 & pi0729;
assign w7715 = pi2868 & w15191;
assign w7716 = (~w2388 & ~w9420) | (~w2388 & w8901) | (~w9420 & w8901);
assign w7717 = pi1531 & w13753;
assign w7718 = ~w3830 & ~w9537;
assign w7719 = ~w13645 & ~w958;
assign w7720 = ~w11237 & ~w10717;
assign w7721 = ~w17577 & w4478;
assign w7722 = pi2338 & ~w15883;
assign w7723 = w14648 & ~pi2732;
assign w7724 = w11209 & ~w8343;
assign w7725 = w7688 & ~w7212;
assign w7726 = ~pi0854 & w15707;
assign w7727 = ~w3038 & ~w7646;
assign w7728 = (pi0889 & ~w13509) | (pi0889 & w18539) | (~w13509 & w18539);
assign w7729 = ~w17010 & ~w16368;
assign w7730 = ~pi3350 & w17935;
assign w7731 = ~w5224 & ~w4305;
assign w7732 = w10818 & ~w10831;
assign w7733 = ~w9166 & ~w11785;
assign w7734 = ~w13220 & ~w12889;
assign w7735 = ~pi3382 & w7793;
assign w7736 = pi3068 & ~pi3159;
assign w7737 = ~w12788 & ~w17670;
assign w7738 = (pi0666 & ~w13509) | (pi0666 & w8411) | (~w13509 & w8411);
assign w7739 = ~pi3056 & w15235;
assign w7740 = w13509 & w17366;
assign w7741 = w4347 & w7734;
assign w7742 = ~w5064 & ~w10164;
assign w7743 = w15705 & w6069;
assign w7744 = w14560 & pi0349;
assign w7745 = (~w3651 & w3409) | (~w3651 & w6142) | (w3409 & w6142);
assign w7746 = w13509 & w1070;
assign w7747 = ~w9437 & ~w7475;
assign w7748 = (pi1114 & ~w13509) | (pi1114 & w16209) | (~w13509 & w16209);
assign w7749 = ~w7844 & pi0603;
assign w7750 = (pi1074 & ~w13509) | (pi1074 & w10832) | (~w13509 & w10832);
assign w7751 = ~w15236 & ~w8884;
assign w7752 = ~pi0853 & w15707;
assign w7753 = ~pi0679 & w9110;
assign w7754 = ~w11667 & ~w3475;
assign w7755 = (pi0700 & ~w13509) | (pi0700 & w16471) | (~w13509 & w16471);
assign w7756 = w16278 & ~w10947;
assign w7757 = ~pi2946 & w261;
assign w7758 = w11106 & w303;
assign w7759 = ~w16695 & ~w15603;
assign w7760 = ~w6381 & ~w9892;
assign w7761 = ~w1545 & ~w6470;
assign w7762 = ~pi3343 & w6072;
assign w7763 = ~w10963 & ~w4321;
assign w7764 = pi2097 & ~w4420;
assign w7765 = w4508 & w2753;
assign w7766 = w10209 & w8632;
assign w7767 = ~pi2906 & ~w8304;
assign w7768 = ~w5091 & ~w4360;
assign w7769 = ~w5864 & w5158;
assign w7770 = w13509 & w321;
assign w7771 = ~w9450 & ~w10214;
assign w7772 = ~w6462 & w470;
assign w7773 = ~w2061 & w5436;
assign w7774 = w17562 & pi1819;
assign w7775 = ~pi1007 & w14641;
assign w7776 = ~pi1017 & w9110;
assign w7777 = w10818 & ~w2554;
assign w7778 = ~w76 & ~w13872;
assign w7779 = ~pi2152 & w13065;
assign w7780 = ~w14228 & pi0629;
assign w7781 = pi1163 & pi3180;
assign w7782 = ~pi2260 & w13065;
assign w7783 = ~w6109 & pi1241;
assign w7784 = ~w2078 & ~w14010;
assign w7785 = w384 & w5295;
assign w7786 = ~w14628 & w14917;
assign w7787 = w13509 & w7756;
assign w7788 = ~pi3336 & w9781;
assign w7789 = ~w11204 & ~w4577;
assign w7790 = (pi0613 & ~w13509) | (pi0613 & w10814) | (~w13509 & w10814);
assign w7791 = ~pi2054 & w13204;
assign w7792 = ~w17382 & ~w16529;
assign w7793 = ~pi3380 & ~pi3381;
assign w7794 = ~w4095 & ~w12686;
assign w7795 = ~pi0585 & w795;
assign w7796 = w12460 & w3920;
assign w7797 = ~w15122 & ~pi2745;
assign w7798 = (pi1264 & ~w5437) | (pi1264 & w4485) | (~w5437 & w4485);
assign w7799 = w9720 & w11637;
assign w7800 = pi3143 & w10389;
assign w7801 = ~w8359 & ~w15094;
assign w7802 = w1368 & pi0389;
assign w7803 = w15092 & w8982;
assign w7804 = ~w8324 & ~w16742;
assign w7805 = pi2547 & w14148;
assign w7806 = pi1771 & pi1792;
assign w7807 = w914 & w2786;
assign w7808 = w10647 & ~w5027;
assign w7809 = ~w17932 & ~w16298;
assign w7810 = ~pi3341 & w6072;
assign w7811 = pi3153 & w18497;
assign w7812 = w13509 & w3824;
assign w7813 = ~w5189 & pi0731;
assign w7814 = ~w7215 & ~w8658;
assign w7815 = ~pi2975 & w17683;
assign w7816 = ~w4847 & ~w10363;
assign w7817 = ~w3254 & ~w9058;
assign w7818 = w15808 & ~w2741;
assign w7819 = ~pi3316 & w6072;
assign w7820 = pi2966 & pi2895;
assign w7821 = w13509 & w5178;
assign w7822 = w13509 & w7861;
assign w7823 = w13509 & w7862;
assign w7824 = w4787 & w4370;
assign w7825 = pi2770 & ~w6463;
assign w7826 = pi1512 & ~w13753;
assign w7827 = ~pi1015 & w12197;
assign w7828 = ~w2341 & pi0838;
assign w7829 = pi1983 & ~w2247;
assign w7830 = ~w8115 & ~w610;
assign w7831 = ~pi1090 & w11739;
assign w7832 = w15808 & ~w13195;
assign w7833 = ~w12855 & ~w11499;
assign w7834 = ~pi2071 & w8617;
assign w7835 = ~w2990 & ~w693;
assign w7836 = pi2484 & ~w15235;
assign w7837 = ~pi0136 & pi1878;
assign w7838 = w11010 & ~w6625;
assign w7839 = ~pi2982 & w5453;
assign w7840 = ~pi2065 & w8617;
assign w7841 = ~w16466 & ~w18211;
assign w7842 = w10689 & w9636;
assign w7843 = ~w13380 & w4593;
assign w7844 = w2613 & w15907;
assign w7845 = pi1524 & ~w14918;
assign w7846 = ~pi3145 & w12427;
assign w7847 = ~w6720 & ~w7535;
assign w7848 = pi2189 & ~w11735;
assign w7849 = ~w16267 & ~w11419;
assign w7850 = (~pi0487 & w17577) | (~pi0487 & w16012) | (w17577 & w16012);
assign w7851 = ~pi3013 & pi3134;
assign w7852 = ~w12679 & ~w9558;
assign w7853 = w15121 & w15432;
assign w7854 = pi3163 & w8088;
assign w7855 = pi2717 & ~w16815;
assign w7856 = ~pi1956 & w11688;
assign w7857 = ~w3575 & ~w12019;
assign w7858 = pi1337 & ~w16598;
assign w7859 = w13193 & ~w3435;
assign w7860 = pi2841 & w605;
assign w7861 = w5189 & ~w14143;
assign w7862 = w5189 & ~w13195;
assign w7863 = ~pi3045 & w16815;
assign w7864 = w5349 & w15786;
assign w7865 = w13509 & w8500;
assign w7866 = ~w12040 & pi0686;
assign w7867 = ~w8423 & ~w14690;
assign w7868 = ~pi3155 & ~pi3160;
assign w7869 = ~pi1964 & w11688;
assign w7870 = w6785 & ~w7449;
assign w7871 = ~w5560 & w16613;
assign w7872 = ~w17248 & ~pi0973;
assign w7873 = w7307 & w15444;
assign w7874 = ~w9667 & ~w5922;
assign w7875 = ~w15808 & ~pi0972;
assign w7876 = ~w2891 & ~w2116;
assign w7877 = ~w12131 & ~w12860;
assign w7878 = pi2784 & ~w261;
assign w7879 = ~w4969 & w3238;
assign w7880 = ~pi3157 & w13570;
assign w7881 = ~pi3146 & w3805;
assign w7882 = w12460 & w8452;
assign w7883 = pi0205 & w9021;
assign w7884 = pi2136 & ~w15883;
assign w7885 = ~pi3128 & w15235;
assign w7886 = w7498 & w762;
assign w7887 = ~w8479 & w8071;
assign w7888 = w13509 & w2285;
assign w7889 = ~w15122 & ~pi2810;
assign w7890 = ~w17248 & pi0878;
assign w7891 = (~w3744 & ~w5517) | (~w3744 & w17148) | (~w5517 & w17148);
assign w7892 = ~pi3135 & w15839;
assign w7893 = w10189 & pi0377;
assign w7894 = ~pi0494 & ~pi1158;
assign w7895 = w13509 & w3882;
assign w7896 = pi0495 & pi0510;
assign w7897 = pi2284 & ~w16815;
assign w7898 = ~pi3135 & w14753;
assign w7899 = ~w17337 & ~w16109;
assign w7900 = ~w12987 & w14405;
assign w7901 = ~pi2110 & w12755;
assign w7902 = w12460 & w12220;
assign w7903 = ~pi2090 & w12724;
assign w7904 = pi1728 & w1924;
assign w7905 = ~w18130 & ~w14717;
assign w7906 = ~w315 & w6756;
assign w7907 = (pi1174 & ~w13509) | (pi1174 & w14256) | (~w13509 & w14256);
assign w7908 = ~w13470 & w8041;
assign w7909 = ~w16686 & ~w178;
assign w7910 = pi1483 & ~w9781;
assign w7911 = ~pi0600 & w12825;
assign w7912 = ~pi2923 & w2276;
assign w7913 = ~w17465 & ~w8560;
assign w7914 = pi2615 & ~w261;
assign w7915 = w1368 & pi0379;
assign w7916 = pi1546 & w13753;
assign w7917 = pi2515 & ~w261;
assign w7918 = w6857 & w7055;
assign w7919 = ~pi2121 & w12755;
assign w7920 = ~w5189 & pi0733;
assign w7921 = pi0506 & pi1149;
assign w7922 = w7703 & w12920;
assign w7923 = (pi1026 & ~w13509) | (pi1026 & w3354) | (~w13509 & w3354);
assign w7924 = pi1236 & pi1237;
assign w7925 = (~pi0289 & ~w6857) | (~pi0289 & w8850) | (~w6857 & w8850);
assign w7926 = ~w11356 & ~w14620;
assign w7927 = ~w5373 & ~w17850;
assign w7928 = ~w14599 & ~w13673;
assign w7929 = ~pi2298 & w12941;
assign w7930 = ~w6528 & ~w4612;
assign w7931 = ~w6047 & ~w8686;
assign w7932 = ~pi0979 & w9110;
assign w7933 = ~w15130 & ~w15189;
assign w7934 = pi2268 & ~w9414;
assign w7935 = w17562 & w384;
assign w7936 = w6617 & ~w9527;
assign w7937 = pi2197 & ~w10299;
assign w7938 = ~pi2914 & pi3205;
assign w7939 = ~w17100 & ~w7140;
assign w7940 = ~w13315 & ~w11962;
assign w7941 = (pi0984 & ~w13509) | (pi0984 & w16568) | (~w13509 & w16568);
assign w7942 = ~w10489 & ~w13839;
assign w7943 = ~pi1932 & w11313;
assign w7944 = pi1527 & w13753;
assign w7945 = w2046 & ~w727;
assign w7946 = w4683 & w876;
assign w7947 = w17562 & pi1855;
assign w7948 = (pi0944 & ~w13509) | (pi0944 & w13531) | (~w13509 & w13531);
assign w7949 = pi2105 & ~w4420;
assign w7950 = ~w7844 & pi1002;
assign w7951 = pi2304 & ~w4508;
assign w7952 = ~w12973 & ~w14140;
assign w7953 = w1962 & ~w17513;
assign w7954 = ~pi3353 & w17935;
assign w7955 = ~w5160 & pi1206;
assign w7956 = ~pi0734 & w17899;
assign w7957 = pi0191 & w5274;
assign w7958 = pi3001 & w12689;
assign w7959 = w10726 & w6645;
assign w7960 = w13509 & w4707;
assign w7961 = ~w7027 & ~w10100;
assign w7962 = ~w12796 & ~w2538;
assign w7963 = ~pi2287 & w8617;
assign w7964 = ~w3477 & ~w2242;
assign w7965 = w16893 & w6827;
assign w7966 = ~w14228 & pi0946;
assign w7967 = ~w15122 & ~pi2754;
assign w7968 = ~w13062 & ~w9415;
assign w7969 = pi1926 & ~w10299;
assign w7970 = ~w11782 & ~w14915;
assign w7971 = pi2410 & ~w14524;
assign w7972 = pi0270 & w5274;
assign w7973 = pi1707 & ~pi3147;
assign w7974 = ~pi0842 & w93;
assign w7975 = w17248 & ~w7449;
assign w7976 = ~pi2228 & w11313;
assign w7977 = pi0136 & w5274;
assign w7978 = ~w15831 & ~w11983;
assign w7979 = ~w12980 & ~w17453;
assign w7980 = ~pi3314 & w17935;
assign w7981 = ~pi2988 & w3555;
assign w7982 = ~w1216 & ~w14808;
assign w7983 = ~pi0955 & w12825;
assign w7984 = ~w1391 & pi1036;
assign w7985 = ~pi3321 & w7090;
assign w7986 = pi2644 & ~w261;
assign w7987 = ~w11655 & w18562;
assign w7988 = pi3160 & ~pi3494;
assign w7989 = w8308 & w2152;
assign w7990 = w16278 & ~w14465;
assign w7991 = pi0192 & w5274;
assign w7992 = (pi1120 & ~w13509) | (pi1120 & w7567) | (~w13509 & w7567);
assign w7993 = w17562 & pi2560;
assign w7994 = pi2176 & ~w14524;
assign w7995 = ~w17938 & w10935;
assign w7996 = ~pi1985 & w4254;
assign w7997 = ~w3055 & w18390;
assign w7998 = ~pi3133 & w11701;
assign w7999 = ~w16765 & ~w2470;
assign w8000 = w2648 & w13856;
assign w8001 = w14216 & w1611;
assign w8002 = ~w3203 & pi0909;
assign w8003 = pi2970 & w12458;
assign w8004 = ~w2155 & w363;
assign w8005 = ~w5189 & pi0735;
assign w8006 = w11383 & w2714;
assign w8007 = w12460 & w17177;
assign w8008 = w8337 & pi3279;
assign w8009 = ~w10618 & ~w14764;
assign w8010 = w13509 & w7666;
assign w8011 = (pi0306 & ~w325) | (pi0306 & w15245) | (~w325 & w15245);
assign w8012 = pi1358 & w17413;
assign w8013 = (pi0550 & ~w13509) | (pi0550 & w9851) | (~w13509 & w9851);
assign w8014 = ~w6421 & ~w7594;
assign w8015 = pi0053 & ~w14148;
assign w8016 = ~pi1911 & w5384;
assign w8017 = w14648 & ~pi2644;
assign w8018 = w10647 & ~w9267;
assign w8019 = pi1430 & ~w6448;
assign w8020 = ~w15967 & ~w6784;
assign w8021 = ~w11940 & ~w17008;
assign w8022 = ~w9548 & ~w12715;
assign w8023 = w14560 & pi0367;
assign w8024 = (pi0999 & ~w13509) | (pi0999 & w10980) | (~w13509 & w10980);
assign w8025 = ~w3259 & ~w7617;
assign w8026 = pi1776 & ~w10389;
assign w8027 = w11345 & w14629;
assign w8028 = pi1465 & ~w7090;
assign w8029 = w5494 & w8837;
assign w8030 = w4886 & w519;
assign w8031 = w11209 & ~w6661;
assign w8032 = ~w9836 & ~w14697;
assign w8033 = (pi1061 & ~w13509) | (pi1061 & w6266) | (~w13509 & w6266);
assign w8034 = ~pi3158 & w15048;
assign w8035 = ~w7191 & ~w9229;
assign w8036 = ~w7491 & ~w16444;
assign w8037 = ~w15382 & w10952;
assign w8038 = pi2198 & ~w11735;
assign w8039 = ~w16832 & ~w4071;
assign w8040 = ~w16056 & ~w12829;
assign w8041 = ~w4515 & ~w12671;
assign w8042 = ~pi1685 & ~pi2908;
assign w8043 = ~pi2198 & w2151;
assign w8044 = pi1526 & w13753;
assign w8045 = w14648 & ~pi2615;
assign w8046 = (~pi1773 & ~w7799) | (~pi1773 & w11171) | (~w7799 & w11171);
assign w8047 = ~w4839 & ~w12043;
assign w8048 = pi3154 & w653;
assign w8049 = ~pi1041 & w543;
assign w8050 = (pi0847 & ~w13509) | (pi0847 & w12548) | (~w13509 & w12548);
assign w8051 = w1368 & pi0406;
assign w8052 = ~w9132 & ~w1125;
assign w8053 = w13231 & ~w17513;
assign w8054 = ~w5451 & ~w17145;
assign w8055 = w6857 & w13404;
assign w8056 = (pi0383 & w5560) | (pi0383 & w2495) | (w5560 & w2495);
assign w8057 = ~pi0808 & w1147;
assign w8058 = ~pi3056 & w6463;
assign w8059 = (pi1077 & ~w13509) | (pi1077 & w10913) | (~w13509 & w10913);
assign w8060 = pi3019 & ~w3987;
assign w8061 = ~w9992 & ~w7740;
assign w8062 = ~w12833 & ~w13994;
assign w8063 = pi2963 & ~w3987;
assign w8064 = ~pi2832 & w13343;
assign w8065 = pi1308 & pi1345;
assign w8066 = w7703 & w4213;
assign w8067 = ~w5657 & ~w11446;
assign w8068 = ~pi2987 & w226;
assign w8069 = ~w6491 & ~w7172;
assign w8070 = ~w10567 & ~w2429;
assign w8071 = pi1786 & ~w2508;
assign w8072 = ~w17248 & pi0887;
assign w8073 = ~w10967 & ~w3461;
assign w8074 = (~pi0297 & ~w6857) | (~pi0297 & w13064) | (~w6857 & w13064);
assign w8075 = pi2167 & ~w15271;
assign w8076 = ~w4249 & w9015;
assign w8077 = ~w13607 & ~w11407;
assign w8078 = w13676 & w4652;
assign w8079 = w11010 & w11942;
assign w8080 = ~w13231 & pi0565;
assign w8081 = ~w16998 & w18380;
assign w8082 = ~w12939 & ~w9325;
assign w8083 = pi1713 & pi3134;
assign w8084 = (pi0342 & w6195) | (pi0342 & w11481) | (w6195 & w11481);
assign w8085 = ~pi0909 & w795;
assign w8086 = pi3143 & w12558;
assign w8087 = ~w14705 & w7692;
assign w8088 = w9332 & w876;
assign w8089 = pi1766 & ~pi3162;
assign w8090 = (pi0609 & ~w13509) | (pi0609 & w7502) | (~w13509 & w7502);
assign w8091 = w5383 & pi2864;
assign w8092 = (~pi0494 & ~w11345) | (~pi0494 & w11447) | (~w11345 & w11447);
assign w8093 = ~pi3098 & w9504;
assign w8094 = ~w14152 & w9066;
assign w8095 = ~pi0867 & w15707;
assign w8096 = ~pi0765 & w6200;
assign w8097 = ~w12752 & ~w3612;
assign w8098 = w18047 & w3481;
assign w8099 = pi1482 & w13753;
assign w8100 = ~w15388 & ~w14683;
assign w8101 = ~w8669 & ~w10003;
assign w8102 = ~w2688 & ~w3578;
assign w8103 = ~pi1005 & w14641;
assign w8104 = w16278 & ~w7449;
assign w8105 = w11209 & ~w10294;
assign w8106 = ~pi2270 & w17439;
assign w8107 = ~w2725 & pi0788;
assign w8108 = ~w2725 & pi0799;
assign w8109 = ~w1671 & ~w17876;
assign w8110 = w4711 & w1800;
assign w8111 = w539 & ~w10969;
assign w8112 = ~pi2946 & w9504;
assign w8113 = w9227 & w16345;
assign w8114 = ~w15524 & ~w9517;
assign w8115 = pi1232 & w15084;
assign w8116 = ~w12158 & ~w12295;
assign w8117 = ~w5189 & pi0737;
assign w8118 = ~pi2217 & w2151;
assign w8119 = pi1628 & ~w13753;
assign w8120 = ~w7873 & ~w10385;
assign w8121 = ~w16506 & pi1151;
assign w8122 = ~w9125 & ~w15462;
assign w8123 = (pi2913 & ~w16679) | (pi2913 & w3893) | (~w16679 & w3893);
assign w8124 = pi2451 & ~w10299;
assign w8125 = ~w18406 & w11621;
assign w8126 = (~w8801 & ~w11743) | (~w8801 & w16622) | (~w11743 & w16622);
assign w8127 = ~w15005 & ~w11935;
assign w8128 = (pi0853 & ~w13509) | (pi0853 & w7352) | (~w13509 & w7352);
assign w8129 = ~w13777 & ~w2887;
assign w8130 = ~w2970 & ~w2759;
assign w8131 = w12771 & w8959;
assign w8132 = ~pi2936 & pi3208;
assign w8133 = w12460 & w5777;
assign w8134 = pi2965 & w16502;
assign w8135 = ~pi3105 & pi3169;
assign w8136 = pi1677 & ~w14980;
assign w8137 = ~pi2264 & w13065;
assign w8138 = ~pi2965 & ~pi3207;
assign w8139 = pi3383 & pi3517;
assign w8140 = ~w2247 & ~w6458;
assign w8141 = pi2043 & ~w10158;
assign w8142 = pi1431 & ~w6448;
assign w8143 = ~pi3330 & w14918;
assign w8144 = ~w13231 & ~pi0952;
assign w8145 = w1869 & w14252;
assign w8146 = ~pi2363 & w16041;
assign w8147 = ~pi0452 & pi1686;
assign w8148 = w8956 & w17156;
assign w8149 = w8658 & pi1808;
assign w8150 = w11345 & w3636;
assign w8151 = ~w8657 & ~w7764;
assign w8152 = ~w15163 & ~w11497;
assign w8153 = w4146 & w10239;
assign w8154 = pi0299 & w5113;
assign w8155 = ~w967 & w15782;
assign w8156 = pi1938 & ~w14833;
assign w8157 = ~w10444 & ~w12210;
assign w8158 = ~w2345 & ~w5799;
assign w8159 = ~pi3060 & w11406;
assign w8160 = pi3151 & w5457;
assign w8161 = w539 & ~w1393;
assign w8162 = pi2834 & w14148;
assign w8163 = ~w17252 & ~w18524;
assign w8164 = ~pi3333 & w6448;
assign w8165 = ~pi1987 & w3019;
assign w8166 = pi0253 & w11247;
assign w8167 = (pi0874 & ~w13509) | (pi0874 & w5705) | (~w13509 & w5705);
assign w8168 = ~w16991 & ~w1037;
assign w8169 = ~w12551 & w10593;
assign w8170 = ~w5746 & w7447;
assign w8171 = w13509 & w3203;
assign w8172 = pi2497 & ~w15235;
assign w8173 = ~pi2975 & w15883;
assign w8174 = ~w7034 & ~w2582;
assign w8175 = pi2172 & ~w15271;
assign w8176 = ~pi3145 & w1843;
assign w8177 = (pi1118 & ~w13509) | (pi1118 & w14390) | (~w13509 & w14390);
assign w8178 = pi1603 & ~w9781;
assign w8179 = pi1940 & ~w17683;
assign w8180 = pi0300 & w5274;
assign w8181 = (pi0750 & ~w13509) | (pi0750 & w3684) | (~w13509 & w3684);
assign w8182 = pi0068 & w5642;
assign w8183 = ~pi2075 & w17439;
assign w8184 = (pi0627 & ~w13509) | (pi0627 & w11803) | (~w13509 & w11803);
assign w8185 = pi0007 & ~w14148;
assign w8186 = (pi1787 & w7215) | (pi1787 & w17211) | (w7215 & w17211);
assign w8187 = ~w692 & ~w259;
assign w8188 = ~pi2420 & w13204;
assign w8189 = ~w18405 & ~w18081;
assign w8190 = w3203 & ~w14465;
assign w8191 = ~w13231 & pi0916;
assign w8192 = w13509 & w15898;
assign w8193 = pi2073 & ~w17683;
assign w8194 = w5453 & pi1970;
assign w8195 = ~w8550 & ~w12074;
assign w8196 = ~w13231 & pi1078;
assign w8197 = ~pi2230 & w2151;
assign w8198 = pi0340 & pi3364;
assign w8199 = ~w3734 & ~w18229;
assign w8200 = ~w10261 & w13602;
assign w8201 = w12460 & w4546;
assign w8202 = pi0179 & w5274;
assign w8203 = ~pi1172 & ~pi3192;
assign w8204 = pi2995 & pi1350;
assign w8205 = w9421 & w4666;
assign w8206 = pi1212 & ~pi1213;
assign w8207 = (~pi0258 & ~w325) | (~pi0258 & w18160) | (~w325 & w18160);
assign w8208 = (pi0259 & ~w325) | (pi0259 & w18161) | (~w325 & w18161);
assign w8209 = ~w13038 & ~w9126;
assign w8210 = w13509 & w6817;
assign w8211 = w15842 & w384;
assign w8212 = pi1652 & ~w6072;
assign w8213 = pi1739 & w1924;
assign w8214 = pi2553 & pi2963;
assign w8215 = pi3009 & ~w3987;
assign w8216 = ~w12507 & ~pi2920;
assign w8217 = w3203 & ~w14978;
assign w8218 = ~w10262 & ~w268;
assign w8219 = ~pi3104 & ~pi3207;
assign w8220 = (pi1035 & ~w13509) | (pi1035 & w13890) | (~w13509 & w13890);
assign w8221 = pi0256 & w5113;
assign w8222 = ~pi2975 & w18123;
assign w8223 = ~w12900 & ~w10800;
assign w8224 = ~w3940 & ~w6540;
assign w8225 = (pi0400 & w5560) | (pi0400 & w2635) | (w5560 & w2635);
assign w8226 = ~w5189 & pi0739;
assign w8227 = pi0099 & w3748;
assign w8228 = pi1826 & ~w12558;
assign w8229 = pi2983 & w14742;
assign w8230 = pi0079 & pi0082;
assign w8231 = ~pi0078 & ~pi0081;
assign w8232 = ~w14648 & ~pi2780;
assign w8233 = ~w12388 & ~w3429;
assign w8234 = ~w5903 & ~w1728;
assign w8235 = ~w13008 & ~w5859;
assign w8236 = ~w11679 & ~w9607;
assign w8237 = ~w14385 & ~w5896;
assign w8238 = w5383 & w15842;
assign w8239 = ~pi3080 & pi3141;
assign w8240 = ~w3054 & w4303;
assign w8241 = ~w5387 & ~w3378;
assign w8242 = ~w1791 & w3576;
assign w8243 = ~w7012 & ~w2477;
assign w8244 = ~w13253 & ~w17143;
assign w8245 = ~w15305 & ~w16936;
assign w8246 = pi3168 & w12558;
assign w8247 = ~pi1250 & w11655;
assign w8248 = w4508 & w6320;
assign w8249 = pi2413 & ~w10299;
assign w8250 = w16824 & w3758;
assign w8251 = pi3160 & ~pi3487;
assign w8252 = pi2936 & ~pi3208;
assign w8253 = ~pi3299 & w6448;
assign w8254 = ~pi3165 & w15839;
assign w8255 = w9891 & w11318;
assign w8256 = (~w12775 & w18153) | (~w12775 & w18233) | (w18153 & w18233);
assign w8257 = ~w7606 & ~w15834;
assign w8258 = ~w17281 & ~w13247;
assign w8259 = (~pi0064 & ~w5642) | (~pi0064 & w8330) | (~w5642 & w8330);
assign w8260 = w13509 & w17280;
assign w8261 = ~pi0483 & ~pi3408;
assign w8262 = ~pi0483 & pi3409;
assign w8263 = w7077 & ~w2587;
assign w8264 = pi2951 & ~w6045;
assign w8265 = ~w2646 & w13675;
assign w8266 = w13509 & w7870;
assign w8267 = pi1728 & ~w4058;
assign w8268 = ~w7368 & ~w16463;
assign w8269 = ~pi0834 & w93;
assign w8270 = w5437 & w78;
assign w8271 = ~w3000 & ~pi2802;
assign w8272 = ~w1368 & ~pi0479;
assign w8273 = ~pi0860 & w15707;
assign w8274 = ~w1391 & pi0767;
assign w8275 = w5580 & w16658;
assign w8276 = ~w15063 & w11649;
assign w8277 = pi1316 & w2325;
assign w8278 = pi2779 & w14148;
assign w8279 = ~w13231 & pi0544;
assign w8280 = ~w14650 & ~w2900;
assign w8281 = w9440 & pi0139;
assign w8282 = ~w14761 & ~w11560;
assign w8283 = ~w16575 & w7639;
assign w8284 = ~w16278 & pi1023;
assign w8285 = pi3017 & ~w3987;
assign w8286 = ~w16432 & w4167;
assign w8287 = ~w13529 & w4588;
assign w8288 = w14109 & pi0432;
assign w8289 = ~pi1835 & w8617;
assign w8290 = pi0119 & w3748;
assign w8291 = ~w17549 & ~w17446;
assign w8292 = ~w5830 & ~w14159;
assign w8293 = pi2701 & ~w3555;
assign w8294 = ~w2382 & ~w6893;
assign w8295 = w1962 & ~w13028;
assign w8296 = ~w15700 & ~w2498;
assign w8297 = w7504 & ~w12650;
assign w8298 = w7844 & ~w3430;
assign w8299 = ~pi3107 & ~w3987;
assign w8300 = w18123 & w3515;
assign w8301 = ~w8723 & ~w4816;
assign w8302 = pi3022 & ~w3987;
assign w8303 = w13569 & w11637;
assign w8304 = ~pi3082 & w6045;
assign w8305 = pi1791 & ~w48;
assign w8306 = ~w2208 & ~w12151;
assign w8307 = ~pi0750 & w17490;
assign w8308 = ~w7163 & ~w9443;
assign w8309 = ~pi3133 & w17669;
assign w8310 = ~w9616 & ~w3179;
assign w8311 = ~w11004 & ~w7934;
assign w8312 = ~w16817 & ~w6118;
assign w8313 = w9440 & pi0171;
assign w8314 = pi3114 & ~pi3164;
assign w8315 = ~w15808 & pi0758;
assign w8316 = w13446 & w5238;
assign w8317 = ~w6681 & ~w14348;
assign w8318 = ~pi0673 & w12197;
assign w8319 = ~pi3333 & w6072;
assign w8320 = ~w18567 & ~w5061;
assign w8321 = ~w4684 & w6649;
assign w8322 = pi1768 & pi1790;
assign w8323 = pi1416 & ~w13753;
assign w8324 = ~w5517 & ~w5312;
assign w8325 = ~w16791 & ~w2908;
assign w8326 = pi2911 & w16598;
assign w8327 = ~pi1831 & w7455;
assign w8328 = ~w1391 & pi0770;
assign w8329 = pi1349 & ~w11272;
assign w8330 = ~w13318 & ~pi0064;
assign w8331 = pi3135 & w3987;
assign w8332 = w3243 & ~pi0314;
assign w8333 = ~pi0666 & w12197;
assign w8334 = w16278 & w1217;
assign w8335 = ~w10697 & ~w4357;
assign w8336 = w1206 & w5577;
assign w8337 = ~w968 & pi2486;
assign w8338 = ~w1962 & pi0646;
assign w8339 = (~w17391 & ~w9420) | (~w17391 & w5166) | (~w9420 & w5166);
assign w8340 = pi1610 & w13753;
assign w8341 = w3546 & w1854;
assign w8342 = ~w10545 & ~w16642;
assign w8343 = w4491 & w6437;
assign w8344 = ~pi0950 & w15707;
assign w8345 = ~w8206 & ~w17438;
assign w8346 = ~pi3007 & pi3057;
assign w8347 = w14228 & ~w13028;
assign w8348 = ~w2005 & ~w17979;
assign w8349 = pi1252 & ~pi3228;
assign w8350 = ~w4667 & ~w8115;
assign w8351 = pi1191 & w9420;
assign w8352 = w10647 & ~w4990;
assign w8353 = ~w15162 & ~w17560;
assign w8354 = pi1450 & ~w13753;
assign w8355 = ~w186 & ~w13916;
assign w8356 = w17378 & pi0255;
assign w8357 = ~w9021 & w4399;
assign w8358 = (pi0596 & ~w13509) | (pi0596 & w8690) | (~w13509 & w8690);
assign w8359 = pi1442 & ~w6448;
assign w8360 = w9985 & w16122;
assign w8361 = ~w5249 & ~w18324;
assign w8362 = w13509 & w4602;
assign w8363 = ~pi2967 & ~pi3033;
assign w8364 = pi1720 & ~w8113;
assign w8365 = ~w6327 & ~w5889;
assign w8366 = pi0896 & ~w3452;
assign w8367 = ~pi1943 & w7455;
assign w8368 = ~pi3347 & w6448;
assign w8369 = (pi1028 & ~w13509) | (pi1028 & w14429) | (~w13509 & w14429);
assign w8370 = pi1983 & w4841;
assign w8371 = ~pi3062 & w9504;
assign w8372 = w13509 & w5601;
assign w8373 = ~pi3288 & w14918;
assign w8374 = ~w12230 & w8375;
assign w8375 = (~pi0271 & ~w325) | (~pi0271 & w2861) | (~w325 & w2861);
assign w8376 = ~w5968 & pi1676;
assign w8377 = w6652 & w1150;
assign w8378 = pi0021 & ~w14148;
assign w8379 = w979 & w10713;
assign w8380 = w10666 & w16213;
assign w8381 = ~pi1229 & w11655;
assign w8382 = pi2233 & ~w11735;
assign w8383 = pi0452 & ~pi1687;
assign w8384 = w13509 & w8494;
assign w8385 = ~pi2967 & ~pi3037;
assign w8386 = ~pi3417 & w15036;
assign w8387 = pi2528 & w14148;
assign w8388 = ~w3243 & pi0320;
assign w8389 = ~pi1353 & w12365;
assign w8390 = ~w8640 & ~w9825;
assign w8391 = ~w5741 & ~w16628;
assign w8392 = w1391 & ~w15296;
assign w8393 = pi3057 & ~w9243;
assign w8394 = w14560 & pi0345;
assign w8395 = (~pi0955 & ~w13509) | (~pi0955 & w13798) | (~w13509 & w13798);
assign w8396 = pi2949 & w1804;
assign w8397 = ~w16895 & ~w9973;
assign w8398 = pi2345 & ~w17683;
assign w8399 = pi1661 & ~w13753;
assign w8400 = w13509 & w2357;
assign w8401 = ~w11692 & ~w9083;
assign w8402 = ~pi2337 & w17439;
assign w8403 = pi2368 & ~w15883;
assign w8404 = ~w15942 & ~w14243;
assign w8405 = ~pi2010 & w11688;
assign w8406 = w13509 & w7340;
assign w8407 = pi3132 & w14951;
assign w8408 = (~w17367 & ~w15717) | (~w17367 & w4585) | (~w15717 & w4585);
assign w8409 = w7703 & w5057;
assign w8410 = pi1337 & ~w446;
assign w8411 = ~w6697 & pi0666;
assign w8412 = (pi0723 & ~w13509) | (pi0723 & w15680) | (~w13509 & w15680);
assign w8413 = pi2631 & ~w9504;
assign w8414 = ~pi2422 & w5075;
assign w8415 = ~pi3077 & ~pi3207;
assign w8416 = w14524 & w614;
assign w8417 = w6857 & w1921;
assign w8418 = pi1584 & ~w13753;
assign w8419 = ~w14560 & pi0236;
assign w8420 = ~w10835 & w1371;
assign w8421 = ~w16476 & w1419;
assign w8422 = w14859 & w7269;
assign w8423 = ~pi0144 & ~pi0150;
assign w8424 = ~w10922 & ~w622;
assign w8425 = w5802 & w14396;
assign w8426 = w13509 & w16328;
assign w8427 = ~w8028 & ~w4873;
assign w8428 = pi3159 & w7946;
assign w8429 = ~pi3041 & ~pi3207;
assign w8430 = ~w16679 & ~w5790;
assign w8431 = w3177 & w3372;
assign w8432 = ~w4855 & ~w13644;
assign w8433 = ~w12226 & ~w14085;
assign w8434 = ~pi3145 & w15839;
assign w8435 = ~pi0276 & w2196;
assign w8436 = ~w3485 & w15638;
assign w8437 = ~w17026 & ~w6903;
assign w8438 = w968 & ~pi0332;
assign w8439 = ~pi2436 & w17213;
assign w8440 = ~pi3133 & w17387;
assign w8441 = pi0126 & ~pi0128;
assign w8442 = ~pi0566 & w11739;
assign w8443 = w539 & ~w6539;
assign w8444 = ~pi0483 & pi3399;
assign w8445 = pi1367 & ~w5043;
assign w8446 = w13143 & w11412;
assign w8447 = pi0060 & w922;
assign w8448 = ~pi0910 & w6200;
assign w8449 = ~w187 & ~w9116;
assign w8450 = pi2914 & ~w6045;
assign w8451 = ~w16620 & ~w13367;
assign w8452 = w9440 & pi0198;
assign w8453 = ~w6388 & ~w9105;
assign w8454 = ~w17595 & ~w5325;
assign w8455 = w709 & pi1876;
assign w8456 = ~w2437 & w12211;
assign w8457 = ~w6972 & ~w14938;
assign w8458 = w16893 & w16560;
assign w8459 = ~w4765 & ~w3064;
assign w8460 = w2341 & ~w15173;
assign w8461 = w62 & w10359;
assign w8462 = ~w18417 & w18326;
assign w8463 = w14648 & ~pi2630;
assign w8464 = ~w14999 & ~w1936;
assign w8465 = ~w16063 & ~w9760;
assign w8466 = ~w2341 & pi0837;
assign w8467 = ~w8701 & ~w16966;
assign w8468 = ~pi3287 & w14918;
assign w8469 = ~pi2972 & w16502;
assign w8470 = (pi0932 & ~w13509) | (pi0932 & w5850) | (~w13509 & w5850);
assign w8471 = ~w1664 & ~w4849;
assign w8472 = ~w6259 & ~w780;
assign w8473 = ~w621 & ~w8350;
assign w8474 = pi1410 & ~w5043;
assign w8475 = ~w2014 & w10758;
assign w8476 = ~pi0913 & w11739;
assign w8477 = ~w13970 & ~w17303;
assign w8478 = pi1863 & ~w15036;
assign w8479 = pi1765 & pi3155;
assign w8480 = ~w7888 & ~w5897;
assign w8481 = pi1337 & pi0252;
assign w8482 = ~pi1224 & ~w16679;
assign w8483 = pi2587 & ~w5274;
assign w8484 = ~w3203 & pi0906;
assign w8485 = pi2879 & ~w16815;
assign w8486 = ~w2994 & w18149;
assign w8487 = w10818 & ~w15440;
assign w8488 = ~w17321 & ~w44;
assign w8489 = ~pi0510 & ~pi1184;
assign w8490 = ~pi3096 & w11406;
assign w8491 = w7703 & w5497;
assign w8492 = ~w5540 & ~w13379;
assign w8493 = ~w5684 & ~w9182;
assign w8494 = w1962 & ~w15296;
assign w8495 = pi1936 & ~w18123;
assign w8496 = ~pi2232 & w2151;
assign w8497 = ~w2014 & w16050;
assign w8498 = ~w2014 & w16051;
assign w8499 = ~w366 & ~w12077;
assign w8500 = w3203 & ~w13028;
assign w8501 = pi1479 & w13753;
assign w8502 = pi1409 & ~w5043;
assign w8503 = ~w7077 & pi0808;
assign w8504 = pi1240 & ~w11655;
assign w8505 = w15122 & ~pi2598;
assign w8506 = ~w11702 & ~w7612;
assign w8507 = w934 & pi0430;
assign w8508 = w6611 & w8250;
assign w8509 = pi2752 & w14148;
assign w8510 = ~w16738 & ~w6151;
assign w8511 = pi2656 & ~w15235;
assign w8512 = ~w12101 & ~w8387;
assign w8513 = ~w16939 & pi0006;
assign w8514 = w1472 & w2157;
assign w8515 = ~w4020 & w15883;
assign w8516 = ~w2577 & ~w6798;
assign w8517 = ~pi2986 & ~w3067;
assign w8518 = ~w16278 & pi0714;
assign w8519 = ~pi0072 & w922;
assign w8520 = ~w8765 & ~w4998;
assign w8521 = ~w13655 & ~w2734;
assign w8522 = ~w6684 & ~w14790;
assign w8523 = w16575 & w16664;
assign w8524 = ~w4729 & ~w7446;
assign w8525 = w4067 & w3678;
assign w8526 = ~w16739 & ~w4280;
assign w8527 = ~pi3326 & w18259;
assign w8528 = w7434 & w8255;
assign w8529 = ~w11559 & ~w13608;
assign w8530 = ~pi0951 & w11739;
assign w8531 = w13231 & ~w2741;
assign w8532 = ~pi2851 & w14148;
assign w8533 = ~w3000 & ~pi2746;
assign w8534 = ~w18354 & ~w4788;
assign w8535 = ~pi3355 & w16922;
assign w8536 = ~w709 & pi1274;
assign w8537 = ~pi2975 & w17646;
assign w8538 = w13509 & w13706;
assign w8539 = pi3118 & ~pi3124;
assign w8540 = ~w2784 & ~w7976;
assign w8541 = ~w13790 & ~w3649;
assign w8542 = w13509 & w18203;
assign w8543 = pi1932 & ~w15271;
assign w8544 = (~pi0972 & ~w13509) | (~pi0972 & w7875) | (~w13509 & w7875);
assign w8545 = pi3165 & w3987;
assign w8546 = ~pi0631 & w14641;
assign w8547 = ~pi1296 & w62;
assign w8548 = w6697 & ~w2741;
assign w8549 = (pi1140 & ~w5437) | (pi1140 & w6500) | (~w5437 & w6500);
assign w8550 = ~pi0555 & w11739;
assign w8551 = pi1447 & ~w13753;
assign w8552 = ~pi2213 & w11313;
assign w8553 = ~w11211 & ~w16155;
assign w8554 = ~w4293 & ~w10785;
assign w8555 = ~w12409 & pi1202;
assign w8556 = w5453 & pi2582;
assign w8557 = w11743 & ~w11365;
assign w8558 = w1391 & ~w1236;
assign w8559 = ~w16506 & pi1193;
assign w8560 = w13509 & w5252;
assign w8561 = w6396 & w1485;
assign w8562 = w8949 & ~w13868;
assign w8563 = ~pi2034 & w7455;
assign w8564 = w13509 & w16643;
assign w8565 = pi1858 & ~pi0332;
assign w8566 = ~w7314 & ~w11273;
assign w8567 = w13509 & w14701;
assign w8568 = ~w2804 & ~pi2920;
assign w8569 = pi2977 & w8229;
assign w8570 = ~w13172 & ~w10396;
assign w8571 = pi2999 & pi3002;
assign w8572 = ~pi2234 & w2151;
assign w8573 = pi0031 & ~w3748;
assign w8574 = ~w6230 & ~w9107;
assign w8575 = pi3506 & w13367;
assign w8576 = ~w14648 & ~pi2710;
assign w8577 = ~w12040 & pi1086;
assign w8578 = pi2552 & w14148;
assign w8579 = ~pi1677 & pi3368;
assign w8580 = ~w15916 & ~w13601;
assign w8581 = ~w15613 & ~w7068;
assign w8582 = w11345 & w14350;
assign w8583 = ~w2725 & pi1089;
assign w8584 = pi1680 & pi1681;
assign w8585 = ~w2233 & ~w14952;
assign w8586 = ~w18282 & ~w156;
assign w8587 = pi1577 & w13753;
assign w8588 = ~w8539 & ~w16360;
assign w8589 = w14020 & w3464;
assign w8590 = ~w4425 & ~w2404;
assign w8591 = pi0046 & ~w14148;
assign w8592 = ~w6556 & ~w10605;
assign w8593 = ~w15808 & pi0745;
assign w8594 = w16575 & w15116;
assign w8595 = w2200 & w2708;
assign w8596 = ~w12995 & w1442;
assign w8597 = pi2321 & ~w4420;
assign w8598 = w13546 & w7010;
assign w8599 = w5874 & w11952;
assign w8600 = pi1391 & w13753;
assign w8601 = w14833 & w2753;
assign w8602 = w1962 & w11010;
assign w8603 = ~w8784 & ~w636;
assign w8604 = (pi1079 & ~w13509) | (pi1079 & w7106) | (~w13509 & w7106);
assign w8605 = w11247 & w5874;
assign w8606 = pi0206 & w9021;
assign w8607 = ~w16737 & ~w11420;
assign w8608 = ~w9605 & ~w5316;
assign w8609 = w9330 & w9792;
assign w8610 = w9440 & pi0159;
assign w8611 = ~w7856 & ~w12406;
assign w8612 = ~w12327 & ~w10869;
assign w8613 = ~pi3439 & w15036;
assign w8614 = w10647 & ~w16143;
assign w8615 = ~w709 & pi1288;
assign w8616 = ~pi1827 & ~w3567;
assign w8617 = w2425 & w17559;
assign w8618 = w10818 & ~w8044;
assign w8619 = ~pi3153 & w3805;
assign w8620 = (~w3771 & ~w9420) | (~w3771 & w16259) | (~w9420 & w16259);
assign w8621 = ~w13179 & ~w7821;
assign w8622 = (pi0833 & ~w13509) | (pi0833 & w629) | (~w13509 & w629);
assign w8623 = w384 & w14891;
assign w8624 = w17562 & pi2574;
assign w8625 = pi1500 & ~w16922;
assign w8626 = w5718 & w8918;
assign w8627 = ~w7844 & pi1062;
assign w8628 = ~w12460 & w12260;
assign w8629 = ~w6844 & ~w4218;
assign w8630 = pi2029 & ~w17646;
assign w8631 = ~w12572 & ~w11467;
assign w8632 = ~w6051 & ~w3342;
assign w8633 = ~w14648 & ~pi1974;
assign w8634 = w10189 & ~pi0453;
assign w8635 = w13509 & w7410;
assign w8636 = ~w9939 & ~w1780;
assign w8637 = ~pi0576 & w795;
assign w8638 = w4766 & w7212;
assign w8639 = ~pi3422 & w15036;
assign w8640 = w13509 & w15033;
assign w8641 = ~w10012 & ~w17328;
assign w8642 = pi1694 & ~pi1695;
assign w8643 = ~w2702 & w16826;
assign w8644 = w17248 & ~w15296;
assign w8645 = (~pi0269 & ~w325) | (~pi0269 & w10387) | (~w325 & w10387);
assign w8646 = ~w12992 & ~w12734;
assign w8647 = ~w7844 & pi0897;
assign w8648 = ~w8673 & ~w7124;
assign w8649 = w1962 & ~w6033;
assign w8650 = w8609 & w15060;
assign w8651 = ~w13969 & ~w6207;
assign w8652 = pi3158 & w10894;
assign w8653 = ~w8137 & ~w5005;
assign w8654 = pi2433 & ~w17646;
assign w8655 = pi0332 & w14001;
assign w8656 = ~w5892 & ~w12668;
assign w8657 = ~pi3165 & w11132;
assign w8658 = w9720 & w6447;
assign w8659 = w13509 & w1701;
assign w8660 = ~w17014 & w9090;
assign w8661 = w6002 & w17055;
assign w8662 = w11383 & w1570;
assign w8663 = w4835 & w7066;
assign w8664 = ~w11931 & ~w2619;
assign w8665 = w10647 & ~w6987;
assign w8666 = w13509 & w2028;
assign w8667 = ~w16278 & pi0936;
assign w8668 = ~w6195 & w15794;
assign w8669 = ~w1791 & w3256;
assign w8670 = (pi1115 & ~w13509) | (pi1115 & w11017) | (~w13509 & w11017);
assign w8671 = w10676 & w12227;
assign w8672 = ~pi3333 & w7090;
assign w8673 = ~w16575 & w6319;
assign w8674 = pi1793 & ~w9520;
assign w8675 = ~w16278 & pi0699;
assign w8676 = ~w8067 & w15450;
assign w8677 = w14228 & ~w15173;
assign w8678 = ~pi3053 & w261;
assign w8679 = pi1314 & pi1302;
assign w8680 = ~w12880 & ~w10478;
assign w8681 = w384 & w1768;
assign w8682 = w1962 & ~w10947;
assign w8683 = ~pi2459 & w13065;
assign w8684 = w16506 & ~w2587;
assign w8685 = ~w17890 & ~w16906;
assign w8686 = ~pi0835 & w93;
assign w8687 = ~w1151 & ~w13614;
assign w8688 = w7307 & w7037;
assign w8689 = pi1668 & ~pi3141;
assign w8690 = ~w7844 & pi0596;
assign w8691 = ~pi2975 & w9414;
assign w8692 = ~w251 & w12472;
assign w8693 = ~w3055 & w3693;
assign w8694 = ~w3055 & w3694;
assign w8695 = pi1282 & pi1345;
assign w8696 = (pi0784 & ~w13509) | (pi0784 & w16310) | (~w13509 & w16310);
assign w8697 = ~w8495 & ~w7554;
assign w8698 = pi2131 & ~w18123;
assign w8699 = ~w1962 & pi1011;
assign w8700 = pi1521 & w13753;
assign w8701 = pi1758 & ~w9520;
assign w8702 = ~w2690 & w16537;
assign w8703 = w9154 & w6760;
assign w8704 = (pi1137 & ~w5437) | (pi1137 & w14552) | (~w5437 & w14552);
assign w8705 = pi2496 & ~w5274;
assign w8706 = ~pi0948 & w1126;
assign w8707 = pi2114 & ~w412;
assign w8708 = (~pi1235 & ~w5437) | (~pi1235 & w14421) | (~w5437 & w14421);
assign w8709 = (w12775 & w9812) | (w12775 & w9367) | (w9812 & w9367);
assign w8710 = ~w6809 & ~w13668;
assign w8711 = w2725 & ~w3374;
assign w8712 = pi1423 & ~w6072;
assign w8713 = ~w13860 & ~w15623;
assign w8714 = ~w814 & ~w6946;
assign w8715 = (pi0618 & ~w13509) | (pi0618 & w17401) | (~w13509 & w17401);
assign w8716 = (~pi1802 & ~w7799) | (~pi1802 & w4302) | (~w7799 & w4302);
assign w8717 = pi1671 & w1924;
assign w8718 = w11247 & w17378;
assign w8719 = w4157 & w3711;
assign w8720 = ~pi3087 & w3555;
assign w8721 = ~pi2804 & w13343;
assign w8722 = ~w1586 & ~w17024;
assign w8723 = ~pi2908 & ~w14370;
assign w8724 = ~pi2639 & w15122;
assign w8725 = w7799 & w6691;
assign w8726 = ~w2530 & ~w14596;
assign w8727 = ~pi0635 & w3791;
assign w8728 = w7718 & w14994;
assign w8729 = ~w15560 & ~w4967;
assign w8730 = ~w14436 & ~w14086;
assign w8731 = ~w13355 & w3722;
assign w8732 = pi3164 & w653;
assign w8733 = w4667 & pi1259;
assign w8734 = ~pi3052 & w6463;
assign w8735 = ~pi0866 & w15707;
assign w8736 = ~w13231 & pi0566;
assign w8737 = ~pi3138 & w17993;
assign w8738 = (~pi0491 & w17577) | (~pi0491 & w13085) | (w17577 & w13085);
assign w8739 = (pi0845 & ~w13509) | (pi0845 & w13820) | (~w13509 & w13820);
assign w8740 = ~pi0292 & w4058;
assign w8741 = w5984 & w11151;
assign w8742 = ~w12798 & ~w17201;
assign w8743 = ~w10641 & ~w6619;
assign w8744 = w13509 & w10281;
assign w8745 = w369 & w300;
assign w8746 = w539 & ~w12823;
assign w8747 = w10680 & w5733;
assign w8748 = w2341 & ~w17513;
assign w8749 = w10818 & ~w10480;
assign w8750 = w13509 & w7485;
assign w8751 = w709 & pi1865;
assign w8752 = pi1933 & ~w11735;
assign w8753 = w13509 & w8649;
assign w8754 = ~w17071 & ~w6489;
assign w8755 = pi1547 & w13753;
assign w8756 = ~pi0980 & w6200;
assign w8757 = ~w2134 & w12401;
assign w8758 = ~w17121 & ~w1110;
assign w8759 = ~pi0630 & w14641;
assign w8760 = ~pi0780 & w543;
assign w8761 = w1144 & w2977;
assign w8762 = ~w1103 & ~w4359;
assign w8763 = w17117 & w8892;
assign w8764 = ~pi0782 & w543;
assign w8765 = ~w3969 & w3906;
assign w8766 = ~w5512 & w13417;
assign w8767 = ~pi3018 & w858;
assign w8768 = ~w11081 & ~w7043;
assign w8769 = ~pi1122 & w14641;
assign w8770 = (pi0830 & ~w13509) | (pi0830 & w2521) | (~w13509 & w2521);
assign w8771 = w13509 & w3545;
assign w8772 = w11015 & ~pi1312;
assign w8773 = pi1368 & w9653;
assign w8774 = w1368 & pi0398;
assign w8775 = ~w2805 & w2228;
assign w8776 = ~w10659 & ~w13719;
assign w8777 = ~pi2360 & w12755;
assign w8778 = ~w9444 & ~w17686;
assign w8779 = ~w17931 & ~w12378;
assign w8780 = ~w14228 & pi1112;
assign w8781 = pi1706 & ~w7946;
assign w8782 = (~pi0292 & ~w6857) | (~pi0292 & w11724) | (~w6857 & w11724);
assign w8783 = ~w9672 & ~w13665;
assign w8784 = w13509 & w4472;
assign w8785 = pi1738 & ~w4058;
assign w8786 = w10818 & ~w15355;
assign w8787 = ~w4318 & ~w8111;
assign w8788 = w17536 & w3987;
assign w8789 = ~pi1335 & ~pi2984;
assign w8790 = ~w10632 & w4947;
assign w8791 = ~w15336 & ~w8403;
assign w8792 = ~w10140 & ~w17815;
assign w8793 = ~w1418 & ~w16942;
assign w8794 = ~w14286 & w16947;
assign w8795 = ~w14626 & ~w15984;
assign w8796 = pi1624 & ~w6448;
assign w8797 = ~w14491 & ~w10531;
assign w8798 = w16138 & w17757;
assign w8799 = pi1597 & ~w13753;
assign w8800 = ~w12040 & pi1019;
assign w8801 = pi1220 & ~pi2969;
assign w8802 = pi1381 & ~w14918;
assign w8803 = ~pi2314 & w16041;
assign w8804 = w5437 & w16506;
assign w8805 = ~w2014 & w18361;
assign w8806 = ~w4075 & w13705;
assign w8807 = w384 & w17765;
assign w8808 = (~w5768 & ~w15717) | (~w5768 & w15274) | (~w15717 & w15274);
assign w8809 = ~w12624 & ~w17473;
assign w8810 = ~w11520 & ~w171;
assign w8811 = w13509 & w17766;
assign w8812 = pi1420 & ~w13753;
assign w8813 = pi1547 & ~w17935;
assign w8814 = ~w14003 & ~w8817;
assign w8815 = pi1668 & ~w2253;
assign w8816 = pi1149 & w9420;
assign w8817 = ~w12231 & w17358;
assign w8818 = ~w1391 & pi1039;
assign w8819 = ~pi1748 & w15122;
assign w8820 = pi1385 & w13753;
assign w8821 = ~w12084 & ~w14135;
assign w8822 = pi2523 & w16699;
assign w8823 = ~w9968 & ~w13906;
assign w8824 = pi2934 & ~w6045;
assign w8825 = w968 & ~pi0273;
assign w8826 = ~w15264 & ~w4891;
assign w8827 = ~w10350 & ~w15015;
assign w8828 = w1127 & ~w18357;
assign w8829 = w2531 & w11618;
assign w8830 = pi1425 & ~w6072;
assign w8831 = ~pi3089 & w16815;
assign w8832 = ~w5674 & ~w17919;
assign w8833 = ~w15979 & ~w10658;
assign w8834 = ~w11434 & w11504;
assign w8835 = ~pi1200 & w12825;
assign w8836 = ~w2665 & ~w2567;
assign w8837 = ~w1182 & ~w879;
assign w8838 = ~w2725 & pi1082;
assign w8839 = ~w8378 & ~w16526;
assign w8840 = pi2570 & ~w5274;
assign w8841 = w11383 & w9052;
assign w8842 = ~pi1166 & ~w13509;
assign w8843 = ~w14236 & ~w18080;
assign w8844 = pi1171 & ~w13509;
assign w8845 = pi2882 & ~w3555;
assign w8846 = ~w8895 & ~w18078;
assign w8847 = (~pi1765 & ~w7799) | (~pi1765 & w12621) | (~w7799 & w12621);
assign w8848 = pi1243 & ~pi1256;
assign w8849 = (~pi1804 & ~w7799) | (~pi1804 & w4583) | (~w7799 & w4583);
assign w8850 = w968 & ~pi0289;
assign w8851 = (pi0316 & w3055) | (pi0316 & w9890) | (w3055 & w9890);
assign w8852 = ~w16640 & ~w1538;
assign w8853 = ~pi0902 & w1147;
assign w8854 = w17248 & ~w2741;
assign w8855 = ~w15450 & ~w997;
assign w8856 = w2447 & w3956;
assign w8857 = ~w466 & ~w5654;
assign w8858 = ~pi2967 & pi3116;
assign w8859 = ~w17349 & ~pi0077;
assign w8860 = ~pi1229 & ~pi1242;
assign w8861 = ~w6697 & pi0943;
assign w8862 = ~w101 & ~w1626;
assign w8863 = ~w16575 & w7514;
assign w8864 = ~w8212 & ~w6082;
assign w8865 = w7136 & w6881;
assign w8866 = w3243 & w15659;
assign w8867 = ~w3567 & w4599;
assign w8868 = ~pi1752 & ~pi3157;
assign w8869 = ~w968 & w6857;
assign w8870 = pi2319 & ~w9414;
assign w8871 = ~w6785 & pi0989;
assign w8872 = ~w12146 & ~w13940;
assign w8873 = w7077 & w15609;
assign w8874 = pi1971 & ~w10539;
assign w8875 = w412 & w14078;
assign w8876 = ~pi2338 & w12941;
assign w8877 = pi1140 & ~w13564;
assign w8878 = (pi0372 & w6195) | (pi0372 & w9907) | (w6195 & w9907);
assign w8879 = pi1362 & ~w4256;
assign w8880 = pi1559 & ~w18259;
assign w8881 = (~pi0495 & w17577) | (~pi0495 & w11464) | (w17577 & w11464);
assign w8882 = ~w18407 & w6871;
assign w8883 = w8195 & w14382;
assign w8884 = pi2091 & ~w4420;
assign w8885 = ~pi1968 & w13729;
assign w8886 = ~w6697 & pi0663;
assign w8887 = w3168 & w2879;
assign w8888 = pi2937 & pi2969;
assign w8889 = w1391 & ~w14143;
assign w8890 = pi1255 & ~w11655;
assign w8891 = w15122 & ~pi2495;
assign w8892 = ~w12484 & ~w12315;
assign w8893 = ~pi3121 & pi3227;
assign w8894 = ~w18593 & ~w17585;
assign w8895 = ~pi3160 & ~pi3164;
assign w8896 = ~w7678 & ~w18196;
assign w8897 = ~pi3169 & w13570;
assign w8898 = ~w3947 & ~w9310;
assign w8899 = ~pi3155 & w3805;
assign w8900 = (~w13367 & w17577) | (~w13367 & w17343) | (w17577 & w17343);
assign w8901 = pi1235 & ~w2388;
assign w8902 = ~w1368 & ~pi0461;
assign w8903 = ~w1016 & ~w10271;
assign w8904 = ~w12917 & w9463;
assign w8905 = ~w2298 & ~w12075;
assign w8906 = pi1939 & ~w14833;
assign w8907 = ~pi3157 & w17669;
assign w8908 = pi3172 & w9520;
assign w8909 = ~w205 & ~w8681;
assign w8910 = ~w9010 & ~w690;
assign w8911 = pi1896 & ~w458;
assign w8912 = ~w13372 & ~w2954;
assign w8913 = ~pi2371 & w8617;
assign w8914 = ~pi0421 & w17173;
assign w8915 = ~w5627 & ~w11642;
assign w8916 = ~w15170 & w14721;
assign w8917 = ~pi2418 & w5075;
assign w8918 = ~w4466 & ~w13015;
assign w8919 = pi1612 & ~w7090;
assign w8920 = ~w8716 & w2275;
assign w8921 = w13509 & w9913;
assign w8922 = ~w15020 & ~w17798;
assign w8923 = w5189 & ~w6680;
assign w8924 = ~pi2174 & w11313;
assign w8925 = ~pi3171 & w15839;
assign w8926 = ~pi0944 & w3791;
assign w8927 = ~w7077 & pi0825;
assign w8928 = (w3987 & ~w4116) | (w3987 & w5176) | (~w4116 & w5176);
assign w8929 = ~w845 & ~w17061;
assign w8930 = w13509 & w14949;
assign w8931 = (w11743 & w11654) | (w11743 & w3264) | (w11654 & w3264);
assign w8932 = pi1720 & ~pi3172;
assign w8933 = ~pi0710 & w3106;
assign w8934 = (pi0841 & ~w13509) | (pi0841 & w5890) | (~w13509 & w5890);
assign w8935 = w14648 & ~pi2728;
assign w8936 = ~pi2275 & w3019;
assign w8937 = w13509 & w1425;
assign w8938 = w1465 & w7699;
assign w8939 = w16849 & w13541;
assign w8940 = ~w2491 & w12175;
assign w8941 = pi3166 & w6853;
assign w8942 = w7844 & ~w13028;
assign w8943 = ~pi3084 & w261;
assign w8944 = (~pi0958 & ~w13509) | (~pi0958 & w1926) | (~w13509 & w1926);
assign w8945 = pi3139 & w3987;
assign w8946 = ~pi0922 & w17899;
assign w8947 = w2770 & w8929;
assign w8948 = pi2557 & ~w5274;
assign w8949 = w7212 & ~w4766;
assign w8950 = w6697 & ~w10947;
assign w8951 = w13509 & w3487;
assign w8952 = w14648 & ~pi2289;
assign w8953 = ~w8254 & ~w9606;
assign w8954 = ~w2355 & w17830;
assign w8955 = ~w5065 & ~w1526;
assign w8956 = ~w12886 & ~w12363;
assign w8957 = pi1987 & ~w9414;
assign w8958 = ~pi1988 & w3019;
assign w8959 = ~w15371 & ~w9247;
assign w8960 = ~pi0135 & pi1878;
assign w8961 = w17954 & w11296;
assign w8962 = ~pi3340 & w18259;
assign w8963 = pi3170 & pi3207;
assign w8964 = ~pi0889 & w1126;
assign w8965 = pi2218 & ~w15271;
assign w8966 = pi1228 & pi3365;
assign w8967 = ~w17412 & ~w13938;
assign w8968 = ~pi3146 & w1843;
assign w8969 = ~w17447 & ~w16241;
assign w8970 = ~w10625 & ~w285;
assign w8971 = ~w3 & ~w2516;
assign w8972 = ~w2997 & ~w9427;
assign w8973 = ~w5650 & w15450;
assign w8974 = ~w17248 & pi1053;
assign w8975 = ~w15748 & ~w11563;
assign w8976 = pi2580 & ~w5274;
assign w8977 = w5189 & ~w2587;
assign w8978 = w6857 & w1012;
assign w8979 = pi1279 & pi1345;
assign w8980 = w13509 & w13007;
assign w8981 = ~w1515 & ~w13863;
assign w8982 = ~w1546 & ~w7251;
assign w8983 = ~w14250 & ~w17400;
assign w8984 = ~w12787 & ~w7372;
assign w8985 = ~w18581 & ~w1298;
assign w8986 = pi0104 & w3748;
assign w8987 = ~w2092 & ~w17865;
assign w8988 = w12081 & w1028;
assign w8989 = ~pi2249 & w12724;
assign w8990 = (~pi0334 & ~w6857) | (~pi0334 & w17431) | (~w6857 & w17431);
assign w8991 = ~w14228 & pi1127;
assign w8992 = w15465 & w9702;
assign w8993 = ~w12317 & ~w11805;
assign w8994 = ~w8822 & w1280;
assign w8995 = w8590 & w218;
assign w8996 = (~w1048 & ~w4903) | (~w1048 & w12522) | (~w4903 & w12522);
assign w8997 = (pi0578 & ~w13509) | (pi0578 & w5578) | (~w13509 & w5578);
assign w8998 = ~w5281 & ~w11192;
assign w8999 = ~pi3330 & w7090;
assign w9000 = pi1808 & ~w8829;
assign w9001 = ~w17822 & ~w11240;
assign w9002 = (pi1057 & ~w13509) | (pi1057 & w11821) | (~w13509 & w11821);
assign w9003 = ~pi0779 & w543;
assign w9004 = ~pi1098 & w17490;
assign w9005 = pi3172 & w5457;
assign w9006 = pi1756 & ~w17565;
assign w9007 = ~w12480 & ~w5429;
assign w9008 = ~w7170 & ~w7411;
assign w9009 = pi2816 & ~w11406;
assign w9010 = (pi0840 & ~w13509) | (pi0840 & w6547) | (~w13509 & w6547);
assign w9011 = pi2490 & ~w15235;
assign w9012 = ~w17410 & ~w8249;
assign w9013 = ~w14105 & ~w14403;
assign w9014 = w15122 & ~pi2627;
assign w9015 = ~w10154 & ~w16394;
assign w9016 = (pi0754 & ~w13509) | (pi0754 & w10044) | (~w13509 & w10044);
assign w9017 = ~pi3346 & w7090;
assign w9018 = w13509 & w16231;
assign w9019 = (pi0390 & w5560) | (pi0390 & w9035) | (w5560 & w9035);
assign w9020 = ~pi0296 & w2196;
assign w9021 = (~w12329 & w5855) | (~w12329 & w4693) | (w5855 & w4693);
assign w9022 = w7077 & ~w2776;
assign w9023 = w11383 & w9662;
assign w9024 = w7077 & ~w4179;
assign w9025 = (pi1068 & ~w13509) | (pi1068 & w670) | (~w13509 & w670);
assign w9026 = w13509 & w2604;
assign w9027 = w15169 & w15562;
assign w9028 = ~w13334 & ~w17743;
assign w9029 = w9243 & ~w10604;
assign w9030 = ~w16506 & pi1146;
assign w9031 = pi2607 & ~w261;
assign w9032 = ~pi0839 & w93;
assign w9033 = w15032 & w17614;
assign w9034 = ~w1368 & ~pi0467;
assign w9035 = w1368 & pi0390;
assign w9036 = ~w3000 & ~pi1890;
assign w9037 = w12460 & w6419;
assign w9038 = ~pi3170 & w17993;
assign w9039 = ~w9373 & w16710;
assign w9040 = w13509 & w15395;
assign w9041 = (~w5769 & ~w15717) | (~w5769 & w17407) | (~w15717 & w17407);
assign w9042 = pi2863 & w15191;
assign w9043 = w9788 & w5959;
assign w9044 = (pi0895 & ~w13509) | (pi0895 & w12429) | (~w13509 & w12429);
assign w9045 = pi1996 & ~w9414;
assign w9046 = w6785 & ~w3374;
assign w9047 = ~pi2488 & w15842;
assign w9048 = ~pi3353 & w16922;
assign w9049 = ~w4658 & ~w5899;
assign w9050 = ~pi0642 & w3791;
assign w9051 = pi3016 & ~w16502;
assign w9052 = w14648 & ~pi2616;
assign w9053 = w7799 & w2297;
assign w9054 = ~pi3049 & w9504;
assign w9055 = ~w1516 & w2912;
assign w9056 = (pi0857 & ~w13509) | (pi0857 & w326) | (~w13509 & w326);
assign w9057 = w7844 & ~w14978;
assign w9058 = ~pi2777 & w17213;
assign w9059 = ~pi3164 & w8515;
assign w9060 = w7703 & w4523;
assign w9061 = ~w13018 & ~w13488;
assign w9062 = w16575 & w1276;
assign w9063 = ~pi0509 & pi3363;
assign w9064 = ~w9751 & ~w12564;
assign w9065 = w934 & pi0425;
assign w9066 = pi1808 & ~w15537;
assign w9067 = w18262 & w6573;
assign w9068 = ~pi1778 & pi1332;
assign w9069 = pi3154 & w15767;
assign w9070 = pi1502 & ~w16922;
assign w9071 = pi0054 & ~w14148;
assign w9072 = (pi1071 & ~w13509) | (pi1071 & w6043) | (~w13509 & w6043);
assign w9073 = (~w10080 & ~w5517) | (~w10080 & w10066) | (~w5517 & w10066);
assign w9074 = w11668 & w14493;
assign w9075 = ~w6195 & w13081;
assign w9076 = w17562 & pi2563;
assign w9077 = pi1560 & ~w13753;
assign w9078 = w14161 & w18502;
assign w9079 = ~w12265 & ~w2885;
assign w9080 = ~pi3162 & w3982;
assign w9081 = ~w9693 & ~w4526;
assign w9082 = ~pi2244 & w17439;
assign w9083 = pi2552 & w605;
assign w9084 = pi0504 & pi0505;
assign w9085 = ~w12721 & ~w4172;
assign w9086 = ~w4671 & ~w5774;
assign w9087 = ~pi1839 & w12941;
assign w9088 = w5437 & w5089;
assign w9089 = ~w15431 & ~w5351;
assign w9090 = ~w1991 & ~w10556;
assign w9091 = pi2090 & ~w4420;
assign w9092 = w3345 & w5348;
assign w9093 = w3029 & w8324;
assign w9094 = pi0107 & w3748;
assign w9095 = ~pi0855 & w15707;
assign w9096 = w8040 & w8789;
assign w9097 = ~pi3286 & w16922;
assign w9098 = ~pi0120 & ~w8441;
assign w9099 = (pi0392 & w5560) | (pi0392 & w11599) | (w5560 & w11599);
assign w9100 = ~pi0841 & w93;
assign w9101 = pi1678 & ~w7177;
assign w9102 = ~w10428 & ~w3624;
assign w9103 = ~pi1802 & ~pi3135;
assign w9104 = ~w1962 & pi0651;
assign w9105 = w13509 & w15234;
assign w9106 = ~w2014 & w6190;
assign w9107 = pi2064 & ~w4508;
assign w9108 = w4599 & ~w16897;
assign w9109 = ~w7096 & ~w18184;
assign w9110 = w10087 & w10724;
assign w9111 = ~w3243 & pi0318;
assign w9112 = ~w9508 & ~w6771;
assign w9113 = ~w14560 & pi0243;
assign w9114 = pi2183 & ~w14524;
assign w9115 = ~w849 & ~w2631;
assign w9116 = pi0325 & w5274;
assign w9117 = ~pi1373 & ~w5144;
assign w9118 = ~pi3053 & w226;
assign w9119 = ~w7178 & ~w9797;
assign w9120 = ~w14228 & pi0899;
assign w9121 = ~w16707 & ~w15791;
assign w9122 = w16575 & w276;
assign w9123 = ~w11014 & ~w5863;
assign w9124 = ~w7431 & ~w13109;
assign w9125 = w13509 & w16140;
assign w9126 = ~pi3101 & w15235;
assign w9127 = ~w7077 & pi1044;
assign w9128 = ~w5189 & pi1100;
assign w9129 = ~pi0877 & pi0896;
assign w9130 = ~w14368 & w14163;
assign w9131 = pi2109 & ~w412;
assign w9132 = (~pi0322 & w3055) | (~pi0322 & w12431) | (w3055 & w12431);
assign w9133 = (pi0323 & w3055) | (pi0323 & w12432) | (w3055 & w12432);
assign w9134 = ~w5093 & ~w6698;
assign w9135 = w1978 & w10446;
assign w9136 = pi1358 & w14565;
assign w9137 = ~pi3052 & w16815;
assign w9138 = ~w6562 & ~w12635;
assign w9139 = ~w11214 & ~w6144;
assign w9140 = pi3153 & w10389;
assign w9141 = pi3160 & ~pi3488;
assign w9142 = ~pi2839 & w13343;
assign w9143 = pi1640 & ~w13753;
assign w9144 = ~pi3131 & w17387;
assign w9145 = ~w7657 & ~w17963;
assign w9146 = pi3113 & ~pi3150;
assign w9147 = ~w1058 & ~w577;
assign w9148 = ~w10627 & ~w3772;
assign w9149 = ~pi3107 & w6225;
assign w9150 = pi2121 & ~w412;
assign w9151 = ~w11200 & ~w9256;
assign w9152 = ~pi2460 & w13065;
assign w9153 = (~w13367 & w17577) | (~w13367 & w16332) | (w17577 & w16332);
assign w9154 = (w14269 & w16452) | (w14269 & w10575) | (w16452 & w10575);
assign w9155 = ~w9935 & ~w7122;
assign w9156 = pi2840 & w14148;
assign w9157 = w15808 & ~w14978;
assign w9158 = w8789 & w8888;
assign w9159 = pi1444 & ~w6448;
assign w9160 = pi2039 & ~w10158;
assign w9161 = ~w9289 & ~w3057;
assign w9162 = w550 & w6755;
assign w9163 = w13509 & w2808;
assign w9164 = ~w1640 & ~w9136;
assign w9165 = pi1984 & w7858;
assign w9166 = ~pi1983 & w7858;
assign w9167 = w13840 & pi1370;
assign w9168 = w539 & ~w12029;
assign w9169 = pi0483 & pi0493;
assign w9170 = w11345 & w10989;
assign w9171 = pi1355 & ~w11272;
assign w9172 = w11630 & w12273;
assign w9173 = ~w3054 & w9909;
assign w9174 = w2725 & ~w6647;
assign w9175 = ~w16331 & ~w8416;
assign w9176 = ~w9998 & w10807;
assign w9177 = pi2909 & ~w9687;
assign w9178 = ~w15221 & ~w5088;
assign w9179 = ~w744 & ~w8175;
assign w9180 = w12460 & w1533;
assign w9181 = pi1812 & ~w12558;
assign w9182 = ~pi2321 & w12724;
assign w9183 = ~w4893 & ~w9752;
assign w9184 = w6785 & ~w6647;
assign w9185 = ~w8181 & ~w5103;
assign w9186 = (pi0918 & ~w13509) | (pi0918 & w18113) | (~w13509 & w18113);
assign w9187 = w8658 & pi1809;
assign w9188 = ~pi2196 & w9340;
assign w9189 = w13509 & w13528;
assign w9190 = pi1556 & ~w18259;
assign w9191 = pi0018 & ~w14148;
assign w9192 = w7499 & w18584;
assign w9193 = ~pi1115 & w12197;
assign w9194 = pi1272 & pi1345;
assign w9195 = ~w13577 & ~w5905;
assign w9196 = w771 & ~w5531;
assign w9197 = pi1576 & w13753;
assign w9198 = ~pi2388 & w13204;
assign w9199 = (pi0837 & ~w13509) | (pi0837 & w8466) | (~w13509 & w8466);
assign w9200 = ~w5678 & ~w10005;
assign w9201 = pi1804 & ~w14951;
assign w9202 = (pi1043 & ~w13509) | (pi1043 & w4082) | (~w13509 & w4082);
assign w9203 = ~pi3153 & w13570;
assign w9204 = w10189 & ~pi0464;
assign w9205 = ~pi1778 & w8147;
assign w9206 = (pi0745 & ~w13509) | (pi0745 & w8593) | (~w13509 & w8593);
assign w9207 = w11735 & w14078;
assign w9208 = w10013 & w4320;
assign w9209 = pi0032 & ~w3748;
assign w9210 = ~w1894 & ~w8006;
assign w9211 = w62 & w15775;
assign w9212 = w5874 & w16033;
assign w9213 = ~w4346 & w7879;
assign w9214 = ~w12439 & ~w13873;
assign w9215 = w15842 & pi1341;
assign w9216 = (pi0501 & ~w11345) | (pi0501 & w5734) | (~w11345 & w5734);
assign w9217 = ~w9216 & ~w6843;
assign w9218 = ~w2725 & pi0790;
assign w9219 = ~w1408 & ~w14295;
assign w9220 = w2254 & w5058;
assign w9221 = ~w13810 & ~w11337;
assign w9222 = ~pi2882 & w15122;
assign w9223 = ~pi1004 & w14641;
assign w9224 = ~pi1251 & ~pi3237;
assign w9225 = ~w14560 & pi0231;
assign w9226 = pi3017 & w16502;
assign w9227 = w13569 & w6584;
assign w9228 = ~w5100 & ~w9481;
assign w9229 = pi1735 & w1924;
assign w9230 = ~pi0514 & ~pi1187;
assign w9231 = w12189 & w5550;
assign w9232 = ~pi0119 & w9284;
assign w9233 = pi2685 & ~w15235;
assign w9234 = ~w5526 & ~w181;
assign w9235 = pi2551 & w605;
assign w9236 = (pi0563 & ~w13509) | (pi0563 & w6743) | (~w13509 & w6743);
assign w9237 = w13509 & w15103;
assign w9238 = (pi0356 & w6195) | (pi0356 & w4006) | (w6195 & w4006);
assign w9239 = ~w4478 & ~pi0490;
assign w9240 = w14782 & w10364;
assign w9241 = ~w9540 & ~w10793;
assign w9242 = ~w2541 & ~w13803;
assign w9243 = ~w18563 & ~w13071;
assign w9244 = ~w2112 & ~w12129;
assign w9245 = ~pi0562 & w11739;
assign w9246 = ~w14311 & ~w13666;
assign w9247 = ~pi1059 & w93;
assign w9248 = pi3026 & ~w16502;
assign w9249 = (~w13367 & w17577) | (~w13367 & w3835) | (w17577 & w3835);
assign w9250 = ~pi3244 & ~pi3245;
assign w9251 = ~pi0769 & w6200;
assign w9252 = w10189 & pi0408;
assign w9253 = ~w8402 & ~w15629;
assign w9254 = w8970 & w11811;
assign w9255 = ~w8476 & ~w2843;
assign w9256 = ~pi0636 & w3791;
assign w9257 = ~w9633 & ~w17831;
assign w9258 = pi0491 & pi1138;
assign w9259 = ~pi0490 & ~pi1137;
assign w9260 = pi1478 & w13753;
assign w9261 = pi1788 & ~w6120;
assign w9262 = pi2042 & ~w10158;
assign w9263 = ~pi2419 & w13204;
assign w9264 = ~w6527 & w15101;
assign w9265 = ~w9991 & w7016;
assign w9266 = ~pi0311 & w13184;
assign w9267 = pi1476 & w13753;
assign w9268 = w11232 & ~w16279;
assign w9269 = w8337 & pi3294;
assign w9270 = ~w11796 & ~w12944;
assign w9271 = ~w11294 & ~w14720;
assign w9272 = w6824 & w11422;
assign w9273 = w2341 & ~w13195;
assign w9274 = ~w3055 & w357;
assign w9275 = pi2269 & ~w11671;
assign w9276 = ~w16369 & ~w3725;
assign w9277 = ~w16005 & ~w8683;
assign w9278 = ~w16278 & pi0709;
assign w9279 = ~w9224 & ~w2084;
assign w9280 = w7703 & w13909;
assign w9281 = ~w3124 & ~w2100;
assign w9282 = ~w3333 & ~pi0506;
assign w9283 = ~w17297 & ~w382;
assign w9284 = w236 & w12057;
assign w9285 = ~w5775 & ~w13774;
assign w9286 = ~pi2000 & w3019;
assign w9287 = ~pi2977 & ~w8229;
assign w9288 = w6785 & ~w1340;
assign w9289 = ~pi0814 & w1147;
assign w9290 = ~w6711 & ~w1015;
assign w9291 = ~w2352 & ~w1087;
assign w9292 = w1767 & w5565;
assign w9293 = pi1381 & w13753;
assign w9294 = w13509 & w14312;
assign w9295 = w16506 & ~w1236;
assign w9296 = w1368 & pi0407;
assign w9297 = ~w14481 & ~w7972;
assign w9298 = ~w4908 & ~w8400;
assign w9299 = pi1732 & ~w4058;
assign w9300 = (~w2913 & ~w1516) | (~w2913 & w1359) | (~w1516 & w1359);
assign w9301 = ~w3203 & pi0576;
assign w9302 = ~w18422 & w3416;
assign w9303 = w15450 & ~w6497;
assign w9304 = pi1587 & ~w16922;
assign w9305 = w9440 & pi0164;
assign w9306 = ~pi1929 & w9340;
assign w9307 = ~w14648 & ~pi2699;
assign w9308 = pi2270 & ~w17683;
assign w9309 = ~w12460 & w4657;
assign w9310 = pi1375 & ~w5043;
assign w9311 = pi1564 & ~w18259;
assign w9312 = ~w3466 & w10560;
assign w9313 = pi1989 & ~w9414;
assign w9314 = ~pi2411 & w7455;
assign w9315 = w6785 & ~w4179;
assign w9316 = ~w14349 & ~w9003;
assign w9317 = pi2712 & ~w261;
assign w9318 = ~w3827 & ~w14868;
assign w9319 = ~w6206 & ~w15855;
assign w9320 = w3509 & w2465;
assign w9321 = ~w3930 & w12358;
assign w9322 = ~w13576 & ~w4826;
assign w9323 = w4240 & ~w2238;
assign w9324 = pi3073 & ~w16502;
assign w9325 = pi2532 & w14148;
assign w9326 = ~w17637 & ~w18310;
assign w9327 = ~w14959 & ~w13151;
assign w9328 = w13509 & w17551;
assign w9329 = w9440 & pi0203;
assign w9330 = w9244 & w9281;
assign w9331 = w6857 & w6819;
assign w9332 = w735 & w657;
assign w9333 = ~w16103 & ~w15252;
assign w9334 = w12775 & ~w13219;
assign w9335 = ~w7242 & w12130;
assign w9336 = ~w7334 & w1389;
assign w9337 = pi1676 & ~w13203;
assign w9338 = pi0419 & w17173;
assign w9339 = w14833 & w17115;
assign w9340 = w5767 & w5410;
assign w9341 = ~w2841 & ~w18475;
assign w9342 = pi1577 & ~w14918;
assign w9343 = ~w6785 & pi0868;
assign w9344 = pi3105 & ~w16502;
assign w9345 = ~w5313 & ~w12334;
assign w9346 = ~pi0277 & w4058;
assign w9347 = pi3203 & ~w14054;
assign w9348 = (w13563 & ~w7807) | (w13563 & w2769) | (~w7807 & w2769);
assign w9349 = w14109 & pi0412;
assign w9350 = ~w3251 & ~w8941;
assign w9351 = (pi0658 & ~w13509) | (pi0658 & w12503) | (~w13509 & w12503);
assign w9352 = pi3043 & w16502;
assign w9353 = w1512 & w8380;
assign w9354 = ~pi0812 & w1147;
assign w9355 = (pi0566 & ~w13509) | (pi0566 & w8736) | (~w13509 & w8736);
assign w9356 = ~w12460 & w13092;
assign w9357 = pi2609 & ~w261;
assign w9358 = ~w13921 & ~w5263;
assign w9359 = ~pi0851 & w15707;
assign w9360 = w17706 & w3993;
assign w9361 = ~w14636 & ~w9995;
assign w9362 = ~w553 & pi1303;
assign w9363 = ~w10349 & ~w12954;
assign w9364 = ~w3427 & ~w566;
assign w9365 = pi2209 & ~w3223;
assign w9366 = ~w6141 & ~w2324;
assign w9367 = w131 & w12775;
assign w9368 = ~pi1955 & w11688;
assign w9369 = w16720 & w11196;
assign w9370 = w15808 & ~w6680;
assign w9371 = w13840 & pi1701;
assign w9372 = ~w6315 & ~w7598;
assign w9373 = (~pi1767 & ~w7799) | (~pi1767 & w12824) | (~w7799 & w12824);
assign w9374 = w10473 & w17084;
assign w9375 = pi2320 & ~w18123;
assign w9376 = ~w14684 & ~w17617;
assign w9377 = ~pi3101 & w3555;
assign w9378 = (pi0887 & ~w13509) | (pi0887 & w8072) | (~w13509 & w8072);
assign w9379 = ~w16329 & ~w14922;
assign w9380 = w14241 & w13671;
assign w9381 = (pi0813 & ~w13509) | (pi0813 & w11620) | (~w13509 & w11620);
assign w9382 = pi2958 & ~w13367;
assign w9383 = w384 & w1365;
assign w9384 = ~w1516 & ~w2555;
assign w9385 = pi2939 & w1326;
assign w9386 = ~w11862 & ~w13079;
assign w9387 = ~w1368 & ~pi0470;
assign w9388 = pi2506 & ~w5274;
assign w9389 = ~w159 & ~w17687;
assign w9390 = pi2396 & ~w10158;
assign w9391 = ~pi3160 & ~pi3161;
assign w9392 = ~w8851 & ~w16434;
assign w9393 = ~pi0989 & w15707;
assign w9394 = pi0506 & pi0512;
assign w9395 = ~pi3150 & w13730;
assign w9396 = w11793 & w4978;
assign w9397 = w13509 & w1965;
assign w9398 = ~w709 & pi1284;
assign w9399 = w15071 & w18021;
assign w9400 = ~w6147 & w1326;
assign w9401 = ~pi1916 & w9340;
assign w9402 = ~pi0515 & w17577;
assign w9403 = (pi1218 & ~w5437) | (pi1218 & w5181) | (~w5437 & w5181);
assign w9404 = ~w1918 & ~w7042;
assign w9405 = ~pi3052 & w9504;
assign w9406 = pi3134 & pi3142;
assign w9407 = ~pi3132 & ~w4020;
assign w9408 = pi0303 & w5113;
assign w9409 = ~w12460 & w3444;
assign w9410 = ~w6697 & pi0660;
assign w9411 = ~w173 & w5018;
assign w9412 = ~pi3160 & ~pi3172;
assign w9413 = pi1803 & pi3138;
assign w9414 = w14342 & w13605;
assign w9415 = pi3155 & w653;
assign w9416 = pi2263 & ~w11671;
assign w9417 = pi2746 & ~w6463;
assign w9418 = (w12436 & w12174) | (w12436 & w17885) | (w12174 & w17885);
assign w9419 = w5113 & w764;
assign w9420 = (w7212 & ~w8616) | (w7212 & w8638) | (~w8616 & w8638);
assign w9421 = ~w16142 & ~w5296;
assign w9422 = w18183 & w10673;
assign w9423 = ~w3203 & pi0586;
assign w9424 = ~w2027 & ~w1743;
assign w9425 = w9543 & pi0510;
assign w9426 = pi3160 & ~pi3501;
assign w9427 = ~pi3085 & w6463;
assign w9428 = ~pi3335 & w7090;
assign w9429 = ~w16730 & ~w13227;
assign w9430 = ~pi3353 & w14918;
assign w9431 = ~w13231 & pi0990;
assign w9432 = ~w3698 & ~w16694;
assign w9433 = w7844 & ~w16498;
assign w9434 = pi2051 & ~w10158;
assign w9435 = pi1802 & pi3135;
assign w9436 = w10103 & w11254;
assign w9437 = pi2290 & ~w9414;
assign w9438 = pi2687 & ~w11406;
assign w9439 = ~w13838 & ~w8475;
assign w9440 = ~w12975 & ~w17534;
assign w9441 = ~w8588 & w10158;
assign w9442 = ~pi3099 & w11406;
assign w9443 = ~w1736 & w14113;
assign w9444 = pi2637 & ~w3555;
assign w9445 = ~w1920 & w2446;
assign w9446 = w10189 & pi0386;
assign w9447 = ~w14508 & ~w14811;
assign w9448 = ~w13014 & ~w12309;
assign w9449 = ~pi3421 & w15036;
assign w9450 = pi2589 & ~w5274;
assign w9451 = pi1275 & pi1345;
assign w9452 = ~pi1305 & ~pi1266;
assign w9453 = ~w2341 & pi0898;
assign w9454 = ~w1042 & ~w14857;
assign w9455 = ~w6992 & ~w11304;
assign w9456 = pi1875 & ~w15036;
assign w9457 = ~w16603 & ~w3136;
assign w9458 = pi2030 & ~w17646;
assign w9459 = ~pi1776 & ~pi3147;
assign w9460 = w13509 & w1551;
assign w9461 = ~w6195 & w12325;
assign w9462 = w7324 & w17904;
assign w9463 = ~w14112 & ~w17271;
assign w9464 = (pi0685 & ~w13509) | (pi0685 & w18522) | (~w13509 & w18522);
assign w9465 = w1007 & w11567;
assign w9466 = pi2054 & ~w10158;
assign w9467 = w5517 & w2458;
assign w9468 = w11383 & w9586;
assign w9469 = w7844 & ~w3374;
assign w9470 = ~pi2455 & w5384;
assign w9471 = ~w2855 & ~w189;
assign w9472 = pi0262 & w5274;
assign w9473 = pi1361 & pi3020;
assign w9474 = pi2996 & ~pi3001;
assign w9475 = ~w1633 & w11489;
assign w9476 = w9394 & w4469;
assign w9477 = pi1623 & w13753;
assign w9478 = ~w11867 & ~w14168;
assign w9479 = pi2606 & ~w261;
assign w9480 = ~w15394 & ~w7418;
assign w9481 = ~pi2086 & w17439;
assign w9482 = ~pi3172 & w4310;
assign w9483 = ~w9543 & ~pi0510;
assign w9484 = ~w9955 & ~w15361;
assign w9485 = ~w16671 & ~w12085;
assign w9486 = w10302 & w8826;
assign w9487 = pi1448 & ~w6448;
assign w9488 = w525 & w6950;
assign w9489 = w13509 & w9288;
assign w9490 = ~w11502 & w17096;
assign w9491 = ~w12963 & ~w16639;
assign w9492 = w709 & pi1886;
assign w9493 = ~pi1178 & ~pi3219;
assign w9494 = (pi1017 & ~w13509) | (pi1017 & w10700) | (~w13509 & w10700);
assign w9495 = pi2236 & ~w11735;
assign w9496 = w12390 & w10328;
assign w9497 = ~w8874 & ~w16611;
assign w9498 = w1127 & ~w2241;
assign w9499 = ~w4598 & ~w13930;
assign w9500 = ~w13148 & w5557;
assign w9501 = ~w4680 & ~w14877;
assign w9502 = w11209 & ~w6966;
assign w9503 = pi1489 & ~w9781;
assign w9504 = pi2949 & w6641;
assign w9505 = ~w7077 & pi1042;
assign w9506 = pi2865 & w15191;
assign w9507 = pi0072 & ~w14148;
assign w9508 = (pi1050 & ~w13509) | (pi1050 & w12781) | (~w13509 & w12781);
assign w9509 = ~pi0550 & w3791;
assign w9510 = ~w13942 & w12452;
assign w9511 = ~w4772 & ~w9981;
assign w9512 = pi1523 & ~w14918;
assign w9513 = ~pi2113 & w12755;
assign w9514 = ~w10476 & ~w347;
assign w9515 = w17709 & w8783;
assign w9516 = w18506 & w1578;
assign w9517 = ~w6195 & w9113;
assign w9518 = ~w2150 & ~w12578;
assign w9519 = w8337 & pi3272;
assign w9520 = w2531 & w17016;
assign w9521 = ~w16087 & ~w13305;
assign w9522 = ~w11763 & ~w843;
assign w9523 = w14109 & pi0416;
assign w9524 = ~pi3145 & w14753;
assign w9525 = w14560 & pi0354;
assign w9526 = ~w13141 & ~w7463;
assign w9527 = pi3042 & pi3124;
assign w9528 = w6697 & ~w1340;
assign w9529 = ~pi1065 & w12825;
assign w9530 = ~pi0483 & pi3385;
assign w9531 = ~w3683 & ~w13222;
assign w9532 = ~w8849 & w14517;
assign w9533 = ~w4124 & w9647;
assign w9534 = ~pi0339 & ~w16205;
assign w9535 = pi2232 & ~w11735;
assign w9536 = w7703 & w3232;
assign w9537 = ~pi0983 & w3106;
assign w9538 = w2029 & w8030;
assign w9539 = pi1305 & pi1311;
assign w9540 = ~w1791 & w12159;
assign w9541 = ~pi2836 & w13343;
assign w9542 = ~w3762 & ~w4507;
assign w9543 = w4936 & w1639;
assign w9544 = ~pi3163 & w15048;
assign w9545 = pi2973 & w8569;
assign w9546 = w14648 & ~pi2831;
assign w9547 = w16575 & w1495;
assign w9548 = pi1797 & ~w5457;
assign w9549 = pi2608 & ~w261;
assign w9550 = (pi1213 & w5560) | (pi1213 & w2780) | (w5560 & w2780);
assign w9551 = ~w6697 & pi1015;
assign w9552 = ~w15499 & ~w414;
assign w9553 = w7703 & w7412;
assign w9554 = ~w8599 & w8207;
assign w9555 = w13231 & ~w1340;
assign w9556 = ~w1324 & ~w13016;
assign w9557 = pi2175 & ~w14524;
assign w9558 = pi3378 & w13367;
assign w9559 = ~w11746 & ~w5215;
assign w9560 = (pi0409 & w5560) | (pi0409 & w11894) | (w5560 & w11894);
assign w9561 = pi0896 & ~w4417;
assign w9562 = ~w1699 & ~w819;
assign w9563 = ~pi3089 & w15235;
assign w9564 = ~w12460 & w4204;
assign w9565 = w16596 & w10457;
assign w9566 = ~w8737 & ~w3729;
assign w9567 = w16893 & w14624;
assign w9568 = ~w9279 & w2273;
assign w9569 = ~w17959 & pi1337;
assign w9570 = ~pi1843 & w16041;
assign w9571 = w10406 & w13209;
assign w9572 = ~w13181 & ~w14747;
assign w9573 = w6857 & w6039;
assign w9574 = ~pi2920 & ~w16893;
assign w9575 = ~w7367 & w4438;
assign w9576 = ~w15792 & ~w14230;
assign w9577 = ~w6998 & ~w7983;
assign w9578 = ~w10539 & ~w7281;
assign w9579 = ~w11056 & ~w16078;
assign w9580 = (pi1084 & ~w13509) | (pi1084 & w17728) | (~w13509 & w17728);
assign w9581 = w13509 & w16052;
assign w9582 = ~w3068 & ~w14674;
assign w9583 = ~w3302 & ~w8597;
assign w9584 = (pi0652 & ~w13509) | (pi0652 & w13023) | (~w13509 & w13023);
assign w9585 = ~pi3018 & pi3102;
assign w9586 = w14648 & ~pi1688;
assign w9587 = ~w8119 & w8749;
assign w9588 = w13509 & w4878;
assign w9589 = ~w7019 & ~w5364;
assign w9590 = w3730 & w16107;
assign w9591 = ~pi1904 & w17213;
assign w9592 = w13509 & w18225;
assign w9593 = ~pi1163 & ~pi3180;
assign w9594 = w14482 & w10613;
assign w9595 = w539 & ~w11971;
assign w9596 = ~pi1750 & w7212;
assign w9597 = pi1905 & ~w11735;
assign w9598 = ~w11655 & w15292;
assign w9599 = pi3171 & w15767;
assign w9600 = w11716 & w4525;
assign w9601 = w16506 & w15609;
assign w9602 = ~w14040 & ~w8371;
assign w9603 = w5453 & pi2583;
assign w9604 = ~w12663 & ~w7173;
assign w9605 = ~pi3155 & w8515;
assign w9606 = pi2047 & ~w10158;
assign w9607 = ~w2014 & w16645;
assign w9608 = ~w1233 & ~w4784;
assign w9609 = pi1607 & ~w7090;
assign w9610 = ~w9660 & ~w9690;
assign w9611 = ~w5853 & ~w1227;
assign w9612 = ~pi3166 & w11701;
assign w9613 = ~w17485 & ~w16927;
assign w9614 = (pi0892 & ~w13509) | (pi0892 & w6108) | (~w13509 & w6108);
assign w9615 = ~w16575 & w6073;
assign w9616 = ~pi2816 & w13343;
assign w9617 = ~pi3288 & w7090;
assign w9618 = ~pi3172 & w15839;
assign w9619 = w2431 & ~w1875;
assign w9620 = pi2066 & ~w4508;
assign w9621 = ~w16145 & w16297;
assign w9622 = pi1337 & pi0305;
assign w9623 = pi3165 & w619;
assign w9624 = (pi0831 & ~w13509) | (pi0831 & w1860) | (~w13509 & w1860);
assign w9625 = w13509 & w497;
assign w9626 = w9720 & pi1714;
assign w9627 = ~w9152 & ~w12698;
assign w9628 = w13509 & w6808;
assign w9629 = w13509 & w10815;
assign w9630 = w13509 & w10816;
assign w9631 = ~w16577 & ~w2117;
assign w9632 = w18139 & w12835;
assign w9633 = w6857 & w15760;
assign w9634 = pi2180 & ~w14524;
assign w9635 = ~pi1124 & w1126;
assign w9636 = w16055 & ~w683;
assign w9637 = ~w11040 & w18520;
assign w9638 = ~w2814 & ~w4477;
assign w9639 = w15842 & pi1349;
assign w9640 = ~w9947 & ~w9258;
assign w9641 = ~w1414 & ~w14309;
assign w9642 = pi1769 & pi1807;
assign w9643 = ~w11299 & ~w17196;
assign w9644 = ~w1121 & ~w10434;
assign w9645 = ~w12192 & w8529;
assign w9646 = ~w16021 & w488;
assign w9647 = (~w4360 & ~w5517) | (~w4360 & w7768) | (~w5517 & w7768);
assign w9648 = ~pi2967 & pi3072;
assign w9649 = ~w14648 & ~pi2625;
assign w9650 = pi0499 & pi1183;
assign w9651 = ~w10130 & ~w10616;
assign w9652 = ~pi3160 & ~pi3165;
assign w9653 = w17741 & w5673;
assign w9654 = ~w13367 & w7513;
assign w9655 = ~pi3162 & w4310;
assign w9656 = pi3160 & w9473;
assign w9657 = ~w12426 & ~w5935;
assign w9658 = ~pi2173 & w11313;
assign w9659 = ~w11819 & ~w13450;
assign w9660 = pi2688 & ~w11406;
assign w9661 = pi1689 & ~w9504;
assign w9662 = w14648 & ~pi2295;
assign w9663 = ~w2014 & w17502;
assign w9664 = w934 & pi0420;
assign w9665 = ~w14073 & w12109;
assign w9666 = ~w11633 & w18436;
assign w9667 = (pi0404 & w5560) | (pi0404 & w15978) | (w5560 & w15978);
assign w9668 = ~w17114 & ~w11986;
assign w9669 = ~w1391 & pi0911;
assign w9670 = w13509 & w14399;
assign w9671 = w8928 & ~w5828;
assign w9672 = w11209 & ~w3707;
assign w9673 = ~pi3350 & w16922;
assign w9674 = pi3018 & ~pi3020;
assign w9675 = w5383 & ~w3432;
assign w9676 = w13509 & w6475;
assign w9677 = pi2850 & w605;
assign w9678 = ~pi3354 & w9781;
assign w9679 = ~w747 & ~w8752;
assign w9680 = ~pi0112 & w3748;
assign w9681 = w11696 & w2599;
assign w9682 = w13509 & w6302;
assign w9683 = (pi0791 & ~w13509) | (pi0791 & w13904) | (~w13509 & w13904);
assign w9684 = ~pi1260 & ~pi2969;
assign w9685 = ~w17315 & ~w8428;
assign w9686 = ~w6237 & ~w7329;
assign w9687 = ~pi2919 & ~pi2925;
assign w9688 = ~pi2708 & w15122;
assign w9689 = ~pi0974 & w6200;
assign w9690 = ~pi3059 & w11406;
assign w9691 = (pi0350 & w6195) | (pi0350 & w10157) | (w6195 & w10157);
assign w9692 = ~pi1153 & pi3194;
assign w9693 = ~pi3022 & ~pi3207;
assign w9694 = ~w4396 & w2221;
assign w9695 = ~pi2439 & w5075;
assign w9696 = ~w2403 & ~w13348;
assign w9697 = w10647 & ~w6042;
assign w9698 = ~pi3099 & w9504;
assign w9699 = ~w14125 & ~w1321;
assign w9700 = ~pi3187 & ~w12114;
assign w9701 = ~w2044 & ~w5130;
assign w9702 = ~w3308 & w4272;
assign w9703 = ~w6410 & ~w16772;
assign w9704 = w15041 & w2406;
assign w9705 = ~w4755 & ~w13006;
assign w9706 = w17562 & pi2506;
assign w9707 = pi1130 & ~pi1131;
assign w9708 = (pi0319 & w3055) | (pi0319 & w13990) | (w3055 & w13990);
assign w9709 = ~w3787 & ~w4223;
assign w9710 = pi3163 & w6853;
assign w9711 = w6857 & w1342;
assign w9712 = ~w6671 & ~w16085;
assign w9713 = ~w18406 & ~w2986;
assign w9714 = pi0444 & pi1827;
assign w9715 = pi2829 & ~w3555;
assign w9716 = ~w12460 & w977;
assign w9717 = ~pi0446 & w17173;
assign w9718 = ~w7880 & ~w5898;
assign w9719 = w5620 & w9078;
assign w9720 = ~pi3001 & w12689;
assign w9721 = ~w13620 & ~w9516;
assign w9722 = ~w4464 & ~w15592;
assign w9723 = (w12580 & ~w1206) | (w12580 & w15275) | (~w1206 & w15275);
assign w9724 = ~w6010 & w14873;
assign w9725 = ~w4384 & ~w7107;
assign w9726 = pi1217 & ~w4921;
assign w9727 = ~w5717 & ~w1941;
assign w9728 = w6857 & w15073;
assign w9729 = (pi0687 & ~w13509) | (pi0687 & w15947) | (~w13509 & w15947);
assign w9730 = w4229 & w16046;
assign w9731 = ~pi0927 & w3106;
assign w9732 = ~w7077 & pi0823;
assign w9733 = pi1337 & pi0268;
assign w9734 = ~pi1360 & w15842;
assign w9735 = ~w8881 & w3107;
assign w9736 = pi2151 & ~w11671;
assign w9737 = ~pi1877 & ~w15450;
assign w9738 = ~pi2401 & w5384;
assign w9739 = (pi0919 & ~w13509) | (pi0919 & w15164) | (~w13509 & w15164);
assign w9740 = pi0035 & ~w14148;
assign w9741 = ~w4751 & ~w18187;
assign w9742 = w2788 & w5596;
assign w9743 = ~w3208 & ~w8933;
assign w9744 = ~w8917 & ~w15835;
assign w9745 = pi2723 & ~w16815;
assign w9746 = w1516 & w15951;
assign w9747 = ~pi3242 & w18267;
assign w9748 = ~w1636 & ~w10491;
assign w9749 = ~pi3311 & w7090;
assign w9750 = ~w8551 & w8352;
assign w9751 = pi0044 & ~w14148;
assign w9752 = w13509 & w5272;
assign w9753 = ~pi3172 & w17993;
assign w9754 = ~pi3286 & w7090;
assign w9755 = ~w4440 & ~w17144;
assign w9756 = (pi0562 & ~w13509) | (pi0562 & w6032) | (~w13509 & w6032);
assign w9757 = ~w7748 & ~w10011;
assign w9758 = w9414 & w3515;
assign w9759 = ~pi3145 & w4310;
assign w9760 = ~pi3438 & w15036;
assign w9761 = w1127 & ~w13609;
assign w9762 = w2414 & w6145;
assign w9763 = ~w14228 & pi0628;
assign w9764 = w6857 & w18434;
assign w9765 = pi2402 & ~w10158;
assign w9766 = ~pi0331 & w2196;
assign w9767 = ~w5182 & ~w12947;
assign w9768 = ~pi3146 & w14753;
assign w9769 = ~w7855 & ~w3986;
assign w9770 = ~pi3350 & w6448;
assign w9771 = pi0509 & ~w17537;
assign w9772 = ~w8421 & ~w15218;
assign w9773 = ~w3156 & ~w4600;
assign w9774 = ~pi2346 & w12755;
assign w9775 = ~pi1994 & w3019;
assign w9776 = pi1968 & ~w7177;
assign w9777 = ~w11531 & ~w83;
assign w9778 = ~w1568 & ~w11113;
assign w9779 = ~pi0427 & w17173;
assign w9780 = w13509 & w6048;
assign w9781 = w1598 & w11747;
assign w9782 = ~pi0547 & w17899;
assign w9783 = pi2342 & ~w4420;
assign w9784 = w7177 & w14379;
assign w9785 = pi0310 & ~pi3218;
assign w9786 = w8163 & w3961;
assign w9787 = ~pi0963 & w543;
assign w9788 = w15075 & w5918;
assign w9789 = w11671 & w614;
assign w9790 = ~w8598 & ~w11546;
assign w9791 = pi2880 & ~w3555;
assign w9792 = w10825 & w1670;
assign w9793 = pi2426 & ~w10158;
assign w9794 = ~w15454 & w1184;
assign w9795 = ~w8172 & ~w15899;
assign w9796 = pi1614 & w13753;
assign w9797 = w13509 & w8190;
assign w9798 = ~w17561 & ~w8068;
assign w9799 = w11247 & w8599;
assign w9800 = ~w15968 & ~w6738;
assign w9801 = ~pi3139 & w14753;
assign w9802 = w13509 & w15135;
assign w9803 = ~pi3330 & w9781;
assign w9804 = w13509 & w2950;
assign w9805 = pi1435 & ~w6448;
assign w9806 = pi1736 & ~w4058;
assign w9807 = ~pi0692 & w9110;
assign w9808 = w13509 & w11575;
assign w9809 = ~pi0326 & ~w291;
assign w9810 = w17741 & w14434;
assign w9811 = ~w2979 & ~w15508;
assign w9812 = (w6228 & w8996) | (w6228 & w10255) | (w8996 & w10255);
assign w9813 = ~pi3326 & w14918;
assign w9814 = ~pi2149 & w13065;
assign w9815 = ~w15445 & ~w3093;
assign w9816 = ~w2710 & ~w15545;
assign w9817 = w9720 & pi1751;
assign w9818 = (pi0553 & ~w13509) | (pi0553 & w16490) | (~w13509 & w16490);
assign w9819 = pi2899 & ~w15235;
assign w9820 = ~pi3057 & ~pi3160;
assign w9821 = w3293 & w308;
assign w9822 = ~w3203 & pi1076;
assign w9823 = ~w14673 & ~w11078;
assign w9824 = (~pi0971 & ~w13509) | (~pi0971 & w331) | (~w13509 & w331);
assign w9825 = (pi0543 & ~w13509) | (pi0543 & w5815) | (~w13509 & w5815);
assign w9826 = ~w1880 & ~w17087;
assign w9827 = w13509 & w18284;
assign w9828 = ~pi2062 & w8617;
assign w9829 = w11209 & ~w9320;
assign w9830 = ~pi3156 & pi3249;
assign w9831 = ~pi0901 & w12825;
assign w9832 = ~pi1821 & w17562;
assign w9833 = w17248 & ~w11978;
assign w9834 = pi0118 & w9284;
assign w9835 = ~w12428 & ~w17309;
assign w9836 = (pi1027 & ~w13509) | (pi1027 & w11435) | (~w13509 & w11435);
assign w9837 = ~w13763 & ~pi0046;
assign w9838 = (pi0085 & ~w10335) | (pi0085 & w15250) | (~w10335 & w15250);
assign w9839 = w13509 & w5819;
assign w9840 = ~w3005 & ~w2680;
assign w9841 = w5437 & w7525;
assign w9842 = pi1588 & ~w9781;
assign w9843 = ~pi3099 & w15235;
assign w9844 = ~w17577 & w5015;
assign w9845 = ~w18148 & ~w16972;
assign w9846 = pi1772 & ~w5457;
assign w9847 = ~w7095 & ~w760;
assign w9848 = ~w3055 & w8866;
assign w9849 = (pi1063 & ~w13509) | (pi1063 & w10859) | (~w13509 & w10859);
assign w9850 = ~w16559 & ~w6136;
assign w9851 = ~w1962 & pi0550;
assign w9852 = ~w1503 & ~w18535;
assign w9853 = pi0248 & pi0260;
assign w9854 = ~w1554 & ~w630;
assign w9855 = w968 & ~pi0330;
assign w9856 = ~pi2391 & w16041;
assign w9857 = ~w13277 & ~w16626;
assign w9858 = (pi1113 & ~w13509) | (pi1113 & w11231) | (~w13509 & w11231);
assign w9859 = ~w2685 & ~w675;
assign w9860 = ~pi3023 & ~pi3207;
assign w9861 = ~w2450 & ~w7087;
assign w9862 = ~w13667 & ~w13114;
assign w9863 = ~w17665 & ~w4894;
assign w9864 = w15774 & w15992;
assign w9865 = ~pi3061 & w16815;
assign w9866 = ~w10343 & ~w3253;
assign w9867 = pi1705 & w4683;
assign w9868 = pi3166 & w4256;
assign w9869 = ~pi1829 & w11688;
assign w9870 = ~w15285 & ~w3898;
assign w9871 = pi2119 & ~w412;
assign w9872 = pi2179 & ~w11735;
assign w9873 = ~w10339 & ~w18232;
assign w9874 = ~w16270 & ~w13505;
assign w9875 = pi0302 & w5113;
assign w9876 = ~w13051 & ~w7386;
assign w9877 = ~pi3143 & pi3157;
assign w9878 = w272 & w1336;
assign w9879 = ~w11118 & ~w10376;
assign w9880 = ~w3763 & ~w1284;
assign w9881 = ~w6330 & ~w14090;
assign w9882 = ~w9545 & w1326;
assign w9883 = ~pi2892 & w15122;
assign w9884 = w4039 & w11798;
assign w9885 = w12040 & ~w6680;
assign w9886 = pi2641 & ~w3555;
assign w9887 = pi0307 & w18583;
assign w9888 = ~w9266 & ~w2862;
assign w9889 = ~w12108 & ~w15683;
assign w9890 = ~w3243 & pi0316;
assign w9891 = ~w7301 & w13352;
assign w9892 = ~w13683 & w9485;
assign w9893 = ~pi2182 & w5384;
assign w9894 = w11383 & w16133;
assign w9895 = ~pi0577 & w795;
assign w9896 = ~w17673 & w10481;
assign w9897 = ~w8367 & ~w4045;
assign w9898 = ~w7337 & ~w9789;
assign w9899 = pi2548 & w605;
assign w9900 = ~pi2043 & w13204;
assign w9901 = pi2710 & ~w16815;
assign w9902 = w8337 & pi3277;
assign w9903 = ~w8876 & ~w16343;
assign w9904 = pi2265 & ~w11671;
assign w9905 = w3255 & w5214;
assign w9906 = pi2374 & ~w3223;
assign w9907 = w14560 & pi0372;
assign w9908 = ~w3757 & ~w18201;
assign w9909 = w9720 & pi1719;
assign w9910 = ~w3039 & ~w14306;
assign w9911 = pi0062 & ~w14148;
assign w9912 = w10189 & ~pi0475;
assign w9913 = w6785 & ~w10947;
assign w9914 = ~pi0608 & w12825;
assign w9915 = pi2765 & w605;
assign w9916 = ~w1368 & ~pi0449;
assign w9917 = pi2694 & ~w16815;
assign w9918 = ~pi3101 & w11406;
assign w9919 = ~w7408 & ~w4737;
assign w9920 = pi1387 & ~w17935;
assign w9921 = ~w5174 & ~w4702;
assign w9922 = ~w12045 & ~w12523;
assign w9923 = ~pi1168 & pi3194;
assign w9924 = w16575 & w3423;
assign w9925 = ~pi0708 & w3106;
assign w9926 = ~w10766 & ~w13354;
assign w9927 = ~w6195 & w11091;
assign w9928 = ~pi2481 & w17213;
assign w9929 = ~pi3286 & w14918;
assign w9930 = w539 & ~w17197;
assign w9931 = pi0039 & ~w14148;
assign w9932 = w13509 & w2218;
assign w9933 = ~w14515 & ~w1541;
assign w9934 = ~pi2160 & w12755;
assign w9935 = pi0141 & ~pi0189;
assign w9936 = (pi1106 & ~w13509) | (pi1106 & w13656) | (~w13509 & w13656);
assign w9937 = ~w12025 & ~w16883;
assign w9938 = ~w4667 & ~w15974;
assign w9939 = pi1802 & ~w5457;
assign w9940 = pi0176 & w5274;
assign w9941 = w7698 & w18472;
assign w9942 = ~w14870 & ~w421;
assign w9943 = ~w12460 & w10529;
assign w9944 = w7703 & w1360;
assign w9945 = ~w1962 & pi0656;
assign w9946 = w2863 & w15626;
assign w9947 = pi0488 & pi1193;
assign w9948 = pi1846 & ~w12558;
assign w9949 = (w12719 & ~w11932) | (w12719 & w2424) | (~w11932 & w2424);
assign w9950 = ~w5189 & pi1102;
assign w9951 = ~w8795 & ~w7274;
assign w9952 = ~w5672 & ~w17406;
assign w9953 = ~w4452 & ~w8875;
assign w9954 = w659 & w18119;
assign w9955 = pi1471 & ~w7090;
assign w9956 = ~w3000 & ~pi2806;
assign w9957 = ~pi1410 & pi3240;
assign w9958 = w5189 & ~w4179;
assign w9959 = w3203 & ~w6680;
assign w9960 = ~pi1262 & w4880;
assign w9961 = ~pi2135 & w12941;
assign w9962 = pi1726 & ~w4058;
assign w9963 = pi2070 & ~w4508;
assign w9964 = w384 & w1122;
assign w9965 = pi2852 & w4140;
assign w9966 = ~w16218 & ~w6308;
assign w9967 = ~pi2058 & w13204;
assign w9968 = pi0172 & ~pi0192;
assign w9969 = pi1481 & ~w9781;
assign w9970 = ~pi1844 & ~w10299;
assign w9971 = w13509 & w2937;
assign w9972 = w13509 & w2938;
assign w9973 = ~pi3097 & w11406;
assign w9974 = ~pi2374 & w5075;
assign w9975 = ~w17248 & pi0882;
assign w9976 = ~pi2003 & w3019;
assign w9977 = ~pi3047 & w9504;
assign w9978 = w6697 & ~w14465;
assign w9979 = ~w4188 & ~w14802;
assign w9980 = ~w17577 & w10217;
assign w9981 = pi0337 & pi0338;
assign w9982 = ~w1962 & pi1117;
assign w9983 = ~w8184 & ~w10612;
assign w9984 = ~w13678 & ~w17792;
assign w9985 = ~w15510 & ~w6633;
assign w9986 = (pi0719 & ~w13509) | (pi0719 & w15509) | (~w13509 & w15509);
assign w9987 = ~pi3158 & w14753;
assign w9988 = w15450 & pi1163;
assign w9989 = ~w14129 & ~w7241;
assign w9990 = ~w16506 & pi1141;
assign w9991 = w5517 & w12983;
assign w9992 = (pi1085 & ~w13509) | (pi1085 & w15594) | (~w13509 & w15594);
assign w9993 = w1027 & ~w10631;
assign w9994 = ~pi1670 & w4667;
assign w9995 = ~w7807 & w961;
assign w9996 = pi2010 & ~w14833;
assign w9997 = ~pi3132 & ~pi3146;
assign w9998 = pi1507 & ~w13753;
assign w9999 = (~pi0282 & ~w6857) | (~pi0282 & w17397) | (~w6857 & w17397);
assign w10000 = ~pi1694 & ~pi1695;
assign w10001 = ~pi0740 & w17490;
assign w10002 = ~w3587 & ~w191;
assign w10003 = ~pi2817 & w17213;
assign w10004 = ~pi3000 & w16502;
assign w10005 = ~w8738 & w8900;
assign w10006 = ~pi3420 & w15036;
assign w10007 = ~w7478 & ~w3885;
assign w10008 = ~w10566 & ~w13738;
assign w10009 = ~w15450 & ~w5568;
assign w10010 = ~w5560 & w483;
assign w10011 = w13509 & w14144;
assign w10012 = pi0025 & ~w3748;
assign w10013 = w15474 & w7101;
assign w10014 = ~w16871 & ~w3863;
assign w10015 = w17581 & ~w5974;
assign w10016 = pi1752 & ~w8113;
assign w10017 = w15271 & w2753;
assign w10018 = ~pi2139 & w12941;
assign w10019 = w4137 & w7469;
assign w10020 = pi1242 & ~w11655;
assign w10021 = w13509 & w1163;
assign w10022 = ~pi3155 & w11132;
assign w10023 = ~w1821 & ~w16607;
assign w10024 = ~w15175 & ~w12442;
assign w10025 = ~pi1028 & w17899;
assign w10026 = pi2975 & ~w5855;
assign w10027 = pi2312 & ~w18123;
assign w10028 = ~pi3354 & w16922;
assign w10029 = ~pi3159 & w1843;
assign w10030 = ~w12254 & ~w16381;
assign w10031 = ~pi0492 & ~pi1139;
assign w10032 = (pi0948 & ~w13509) | (pi0948 & w1174) | (~w13509 & w1174);
assign w10033 = ~pi3347 & w6072;
assign w10034 = w934 & pi0439;
assign w10035 = ~w16506 & pi1183;
assign w10036 = ~w13068 & ~w13826;
assign w10037 = w9440 & pi0169;
assign w10038 = pi0261 & pi0268;
assign w10039 = ~pi0596 & w12825;
assign w10040 = w11077 & w3298;
assign w10041 = w13509 & w999;
assign w10042 = ~w12040 & ~pi0962;
assign w10043 = ~w16337 & ~w4591;
assign w10044 = ~w15808 & pi0754;
assign w10045 = ~pi2229 & w11313;
assign w10046 = pi1643 & ~w18259;
assign w10047 = ~pi3139 & w11701;
assign w10048 = ~w9173 & ~w13594;
assign w10049 = ~w5240 & ~w7551;
assign w10050 = ~w10923 & w11258;
assign w10051 = ~w12978 & ~w1873;
assign w10052 = pi3159 & w13786;
assign w10053 = w11247 & w918;
assign w10054 = (pi0663 & ~w13509) | (pi0663 & w8886) | (~w13509 & w8886);
assign w10055 = ~pi3155 & w17669;
assign w10056 = w384 & w9603;
assign w10057 = pi0896 & ~w2736;
assign w10058 = ~pi2980 & ~pi3109;
assign w10059 = pi1170 & ~w13509;
assign w10060 = ~w2699 & ~w10169;
assign w10061 = w4244 & w7564;
assign w10062 = ~w14588 & ~w9904;
assign w10063 = ~w13449 & ~w2089;
assign w10064 = ~w17090 & ~w9623;
assign w10065 = pi2272 & ~w17683;
assign w10066 = ~w1712 & ~w10080;
assign w10067 = ~w6726 & ~w15526;
assign w10068 = w14228 & ~w14978;
assign w10069 = w5589 & w17357;
assign w10070 = ~w13861 & w6078;
assign w10071 = ~w9019 & ~w12310;
assign w10072 = ~pi3163 & w11701;
assign w10073 = pi2254 & ~w15883;
assign w10074 = ~w16571 & ~w18426;
assign w10075 = ~w6326 & ~w13684;
assign w10076 = ~w5994 & ~w3999;
assign w10077 = w2460 & ~w7860;
assign w10078 = pi1382 & ~w17935;
assign w10079 = (pi1095 & ~w13509) | (pi1095 & w3929) | (~w13509 & w3929);
assign w10080 = ~pi0116 & w9284;
assign w10081 = pi0117 & w9284;
assign w10082 = ~w4670 & ~w1917;
assign w10083 = ~w5128 & ~w17182;
assign w10084 = ~w482 & ~w12250;
assign w10085 = ~pi2124 & w12755;
assign w10086 = pi2645 & ~w3555;
assign w10087 = ~w17666 & ~w1659;
assign w10088 = ~pi0965 & w93;
assign w10089 = ~w17019 & ~w10465;
assign w10090 = ~pi3343 & w14918;
assign w10091 = ~w9711 & w14534;
assign w10092 = ~w4575 & ~w7046;
assign w10093 = ~pi2052 & w13204;
assign w10094 = (pi0003 & ~w1766) | (pi0003 & w17990) | (~w1766 & w17990);
assign w10095 = pi0028 & ~w14148;
assign w10096 = ~w12040 & pi0692;
assign w10097 = pi1928 & ~w15271;
assign w10098 = ~w3491 & ~w15535;
assign w10099 = w7807 & w14738;
assign w10100 = ~pi2334 & w8617;
assign w10101 = w10818 & ~w1508;
assign w10102 = ~w17660 & ~w7474;
assign w10103 = w15749 & w12061;
assign w10104 = w13509 & w17526;
assign w10105 = ~w8087 & w4486;
assign w10106 = ~pi3293 & w9781;
assign w10107 = ~w16912 & ~w16326;
assign w10108 = w13509 & w12040;
assign w10109 = ~pi1828 & ~pi1984;
assign w10110 = ~pi0071 & ~pi0202;
assign w10111 = ~w11264 & ~w5894;
assign w10112 = ~w13724 & ~w15948;
assign w10113 = pi0261 & w5113;
assign w10114 = w16575 & w17627;
assign w10115 = w6649 & ~w4875;
assign w10116 = ~w2700 & ~w6581;
assign w10117 = w8626 & w2723;
assign w10118 = ~w4617 & ~w6750;
assign w10119 = ~w14228 & pi0633;
assign w10120 = w10189 & ~pi0456;
assign w10121 = ~pi2060 & w8617;
assign w10122 = pi3166 & w4324;
assign w10123 = w13509 & w8392;
assign w10124 = w13509 & w14799;
assign w10125 = w8928 & w12524;
assign w10126 = ~pi3314 & w9781;
assign w10127 = ~pi1305 & w14094;
assign w10128 = ~w15122 & ~pi2900;
assign w10129 = ~w17534 & pi0140;
assign w10130 = ~pi3163 & w3805;
assign w10131 = pi2719 & ~w9504;
assign w10132 = w6785 & ~w9852;
assign w10133 = w9440 & pi0196;
assign w10134 = pi3115 & ~pi3136;
assign w10135 = ~w3000 & ~pi2782;
assign w10136 = ~w5609 & ~w7929;
assign w10137 = ~w4274 & ~w14415;
assign w10138 = ~pi2966 & ~w1519;
assign w10139 = ~w8228 & ~w6876;
assign w10140 = w11345 & w891;
assign w10141 = pi3141 & w12558;
assign w10142 = w16278 & ~w16498;
assign w10143 = w6045 & ~w429;
assign w10144 = ~w14607 & ~w2812;
assign w10145 = ~pi3162 & w17669;
assign w10146 = ~w4556 & ~w8630;
assign w10147 = ~w255 & w3050;
assign w10148 = ~w11270 & ~w11658;
assign w10149 = w968 & ~pi0294;
assign w10150 = ~w7941 & ~w5030;
assign w10151 = w15122 & ~pi2597;
assign w10152 = pi3114 & ~w16502;
assign w10153 = ~w1647 & ~w14028;
assign w10154 = ~pi1133 & w9420;
assign w10155 = pi1134 & w9420;
assign w10156 = ~w15178 & ~w3937;
assign w10157 = w14560 & pi0350;
assign w10158 = w4841 & w3167;
assign w10159 = pi3160 & ~pi3480;
assign w10160 = (pi0582 & ~w13509) | (pi0582 & w16875) | (~w13509 & w16875);
assign w10161 = pi2365 & ~w15883;
assign w10162 = ~w12083 & ~w15040;
assign w10163 = ~w11614 & ~w12981;
assign w10164 = ~pi0809 & w1147;
assign w10165 = w9162 & w3227;
assign w10166 = pi0483 & pi0492;
assign w10167 = pi1666 & ~w4058;
assign w10168 = pi3160 & ~pi3490;
assign w10169 = ~w5560 & w16843;
assign w10170 = ~w3924 & ~w5501;
assign w10171 = w11077 & w6245;
assign w10172 = pi3146 & w8829;
assign w10173 = ~w11241 & ~w10797;
assign w10174 = pi3041 & ~w3987;
assign w10175 = w18123 & w14078;
assign w10176 = ~w14648 & ~pi2602;
assign w10177 = (~w18374 & ~w7807) | (~w18374 & w13954) | (~w7807 & w13954);
assign w10178 = ~w14407 & ~w583;
assign w10179 = ~w14473 & ~w12932;
assign w10180 = pi1334 & pi2966;
assign w10181 = w11766 & w17386;
assign w10182 = ~w5669 & ~w10773;
assign w10183 = w12436 & ~w3590;
assign w10184 = ~w13988 & ~w1212;
assign w10185 = w709 & pi2952;
assign w10186 = ~w9934 & ~w8118;
assign w10187 = ~pi3336 & w14918;
assign w10188 = ~pi3061 & w15235;
assign w10189 = w8789 & ~pi0896;
assign w10190 = ~w5189 & pi0718;
assign w10191 = (pi1121 & ~w13509) | (pi1121 & w3628) | (~w13509 & w3628);
assign w10192 = ~w6195 & w17146;
assign w10193 = ~w396 & ~w4532;
assign w10194 = ~w14648 & ~pi2879;
assign w10195 = ~pi1952 & w7455;
assign w10196 = ~w9230 & ~w10031;
assign w10197 = w15883 & w6320;
assign w10198 = ~pi0571 & w11739;
assign w10199 = ~w4077 & w10297;
assign w10200 = w16898 & w3945;
assign w10201 = ~w11484 & ~w11325;
assign w10202 = w11209 & ~w8148;
assign w10203 = w5437 & w10310;
assign w10204 = ~w17248 & pi0891;
assign w10205 = ~w13231 & pi0556;
assign w10206 = w8985 & w18528;
assign w10207 = w17562 & pi2566;
assign w10208 = ~pi0279 & w2196;
assign w10209 = ~w3570 & ~w868;
assign w10210 = ~w11933 & ~w9380;
assign w10211 = w7958 & w3977;
assign w10212 = (~pi0970 & ~w13509) | (~pi0970 & w7569) | (~w13509 & w7569);
assign w10213 = ~pi0259 & w5274;
assign w10214 = pi0260 & w5274;
assign w10215 = pi1514 & ~w14918;
assign w10216 = ~w13473 & ~w9354;
assign w10217 = w15146 & pi0513;
assign w10218 = w8789 & pi0477;
assign w10219 = w1308 & w2505;
assign w10220 = (pi0642 & ~w13509) | (pi0642 & w11394) | (~w13509 & w11394);
assign w10221 = ~w11775 & ~w16910;
assign w10222 = (~pi2920 & ~w384) | (~pi2920 & w111) | (~w384 & w111);
assign w10223 = w13509 & w11814;
assign w10224 = w11209 & ~w3249;
assign w10225 = ~w16210 & w3340;
assign w10226 = ~w16120 & ~w12565;
assign w10227 = ~pi0504 & ~pi1345;
assign w10228 = ~w16249 & ~w1974;
assign w10229 = ~w12852 & ~w12418;
assign w10230 = ~pi2313 & w12724;
assign w10231 = ~pi2381 & w12941;
assign w10232 = w14617 & w12164;
assign w10233 = ~pi0966 & w15707;
assign w10234 = ~w6780 & ~w9736;
assign w10235 = ~w5704 & ~w15939;
assign w10236 = ~w10138 & w13174;
assign w10237 = ~w3203 & pi0994;
assign w10238 = ~w15425 & w8855;
assign w10239 = w3020 & w784;
assign w10240 = pi2328 & ~w15883;
assign w10241 = ~w110 & ~w17905;
assign w10242 = ~w9965 & ~w5271;
assign w10243 = ~w8989 & ~w6648;
assign w10244 = pi1502 & ~w13753;
assign w10245 = ~pi3059 & w3555;
assign w10246 = ~w6071 & ~w9809;
assign w10247 = w3200 & w4686;
assign w10248 = ~pi1905 & w2151;
assign w10249 = pi2995 & w11232;
assign w10250 = (pi0927 & ~w13509) | (pi0927 & w5525) | (~w13509 & w5525);
assign w10251 = pi0087 & w9284;
assign w10252 = pi2782 & ~w6463;
assign w10253 = w8155 & w1528;
assign w10254 = pi2956 & ~pi3205;
assign w10255 = pi2969 & w6228;
assign w10256 = w15232 & w5192;
assign w10257 = pi1665 & ~w4058;
assign w10258 = pi2632 & ~w9504;
assign w10259 = w13509 & w350;
assign w10260 = ~pi3145 & w17993;
assign w10261 = (pi0133 & ~w10992) | (pi0133 & w1078) | (~w10992 & w1078);
assign w10262 = pi2954 & ~w6045;
assign w10263 = w11247 & w9212;
assign w10264 = w8337 & pi3304;
assign w10265 = ~pi0936 & w3106;
assign w10266 = (pi1056 & ~w13509) | (pi1056 & w15838) | (~w13509 & w15838);
assign w10267 = pi1635 & ~w6448;
assign w10268 = w5604 & w15529;
assign w10269 = pi1627 & ~w13753;
assign w10270 = ~w1391 & pi0771;
assign w10271 = (~pi0965 & ~w13509) | (~pi0965 & w2475) | (~w13509 & w2475);
assign w10272 = w7970 & w2313;
assign w10273 = w13177 & w18280;
assign w10274 = ~pi3139 & w12427;
assign w10275 = pi2363 & ~w18123;
assign w10276 = w3953 & w7743;
assign w10277 = pi2732 & ~w261;
assign w10278 = ~w17999 & w8339;
assign w10279 = (pi0858 & ~w13509) | (pi0858 & w17732) | (~w13509 & w17732);
assign w10280 = ~pi3290 & w14918;
assign w10281 = w16278 & ~w305;
assign w10282 = pi0501 & ~pi1147;
assign w10283 = w13509 & w3850;
assign w10284 = ~w13367 & w10447;
assign w10285 = ~w4155 & ~w18510;
assign w10286 = pi2541 & w605;
assign w10287 = pi2714 & ~w3555;
assign w10288 = ~w582 & ~w17069;
assign w10289 = ~w13183 & ~w10949;
assign w10290 = w5650 & ~pi1162;
assign w10291 = w17741 & w2047;
assign w10292 = pi1175 & ~w13509;
assign w10293 = w3132 & w9436;
assign w10294 = w17748 & w475;
assign w10295 = ~pi0587 & w795;
assign w10296 = pi1304 & w17477;
assign w10297 = ~pi3027 & ~w15276;
assign w10298 = pi1699 & ~w18497;
assign w10299 = pi1983 & w2247;
assign w10300 = (pi0744 & ~w13509) | (pi0744 & w11665) | (~w13509 & w11665);
assign w10301 = ~pi3158 & w1843;
assign w10302 = ~w2949 & ~w16748;
assign w10303 = w13231 & ~w4179;
assign w10304 = pi2617 & ~w261;
assign w10305 = ~w1562 & ~w11185;
assign w10306 = w1368 & pi0391;
assign w10307 = w7844 & ~w1340;
assign w10308 = (w8375 & ~w11247) | (w8375 & w8374) | (~w11247 & w8374);
assign w10309 = w8337 & pi3282;
assign w10310 = w16506 & ~w9852;
assign w10311 = ~w5453 & ~pi1776;
assign w10312 = ~w15225 & ~w16187;
assign w10313 = ~w17217 & ~w10999;
assign w10314 = ~w8789 & ~w4084;
assign w10315 = ~pi2339 & w17439;
assign w10316 = ~w13499 & ~w12383;
assign w10317 = ~pi2316 & w3019;
assign w10318 = ~w6564 & ~w12802;
assign w10319 = pi0505 & pi1192;
assign w10320 = ~pi3170 & w13730;
assign w10321 = ~w6195 & w13814;
assign w10322 = w11064 & w277;
assign w10323 = ~pi2400 & w17439;
assign w10324 = w7703 & w12350;
assign w10325 = ~pi1759 & ~pi3168;
assign w10326 = ~w14743 & ~w15926;
assign w10327 = ~w2276 & ~w6673;
assign w10328 = ~w3955 & ~w14561;
assign w10329 = w384 & w9706;
assign w10330 = ~w16842 & w16225;
assign w10331 = w7844 & ~w14143;
assign w10332 = pi1427 & ~w6072;
assign w10333 = ~w10368 & ~w5038;
assign w10334 = pi2202 & ~w10158;
assign w10335 = ~pi0452 & ~pi1687;
assign w10336 = pi1429 & ~w6072;
assign w10337 = ~w7702 & ~w199;
assign w10338 = ~w14678 & ~w796;
assign w10339 = pi3076 & ~pi3142;
assign w10340 = pi1604 & ~w9781;
assign w10341 = pi0039 & w922;
assign w10342 = (pi0601 & ~w13509) | (pi0601 & w905) | (~w13509 & w905);
assign w10343 = ~pi3138 & w13570;
assign w10344 = pi1683 & w18583;
assign w10345 = pi1563 & ~w18259;
assign w10346 = pi1903 & ~w226;
assign w10347 = w735 & pi1339;
assign w10348 = ~w1391 & pi0774;
assign w10349 = pi2516 & ~w16815;
assign w10350 = pi3008 & ~w3987;
assign w10351 = w15323 & w18152;
assign w10352 = w7799 & w735;
assign w10353 = pi3038 & ~w3987;
assign w10354 = ~w2733 & ~w15752;
assign w10355 = pi2551 & w14148;
assign w10356 = ~pi2402 & w13204;
assign w10357 = pi0036 & ~w3748;
assign w10358 = ~pi3330 & w16922;
assign w10359 = w4964 & w16228;
assign w10360 = ~w1158 & w4568;
assign w10361 = pi2563 & ~w5274;
assign w10362 = w11383 & w4298;
assign w10363 = w539 & ~w10853;
assign w10364 = w16836 & w9374;
assign w10365 = ~w13389 & ~w7531;
assign w10366 = ~w10548 & w11708;
assign w10367 = ~w3437 & ~w5698;
assign w10368 = pi1583 & ~w14918;
assign w10369 = pi2961 & ~w6617;
assign w10370 = ~w7523 & ~w14418;
assign w10371 = pi1921 & ~w15271;
assign w10372 = ~w3126 & ~w948;
assign w10373 = (pi0338 & w3055) | (pi0338 & w12011) | (w3055 & w12011);
assign w10374 = ~w8588 & w412;
assign w10375 = pi1590 & ~w16922;
assign w10376 = pi2219 & ~w11735;
assign w10377 = pi0120 & w10784;
assign w10378 = ~w10755 & ~w13931;
assign w10379 = w7703 & w8891;
assign w10380 = ~w2725 & pi0792;
assign w10381 = ~w709 & pi1294;
assign w10382 = ~w17612 & ~w17863;
assign w10383 = (pi0747 & ~w13509) | (pi0747 & w2471) | (~w13509 & w2471);
assign w10384 = ~w6499 & ~w4905;
assign w10385 = w7703 & w3292;
assign w10386 = ~w14648 & ~pi2626;
assign w10387 = pi1337 & ~pi0269;
assign w10388 = pi1776 & pi3147;
assign w10389 = w8658 & w4304;
assign w10390 = ~pi3050 & w6463;
assign w10391 = ~w16210 & ~w10609;
assign w10392 = ~w12040 & pi0684;
assign w10393 = w13509 & w1733;
assign w10394 = ~w2310 & ~w7057;
assign w10395 = ~w17408 & ~w13115;
assign w10396 = ~pi3088 & w3555;
assign w10397 = ~pi2988 & w16815;
assign w10398 = pi1480 & w13753;
assign w10399 = pi2041 & ~w10158;
assign w10400 = w17683 & w17115;
assign w10401 = ~pi2409 & w7455;
assign w10402 = pi1770 & ~w5457;
assign w10403 = ~pi3335 & w9781;
assign w10404 = ~w6963 & ~w9588;
assign w10405 = w9440 & pi0157;
assign w10406 = ~w7726 & ~w12155;
assign w10407 = w11209 & ~w5368;
assign w10408 = w16575 & w10782;
assign w10409 = pi0106 & w3748;
assign w10410 = (pi1167 & ~w13509) | (pi1167 & w11660) | (~w13509 & w11660);
assign w10411 = ~pi2549 & w5453;
assign w10412 = ~w3604 & ~w8563;
assign w10413 = w13509 & w12827;
assign w10414 = ~w17538 & ~w11180;
assign w10415 = ~w2341 & pi1064;
assign w10416 = w15118 & ~w2745;
assign w10417 = ~w12895 & ~w9615;
assign w10418 = ~pi2238 & w2151;
assign w10419 = ~w8056 & ~w18034;
assign w10420 = ~w14310 & ~w15589;
assign w10421 = ~w7791 & ~w916;
assign w10422 = ~pi3288 & w16922;
assign w10423 = pi0091 & w3748;
assign w10424 = pi1709 & w4683;
assign w10425 = ~pi2721 & w15122;
assign w10426 = w968 & ~pi0287;
assign w10427 = w13867 & w4333;
assign w10428 = pi3164 & ~w17800;
assign w10429 = w7396 & w2456;
assign w10430 = pi2522 & w4140;
assign w10431 = ~w9739 & ~w6204;
assign w10432 = ~pi2271 & w17439;
assign w10433 = w13509 & w12842;
assign w10434 = ~w6195 & w14246;
assign w10435 = ~pi3062 & w11406;
assign w10436 = w13231 & ~w2587;
assign w10437 = ~pi2433 & w7455;
assign w10438 = pi2382 & ~w18123;
assign w10439 = w6442 & w13561;
assign w10440 = ~pi1410 & w5043;
assign w10441 = ~w17481 & ~w5582;
assign w10442 = ~w7271 & ~w4206;
assign w10443 = ~w15314 & ~w5682;
assign w10444 = pi2128 & ~w18123;
assign w10445 = (pi0364 & w6195) | (pi0364 & w11072) | (w6195 & w11072);
assign w10446 = ~w14964 & ~w3366;
assign w10447 = (pi0496 & ~w5754) | (pi0496 & ~w17577) | (~w5754 & ~w17577);
assign w10448 = ~pi2771 & w13343;
assign w10449 = ~w4253 & ~w2284;
assign w10450 = ~w14725 & ~w15724;
assign w10451 = ~pi0771 & w6200;
assign w10452 = ~w2725 & pi0781;
assign w10453 = w13509 & w9273;
assign w10454 = ~w15256 & ~w12191;
assign w10455 = ~pi1367 & ~pi1407;
assign w10456 = ~w1368 & ~pi0481;
assign w10457 = ~w10295 & ~w665;
assign w10458 = (pi1212 & w5560) | (pi1212 & w6748) | (w5560 & w6748);
assign w10459 = ~w10244 & w5624;
assign w10460 = (pi1032 & ~w13509) | (pi1032 & w16430) | (~w13509 & w16430);
assign w10461 = pi1537 & w13753;
assign w10462 = ~pi0549 & w14641;
assign w10463 = pi0102 & w9284;
assign w10464 = w14560 & pi0368;
assign w10465 = w13509 & w4811;
assign w10466 = ~w9440 & ~w17160;
assign w10467 = ~w9665 & w4832;
assign w10468 = w13467 & w12127;
assign w10469 = pi2542 & w7965;
assign w10470 = w16506 & ~w10235;
assign w10471 = ~w2187 & ~w91;
assign w10472 = ~w4639 & ~w13881;
assign w10473 = pi0043 & pi0047;
assign w10474 = ~pi3150 & w11701;
assign w10475 = ~w2286 & ~w17095;
assign w10476 = pi3037 & ~pi3131;
assign w10477 = (pi1052 & ~w13509) | (pi1052 & w10909) | (~w13509 & w10909);
assign w10478 = (w8562 & w1682) | (w8562 & w3978) | (w1682 & w3978);
assign w10479 = ~w1791 & w1657;
assign w10480 = pi1581 & w13753;
assign w10481 = (pi1376 & ~w2235) | (pi1376 & w11512) | (~w2235 & w11512);
assign w10482 = ~w15010 & ~w481;
assign w10483 = pi2231 & ~w15271;
assign w10484 = ~pi2205 & w5075;
assign w10485 = w2341 & ~w11978;
assign w10486 = pi2720 & ~w16815;
assign w10487 = ~pi1991 & w11688;
assign w10488 = ~w16795 & ~w3736;
assign w10489 = ~pi3165 & w17993;
assign w10490 = ~pi0068 & ~w5642;
assign w10491 = ~w16438 & ~w16974;
assign w10492 = pi1456 & w13753;
assign w10493 = ~pi0514 & ~pi1345;
assign w10494 = w4653 & w3330;
assign w10495 = ~pi3343 & w16922;
assign w10496 = ~w11640 & ~w12737;
assign w10497 = w2341 & ~w12800;
assign w10498 = ~w11864 & w11516;
assign w10499 = pi1404 & ~w7946;
assign w10500 = ~w18391 & ~w5998;
assign w10501 = ~pi3157 & w11701;
assign w10502 = (pi0586 & ~w13509) | (pi0586 & w9423) | (~w13509 & w9423);
assign w10503 = pi0013 & ~w14148;
assign w10504 = ~w388 & ~w17826;
assign w10505 = (pi1176 & ~w13509) | (pi1176 & w4051) | (~w13509 & w4051);
assign w10506 = ~w12675 & ~w6376;
assign w10507 = ~w16366 & ~w5629;
assign w10508 = ~w12104 & ~w14156;
assign w10509 = ~w2203 & ~w6589;
assign w10510 = (pi0908 & ~w13509) | (pi0908 & w3155) | (~w13509 & w3155);
assign w10511 = ~pi3060 & w6463;
assign w10512 = ~w2014 & w13340;
assign w10513 = ~pi3340 & w17935;
assign w10514 = w13509 & w1996;
assign w10515 = ~w14228 & pi1126;
assign w10516 = ~w6375 & ~w8740;
assign w10517 = ~w3000 & ~pi2665;
assign w10518 = ~w15616 & ~w9176;
assign w10519 = ~w14204 & w17543;
assign w10520 = ~pi2736 & w15842;
assign w10521 = ~w14991 & w1744;
assign w10522 = w10647 & ~w14897;
assign w10523 = ~w16781 & ~w18008;
assign w10524 = pi2339 & ~w17683;
assign w10525 = ~w7578 & ~w10678;
assign w10526 = pi2869 & w14148;
assign w10527 = ~w13986 & ~w5140;
assign w10528 = ~pi0623 & w14641;
assign w10529 = w14109 & pi0427;
assign w10530 = ~pi2794 & w13343;
assign w10531 = w13509 & w8295;
assign w10532 = ~w6785 & pi0867;
assign w10533 = ~w16633 & ~w16708;
assign w10534 = ~w4261 & w15109;
assign w10535 = w5453 & pi2888;
assign w10536 = ~pi2604 & w15122;
assign w10537 = ~w12768 & ~w13383;
assign w10538 = ~w16278 & pi0703;
assign w10539 = ~pi2461 & w7399;
assign w10540 = ~w18104 & ~w11830;
assign w10541 = ~pi3138 & w13730;
assign w10542 = (~pi0329 & ~w6857) | (~pi0329 & w5367) | (~w6857 & w5367);
assign w10543 = ~pi2443 & w9340;
assign w10544 = ~w15449 & ~w3658;
assign w10545 = pi1446 & ~w6448;
assign w10546 = ~pi1843 & ~w18123;
assign w10547 = pi2438 & ~w10299;
assign w10548 = w7807 & w7248;
assign w10549 = w5189 & ~w6033;
assign w10550 = pi2146 & ~w11671;
assign w10551 = w9414 & w2753;
assign w10552 = w13868 & w9596;
assign w10553 = (pi0836 & ~w13509) | (pi0836 & w17319) | (~w13509 & w17319);
assign w10554 = ~w17278 & ~w2917;
assign w10555 = ~w14167 & ~w15318;
assign w10556 = w11383 & w13999;
assign w10557 = ~w7422 & w8620;
assign w10558 = w5517 & w8385;
assign w10559 = pi3153 & ~pi3159;
assign w10560 = w62 & ~w11689;
assign w10561 = ~w18249 & ~w2188;
assign w10562 = ~w13617 & ~w17154;
assign w10563 = (w8207 & ~w11247) | (w8207 & w9554) | (~w11247 & w9554);
assign w10564 = pi2004 & ~w9414;
assign w10565 = ~pi3048 & w9504;
assign w10566 = ~w1791 & w4565;
assign w10567 = ~pi0760 & w6200;
assign w10568 = w8814 & w15997;
assign w10569 = ~w7077 & pi0821;
assign w10570 = ~w10898 & ~w16272;
assign w10571 = ~w5687 & ~w17976;
assign w10572 = ~w6210 & w4315;
assign w10573 = ~w8027 & ~w18094;
assign w10574 = pi2995 & w5383;
assign w10575 = w14705 & w14269;
assign w10576 = ~w15140 & ~w14389;
assign w10577 = (pi0559 & ~w13509) | (pi0559 & w12219) | (~w13509 & w12219);
assign w10578 = w13509 & w4797;
assign w10579 = ~w3528 & ~w13518;
assign w10580 = pi1598 & ~w13753;
assign w10581 = (pi0922 & ~w13509) | (pi0922 & w5727) | (~w13509 & w5727);
assign w10582 = w384 & w15863;
assign w10583 = ~w11440 & ~w10975;
assign w10584 = ~pi1286 & pi1345;
assign w10585 = pi1287 & pi1345;
assign w10586 = (~w13367 & w17577) | (~w13367 & w1328) | (w17577 & w1328);
assign w10587 = ~pi3150 & w17387;
assign w10588 = w11652 & w3402;
assign w10589 = ~w14648 & ~pi2717;
assign w10590 = ~w18463 & w10417;
assign w10591 = ~w200 & ~w6840;
assign w10592 = w11033 & w17689;
assign w10593 = ~w17836 & ~w6236;
assign w10594 = ~pi2987 & w11406;
assign w10595 = ~w484 & ~w13367;
assign w10596 = ~w1962 & pi0637;
assign w10597 = pi0145 & pi0195;
assign w10598 = ~w18335 & ~w18235;
assign w10599 = w1368 & pi0408;
assign w10600 = (~w11215 & w5198) | (~w11215 & w18321) | (w5198 & w18321);
assign w10601 = pi3163 & ~w17313;
assign w10602 = w2561 & w4758;
assign w10603 = ~w6785 & pi0862;
assign w10604 = ~w12398 & ~w2294;
assign w10605 = w13509 & w14081;
assign w10606 = ~w3246 & ~w4152;
assign w10607 = ~w7622 & ~w7811;
assign w10608 = ~pi2521 & ~w1975;
assign w10609 = ~w4346 & ~w15026;
assign w10610 = ~w13367 & ~w11981;
assign w10611 = w6785 & w1217;
assign w10612 = w13509 & w8347;
assign w10613 = ~w16800 & ~w9553;
assign w10614 = ~w2277 & ~w10692;
assign w10615 = w5189 & ~w10235;
assign w10616 = pi1994 & ~w9414;
assign w10617 = ~w8739 & ~w1604;
assign w10618 = pi2292 & ~w9504;
assign w10619 = ~w8845 & ~w17509;
assign w10620 = ~pi1166 & ~pi3198;
assign w10621 = ~pi1925 & w11313;
assign w10622 = ~w8323 & w12490;
assign w10623 = ~w17665 & ~w15981;
assign w10624 = ~w16278 & ~pi0968;
assign w10625 = ~pi0696 & w9110;
assign w10626 = ~w8840 & ~w5594;
assign w10627 = w6857 & w4968;
assign w10628 = (pi1073 & ~w13509) | (pi1073 & w16146) | (~w13509 & w16146);
assign w10629 = ~w4092 & ~w6103;
assign w10630 = ~w5560 & w11989;
assign w10631 = pi1796 & ~w11388;
assign w10632 = w14782 & w16703;
assign w10633 = ~w16575 & w15647;
assign w10634 = ~w2090 & ~w6116;
assign w10635 = pi1983 & ~pi1985;
assign w10636 = ~w3383 & ~w11415;
assign w10637 = ~w14730 & ~w9377;
assign w10638 = ~w17248 & pi1124;
assign w10639 = w6649 & ~w9477;
assign w10640 = ~pi3138 & w3805;
assign w10641 = pi2436 & ~w15235;
assign w10642 = pi2972 & ~w17511;
assign w10643 = ~pi2520 & ~w1975;
assign w10644 = (pi0809 & ~w13509) | (pi0809 & w2852) | (~w13509 & w2852);
assign w10645 = pi1999 & ~w9414;
assign w10646 = ~w11502 & w1463;
assign w10647 = ~w8430 & w16095;
assign w10648 = w1962 & ~w9852;
assign w10649 = ~w1047 & ~w12591;
assign w10650 = ~w2847 & ~w8678;
assign w10651 = ~w18133 & ~w17192;
assign w10652 = w10189 & pi0400;
assign w10653 = ~w3235 & w14739;
assign w10654 = w11383 & w8232;
assign w10655 = pi0249 & w5113;
assign w10656 = pi2276 & ~w4420;
assign w10657 = w17248 & w1217;
assign w10658 = ~pi3087 & w16815;
assign w10659 = pi2711 & ~w16815;
assign w10660 = (w16442 & w12276) | (w16442 & w16808) | (w12276 & w16808);
assign w10661 = (pi1757 & w7215) | (pi1757 & w17423) | (w7215 & w17423);
assign w10662 = ~pi0483 & ~pi3397;
assign w10663 = ~pi0483 & pi3398;
assign w10664 = (pi0728 & ~w13509) | (pi0728 & w2448) | (~w13509 & w2448);
assign w10665 = ~w7162 & w17450;
assign w10666 = ~w12873 & ~w307;
assign w10667 = pi1361 & w4638;
assign w10668 = w3203 & ~w3430;
assign w10669 = pi0025 & ~w14148;
assign w10670 = w18262 & w16958;
assign w10671 = ~w15122 & ~pi1746;
assign w10672 = w13704 & w4026;
assign w10673 = ~pi1210 & ~w11335;
assign w10674 = ~pi3036 & ~w3987;
assign w10675 = ~pi3138 & w11701;
assign w10676 = ~pi2995 & w2363;
assign w10677 = pi0078 & ~pi3230;
assign w10678 = ~pi0103 & w9284;
assign w10679 = pi0104 & w9284;
assign w10680 = ~w18064 & ~w11797;
assign w10681 = w13509 & w12255;
assign w10682 = w15122 & ~pi2494;
assign w10683 = ~w16722 & ~w11090;
assign w10684 = w18123 & w9407;
assign w10685 = pi2536 & w14148;
assign w10686 = ~w17307 & ~w5298;
assign w10687 = pi1450 & ~w6448;
assign w10688 = ~w3595 & ~w16456;
assign w10689 = (pi2993 & ~w545) | (pi2993 & w12397) | (~w545 & w12397);
assign w10690 = ~w9848 & ~w1898;
assign w10691 = (pi0654 & ~w13509) | (pi0654 & w2191) | (~w13509 & w2191);
assign w10692 = w12460 & w8313;
assign w10693 = ~w2287 & ~w12132;
assign w10694 = ~pi2463 & w11606;
assign w10695 = ~w4154 & ~w14973;
assign w10696 = w13509 & w2023;
assign w10697 = ~pi3138 & w4310;
assign w10698 = ~w8785 & ~w4578;
assign w10699 = ~w16753 & ~w18017;
assign w10700 = ~w12040 & pi1017;
assign w10701 = pi2972 & ~pi3057;
assign w10702 = ~pi0569 & w11739;
assign w10703 = ~w9077 & w980;
assign w10704 = ~w10114 & ~w6612;
assign w10705 = ~w7844 & pi1000;
assign w10706 = ~w16746 & ~w10213;
assign w10707 = ~pi1198 & w3106;
assign w10708 = ~w2300 & ~w14713;
assign w10709 = w13509 & w1737;
assign w10710 = ~w3243 & pi0314;
assign w10711 = ~w17418 & ~w257;
assign w10712 = w16979 & w6445;
assign w10713 = ~w13997 & w9656;
assign w10714 = ~pi0659 & w12197;
assign w10715 = pi1422 & ~w13753;
assign w10716 = ~w11210 & ~w3574;
assign w10717 = w384 & w5416;
assign w10718 = w6940 & w2432;
assign w10719 = ~w14643 & ~w6482;
assign w10720 = ~w3318 & w3498;
assign w10721 = ~w8095 & ~w16183;
assign w10722 = pi1795 & ~w9520;
assign w10723 = w7307 & w3160;
assign w10724 = ~w10020 & ~w6261;
assign w10725 = (pi0371 & w6195) | (pi0371 & w7487) | (w6195 & w7487);
assign w10726 = w5408 & w6488;
assign w10727 = pi0502 & ~pi1378;
assign w10728 = ~w409 & ~w3799;
assign w10729 = ~pi2053 & w13204;
assign w10730 = ~w16506 & pi1157;
assign w10731 = ~w3733 & ~w6287;
assign w10732 = ~w4648 & ~w6973;
assign w10733 = w13509 & w16411;
assign w10734 = (~pi1759 & ~w7799) | (~pi1759 & w14355) | (~w7799 & w14355);
assign w10735 = w7307 & w7397;
assign w10736 = w13231 & ~w17210;
assign w10737 = ~pi1367 & ~pi2913;
assign w10738 = pi2161 & ~w11671;
assign w10739 = pi1466 & ~w7090;
assign w10740 = w13231 & ~w13195;
assign w10741 = ~w14228 & ~pi0957;
assign w10742 = ~pi1236 & ~w8966;
assign w10743 = pi2513 & ~w226;
assign w10744 = ~w17631 & w12569;
assign w10745 = ~w9543 & ~w13367;
assign w10746 = ~pi0663 & w12197;
assign w10747 = ~w17033 & ~w115;
assign w10748 = ~pi0575 & w795;
assign w10749 = (pi1059 & ~w13509) | (pi1059 & w12488) | (~w13509 & w12488);
assign w10750 = w7703 & w7967;
assign w10751 = ~w14215 & w4806;
assign w10752 = w7844 & ~w14597;
assign w10753 = (pi0696 & ~w13509) | (pi0696 & w5009) | (~w13509 & w5009);
assign w10754 = ~w12040 & ~pi0979;
assign w10755 = pi0064 & ~w14148;
assign w10756 = ~pi1771 & pi3150;
assign w10757 = pi2278 & ~w14524;
assign w10758 = ~w709 & pi1308;
assign w10759 = w13818 & w2380;
assign w10760 = w1531 & w7425;
assign w10761 = ~w3389 & ~w14937;
assign w10762 = ~w9658 & ~w12710;
assign w10763 = ~pi3044 & pi3172;
assign w10764 = ~pi3164 & w3805;
assign w10765 = ~w3054 & w17440;
assign w10766 = ~w4118 & w8618;
assign w10767 = w384 & w18320;
assign w10768 = ~w18272 & ~w5098;
assign w10769 = pi2446 & ~w14524;
assign w10770 = pi3160 & ~pi3372;
assign w10771 = ~w473 & w711;
assign w10772 = ~w5142 & w5921;
assign w10773 = ~pi2245 & w16041;
assign w10774 = w1303 & w4616;
assign w10775 = ~pi1043 & w1147;
assign w10776 = ~pi0286 & w4058;
assign w10777 = ~pi3055 & w15235;
assign w10778 = ~w13708 & w6382;
assign w10779 = (pi0691 & ~w13509) | (pi0691 & w2075) | (~w13509 & w2075);
assign w10780 = ~w10972 & w7452;
assign w10781 = ~w3021 & w11059;
assign w10782 = w10189 & ~pi0467;
assign w10783 = ~pi2975 & w412;
assign w10784 = ~w13312 & ~w8893;
assign w10785 = ~pi0764 & w6200;
assign w10786 = ~w190 & ~w13025;
assign w10787 = ~w10016 & ~w1275;
assign w10788 = ~w5560 & w11617;
assign w10789 = ~w11930 & ~w7994;
assign w10790 = w13509 & w3195;
assign w10791 = pi2158 & ~w16815;
assign w10792 = pi0510 & pi1184;
assign w10793 = ~pi2659 & w17213;
assign w10794 = ~pi1239 & ~pi3223;
assign w10795 = ~w7077 & pi0815;
assign w10796 = ~w12870 & ~w10895;
assign w10797 = pi2408 & ~w10158;
assign w10798 = ~pi3073 & pi3153;
assign w10799 = w14648 & ~pi2612;
assign w10800 = pi0198 & w5274;
assign w10801 = pi2995 & pi1402;
assign w10802 = w10243 & w9376;
assign w10803 = pi2658 & ~w15235;
assign w10804 = ~w14291 & ~w16423;
assign w10805 = ~w13500 & ~w7583;
assign w10806 = ~pi0641 & w3791;
assign w10807 = w1127 & ~w8755;
assign w10808 = ~w8907 & ~w7230;
assign w10809 = ~pi0972 & w17490;
assign w10810 = ~w397 & w722;
assign w10811 = ~w16367 & ~w6644;
assign w10812 = w10647 & ~w8501;
assign w10813 = ~pi1668 & pi3141;
assign w10814 = ~w7844 & pi0613;
assign w10815 = w2725 & ~w10235;
assign w10816 = w6697 & ~w7449;
assign w10817 = ~w13103 & ~w13442;
assign w10818 = w8430 & ~w16095;
assign w10819 = pi1414 & ~w6072;
assign w10820 = ~pi1254 & ~pi3232;
assign w10821 = pi1958 & ~w14833;
assign w10822 = w14109 & pi0431;
assign w10823 = w6797 & w15866;
assign w10824 = w12864 & w17978;
assign w10825 = ~w298 & ~w11395;
assign w10826 = ~pi3142 & w15839;
assign w10827 = ~pi3099 & w3555;
assign w10828 = w15808 & ~w14597;
assign w10829 = w709 & pi1885;
assign w10830 = w15122 & ~pi2932;
assign w10831 = pi1580 & w13753;
assign w10832 = ~w7077 & pi1074;
assign w10833 = ~pi1099 & w17899;
assign w10834 = w14560 & pi0346;
assign w10835 = pi1415 & ~w13753;
assign w10836 = ~w4407 & ~w6283;
assign w10837 = w14228 & ~w10235;
assign w10838 = pi3019 & w16502;
assign w10839 = ~pi3018 & w16502;
assign w10840 = pi2107 & ~w412;
assign w10841 = w9284 & ~pi0975;
assign w10842 = ~w10664 & ~w15763;
assign w10843 = ~w510 & w4965;
assign w10844 = ~pi3288 & w17935;
assign w10845 = ~w5189 & pi1104;
assign w10846 = pi1129 & w15450;
assign w10847 = (pi0856 & ~w13509) | (pi0856 & w11904) | (~w13509 & w11904);
assign w10848 = ~w2325 & ~w2125;
assign w10849 = pi2737 & ~w5274;
assign w10850 = ~pi3166 & w14753;
assign w10851 = ~w3433 & ~w6888;
assign w10852 = pi2503 & w7498;
assign w10853 = w1709 & w10316;
assign w10854 = ~w12976 & ~w13506;
assign w10855 = ~w11525 & ~w2383;
assign w10856 = ~w10734 & w4142;
assign w10857 = ~pi1901 & w13343;
assign w10858 = w15122 & ~pi2507;
assign w10859 = ~w2341 & pi1063;
assign w10860 = ~w11589 & ~w17216;
assign w10861 = pi1337 & pi0300;
assign w10862 = ~pi1971 & ~pi2461;
assign w10863 = (pi0621 & ~w13509) | (pi0621 & w3061) | (~w13509 & w3061);
assign w10864 = w11383 & w4105;
assign w10865 = ~pi0713 & w3106;
assign w10866 = ~pi0279 & w4058;
assign w10867 = ~w3209 & ~w2896;
assign w10868 = w8589 & w3565;
assign w10869 = w13509 & w17939;
assign w10870 = pi1172 & w13509;
assign w10871 = w16652 & w17744;
assign w10872 = (pi0879 & ~w13509) | (pi0879 & w3727) | (~w13509 & w3727);
assign w10873 = w13509 & w6318;
assign w10874 = ~pi1250 & ~pi3226;
assign w10875 = w13231 & ~w10235;
assign w10876 = w13509 & w580;
assign w10877 = ~pi3343 & w7090;
assign w10878 = w11010 & ~w2270;
assign w10879 = ~w15287 & ~w5761;
assign w10880 = ~pi3093 & w15235;
assign w10881 = w14648 & ~pi2706;
assign w10882 = ~pi0824 & w1147;
assign w10883 = ~w8812 & w12810;
assign w10884 = (~pi0505 & w17577) | (~pi0505 & w16505) | (w17577 & w16505);
assign w10885 = w13509 & w7146;
assign w10886 = ~w13884 & ~w1757;
assign w10887 = ~w13712 & w14974;
assign w10888 = ~w8085 & ~w5003;
assign w10889 = w13509 & w8923;
assign w10890 = w1391 & ~w16498;
assign w10891 = (pi0993 & ~w13509) | (pi0993 & w4555) | (~w13509 & w4555);
assign w10892 = w11383 & w8576;
assign w10893 = w9721 & w5094;
assign w10894 = w14216 & w2531;
assign w10895 = w13509 & w2614;
assign w10896 = ~w10670 & w3352;
assign w10897 = ~w8297 & ~w2962;
assign w10898 = pi2332 & ~w18123;
assign w10899 = ~pi0785 & w543;
assign w10900 = ~pi2141 & w12941;
assign w10901 = ~pi2087 & w17439;
assign w10902 = pi1516 & ~w14918;
assign w10903 = ~pi2031 & w7455;
assign w10904 = ~w17888 & ~w10931;
assign w10905 = ~w3000 & ~pi2808;
assign w10906 = ~pi3326 & w6072;
assign w10907 = ~w9044 & ~w5146;
assign w10908 = pi1558 & ~w18259;
assign w10909 = ~w15808 & pi1052;
assign w10910 = w4009 & ~w1595;
assign w10911 = ~pi0515 & ~pi1345;
assign w10912 = ~w15254 & ~w8414;
assign w10913 = ~w2725 & pi1077;
assign w10914 = w7799 & w7125;
assign w10915 = ~w6699 & w5047;
assign w10916 = ~w9201 & ~w8407;
assign w10917 = pi2329 & ~w9414;
assign w10918 = ~w11892 & ~w15464;
assign w10919 = (pi0727 & ~w13509) | (pi0727 & w15848) | (~w13509 & w15848);
assign w10920 = ~w17896 & ~w12926;
assign w10921 = ~w1206 & ~w383;
assign w10922 = pi3115 & ~w16502;
assign w10923 = w3546 & w13933;
assign w10924 = ~pi2820 & w17213;
assign w10925 = ~w3673 & ~w4706;
assign w10926 = ~w3203 & pi0583;
assign w10927 = ~w13231 & pi0557;
assign w10928 = ~w6767 & ~w14714;
assign w10929 = w384 & w8624;
assign w10930 = ~w14071 & ~w18194;
assign w10931 = ~pi0656 & w3791;
assign w10932 = pi2823 & ~w15235;
assign w10933 = ~w5175 & ~w16957;
assign w10934 = ~w5797 & ~w11227;
assign w10935 = ~w10868 & w4381;
assign w10936 = ~w11098 & w500;
assign w10937 = w13231 & w11302;
assign w10938 = ~w16278 & pi0546;
assign w10939 = pi1534 & ~w17935;
assign w10940 = ~pi3160 & ~pi3241;
assign w10941 = pi1924 & ~w14833;
assign w10942 = ~pi3172 & w17669;
assign w10943 = w8658 & pi1791;
assign w10944 = ~w11550 & w7003;
assign w10945 = pi0249 & w5274;
assign w10946 = ~w15500 & ~w10526;
assign w10947 = ~w8979 & ~w6935;
assign w10948 = ~w16602 & ~w6058;
assign w10949 = w13509 & w11669;
assign w10950 = ~w3203 & ~pi0953;
assign w10951 = (pi1808 & w7215) | (pi1808 & w8149) | (w7215 & w8149);
assign w10952 = ~w11259 & ~w4779;
assign w10953 = ~w2636 & ~w10067;
assign w10954 = ~w7844 & pi1069;
assign w10955 = ~pi1813 & ~w11388;
assign w10956 = ~w18544 & ~w15637;
assign w10957 = pi2132 & ~w18123;
assign w10958 = ~pi0767 & w6200;
assign w10959 = ~pi1676 & ~pi1698;
assign w10960 = ~w18079 & ~w2785;
assign w10961 = ~w709 & pi1275;
assign w10962 = ~pi3147 & w12427;
assign w10963 = ~pi2398 & w5075;
assign w10964 = pi1593 & ~w16922;
assign w10965 = ~w13469 & ~w8537;
assign w10966 = ~w9209 & ~w2110;
assign w10967 = ~pi1804 & pi3132;
assign w10968 = ~w4740 & ~w10321;
assign w10969 = w9743 & w12261;
assign w10970 = ~w12988 & ~w9824;
assign w10971 = ~w6397 & ~w14645;
assign w10972 = ~pi2960 & ~w15756;
assign w10973 = ~w7060 & w13546;
assign w10974 = ~w14400 & ~w4824;
assign w10975 = ~w13458 & w10586;
assign w10976 = ~w2014 & w8615;
assign w10977 = w13231 & ~w13028;
assign w10978 = ~pi3162 & w17387;
assign w10979 = ~w3512 & ~w6880;
assign w10980 = ~w7844 & pi0999;
assign w10981 = pi3020 & w3987;
assign w10982 = pi3139 & w18497;
assign w10983 = ~w6915 & ~w13596;
assign w10984 = pi0205 & pi1902;
assign w10985 = ~w11712 & w12091;
assign w10986 = ~w15404 & ~w14777;
assign w10987 = ~w14228 & pi0616;
assign w10988 = w1199 & w7056;
assign w10989 = ~pi0483 & pi3388;
assign w10990 = w255 & pi0272;
assign w10991 = ~pi3166 & w3982;
assign w10992 = w9227 & w9653;
assign w10993 = w7703 & w16449;
assign w10994 = w15271 & w3515;
assign w10995 = ~w7625 & ~w7796;
assign w10996 = pi1818 & ~w653;
assign w10997 = (pi0795 & ~w13509) | (pi0795 & w16265) | (~w13509 & w16265);
assign w10998 = (~w4455 & ~w5517) | (~w4455 & w403) | (~w5517 & w403);
assign w10999 = ~pi2082 & w17439;
assign w11000 = ~pi3298 & w17935;
assign w11001 = pi0149 & w5274;
assign w11002 = ~pi2364 & w5075;
assign w11003 = pi1700 & ~w18497;
assign w11004 = ~pi3142 & w3805;
assign w11005 = ~w12940 & ~w14145;
assign w11006 = ~w13682 & ~w2412;
assign w11007 = ~w726 & w8645;
assign w11008 = ~w547 & ~w15962;
assign w11009 = ~w14648 & ~pi2689;
assign w11010 = ~w18532 & w785;
assign w11011 = ~w11114 & ~w9784;
assign w11012 = ~w16197 & ~w18023;
assign w11013 = ~w6171 & ~w13165;
assign w11014 = w11209 & ~w8747;
assign w11015 = ~w9721 & w8598;
assign w11016 = ~pi1830 & ~w15271;
assign w11017 = ~w6697 & pi1115;
assign w11018 = ~pi0755 & w17490;
assign w11019 = ~w12414 & ~w10679;
assign w11020 = (pi0252 & ~w325) | (pi0252 & w8481) | (~w325 & w8481);
assign w11021 = pi1177 & ~w14073;
assign w11022 = ~w7462 & ~w4597;
assign w11023 = ~w12711 & ~w4183;
assign w11024 = ~w15938 & ~w17036;
assign w11025 = pi1740 & w1924;
assign w11026 = ~w17035 & ~w12341;
assign w11027 = ~w5642 & ~w7843;
assign w11028 = w10647 & ~w5558;
assign w11029 = w17179 & w11349;
assign w11030 = w13509 & w1740;
assign w11031 = ~w4264 & ~w13164;
assign w11032 = ~pi3084 & w16815;
assign w11033 = ~w18092 & ~w11015;
assign w11034 = ~w3567 & w8949;
assign w11035 = w13509 & w6672;
assign w11036 = pi1434 & ~w13753;
assign w11037 = ~w1826 & ~w7560;
assign w11038 = ~pi2143 & w12941;
assign w11039 = ~pi2830 & w14325;
assign w11040 = pi1215 & w5566;
assign w11041 = ~w10025 & ~w1169;
assign w11042 = w1127 & ~w15442;
assign w11043 = ~pi3124 & ~pi3160;
assign w11044 = ~w5136 & ~w7131;
assign w11045 = (pi1047 & ~w13509) | (pi1047 & w15332) | (~w13509 & w15332);
assign w11046 = ~w8409 & w3806;
assign w11047 = ~w16506 & pi1136;
assign w11048 = w9440 & pi0189;
assign w11049 = ~w4408 & ~w3212;
assign w11050 = pi2344 & ~w18123;
assign w11051 = w6785 & ~w14597;
assign w11052 = ~w15822 & ~w13134;
assign w11053 = ~w12460 & w13349;
assign w11054 = ~pi1926 & w9340;
assign w11055 = pi2700 & ~w9504;
assign w11056 = (w14403 & ~w14705) | (w14403 & w2973) | (~w14705 & w2973);
assign w11057 = ~w1791 & w11430;
assign w11058 = ~w3203 & pi0907;
assign w11059 = w6981 & w2380;
assign w11060 = w13840 & w17562;
assign w11061 = ~w4719 & ~w11377;
assign w11062 = (w6928 & ~w17173) | (w6928 & w14847) | (~w17173 & w14847);
assign w11063 = w13509 & w10485;
assign w11064 = ~w11648 & ~w15577;
assign w11065 = ~w7844 & pi0607;
assign w11066 = ~w16278 & pi0929;
assign w11067 = w709 & pi1874;
assign w11068 = ~w7220 & w5148;
assign w11069 = ~pi3135 & ~pi3160;
assign w11070 = pi0247 & pi0255;
assign w11071 = ~pi1003 & w12825;
assign w11072 = w14560 & pi0364;
assign w11073 = ~w254 & ~w6848;
assign w11074 = ~w143 & w13764;
assign w11075 = pi1445 & ~w6448;
assign w11076 = w13509 & w13059;
assign w11077 = ~w16055 & w10058;
assign w11078 = ~w12985 & w17414;
assign w11079 = ~w4208 & ~w9163;
assign w11080 = w13509 & w13398;
assign w11081 = ~pi1924 & w11688;
assign w11082 = ~w5947 & ~w18186;
assign w11083 = ~pi2215 & w11313;
assign w11084 = ~pi2146 & w13065;
assign w11085 = pi2330 & ~w17646;
assign w11086 = w9440 & pi0201;
assign w11087 = pi2568 & ~w5274;
assign w11088 = ~pi0624 & w14641;
assign w11089 = (pi0742 & ~w13509) | (pi0742 & w17861) | (~w13509 & w17861);
assign w11090 = ~pi3316 & w17935;
assign w11091 = ~w14560 & pi0244;
assign w11092 = ~w17675 & ~w13532;
assign w11093 = w17577 & ~w17370;
assign w11094 = pi2123 & ~w15271;
assign w11095 = ~pi0110 & w3748;
assign w11096 = w10818 & ~w5327;
assign w11097 = ~w8364 & ~w2865;
assign w11098 = pi1770 & pi3172;
assign w11099 = ~pi3097 & w15235;
assign w11100 = ~pi2426 & w13204;
assign w11101 = ~pi0828 & w93;
assign w11102 = ~w5399 & ~w1685;
assign w11103 = ~w1594 & ~w6778;
assign w11104 = w6857 & w15133;
assign w11105 = w6785 & ~w11978;
assign w11106 = w3864 & w7662;
assign w11107 = ~w8715 & ~w3517;
assign w11108 = w13509 & w4130;
assign w11109 = w5437 & w13894;
assign w11110 = pi2706 & ~w261;
assign w11111 = (pi0710 & ~w13509) | (pi0710 & w6609) | (~w13509 & w6609);
assign w11112 = w12460 & w13661;
assign w11113 = pi1952 & ~w17646;
assign w11114 = pi1679 & ~w7177;
assign w11115 = w539 & ~w13747;
assign w11116 = pi0109 & ~w2632;
assign w11117 = ~pi3349 & w7090;
assign w11118 = ~pi3163 & w17387;
assign w11119 = ~pi1128 & pi1130;
assign w11120 = (~w5967 & ~w5517) | (~w5967 & w11226) | (~w5517 & w11226);
assign w11121 = ~w18462 & w8321;
assign w11122 = w3194 & w16823;
assign w11123 = w2725 & ~w10947;
assign w11124 = w6697 & ~w14143;
assign w11125 = ~w1269 & ~w16201;
assign w11126 = ~w1143 & ~w336;
assign w11127 = pi1977 & ~w6463;
assign w11128 = ~w16402 & ~w12282;
assign w11129 = ~w3054 & w7553;
assign w11130 = ~w15514 & ~w18507;
assign w11131 = ~w2725 & pi1190;
assign w11132 = ~w4020 & w4420;
assign w11133 = ~pi0620 & w14641;
assign w11134 = pi1509 & ~w16922;
assign w11135 = w6649 & ~w12396;
assign w11136 = ~w15711 & ~w9872;
assign w11137 = pi1793 & ~w15297;
assign w11138 = w7703 & w378;
assign w11139 = ~w4145 & w8909;
assign w11140 = pi1394 & ~w17935;
assign w11141 = ~w15808 & pi0924;
assign w11142 = ~w6849 & ~w3732;
assign w11143 = (pi0655 & ~w13509) | (pi0655 & w6065) | (~w13509 & w6065);
assign w11144 = ~w12952 & ~w4679;
assign w11145 = ~w17480 & ~w9698;
assign w11146 = ~pi0971 & w17490;
assign w11147 = pi1777 & pi3134;
assign w11148 = w9440 & pi0162;
assign w11149 = w13509 & w4884;
assign w11150 = ~w458 & w14773;
assign w11151 = ~w18202 & ~w3291;
assign w11152 = ~w6826 & w5334;
assign w11153 = ~w3000 & ~pi2667;
assign w11154 = w7703 & w16166;
assign w11155 = ~w7077 & pi1072;
assign w11156 = ~w5563 & ~w13507;
assign w11157 = ~w1691 & ~w10564;
assign w11158 = pi2530 & w14148;
assign w11159 = ~pi1219 & w9284;
assign w11160 = pi3081 & ~w16502;
assign w11161 = pi0515 & pi0503;
assign w11162 = ~w12120 & ~w5242;
assign w11163 = (pi1180 & w5560) | (pi1180 & w7302) | (w5560 & w7302);
assign w11164 = w7703 & w10671;
assign w11165 = ~w10053 & w1856;
assign w11166 = ~w6444 & ~w3193;
assign w11167 = pi1337 & ~pi0262;
assign w11168 = w7703 & w15811;
assign w11169 = pi1169 & ~w13509;
assign w11170 = pi1256 & ~w11655;
assign w11171 = ~w5453 & ~pi1773;
assign w11172 = pi1736 & w1924;
assign w11173 = w6086 & w2436;
assign w11174 = ~w17482 & ~w4687;
assign w11175 = ~w10356 & ~w15690;
assign w11176 = ~pi3169 & w1843;
assign w11177 = w17475 & w17428;
assign w11178 = ~pi3318 & w7090;
assign w11179 = ~w5560 & w12733;
assign w11180 = pi0307 & w5274;
assign w11181 = w13509 & w7257;
assign w11182 = (pi1692 & ~w3023) | (pi1692 & ~w5855) | (~w3023 & ~w5855);
assign w11183 = ~pi2430 & w5075;
assign w11184 = ~w2540 & ~w9932;
assign w11185 = ~pi1711 & pi3132;
assign w11186 = ~w12830 & ~w7543;
assign w11187 = ~w3935 & ~w1378;
assign w11188 = ~w14560 & pi0232;
assign w11189 = w934 & pi0429;
assign w11190 = pi2234 & ~w11735;
assign w11191 = w2341 & ~w10235;
assign w11192 = w13509 & w5315;
assign w11193 = ~pi2195 & w9340;
assign w11194 = (~w10251 & ~w5517) | (~w10251 & w15430) | (~w5517 & w15430);
assign w11195 = (pi0906 & ~w13509) | (pi0906 & w8484) | (~w13509 & w8484);
assign w11196 = ~w2871 & ~w2177;
assign w11197 = (pi1143 & ~w5437) | (pi1143 & w17134) | (~w5437 & w17134);
assign w11198 = ~pi1824 & w17562;
assign w11199 = ~w11577 & ~w12314;
assign w11200 = ~pi0924 & w17490;
assign w11201 = ~w8399 & w6753;
assign w11202 = w10647 & ~w2821;
assign w11203 = pi1729 & w1924;
assign w11204 = ~pi0947 & w1126;
assign w11205 = (pi1022 & ~w13509) | (pi1022 & w15326) | (~w13509 & w15326);
assign w11206 = ~w8853 & ~w5049;
assign w11207 = ~pi2975 & w3223;
assign w11208 = ~w1445 & ~w16649;
assign w11209 = w10087 & ~w6575;
assign w11210 = ~pi0996 & w795;
assign w11211 = ~pi3169 & w12427;
assign w11212 = ~w3000 & ~pi2769;
assign w11213 = (pi1203 & ~w13509) | (pi1203 & w14635) | (~w13509 & w14635);
assign w11214 = ~pi0669 & w12197;
assign w11215 = w8795 & ~w12126;
assign w11216 = ~w18224 & w4025;
assign w11217 = ~pi3085 & w9504;
assign w11218 = w8337 & pi3292;
assign w11219 = ~pi3165 & w13730;
assign w11220 = ~pi3131 & w13730;
assign w11221 = ~w10340 & ~w11677;
assign w11222 = (pi0076 & w5421) | (pi0076 & w15417) | (w5421 & w15417);
assign w11223 = w539 & ~w1245;
assign w11224 = w13509 & w10132;
assign w11225 = ~pi3355 & w7090;
assign w11226 = ~w8858 & ~w5967;
assign w11227 = pi2168 & ~w15271;
assign w11228 = pi2573 & ~w5274;
assign w11229 = ~w995 & ~w14119;
assign w11230 = ~pi0732 & w17899;
assign w11231 = ~w1962 & pi1113;
assign w11232 = w7958 & w11060;
assign w11233 = ~w11786 & ~w18173;
assign w11234 = pi3063 & ~w3987;
assign w11235 = ~pi0088 & w9284;
assign w11236 = pi0089 & w9284;
assign w11237 = w7799 & w7774;
assign w11238 = ~w507 & ~w13256;
assign w11239 = ~w1791 & w16542;
assign w11240 = pi3132 & w653;
assign w11241 = ~pi3133 & w15839;
assign w11242 = pi1443 & ~w6448;
assign w11243 = pi2818 & w14148;
assign w11244 = ~pi2147 & w13065;
assign w11245 = ~pi3057 & ~pi3109;
assign w11246 = w13509 & w2600;
assign w11247 = w1516 & w12312;
assign w11248 = w9345 & w15241;
assign w11249 = ~pi3328 & w18259;
assign w11250 = ~w14692 & ~w20;
assign w11251 = w14768 & w11199;
assign w11252 = pi1789 & ~w15767;
assign w11253 = ~w17527 & ~w4048;
assign w11254 = w10312 & w12586;
assign w11255 = ~pi1073 & w12825;
assign w11256 = ~w3277 & ~w15461;
assign w11257 = ~w125 & ~w3865;
assign w11258 = ~pi1706 & ~pi1708;
assign w11259 = ~pi1269 & w9420;
assign w11260 = ~w14782 & w10998;
assign w11261 = ~w11770 & w5697;
assign w11262 = ~pi2319 & w3019;
assign w11263 = ~w14124 & w12761;
assign w11264 = pi0030 & ~w3748;
assign w11265 = ~w6172 & ~w11507;
assign w11266 = w16761 & w685;
assign w11267 = ~pi1773 & pi3139;
assign w11268 = w16575 & w1882;
assign w11269 = w13231 & ~w3374;
assign w11270 = pi3158 & w3615;
assign w11271 = ~pi3128 & w261;
assign w11272 = w3774 & w876;
assign w11273 = ~pi1037 & w6200;
assign w11274 = (pi1006 & ~w13509) | (pi1006 & w2488) | (~w13509 & w2488);
assign w11275 = pi3082 & w11406;
assign w11276 = ~w11338 & ~w7437;
assign w11277 = ~pi1717 & pi3153;
assign w11278 = w2341 & ~w14143;
assign w11279 = pi1816 & ~w3709;
assign w11280 = pi2777 & ~w15235;
assign w11281 = ~pi2974 & ~w12881;
assign w11282 = ~pi1957 & w12941;
assign w11283 = w15122 & ~pi2632;
assign w11284 = (pi0629 & ~w13509) | (pi0629 & w7780) | (~w13509 & w7780);
assign w11285 = pi1942 & ~w17683;
assign w11286 = w1306 & w6875;
assign w11287 = w2725 & ~w2776;
assign w11288 = (~pi0299 & ~w7807) | (~pi0299 & w697) | (~w7807 & w697);
assign w11289 = ~w3842 & ~w16755;
assign w11290 = (pi0779 & ~w13509) | (pi0779 & w1204) | (~w13509 & w1204);
assign w11291 = w13116 & ~w9399;
assign w11292 = w10818 & ~w8587;
assign w11293 = ~w6020 & ~w14319;
assign w11294 = pi2572 & ~w5274;
assign w11295 = ~pi0503 & ~pi1345;
assign w11296 = ~w18230 & ~w3582;
assign w11297 = pi1645 & ~w13753;
assign w11298 = w384 & w13688;
assign w11299 = (pi0387 & w5560) | (pi0387 & w15772) | (w5560 & w15772);
assign w11300 = pi1359 & w17413;
assign w11301 = w6857 & w14572;
assign w11302 = ~w7021 & ~w6135;
assign w11303 = ~w8176 & ~w6545;
assign w11304 = ~pi3088 & w9504;
assign w11305 = ~w2341 & pi0849;
assign w11306 = pi2318 & ~w3223;
assign w11307 = (pi0606 & ~w13509) | (pi0606 & w3483) | (~w13509 & w3483);
assign w11308 = ~w99 & ~w17779;
assign w11309 = ~w10252 & ~w16519;
assign w11310 = pi1476 & ~w9781;
assign w11311 = pi2839 & ~w11406;
assign w11312 = ~pi1805 & w16618;
assign w11313 = w5410 & w2246;
assign w11314 = ~w12622 & ~w3013;
assign w11315 = ~w10840 & ~w15484;
assign w11316 = pi2995 & pi1401;
assign w11317 = (pi0814 & ~w13509) | (pi0814 & w16489) | (~w13509 & w16489);
assign w11318 = ~w15096 & ~w16416;
assign w11319 = pi0112 & ~w2632;
assign w11320 = ~w5914 & ~w13205;
assign w11321 = ~w7724 & ~w2975;
assign w11322 = pi1368 & ~w1993;
assign w11323 = w12460 & w11898;
assign w11324 = ~pi2429 & w7455;
assign w11325 = ~pi2331 & w12755;
assign w11326 = ~w116 & ~w13093;
assign w11327 = ~w2341 & pi0829;
assign w11328 = w7030 & w848;
assign w11329 = pi1714 & ~w619;
assign w11330 = ~w4354 & ~w10390;
assign w11331 = ~w16506 & pi1230;
assign w11332 = ~w774 & ~w648;
assign w11333 = ~w9287 & w6746;
assign w11334 = ~w1513 & w15725;
assign w11335 = w2880 & w572;
assign w11336 = ~pi2954 & pi3199;
assign w11337 = w13509 & w17311;
assign w11338 = (pi0849 & ~w13509) | (pi0849 & w11305) | (~w13509 & w11305);
assign w11339 = pi2721 & ~w3555;
assign w11340 = ~w4589 & ~w2825;
assign w11341 = ~pi2191 & w2151;
assign w11342 = ~w3459 & ~w16327;
assign w11343 = w3333 & w9394;
assign w11344 = pi2634 & ~w9504;
assign w11345 = w17857 & w13556;
assign w11346 = ~w16575 & w5169;
assign w11347 = (pi1157 & ~w5437) | (pi1157 & w10730) | (~w5437 & w10730);
assign w11348 = ~w16278 & pi1107;
assign w11349 = ~w9895 & ~w4646;
assign w11350 = ~w7073 & ~w3845;
assign w11351 = w10338 & w3215;
assign w11352 = ~w7912 & w16661;
assign w11353 = ~w1855 & ~w1726;
assign w11354 = w8664 & w14851;
assign w11355 = pi3039 & ~w3987;
assign w11356 = w2325 & w12877;
assign w11357 = pi2087 & ~w17683;
assign w11358 = pi3136 & w11272;
assign w11359 = ~pi3171 & w17993;
assign w11360 = ~pi0077 & ~w10784;
assign w11361 = pi1145 & w9420;
assign w11362 = ~pi0053 & w922;
assign w11363 = pi1340 & ~w7705;
assign w11364 = ~w15122 & ~pi2877;
assign w11365 = ~pi2944 & ~w15587;
assign w11366 = ~pi3151 & ~pi3158;
assign w11367 = w6857 & w9664;
assign w11368 = ~pi0926 & w9110;
assign w11369 = w13509 & w4690;
assign w11370 = w7077 & ~w14465;
assign w11371 = ~w8182 & ~w2901;
assign w11372 = ~pi1944 & w7455;
assign w11373 = w13509 & w15012;
assign w11374 = ~w2014 & w10961;
assign w11375 = pi1531 & ~w14918;
assign w11376 = ~w487 & w660;
assign w11377 = ~pi0328 & w2196;
assign w11378 = ~pi3087 & w261;
assign w11379 = ~w9479 & ~w18397;
assign w11380 = ~pi0905 & w795;
assign w11381 = w11345 & w113;
assign w11382 = ~pi0327 & w4058;
assign w11383 = ~w3000 & w15122;
assign w11384 = ~w8060 & ~w5549;
assign w11385 = ~w12460 & w15710;
assign w11386 = ~pi2379 & w8617;
assign w11387 = (pi1104 & ~w13509) | (pi1104 & w10845) | (~w13509 & w10845);
assign w11388 = pi1778 & w15622;
assign w11389 = w9440 & pi0130;
assign w11390 = w384 & w16916;
assign w11391 = pi3141 & w2253;
assign w11392 = w17562 & pi2569;
assign w11393 = ~w16575 & w100;
assign w11394 = ~w1962 & pi0642;
assign w11395 = ~pi2203 & w12724;
assign w11396 = pi2504 & ~w226;
assign w11397 = (pi0005 & ~w1766) | (pi0005 & w1958) | (~w1766 & w1958);
assign w11398 = w968 & ~pi0328;
assign w11399 = ~pi1407 & w4517;
assign w11400 = ~w16278 & pi0698;
assign w11401 = ~w5820 & ~w3503;
assign w11402 = ~w9715 & ~w4915;
assign w11403 = ~w11247 & w341;
assign w11404 = ~w2758 & ~w1344;
assign w11405 = w10533 & ~w10781;
assign w11406 = ~pi2949 & w5675;
assign w11407 = ~pi3098 & w15235;
assign w11408 = ~pi1902 & pi0205;
assign w11409 = ~w4724 & ~w6173;
assign w11410 = ~pi3100 & w261;
assign w11411 = pi2048 & ~w10158;
assign w11412 = ~w10319 & ~w2141;
assign w11413 = pi1519 & w13753;
assign w11414 = (pi0805 & ~w13509) | (pi0805 & w12727) | (~w13509 & w12727);
assign w11415 = w17683 & w2753;
assign w11416 = ~w1775 & ~w1660;
assign w11417 = ~pi3169 & w14753;
assign w11418 = ~pi3170 & w15839;
assign w11419 = pi2444 & ~w10299;
assign w11420 = ~w7353 & ~w9562;
assign w11421 = w17741 & w16744;
assign w11422 = ~w9502 & ~w15583;
assign w11423 = ~w14494 & ~w10006;
assign w11424 = ~pi3159 & w15839;
assign w11425 = pi2753 & ~w6463;
assign w11426 = pi2034 & ~w17646;
assign w11427 = pi1918 & ~w10299;
assign w11428 = ~pi3085 & w11406;
assign w11429 = w14794 & w9007;
assign w11430 = ~pi2881 & w15122;
assign w11431 = ~pi0706 & w3106;
assign w11432 = ~w13918 & ~w1694;
assign w11433 = ~w1069 & w18516;
assign w11434 = pi1647 & ~w13753;
assign w11435 = ~w16278 & pi1027;
assign w11436 = ~pi0682 & w9110;
assign w11437 = ~w11329 & ~w2815;
assign w11438 = w7799 & w4973;
assign w11439 = w13509 & w4064;
assign w11440 = w11345 & w7330;
assign w11441 = ~w14611 & ~w17255;
assign w11442 = ~w2523 & w11744;
assign w11443 = ~w2615 & ~w7028;
assign w11444 = ~w4330 & ~w5934;
assign w11445 = w12460 & w6515;
assign w11446 = pi1131 & w14073;
assign w11447 = ~w8444 & ~pi0494;
assign w11448 = ~pi0494 & ~pi1345;
assign w11449 = pi1974 & ~w16815;
assign w11450 = (pi0253 & ~w325) | (pi0253 & w14008) | (~w325 & w14008);
assign w11451 = ~w12785 & ~w1507;
assign w11452 = pi2455 & ~w14524;
assign w11453 = ~w15122 & ~pi2887;
assign w11454 = ~w16575 & w6328;
assign w11455 = pi1619 & ~w13753;
assign w11456 = ~pi2949 & w4095;
assign w11457 = ~w2911 & ~w9793;
assign w11458 = pi2911 & ~w16598;
assign w11459 = w18345 & ~w6499;
assign w11460 = ~w11954 & ~w15674;
assign w11461 = w11209 & ~w14057;
assign w11462 = ~w6697 & pi0664;
assign w11463 = ~pi3135 & w1843;
assign w11464 = ~w9425 & ~pi0495;
assign w11465 = ~pi0617 & w14641;
assign w11466 = pi1649 & ~w6072;
assign w11467 = ~pi2186 & w2151;
assign w11468 = ~pi3002 & w1326;
assign w11469 = ~pi2208 & w5075;
assign w11470 = w13509 & w9958;
assign w11471 = w13509 & w9959;
assign w11472 = ~w15228 & ~w10410;
assign w11473 = ~w16670 & ~w16945;
assign w11474 = (~pi0896 & w461) | (~pi0896 & w12695) | (w461 & w12695);
assign w11475 = ~pi0647 & w3791;
assign w11476 = (~pi1763 & ~w7799) | (~pi1763 & w4235) | (~w7799 & w4235);
assign w11477 = (pi1891 & w2014) | (pi1891 & w834) | (w2014 & w834);
assign w11478 = pi2072 & ~w17683;
assign w11479 = ~pi1219 & ~w5652;
assign w11480 = w384 & w14618;
assign w11481 = w14560 & pi0342;
assign w11482 = pi1943 & ~w17646;
assign w11483 = (pi0898 & ~w13509) | (pi0898 & w9453) | (~w13509 & w9453);
assign w11484 = ~pi2251 & w3019;
assign w11485 = ~w4955 & w14982;
assign w11486 = ~w2956 & ~w13585;
assign w11487 = ~w15714 & ~w14055;
assign w11488 = ~w17894 & ~w6884;
assign w11489 = ~w17665 & ~w4698;
assign w11490 = pi2966 & pi2480;
assign w11491 = ~pi0504 & ~pi1186;
assign w11492 = ~w5955 & ~w18318;
assign w11493 = w1127 & ~w16019;
assign w11494 = pi1600 & ~w9781;
assign w11495 = ~pi3166 & w1843;
assign w11496 = w2466 & w9033;
assign w11497 = pi2117 & ~w412;
assign w11498 = ~w3000 & ~pi2927;
assign w11499 = ~pi3052 & w11406;
assign w11500 = ~w12460 & w18279;
assign w11501 = w13509 & w4373;
assign w11502 = w5017 & w4176;
assign w11503 = ~w12153 & ~w11243;
assign w11504 = w6649 & ~w15642;
assign w11505 = w8966 & w7924;
assign w11506 = pi1851 & ~w2732;
assign w11507 = w13509 & w13642;
assign w11508 = ~pi0579 & w795;
assign w11509 = ~pi3037 & pi3131;
assign w11510 = ~w7209 & ~w12491;
assign w11511 = ~w7938 & ~w533;
assign w11512 = pi1376 & ~w8966;
assign w11513 = pi1384 & ~w17935;
assign w11514 = ~w16128 & ~w18409;
assign w11515 = pi1801 & pi3165;
assign w11516 = w62 & ~w4964;
assign w11517 = pi1161 & pi0077;
assign w11518 = w11345 & w4519;
assign w11519 = pi2972 & w3987;
assign w11520 = w15328 & ~w10241;
assign w11521 = ~w8170 & ~w14064;
assign w11522 = ~w6640 & ~w6995;
assign w11523 = ~w807 & ~w7390;
assign w11524 = w10189 & ~pi0478;
assign w11525 = pi1741 & ~w4058;
assign w11526 = ~w17566 & ~w6087;
assign w11527 = ~w3203 & pi0904;
assign w11528 = pi3082 & w15235;
assign w11529 = pi2629 & ~w9504;
assign w11530 = (pi0846 & ~w13509) | (pi0846 & w13167) | (~w13509 & w13167);
assign w11531 = pi2616 & ~w261;
assign w11532 = ~w8341 & ~w17550;
assign w11533 = pi1536 & w13753;
assign w11534 = ~w6768 & ~w14943;
assign w11535 = ~w10277 & ~w4774;
assign w11536 = w7799 & w5545;
assign w11537 = ~pi2144 & w12941;
assign w11538 = ~w8934 & ~w3286;
assign w11539 = (~w1877 & ~w5517) | (~w1877 & w12757) | (~w5517 & w12757);
assign w11540 = pi3157 & w5457;
assign w11541 = ~w9299 & ~w1242;
assign w11542 = ~w14687 & ~w6131;
assign w11543 = ~w7187 & ~w8564;
assign w11544 = ~w14417 & w1326;
assign w11545 = w13569 & w3550;
assign w11546 = ~w15036 & ~w15955;
assign w11547 = ~pi3146 & w15048;
assign w11548 = ~w633 & ~w3105;
assign w11549 = pi3040 & w16502;
assign w11550 = ~w17882 & w17753;
assign w11551 = w2725 & ~w15296;
assign w11552 = ~w14521 & ~w12356;
assign w11553 = ~w3816 & ~w6350;
assign w11554 = pi3024 & w16502;
assign w11555 = ~w18240 & ~w7550;
assign w11556 = ~pi2085 & w16041;
assign w11557 = ~w5044 & w9761;
assign w11558 = pi2418 & ~w3223;
assign w11559 = w6857 & w9902;
assign w11560 = ~pi3091 & w3555;
assign w11561 = w9440 & pi0150;
assign w11562 = ~w2689 & ~w723;
assign w11563 = (~pi0294 & ~w6857) | (~pi0294 & w10149) | (~w6857 & w10149);
assign w11564 = w451 & w8205;
assign w11565 = ~w7374 & w7509;
assign w11566 = ~w3237 & ~w17716;
assign w11567 = w9216 & pi0502;
assign w11568 = ~w13231 & pi0558;
assign w11569 = w12040 & w11302;
assign w11570 = w7228 & w5711;
assign w11571 = ~w16575 & w9446;
assign w11572 = pi1483 & w13753;
assign w11573 = ~pi1914 & w9340;
assign w11574 = pi2677 & ~w226;
assign w11575 = w2725 & ~w11978;
assign w11576 = pi0052 & w922;
assign w11577 = ~pi2440 & w5075;
assign w11578 = ~w16619 & ~w7347;
assign w11579 = ~w7151 & ~w15773;
assign w11580 = (pi0517 & ~w13509) | (pi0517 & w7366) | (~w13509 & w7366);
assign w11581 = (w17577 & w11928) | (w17577 & w6870) | (w11928 & w6870);
assign w11582 = pi2252 & ~w18209;
assign w11583 = ~pi3155 & w11701;
assign w11584 = ~w17481 & ~w2055;
assign w11585 = ~w14792 & w15539;
assign w11586 = w11383 & w14948;
assign w11587 = ~w15628 & ~w9091;
assign w11588 = ~w2397 & ~w15159;
assign w11589 = pi1748 & ~w3555;
assign w11590 = w7703 & w18195;
assign w11591 = pi2757 & ~w4667;
assign w11592 = ~w7956 & ~w6580;
assign w11593 = pi2619 & ~w261;
assign w11594 = ~pi3146 & ~pi3160;
assign w11595 = (pi1756 & w7215) | (pi1756 & w16405) | (w7215 & w16405);
assign w11596 = ~pi0968 & w3106;
assign w11597 = ~w9723 & w1684;
assign w11598 = ~w6638 & ~w15386;
assign w11599 = w1368 & pi0392;
assign w11600 = (pi1177 & w14073) | (pi1177 & w15970) | (w14073 & w15970);
assign w11601 = ~w15808 & pi1098;
assign w11602 = ~w2725 & pi0783;
assign w11603 = ~w5245 & ~w18219;
assign w11604 = w1962 & ~w6922;
assign w11605 = w17665 & ~w10660;
assign w11606 = ~pi2294 & ~w15974;
assign w11607 = ~w5617 & ~w15676;
assign w11608 = w13149 & w8671;
assign w11609 = ~pi1700 & w4667;
assign w11610 = ~w17312 & ~w567;
assign w11611 = ~pi0293 & w4058;
assign w11612 = pi1608 & ~w9781;
assign w11613 = ~w16954 & w7858;
assign w11614 = w11383 & w14511;
assign w11615 = ~w12666 & ~w8753;
assign w11616 = w4002 & w11899;
assign w11617 = ~w1368 & ~pi0472;
assign w11618 = w254 & w2878;
assign w11619 = pi0110 & ~w2632;
assign w11620 = ~w7077 & pi0813;
assign w11621 = ~pi0049 & w922;
assign w11622 = pi0050 & w922;
assign w11623 = ~pi0059 & ~w17103;
assign w11624 = ~pi0964 & w1147;
assign w11625 = (pi0374 & w6195) | (pi0374 & w4427) | (w6195 & w4427);
assign w11626 = w13509 & w15269;
assign w11627 = ~w3614 & ~w18408;
assign w11628 = ~w1262 & ~w11119;
assign w11629 = pi2760 & w14148;
assign w11630 = pi3152 & w545;
assign w11631 = ~w4771 & ~w5714;
assign w11632 = ~w17671 & ~w4351;
assign w11633 = pi2795 & w7965;
assign w11634 = ~w15347 & ~w13135;
assign w11635 = pi1792 & ~w3140;
assign w11636 = ~w2130 & w858;
assign w11637 = pi2981 & w13584;
assign w11638 = ~w15741 & ~w1801;
assign w11639 = w15450 & ~pi1181;
assign w11640 = pi2560 & ~w5274;
assign w11641 = (~pi0967 & ~w13509) | (~pi0967 & w2639) | (~w13509 & w2639);
assign w11642 = ~pi3299 & w6072;
assign w11643 = ~pi0291 & w2196;
assign w11644 = w11822 & w11206;
assign w11645 = ~w700 & w7693;
assign w11646 = w16575 & w5067;
assign w11647 = pi3160 & ~pi3485;
assign w11648 = ~pi0752 & w17490;
assign w11649 = ~w1543 & w3409;
assign w11650 = w13509 & w18571;
assign w11651 = ~w12674 & ~w9150;
assign w11652 = ~w13818 & ~w6981;
assign w11653 = ~w2101 & ~w9547;
assign w11654 = ~w7652 & w12424;
assign w11655 = ~w11034 & ~w3315;
assign w11656 = w5453 & pi2587;
assign w11657 = ~w17986 & ~w5822;
assign w11658 = pi1378 & ~w3615;
assign w11659 = pi3138 & w8113;
assign w11660 = ~w6785 & pi1167;
assign w11661 = ~w5828 & ~w12780;
assign w11662 = ~w10077 & w7069;
assign w11663 = w968 & ~pi0276;
assign w11664 = (pi0408 & w5560) | (pi0408 & w10599) | (w5560 & w10599);
assign w11665 = ~w15808 & pi0744;
assign w11666 = ~w12460 & w14490;
assign w11667 = ~pi3147 & w4310;
assign w11668 = ~w16962 & ~w15210;
assign w11669 = w3203 & ~w16498;
assign w11670 = pi1285 & pi1345;
assign w11671 = ~pi1985 & w8370;
assign w11672 = w922 & pi0048;
assign w11673 = pi1214 & ~pi3193;
assign w11674 = pi2467 & ~w9504;
assign w11675 = ~pi2209 & w5075;
assign w11676 = ~pi2107 & w12755;
assign w11677 = ~pi3326 & w9781;
assign w11678 = ~w16175 & w10661;
assign w11679 = (pi1900 & w2014) | (pi1900 & w3301) | (w2014 & w3301);
assign w11680 = ~w7649 & ~w355;
assign w11681 = ~pi3157 & w3805;
assign w11682 = ~w6646 & w3305;
assign w11683 = w13509 & w58;
assign w11684 = ~pi3164 & w12427;
assign w11685 = pi1334 & ~w17504;
assign w11686 = w2725 & ~w6680;
assign w11687 = ~pi3163 & w3679;
assign w11688 = w17559 & w2246;
assign w11689 = w17477 & w553;
assign w11690 = pi3135 & w9520;
assign w11691 = w13509 & w6850;
assign w11692 = pi1589 & w4683;
assign w11693 = ~w3681 & ~w4608;
assign w11694 = ~w13367 & ~w1300;
assign w11695 = pi0111 & ~w2632;
assign w11696 = ~w13731 & w12018;
assign w11697 = w4923 & w8955;
assign w11698 = w7703 & w10682;
assign w11699 = ~w15255 & ~w6593;
assign w11700 = pi2786 & ~w3555;
assign w11701 = ~w4020 & w14524;
assign w11702 = ~pi3172 & w11132;
assign w11703 = pi2913 & ~w8430;
assign w11704 = pi2885 & ~w5274;
assign w11705 = w7844 & ~w17513;
assign w11706 = ~w12190 & ~w12924;
assign w11707 = pi3172 & w2732;
assign w11708 = ~w10155 & ~w13709;
assign w11709 = ~w6697 & pi0676;
assign w11710 = ~w1387 & ~w1065;
assign w11711 = w532 & w5221;
assign w11712 = pi1652 & ~w13753;
assign w11713 = pi1849 & ~w12558;
assign w11714 = ~pi1827 & w14347;
assign w11715 = ~w16554 & ~w8490;
assign w11716 = ~w9188 & ~w12;
assign w11717 = w7844 & w1217;
assign w11718 = w13509 & w5556;
assign w11719 = ~w10872 & ~w4688;
assign w11720 = ~w15915 & ~w14677;
assign w11721 = w17562 & pi1854;
assign w11722 = ~w18399 & ~w18353;
assign w11723 = w13840 & pi1708;
assign w11724 = w968 & ~pi0292;
assign w11725 = w13231 & ~w6033;
assign w11726 = ~pi3314 & w6448;
assign w11727 = ~w3000 & ~pi2669;
assign w11728 = w13308 & ~w2623;
assign w11729 = ~w14781 & ~w9017;
assign w11730 = ~pi3330 & w6072;
assign w11731 = pi1365 & w15290;
assign w11732 = ~pi3337 & w14918;
assign w11733 = ~w16238 & ~w3362;
assign w11734 = (pi0365 & w6195) | (pi0365 & w13538) | (w6195 & w13538);
assign w11735 = w14651 & w14245;
assign w11736 = ~w7332 & ~w11217;
assign w11737 = (pi0712 & ~w13509) | (pi0712 & w3447) | (~w13509 & w3447);
assign w11738 = w13509 & w14504;
assign w11739 = w134 & w17899;
assign w11740 = w13184 & w1493;
assign w11741 = ~w2790 & ~w5008;
assign w11742 = w7703 & w7683;
assign w11743 = w10000 & w18002;
assign w11744 = (pi1788 & w7215) | (pi1788 & w18290) | (w7215 & w18290);
assign w11745 = ~w1492 & ~w15406;
assign w11746 = ~pi1918 & w9340;
assign w11747 = pi1407 & w5043;
assign w11748 = pi2177 & ~w14524;
assign w11749 = w13231 & ~w12800;
assign w11750 = pi1589 & ~w7946;
assign w11751 = ~pi2522 & w14148;
assign w11752 = ~w16223 & ~w15658;
assign w11753 = w7844 & ~w13195;
assign w11754 = ~w1348 & ~w6833;
assign w11755 = ~w13742 & w13846;
assign w11756 = w12460 & w1999;
assign w11757 = w4508 & w614;
assign w11758 = w15808 & ~w6647;
assign w11759 = pi3153 & w12558;
assign w11760 = w10000 & w18403;
assign w11761 = ~pi3155 & pi3207;
assign w11762 = ~pi0888 & w1126;
assign w11763 = ~pi3165 & w13570;
assign w11764 = ~pi1114 & w12197;
assign w11765 = (pi0686 & ~w13509) | (pi0686 & w7866) | (~w13509 & w7866);
assign w11766 = ~w3878 & ~w12027;
assign w11767 = ~pi1026 & w3106;
assign w11768 = ~w13882 & ~w3605;
assign w11769 = ~pi3299 & w18259;
assign w11770 = w14322 & w15663;
assign w11771 = ~w18126 & ~w7863;
assign w11772 = pi1782 & ~w8829;
assign w11773 = ~w14560 & pi0208;
assign w11774 = ~w8486 & ~w9621;
assign w11775 = pi3043 & ~w3987;
assign w11776 = w5383 & ~pi2966;
assign w11777 = ~w17970 & ~w12872;
assign w11778 = (pi0620 & ~w13509) | (pi0620 & w5054) | (~w13509 & w5054);
assign w11779 = ~w10891 & ~w16410;
assign w11780 = ~w17980 & ~w286;
assign w11781 = ~pi0990 & w11739;
assign w11782 = ~pi2237 & w2151;
assign w11783 = ~pi0580 & w795;
assign w11784 = ~w9587 & ~w18468;
assign w11785 = pi1986 & ~w7858;
assign w11786 = (pi0388 & w5560) | (pi0388 & w17015) | (w5560 & w17015);
assign w11787 = ~w9994 & ~w1458;
assign w11788 = ~w1791 & w1588;
assign w11789 = w13509 & w7589;
assign w11790 = ~pi3333 & w16922;
assign w11791 = ~w16798 & ~w9676;
assign w11792 = ~w6785 & pi0861;
assign w11793 = w7369 & w4447;
assign w11794 = ~w11828 & ~w17870;
assign w11795 = w7703 & w13411;
assign w11796 = pi2495 & ~w9504;
assign w11797 = ~pi0655 & w3791;
assign w11798 = ~w3426 & w5212;
assign w11799 = (pi0949 & ~w13509) | (pi0949 & w15769) | (~w13509 & w15769);
assign w11800 = pi0079 & ~pi0082;
assign w11801 = ~pi2425 & w11313;
assign w11802 = ~w18044 & ~w13302;
assign w11803 = ~w14228 & pi0627;
assign w11804 = ~w3992 & ~w18067;
assign w11805 = pi2533 & w15191;
assign w11806 = ~w16163 & w10984;
assign w11807 = pi1222 & w5566;
assign w11808 = w6697 & ~w16498;
assign w11809 = ~pi3147 & ~pi3160;
assign w11810 = ~w14939 & w6600;
assign w11811 = ~w15149 & ~w17231;
assign w11812 = ~w18410 & ~w10865;
assign w11813 = ~w8307 & ~w335;
assign w11814 = w1391 & ~w14597;
assign w11815 = pi2932 & ~w9504;
assign w11816 = ~w709 & pi1285;
assign w11817 = ~w15580 & w4230;
assign w11818 = w8789 & w2184;
assign w11819 = pi2419 & ~w10158;
assign w11820 = w6857 & w14214;
assign w11821 = ~w17248 & pi1057;
assign w11822 = ~w16001 & ~w4462;
assign w11823 = ~w13636 & ~w3031;
assign w11824 = w15122 & ~pi2715;
assign w11825 = ~w13367 & ~w9980;
assign w11826 = pi1475 & ~w9781;
assign w11827 = pi1572 & ~w13753;
assign w11828 = pi2793 & ~w6463;
assign w11829 = ~w17122 & ~w9834;
assign w11830 = pi0322 & pi3229;
assign w11831 = ~pi2772 & w13343;
assign w11832 = ~w18138 & ~w11943;
assign w11833 = w13453 & w16774;
assign w11834 = ~pi3170 & w11132;
assign w11835 = ~w4937 & ~w8227;
assign w11836 = pi3165 & w14951;
assign w11837 = w15122 & ~pi2596;
assign w11838 = pi2599 & ~w16815;
assign w11839 = pi3136 & w5762;
assign w11840 = (pi0324 & w3055) | (pi0324 & w6852) | (w3055 & w6852);
assign w11841 = ~pi0848 & w93;
assign w11842 = pi1560 & ~w18259;
assign w11843 = ~w253 & ~w8146;
assign w11844 = ~pi3337 & w16922;
assign w11845 = ~w14648 & ~pi2723;
assign w11846 = ~pi0731 & w17899;
assign w11847 = ~w185 & ~w12509;
assign w11848 = ~w1426 & w16057;
assign w11849 = ~w9969 & ~w1970;
assign w11850 = pi0124 & w3748;
assign w11851 = ~w11170 & ~w16860;
assign w11852 = ~w11466 & ~w18013;
assign w11853 = w9440 & pi0167;
assign w11854 = ~pi2083 & w17439;
assign w11855 = w10189 & ~pi0454;
assign w11856 = pi0205 & w10959;
assign w11857 = w12460 & w10133;
assign w11858 = w7307 & w1904;
assign w11859 = ~pi0793 & w543;
assign w11860 = ~w15957 & ~w8160;
assign w11861 = ~pi1203 & w93;
assign w11862 = pi2650 & ~w16815;
assign w11863 = (pi1101 & ~w13509) | (pi1101 & w14809) | (~w13509 & w14809);
assign w11864 = pi1315 & ~w13834;
assign w11865 = w8337 & pi3275;
assign w11866 = ~pi0753 & w17490;
assign w11867 = pi2295 & ~w261;
assign w11868 = ~pi0884 & w1126;
assign w11869 = ~w11570 & w14908;
assign w11870 = ~w18245 & ~w9827;
assign w11871 = ~w3171 & ~w10645;
assign w11872 = ~pi3144 & ~w16370;
assign w11873 = w13509 & w6813;
assign w11874 = ~w2602 & ~w16583;
assign w11875 = ~pi2350 & w8617;
assign w11876 = ~w15618 & ~w7029;
assign w11877 = ~w748 & ~w11751;
assign w11878 = ~w17862 & ~w9458;
assign w11879 = ~w18016 & ~w17981;
assign w11880 = ~w9395 & ~w18198;
assign w11881 = w12460 & w13639;
assign w11882 = ~pi2025 & w7455;
assign w11883 = ~pi3039 & ~pi3207;
assign w11884 = ~w1791 & w6106;
assign w11885 = ~w8318 & ~w5895;
assign w11886 = ~w17237 & ~w6518;
assign w11887 = pi0306 & w18583;
assign w11888 = pi3139 & w12558;
assign w11889 = ~pi3171 & w1843;
assign w11890 = pi2996 & ~w3987;
assign w11891 = pi1661 & ~w6072;
assign w11892 = pi1779 & ~w15767;
assign w11893 = ~w11772 & ~w12163;
assign w11894 = w1368 & pi0409;
assign w11895 = ~w10803 & ~w18480;
assign w11896 = (pi0832 & ~w13509) | (pi0832 & w1261) | (~w13509 & w1261);
assign w11897 = ~pi3078 & pi3143;
assign w11898 = w9440 & pi0194;
assign w11899 = ~w16191 & ~w3446;
assign w11900 = ~w5665 & ~w15452;
assign w11901 = ~w10792 & ~w250;
assign w11902 = ~w8267 & ~w9346;
assign w11903 = w7656 & pi0476;
assign w11904 = ~w6785 & pi0856;
assign w11905 = ~pi2990 & ~w3987;
assign w11906 = ~w6624 & ~w628;
assign w11907 = w7703 & w11283;
assign w11908 = w1962 & ~w15173;
assign w11909 = ~pi0746 & w17490;
assign w11910 = ~w13329 & ~pi0486;
assign w11911 = pi0023 & ~w14148;
assign w11912 = w8658 & pi1782;
assign w11913 = ~pi3157 & w17993;
assign w11914 = w13509 & w18496;
assign w11915 = pi2508 & w384;
assign w11916 = w16575 & w15716;
assign w11917 = pi3032 & ~pi3135;
assign w11918 = ~pi2641 & w15122;
assign w11919 = w539 & ~w15953;
assign w11920 = ~pi2188 & w2151;
assign w11921 = w12126 & ~w489;
assign w11922 = (pi0317 & w3055) | (pi0317 & w4269) | (w3055 & w4269);
assign w11923 = (pi0863 & ~w13509) | (pi0863 & w17642) | (~w13509 & w17642);
assign w11924 = ~w1975 & w1473;
assign w11925 = ~w16099 & w13087;
assign w11926 = pi2521 & w4140;
assign w11927 = w17248 & w15609;
assign w11928 = ~pi0492 & ~w13367;
assign w11929 = ~w11406 & ~w18296;
assign w11930 = ~pi3147 & w11701;
assign w11931 = ~pi1931 & w11313;
assign w11932 = ~w3504 & w7341;
assign w11933 = ~pi0896 & ~w2621;
assign w11934 = ~pi3163 & w17313;
assign w11935 = ~pi0875 & w1126;
assign w11936 = w14061 & w12421;
assign w11937 = ~w17534 & ~w14414;
assign w11938 = ~w4866 & ~w17364;
assign w11939 = ~w15019 & w6811;
assign w11940 = ~pi0736 & w17899;
assign w11941 = ~w2341 & pi0848;
assign w11942 = ~pi1209 & ~w2270;
assign w11943 = w13509 & w9024;
assign w11944 = (pi1105 & ~w13509) | (pi1105 & w5455) | (~w13509 & w5455);
assign w11945 = ~w2703 & ~w7120;
assign w11946 = ~w6567 & w16173;
assign w11947 = w12460 & w14529;
assign w11948 = pi2704 & ~w3555;
assign w11949 = ~w11442 & w5042;
assign w11950 = pi1397 & w2925;
assign w11951 = ~w3387 & ~w17901;
assign w11952 = pi0256 & pi0257;
assign w11953 = (pi0766 & ~w13509) | (pi0766 & w14432) | (~w13509 & w14432);
assign w11954 = ~w15450 & w16954;
assign w11955 = w17562 & pi2502;
assign w11956 = pi1168 & ~w13509;
assign w11957 = pi1734 & w1924;
assign w11958 = ~w2378 & ~w4776;
assign w11959 = w17248 & ~w14143;
assign w11960 = pi2745 & ~w226;
assign w11961 = pi0123 & w3748;
assign w11962 = ~w3055 & w16286;
assign w11963 = w9705 & w13548;
assign w11964 = ~w18083 & ~w2401;
assign w11965 = ~pi3090 & w226;
assign w11966 = ~pi2918 & w17770;
assign w11967 = w2341 & ~w2587;
assign w11968 = ~w4247 & ~w17625;
assign w11969 = ~w10978 & ~w18099;
assign w11970 = ~w6697 & pi1013;
assign w11971 = w3295 & w7123;
assign w11972 = ~w12151 & ~w8007;
assign w11973 = ~pi0485 & ~pi1345;
assign w11974 = pi0026 & ~w3748;
assign w11975 = ~w18486 & w7720;
assign w11976 = w6649 & ~w3998;
assign w11977 = ~pi2344 & w16041;
assign w11978 = ~w8695 & ~w4234;
assign w11979 = ~w7844 & pi0600;
assign w11980 = ~w2341 & pi0828;
assign w11981 = ~w17577 & w9425;
assign w11982 = w54 & w9590;
assign w11983 = ~pi3290 & w6448;
assign w11984 = pi0015 & ~w14148;
assign w11985 = ~w10592 & ~w13367;
assign w11986 = w14833 & w614;
assign w11987 = ~w6697 & pi0661;
assign w11988 = w7307 & w3296;
assign w11989 = ~w1368 & ~pi0475;
assign w11990 = ~w11992 & ~w632;
assign w11991 = ~w15087 & ~w18025;
assign w11992 = ~pi1309 & ~pi3214;
assign w11993 = ~pi0619 & w14641;
assign w11994 = ~w16415 & ~w797;
assign w11995 = ~w17869 & ~w10945;
assign w11996 = pi3131 & w7946;
assign w11997 = w9744 & w5111;
assign w11998 = ~w14385 & ~w4069;
assign w11999 = pi1660 & ~w6072;
assign w12000 = w1962 & w15609;
assign w12001 = ~w3033 & ~w12560;
assign w12002 = ~pi2417 & w5075;
assign w12003 = w709 & pi1895;
assign w12004 = pi2662 & ~w15235;
assign w12005 = w8304 & ~w18086;
assign w12006 = pi3141 & w18497;
assign w12007 = ~w2859 & ~w943;
assign w12008 = ~w14036 & w12150;
assign w12009 = ~w13432 & ~w4694;
assign w12010 = ~w17695 & ~w10551;
assign w12011 = ~w3243 & pi0338;
assign w12012 = ~pi2308 & w12941;
assign w12013 = pi2511 & ~w9504;
assign w12014 = pi3150 & w3987;
assign w12015 = w5437 & w2250;
assign w12016 = w13509 & w10740;
assign w12017 = ~pi3089 & w3555;
assign w12018 = ~w1977 & ~w5725;
assign w12019 = ~pi3333 & w17935;
assign w12020 = pi2840 & w605;
assign w12021 = (pi0555 & ~w13509) | (pi0555 & w17807) | (~w13509 & w17807);
assign w12022 = pi2186 & ~w11735;
assign w12023 = pi1569 & ~w13753;
assign w12024 = w12040 & ~w6922;
assign w12025 = w13509 & w3341;
assign w12026 = w13231 & ~w11978;
assign w12027 = ~w10971 & ~w15819;
assign w12028 = (pi0720 & ~w13509) | (pi0720 & w2096) | (~w13509 & w2096);
assign w12029 = w16487 & w3150;
assign w12030 = ~w15880 & w1210;
assign w12031 = ~pi2848 & w14148;
assign w12032 = pi2849 & w14148;
assign w12033 = ~w10919 & ~w17607;
assign w12034 = ~w5576 & ~w17263;
assign w12035 = ~pi3132 & pi3207;
assign w12036 = ~pi3065 & ~pi3207;
assign w12037 = ~w1364 & w4194;
assign w12038 = ~w9860 & ~w2687;
assign w12039 = w9847 & ~w9145;
assign w12040 = w7254 & w15907;
assign w12041 = ~w8890 & ~w15929;
assign w12042 = ~pi1033 & w17490;
assign w12043 = w13509 & w8558;
assign w12044 = ~pi2074 & w17439;
assign w12045 = (pi1000 & ~w13509) | (pi1000 & w10705) | (~w13509 & w10705);
assign w12046 = pi1360 & ~w4256;
assign w12047 = ~pi0838 & w93;
assign w12048 = ~pi3094 & w261;
assign w12049 = w12460 & w11853;
assign w12050 = ~pi2329 & w3019;
assign w12051 = w10544 & w98;
assign w12052 = ~w7350 & ~w7951;
assign w12053 = ~pi2918 & ~pi3231;
assign w12054 = (pi1036 & ~w13509) | (pi1036 & w7984) | (~w13509 & w7984);
assign w12055 = ~w2534 & ~w8535;
assign w12056 = ~w14627 & ~w571;
assign w12057 = ~pi2967 & w13427;
assign w12058 = ~w13765 & w17368;
assign w12059 = pi2836 & ~w11406;
assign w12060 = ~w18515 & w14878;
assign w12061 = ~w10248 & ~w2068;
assign w12062 = pi3113 & ~w16502;
assign w12063 = (pi0764 & ~w13509) | (pi0764 & w122) | (~w13509 & w122);
assign w12064 = ~w12395 & w2893;
assign w12065 = w15808 & ~w14465;
assign w12066 = pi2428 & ~w3223;
assign w12067 = ~w2551 & ~w2050;
assign w12068 = pi3154 & w14951;
assign w12069 = ~w5788 & ~w12464;
assign w12070 = pi2185 & ~w11735;
assign w12071 = ~pi3110 & ~pi3207;
assign w12072 = w1368 & pi0401;
assign w12073 = ~pi1085 & w543;
assign w12074 = ~pi0876 & w1126;
assign w12075 = ~w16575 & w13958;
assign w12076 = ~w14705 & ~w4911;
assign w12077 = ~pi2660 & w17213;
assign w12078 = ~w8830 & ~w3175;
assign w12079 = ~pi3170 & w1843;
assign w12080 = pi3007 & ~w16502;
assign w12081 = w14719 & w15991;
assign w12082 = ~w2341 & pi1060;
assign w12083 = (pi0375 & w6195) | (pi0375 & w6934) | (w6195 & w6934);
assign w12084 = pi1572 & ~w18259;
assign w12085 = ~pi0148 & pi0187;
assign w12086 = pi2388 & ~w10158;
assign w12087 = w16506 & ~w14597;
assign w12088 = w16278 & ~w13028;
assign w12089 = ~w9936 & ~w15496;
assign w12090 = w11286 & w8292;
assign w12091 = w6649 & ~w2143;
assign w12092 = w13509 & w10331;
assign w12093 = ~pi0678 & w9110;
assign w12094 = pi2888 & ~w5274;
assign w12095 = (pi1676 & w5855) | (pi1676 & w8376) | (w5855 & w8376);
assign w12096 = ~pi0483 & pi3401;
assign w12097 = ~w6336 & ~w2522;
assign w12098 = ~w3054 & w4613;
assign w12099 = (pi1100 & ~w13509) | (pi1100 & w9128) | (~w13509 & w9128);
assign w12100 = pi1519 & ~w14918;
assign w12101 = pi0052 & ~w14148;
assign w12102 = ~pi1716 & ~pi3164;
assign w12103 = ~w1256 & ~w17003;
assign w12104 = ~pi3155 & w17993;
assign w12105 = ~w9181 & ~w11888;
assign w12106 = pi2972 & ~pi3111;
assign w12107 = ~w7684 & ~w11271;
assign w12108 = pi2791 & ~w6463;
assign w12109 = w15450 & ~w1466;
assign w12110 = ~pi3288 & w9781;
assign w12111 = ~pi1024 & w3106;
assign w12112 = pi2267 & ~w9414;
assign w12113 = ~pi2280 & w13065;
assign w12114 = ~w4522 & w5763;
assign w12115 = pi2005 & ~w9414;
assign w12116 = pi0515 & pi1185;
assign w12117 = ~w7892 & ~w9434;
assign w12118 = ~pi2645 & w15122;
assign w12119 = ~pi3295 & w6072;
assign w12120 = pi2800 & ~w6463;
assign w12121 = pi2530 & w15191;
assign w12122 = ~w11728 & ~w13180;
assign w12123 = w3203 & ~w4043;
assign w12124 = ~pi3313 & w6448;
assign w12125 = pi1463 & ~w7090;
assign w12126 = ~w17286 & w16618;
assign w12127 = ~w7320 & ~w7436;
assign w12128 = pi1234 & w13142;
assign w12129 = ~pi2161 & w13065;
assign w12130 = ~w17665 & ~w3181;
assign w12131 = ~w16250 & w17242;
assign w12132 = w13509 & w1411;
assign w12133 = pi3151 & w9520;
assign w12134 = ~w502 & ~w6996;
assign w12135 = w13509 & w18360;
assign w12136 = ~w12921 & ~w8990;
assign w12137 = ~w6615 & w10639;
assign w12138 = ~w1716 & ~w8702;
assign w12139 = (pi0345 & w6195) | (pi0345 & w8394) | (w6195 & w8394);
assign w12140 = w16575 & w14793;
assign w12141 = w6785 & ~w17513;
assign w12142 = ~w10541 & ~w1462;
assign w12143 = ~w16575 & w17052;
assign w12144 = pi1438 & ~w6448;
assign w12145 = ~w65 & ~w1973;
assign w12146 = pi2691 & ~w15235;
assign w12147 = ~w4040 & ~w16074;
assign w12148 = ~pi0777 & w6200;
assign w12149 = pi1855 & ~w653;
assign w12150 = (~w4084 & ~w6920) | (~w4084 & w2959) | (~w6920 & w2959);
assign w12151 = ~w746 & w15424;
assign w12152 = pi3159 & w4256;
assign w12153 = pi0022 & ~w14148;
assign w12154 = ~pi0266 & ~w18262;
assign w12155 = ~pi0557 & w11739;
assign w12156 = ~w174 & ~w18234;
assign w12157 = pi2858 & w14148;
assign w12158 = (pi0692 & ~w13509) | (pi0692 & w10096) | (~w13509 & w10096);
assign w12159 = ~pi2828 & w15122;
assign w12160 = ~w10047 & ~w9557;
assign w12161 = ~pi0079 & ~pi1811;
assign w12162 = ~w14228 & pi0632;
assign w12163 = pi3168 & w8829;
assign w12164 = ~w9053 & ~w10329;
assign w12165 = pi2415 & ~w3223;
assign w12166 = (~w9205 & ~w10533) | (~w9205 & w11) | (~w10533 & w11);
assign w12167 = ~pi3290 & w6072;
assign w12168 = ~w1391 & ~pi0974;
assign w12169 = ~pi1257 & pi1376;
assign w12170 = ~w13794 & ~w12071;
assign w12171 = ~w17248 & pi0886;
assign w12172 = ~w7181 & ~w18438;
assign w12173 = ~pi0080 & w3584;
assign w12174 = (w11360 & w10646) | (w11360 & w3870) | (w10646 & w3870);
assign w12175 = ~w17635 & ~w2654;
assign w12176 = ~w18313 & ~w16194;
assign w12177 = ~w993 & ~w1532;
assign w12178 = ~w555 & w18132;
assign w12179 = ~w10528 & ~w4860;
assign w12180 = pi0069 & w922;
assign w12181 = w13509 & w11967;
assign w12182 = ~pi3314 & w6072;
assign w12183 = ~pi3158 & w12427;
assign w12184 = ~w4851 & ~w6758;
assign w12185 = ~w3817 & w11103;
assign w12186 = w17562 & pi1826;
assign w12187 = ~w8605 & w17600;
assign w12188 = ~w9087 & ~w5107;
assign w12189 = ~w8936 & ~w13816;
assign w12190 = pi1747 & ~w6463;
assign w12191 = w12483 & w650;
assign w12192 = w6857 & w8507;
assign w12193 = ~w10530 & w1033;
assign w12194 = ~pi1941 & w7455;
assign w12195 = ~w1962 & pi0647;
assign w12196 = pi1324 & pi1345;
assign w12197 = w134 & w3106;
assign w12198 = pi1653 & ~w6072;
assign w12199 = ~w662 & ~w18018;
assign w12200 = (pi0347 & w6195) | (pi0347 & w13268) | (w6195 & w13268);
assign w12201 = ~w8588 & w14524;
assign w12202 = pi1978 & ~w6463;
assign w12203 = pi2930 & ~w15122;
assign w12204 = ~w17089 & ~w9682;
assign w12205 = pi2947 & w14417;
assign w12206 = ~pi3514 & pi3515;
assign w12207 = (pi0653 & ~w13509) | (pi0653 & w16973) | (~w13509 & w16973);
assign w12208 = ~w16271 & w1183;
assign w12209 = w12051 & w10019;
assign w12210 = ~pi3162 & w14753;
assign w12211 = w6649 & ~w2000;
assign w12212 = pi2294 & pi2463;
assign w12213 = ~w4483 & ~w7295;
assign w12214 = pi2153 & ~w11671;
assign w12215 = (pi0774 & ~w13509) | (pi0774 & w10348) | (~w13509 & w10348);
assign w12216 = pi0485 & pi1134;
assign w12217 = pi2485 & w7965;
assign w12218 = ~w7077 & pi0902;
assign w12219 = ~w13231 & pi0559;
assign w12220 = w9440 & pi0155;
assign w12221 = ~w17259 & ~w13351;
assign w12222 = pi3163 & w13786;
assign w12223 = w11074 & w8120;
assign w12224 = ~pi2008 & w11688;
assign w12225 = (pi0740 & ~w13509) | (pi0740 & w13530) | (~w13509 & w13530);
assign w12226 = (pi1895 & w2014) | (pi1895 & w12003) | (w2014 & w12003);
assign w12227 = w13569 & w5453;
assign w12228 = ~w11583 & ~w6028;
assign w12229 = w16575 & w6706;
assign w12230 = w5874 & w4374;
assign w12231 = pi1508 & ~w13753;
assign w12232 = ~w10078 & ~w18236;
assign w12233 = ~w3303 & ~w18478;
assign w12234 = ~pi2153 & w13065;
assign w12235 = ~pi3335 & w17935;
assign w12236 = ~pi0448 & w17173;
assign w12237 = ~w4085 & ~w3965;
assign w12238 = pi1324 & w458;
assign w12239 = w6056 & w9786;
assign w12240 = ~pi2437 & w5075;
assign w12241 = ~pi3354 & w17935;
assign w12242 = ~w4128 & ~w12653;
assign w12243 = ~pi3103 & w261;
assign w12244 = w8337 & pi3280;
assign w12245 = ~w1010 & ~w11158;
assign w12246 = w7307 & w16356;
assign w12247 = ~pi3093 & w226;
assign w12248 = w13509 & w15194;
assign w12249 = ~w14804 & ~w5143;
assign w12250 = (~pi0291 & ~w6857) | (~pi0291 & w7317) | (~w6857 & w7317);
assign w12251 = pi1520 & w13753;
assign w12252 = w13509 & w6182;
assign w12253 = w16506 & ~w3430;
assign w12254 = (pi0799 & ~w13509) | (pi0799 & w8108) | (~w13509 & w8108);
assign w12255 = w5189 & ~w4043;
assign w12256 = (pi0640 & ~w13509) | (pi0640 & w3591) | (~w13509 & w3591);
assign w12257 = ~pi1927 & w9340;
assign w12258 = ~w8096 & ~w13012;
assign w12259 = ~pi3170 & w14753;
assign w12260 = w14109 & pi0446;
assign w12261 = ~w17701 & ~w5546;
assign w12262 = w13509 & w15679;
assign w12263 = ~w8674 & ~w1357;
assign w12264 = ~w12139 & ~w10192;
assign w12265 = ~pi1709 & w8341;
assign w12266 = w1815 & w3600;
assign w12267 = pi3134 & w619;
assign w12268 = ~w11359 & ~w6383;
assign w12269 = ~w7844 & pi0594;
assign w12270 = ~w13515 & ~w8406;
assign w12271 = (pi0865 & ~w13509) | (pi0865 & w4736) | (~w13509 & w4736);
assign w12272 = ~w1437 & ~w7624;
assign w12273 = w14334 & w10701;
assign w12274 = pi1790 & ~w9520;
assign w12275 = pi0142 & w5274;
assign w12276 = w13428 & w9130;
assign w12277 = w12606 & w12839;
assign w12278 = w8789 & ~pi0460;
assign w12279 = ~w3203 & pi1088;
assign w12280 = pi1550 & w13753;
assign w12281 = w13318 & pi0064;
assign w12282 = ~w12975 & w13555;
assign w12283 = w10818 & ~w7944;
assign w12284 = w9277 & w12676;
assign w12285 = pi1341 & w5274;
assign w12286 = ~w16987 & w2874;
assign w12287 = ~w6098 & ~w10423;
assign w12288 = pi1431 & ~w13753;
assign w12289 = w13509 & w106;
assign w12290 = (w18569 & ~w11247) | (w18569 & w534) | (~w11247 & w534);
assign w12291 = ~pi3021 & ~pi3207;
assign w12292 = ~pi3146 & w11701;
assign w12293 = ~pi0632 & w14641;
assign w12294 = pi0268 & w5274;
assign w12295 = w13509 & w17787;
assign w12296 = w5511 & w13047;
assign w12297 = ~w2641 & ~w15411;
assign w12298 = pi2384 & ~w7858;
assign w12299 = ~pi0447 & w17173;
assign w12300 = w1391 & ~w17210;
assign w12301 = w14782 & w14460;
assign w12302 = ~w16575 & w10189;
assign w12303 = ~pi0618 & w14641;
assign w12304 = ~w1391 & pi0915;
assign w12305 = w3243 & pi0317;
assign w12306 = ~w5658 & ~w1735;
assign w12307 = ~w5247 & ~w16470;
assign w12308 = (pi1810 & w5453) | (pi1810 & w15202) | (w5453 & w15202);
assign w12309 = ~w5560 & w5621;
assign w12310 = ~w5560 & w15263;
assign w12311 = pi2894 & ~w5274;
assign w12312 = w726 & pi0269;
assign w12313 = ~pi0880 & w1126;
assign w12314 = ~pi2072 & w17439;
assign w12315 = pi0254 & w5113;
assign w12316 = ~w10059 & ~w10870;
assign w12317 = ~w3054 & w15634;
assign w12318 = (w16679 & w15009) | (w16679 & w1249) | (w15009 & w1249);
assign w12319 = w7799 & w557;
assign w12320 = pi1586 & w13753;
assign w12321 = pi2381 & ~w15883;
assign w12322 = ~pi2263 & w13065;
assign w12323 = ~pi3354 & w18259;
assign w12324 = w17248 & ~w305;
assign w12325 = ~w14560 & pi0215;
assign w12326 = ~pi1962 & w11313;
assign w12327 = (pi0994 & ~w13509) | (pi0994 & w10237) | (~w13509 & w10237);
assign w12328 = ~w6697 & pi1110;
assign w12329 = (~pi2989 & ~w325) | (~pi2989 & w1596) | (~w325 & w1596);
assign w12330 = ~w15291 & ~w2571;
assign w12331 = ~pi2441 & w8617;
assign w12332 = pi1364 & w17382;
assign w12333 = ~pi2200 & w9340;
assign w12334 = ~pi0674 & w12197;
assign w12335 = w16506 & pi2952;
assign w12336 = ~w12301 & w14027;
assign w12337 = ~pi2253 & w12941;
assign w12338 = ~w14267 & ~w2886;
assign w12339 = ~w3044 & ~w10827;
assign w12340 = ~w17665 & ~w9564;
assign w12341 = pi2762 & w14148;
assign w12342 = pi3132 & w619;
assign w12343 = pi0047 & ~w14148;
assign w12344 = w6009 & ~w7177;
assign w12345 = pi2306 & ~w4420;
assign w12346 = ~pi3145 & w3982;
assign w12347 = pi1962 & ~w15271;
assign w12348 = ~w4827 & ~w4685;
assign w12349 = ~pi3154 & w3805;
assign w12350 = ~w15122 & ~pi2855;
assign w12351 = ~pi3103 & w9504;
assign w12352 = ~pi0762 & w6200;
assign w12353 = w13509 & w14299;
assign w12354 = w4800 & w3667;
assign w12355 = pi1799 & ~w10389;
assign w12356 = ~pi2041 & w13204;
assign w12357 = ~w14082 & ~w6917;
assign w12358 = ~w4120 & w17698;
assign w12359 = ~w6696 & w17229;
assign w12360 = ~w14741 & ~w10125;
assign w12361 = ~w8128 & ~w267;
assign w12362 = ~w6052 & w5393;
assign w12363 = ~pi0650 & w3791;
assign w12364 = ~pi3128 & w3555;
assign w12365 = pi0081 & pi1318;
assign w12366 = pi1645 & ~w6448;
assign w12367 = ~w25 & ~w17601;
assign w12368 = (pi0304 & ~w325) | (pi0304 & w4033) | (~w325 & w4033);
assign w12369 = w6649 & ~w13438;
assign w12370 = pi1666 & w1924;
assign w12371 = w12281 & pi0051;
assign w12372 = pi1141 & ~w11020;
assign w12373 = ~w16749 & w7628;
assign w12374 = w8291 & w11022;
assign w12375 = pi1632 & ~w6448;
assign w12376 = w384 & w5191;
assign w12377 = pi1278 & pi1345;
assign w12378 = pi2767 & w14148;
assign w12379 = ~w8179 & ~w1787;
assign w12380 = w11383 & w3403;
assign w12381 = ~w7234 & ~w13158;
assign w12382 = ~w7256 & ~w15160;
assign w12383 = ~pi0594 & w12825;
assign w12384 = w13509 & w12811;
assign w12385 = ~w3054 & w2223;
assign w12386 = w4181 & w16266;
assign w12387 = w4931 & pi0268;
assign w12388 = (pi0551 & ~w13509) | (pi0551 & w17985) | (~w13509 & w17985);
assign w12389 = ~w13300 & ~w15215;
assign w12390 = ~w1591 & ~w12111;
assign w12391 = w17679 & ~w1229;
assign w12392 = (pi1269 & ~w5437) | (pi1269 & w4107) | (~w5437 & w4107);
assign w12393 = ~pi3355 & w14918;
assign w12394 = ~pi3062 & w261;
assign w12395 = ~pi0129 & pi3377;
assign w12396 = pi1621 & w13753;
assign w12397 = ~pi3130 & pi2993;
assign w12398 = w13207 & w6714;
assign w12399 = ~w14950 & ~w10777;
assign w12400 = ~pi2979 & ~w6147;
assign w12401 = ~w6688 & ~w236;
assign w12402 = ~w1391 & pi0762;
assign w12403 = pi1418 & ~w13753;
assign w12404 = ~w10161 & ~w15919;
assign w12405 = ~pi2664 & w17213;
assign w12406 = ~pi2104 & w12724;
assign w12407 = pi0412 & w17173;
assign w12408 = w16148 & w6440;
assign w12409 = w13509 & w7077;
assign w12410 = ~w4822 & ~w14300;
assign w12411 = ~pi2967 & pi3028;
assign w12412 = ~w17124 & w11165;
assign w12413 = ~w17578 & ~w7384;
assign w12414 = ~pi2967 & pi3032;
assign w12415 = ~w1368 & ~pi0454;
assign w12416 = pi3136 & w6853;
assign w12417 = w15450 & pi1164;
assign w12418 = pi2205 & ~w3223;
assign w12419 = ~w10819 & ~w18032;
assign w12420 = ~w12460 & w10822;
assign w12421 = ~w7887 & ~w11635;
assign w12422 = ~pi0301 & ~w1698;
assign w12423 = ~w8344 & ~w12773;
assign w12424 = pi1858 & w11182;
assign w12425 = ~w17187 & ~w7954;
assign w12426 = ~pi3160 & ~pi3166;
assign w12427 = ~w4020 & w10299;
assign w12428 = ~w11582 & w4941;
assign w12429 = ~w17248 & pi0895;
assign w12430 = ~w9894 & ~w11164;
assign w12431 = ~w3243 & ~pi0322;
assign w12432 = ~w3243 & pi0323;
assign w12433 = ~w559 & w11539;
assign w12434 = ~w1391 & pi0778;
assign w12435 = pi1379 & w9653;
assign w12436 = w4009 & ~w8795;
assign w12437 = ~w12599 & w9148;
assign w12438 = pi2734 & ~w261;
assign w12439 = pi2766 & w605;
assign w12440 = (pi1116 & ~w13509) | (pi1116 & w5626) | (~w13509 & w5626);
assign w12441 = (pi0721 & ~w13509) | (pi0721 & w15598) | (~w13509 & w15598);
assign w12442 = pi2914 & w6045;
assign w12443 = ~w12458 & w1326;
assign w12444 = ~w16278 & pi0707;
assign w12445 = w13509 & w972;
assign w12446 = ~w2137 & w10810;
assign w12447 = w12786 & w8993;
assign w12448 = w1127 & ~w2434;
assign w12449 = w13231 & ~w6647;
assign w12450 = (pi0842 & ~w13509) | (pi0842 & w5200) | (~w13509 & w5200);
assign w12451 = ~w7077 & pi0811;
assign w12452 = w6649 & ~w16032;
assign w12453 = ~w10152 & ~w16520;
assign w12454 = (pi0660 & ~w13509) | (pi0660 & w9410) | (~w13509 & w9410);
assign w12455 = w10189 & ~pi0465;
assign w12456 = ~w3928 & ~w2472;
assign w12457 = ~w2545 & ~w3527;
assign w12458 = pi2978 & w9545;
assign w12459 = ~w4278 & ~w16539;
assign w12460 = ~w12775 & ~w2445;
assign w12461 = pi0007 & ~w3748;
assign w12462 = pi1254 & ~w11655;
assign w12463 = ~pi3033 & ~pi3155;
assign w12464 = ~pi3349 & w6448;
assign w12465 = pi0088 & w3748;
assign w12466 = w3813 & w11588;
assign w12467 = w6697 & ~w15173;
assign w12468 = ~w17155 & ~w12275;
assign w12469 = ~pi3086 & w226;
assign w12470 = pi0271 & w5274;
assign w12471 = w922 & ~w759;
assign w12472 = ~w5764 & ~w13188;
assign w12473 = w15122 & ~pi2512;
assign w12474 = ~pi0773 & w6200;
assign w12475 = pi2846 & w16699;
assign w12476 = w5396 & w4768;
assign w12477 = ~pi3045 & w3555;
assign w12478 = ~pi1375 & pi3224;
assign w12479 = ~w16953 & ~w7375;
assign w12480 = ~w17795 & w15668;
assign w12481 = ~pi2106 & w12724;
assign w12482 = w13509 & w9315;
assign w12483 = w18351 & w1778;
assign w12484 = pi1665 & w1924;
assign w12485 = ~pi2687 & w13343;
assign w12486 = (~w6843 & ~w1007) | (~w6843 & w9217) | (~w1007 & w9217);
assign w12487 = ~w14444 & ~w14176;
assign w12488 = ~w2341 & pi1059;
assign w12489 = ~w644 & ~w10775;
assign w12490 = w6649 & ~w5056;
assign w12491 = ~pi0321 & ~pi3225;
assign w12492 = ~pi2202 & w13204;
assign w12493 = pi2858 & w15191;
assign w12494 = w13509 & w2054;
assign w12495 = ~w6535 & ~w12259;
assign w12496 = ~w6215 & ~w17934;
assign w12497 = pi3166 & w8088;
assign w12498 = ~w4676 & ~w1373;
assign w12499 = ~pi0882 & w1126;
assign w12500 = pi2228 & ~w15271;
assign w12501 = ~w18577 & ~w6974;
assign w12502 = ~w8177 & ~w13010;
assign w12503 = ~w6697 & pi0658;
assign w12504 = w14648 & ~pi2608;
assign w12505 = ~pi1811 & pi2465;
assign w12506 = ~pi0967 & w3106;
assign w12507 = pi2966 & pi2755;
assign w12508 = ~w8188 & ~w3862;
assign w12509 = pi3147 & w8829;
assign w12510 = ~w11778 & ~w11718;
assign w12511 = pi1605 & ~w18259;
assign w12512 = ~w13657 & ~w275;
assign w12513 = ~w11494 & ~w5039;
assign w12514 = ~w13919 & w2672;
assign w12515 = ~w5489 & ~w14892;
assign w12516 = ~w13689 & ~w14463;
assign w12517 = ~w15469 & ~w3606;
assign w12518 = ~w5078 & w14137;
assign w12519 = (pi0646 & ~w13509) | (pi0646 & w8338) | (~w13509 & w8338);
assign w12520 = ~w3654 & ~w3944;
assign w12521 = ~w11399 & w4539;
assign w12522 = ~w3479 & ~w1048;
assign w12523 = w13509 & w13410;
assign w12524 = ~pi2943 & ~pi3123;
assign w12525 = pi3184 & ~pi3239;
assign w12526 = ~pi0597 & w12825;
assign w12527 = ~w18589 & ~w7730;
assign w12528 = ~w7728 & ~w452;
assign w12529 = ~w8141 & ~w15489;
assign w12530 = ~w7526 & ~w5324;
assign w12531 = ~w15383 & ~w16236;
assign w12532 = ~pi3100 & w3555;
assign w12533 = ~pi2755 & ~w5274;
assign w12534 = pi2159 & ~w17683;
assign w12535 = w5383 & w17562;
assign w12536 = w13509 & w7254;
assign w12537 = w13509 & w18159;
assign w12538 = ~pi3054 & w261;
assign w12539 = ~w352 & w8975;
assign w12540 = w6365 & w3078;
assign w12541 = ~w8925 & ~w689;
assign w12542 = ~w14344 & ~w18519;
assign w12543 = ~w10087 & ~w6575;
assign w12544 = pi2143 & ~w15883;
assign w12545 = ~pi3135 & w17669;
assign w12546 = w13961 & w14963;
assign w12547 = ~w4963 & w17047;
assign w12548 = ~w2341 & pi0847;
assign w12549 = ~w14797 & ~w13874;
assign w12550 = (~pi0083 & ~w18005) | (~pi0083 & w16779) | (~w18005 & w16779);
assign w12551 = ~w4862 & ~w10597;
assign w12552 = w12848 & w12749;
assign w12553 = w13509 & w1971;
assign w12554 = w384 & w11656;
assign w12555 = w12040 & ~w15296;
assign w12556 = ~pi2421 & w5075;
assign w12557 = ~w15713 & ~w8283;
assign w12558 = w1611 & w11618;
assign w12559 = pi1991 & ~w14833;
assign w12560 = w7307 & w12813;
assign w12561 = pi2282 & ~w11671;
assign w12562 = ~w2014 & w9398;
assign w12563 = ~w6901 & ~w12241;
assign w12564 = pi2867 & w14148;
assign w12565 = pi3020 & w3384;
assign w12566 = w5437 & w4168;
assign w12567 = ~pi2688 & w13343;
assign w12568 = pi1413 & ~w6072;
assign w12569 = ~w13150 & ~w17241;
assign w12570 = ~pi3295 & w6448;
assign w12571 = (w17562 & ~w384) | (w17562 & w14453) | (~w384 & w14453);
assign w12572 = ~pi2029 & w7455;
assign w12573 = pi0032 & ~w14148;
assign w12574 = ~w13387 & ~w11683;
assign w12575 = ~w16506 & pi1147;
assign w12576 = w5453 & pi2787;
assign w12577 = pi2532 & w15191;
assign w12578 = pi2083 & ~w17683;
assign w12579 = ~pi3160 & ~pi3168;
assign w12580 = (~pi0248 & ~w325) | (~pi0248 & w2360) | (~w325 & w2360);
assign w12581 = (pi0249 & ~w325) | (pi0249 & w2361) | (~w325 & w2361);
assign w12582 = w1391 & ~w305;
assign w12583 = pi3361 & pi3362;
assign w12584 = ~w6929 & ~w16902;
assign w12585 = w14094 & ~w2225;
assign w12586 = ~w564 & ~w16081;
assign w12587 = ~w2961 & ~w8805;
assign w12588 = ~pi2099 & w12724;
assign w12589 = ~w15288 & ~w2334;
assign w12590 = w6697 & ~w11978;
assign w12591 = w5437 & w15779;
assign w12592 = ~w1391 & pi1189;
assign w12593 = ~w11698 & ~w1678;
assign w12594 = pi2062 & ~w4508;
assign w12595 = ~w15122 & ~pi2929;
assign w12596 = ~pi1121 & w1126;
assign w12597 = ~pi3159 & w8515;
assign w12598 = ~pi0266 & pi3217;
assign w12599 = pi0448 & w4643;
assign w12600 = ~w12046 & ~w565;
assign w12601 = ~pi0759 & w6200;
assign w12602 = ~w13744 & ~w16390;
assign w12603 = pi1732 & w1924;
assign w12604 = ~pi3433 & w15036;
assign w12605 = ~pi2274 & w8617;
assign w12606 = ~w4027 & ~w2484;
assign w12607 = ~w6431 & ~w16037;
assign w12608 = ~pi1961 & w11688;
assign w12609 = ~pi0586 & w795;
assign w12610 = w4108 & w5433;
assign w12611 = ~w13922 & ~w8173;
assign w12612 = ~w3701 & ~w13640;
assign w12613 = ~w2341 & pi0827;
assign w12614 = ~w3000 & ~pi2692;
assign w12615 = pi2940 & w6045;
assign w12616 = ~pi1215 & ~pi3220;
assign w12617 = ~pi3157 & w3982;
assign w12618 = pi2169 & ~w15271;
assign w12619 = ~w5561 & ~w8639;
assign w12620 = w10189 & pi0387;
assign w12621 = ~w5453 & ~pi1765;
assign w12622 = ~w10820 & ~w16783;
assign w12623 = (pi0004 & ~w1766) | (pi0004 & w5831) | (~w1766 & w5831);
assign w12624 = ~pi3165 & w3982;
assign w12625 = pi2280 & ~w11671;
assign w12626 = w8508 & w11564;
assign w12627 = pi1336 & w5274;
assign w12628 = w9178 & w15144;
assign w12629 = ~w4350 & ~w13619;
assign w12630 = ~w15122 & ~pi2876;
assign w12631 = ~w9 & ~pi1687;
assign w12632 = ~w2678 & w8408;
assign w12633 = ~w9887 & ~w11856;
assign w12634 = w7844 & ~w1236;
assign w12635 = ~w16575 & w1655;
assign w12636 = ~pi3153 & w17669;
assign w12637 = ~w2731 & ~w10462;
assign w12638 = w14782 & w16836;
assign w12639 = ~w2671 & ~w3436;
assign w12640 = ~pi0146 & w9966;
assign w12641 = pi1396 & ~w6853;
assign w12642 = w14560 & pi0351;
assign w12643 = ~w8588 & w11735;
assign w12644 = ~w15196 & ~w769;
assign w12645 = ~w12183 & ~w14813;
assign w12646 = ~w7006 & w8305;
assign w12647 = ~w2288 & ~w12006;
assign w12648 = (w2460 & ~w7799) | (w2460 & w16018) | (~w7799 & w16018);
assign w12649 = w13509 & w3314;
assign w12650 = ~w6193 & ~w8169;
assign w12651 = ~pi3018 & pi3020;
assign w12652 = ~pi3347 & w7090;
assign w12653 = ~pi2658 & w17213;
assign w12654 = (pi0568 & ~w13509) | (pi0568 & w1923) | (~w13509 & w1923);
assign w12655 = w2359 & w17944;
assign w12656 = ~w7557 & ~w9140;
assign w12657 = w11334 & w6469;
assign w12658 = pi1451 & ~w13753;
assign w12659 = ~pi3313 & w16922;
assign w12660 = ~pi2962 & ~w8003;
assign w12661 = pi2101 & ~w4420;
assign w12662 = (pi0803 & ~w13509) | (pi0803 & w13588) | (~w13509 & w13588);
assign w12663 = (pi1107 & ~w13509) | (pi1107 & w11348) | (~w13509 & w11348);
assign w12664 = pi3151 & w3987;
assign w12665 = (pi1784 & w7215) | (pi1784 & w14014) | (w7215 & w14014);
assign w12666 = (pi0639 & ~w13509) | (pi0639 & w18457) | (~w13509 & w18457);
assign w12667 = pi1845 & w7799;
assign w12668 = w9414 & w17115;
assign w12669 = pi2326 & ~w18123;
assign w12670 = w10804 & w16159;
assign w12671 = (~pi0283 & ~w6857) | (~pi0283 & w3143) | (~w6857 & w3143);
assign w12672 = ~pi0310 & ~w18262;
assign w12673 = ~w9159 & ~w3792;
assign w12674 = ~pi3150 & w4310;
assign w12675 = ~pi3131 & w11132;
assign w12676 = ~w9470 & ~w10432;
assign w12677 = w7799 & w6085;
assign w12678 = (~w6499 & w1225) | (~w6499 & w5426) | (w1225 & w5426);
assign w12679 = pi2938 & ~w13367;
assign w12680 = ~w1755 & ~w4541;
assign w12681 = ~w10065 & ~w16850;
assign w12682 = ~w3000 & ~pi2788;
assign w12683 = pi1153 & ~pi3194;
assign w12684 = ~w13792 & ~w9738;
assign w12685 = ~w11310 & ~w16320;
assign w12686 = ~pi2949 & w6045;
assign w12687 = ~pi2898 & w15122;
assign w12688 = w15113 & w9594;
assign w12689 = ~pi2996 & ~pi2997;
assign w12690 = (pi0682 & ~w13509) | (pi0682 & w12961) | (~w13509 & w12961);
assign w12691 = ~w10121 & ~w2572;
assign w12692 = (pi0758 & ~w13509) | (pi0758 & w8315) | (~w13509 & w8315);
assign w12693 = ~w7395 & ~w18199;
assign w12694 = ~w2289 & ~w8773;
assign w12695 = ~w18215 & ~pi0896;
assign w12696 = w13509 & w15370;
assign w12697 = pi3132 & w3987;
assign w12698 = ~pi2403 & w12755;
assign w12699 = ~pi3145 & w3805;
assign w12700 = pi2727 & ~w261;
assign w12701 = w8337 & pi3307;
assign w12702 = ~w9729 & ~w6290;
assign w12703 = w1225 & w3003;
assign w12704 = ~w15007 & ~w14805;
assign w12705 = ~w6221 & ~w11767;
assign w12706 = (pi0909 & ~w13509) | (pi0909 & w8002) | (~w13509 & w8002);
assign w12707 = ~w12205 & w1326;
assign w12708 = ~w3099 & ~w11088;
assign w12709 = ~w5253 & ~w11411;
assign w12710 = ~pi2448 & w9340;
assign w12711 = pi1532 & ~w14918;
assign w12712 = pi1269 & pi1310;
assign w12713 = ~w17864 & ~w9599;
assign w12714 = w2341 & w1217;
assign w12715 = pi3158 & w5457;
assign w12716 = ~w14648 & ~pi2621;
assign w12717 = w11383 & w13464;
assign w12718 = ~w8059 & ~w12353;
assign w12719 = ~w11887 & ~w16264;
assign w12720 = w934 & pi0438;
assign w12721 = w13509 & w3276;
assign w12722 = ~w17140 & w12340;
assign w12723 = w6857 & w4016;
assign w12724 = w13807 & w14138;
assign w12725 = ~w10791 & ~w59;
assign w12726 = pi2314 & ~w18123;
assign w12727 = ~w7077 & pi0805;
assign w12728 = ~w1721 & ~w15343;
assign w12729 = ~pi1407 & ~pi2913;
assign w12730 = ~w626 & ~w2202;
assign w12731 = pi2369 & ~w17683;
assign w12732 = ~w17843 & ~w1056;
assign w12733 = ~w1368 & ~pi0457;
assign w12734 = pi0176 & pi0201;
assign w12735 = ~w16691 & ~w16061;
assign w12736 = ~pi0616 & w14641;
assign w12737 = pi0141 & w5274;
assign w12738 = w2229 & w9210;
assign w12739 = w7498 & w13876;
assign w12740 = ~w17676 & ~w1527;
assign w12741 = ~pi0943 & w12197;
assign w12742 = ~w5055 & w9041;
assign w12743 = ~pi3087 & w226;
assign w12744 = pi2803 & ~w11406;
assign w12745 = pi3159 & w3987;
assign w12746 = ~w3243 & ~pi0335;
assign w12747 = pi2002 & ~w9414;
assign w12748 = ~w18556 & ~w9294;
assign w12749 = ~w9829 & ~w14104;
assign w12750 = pi1639 & ~w13753;
assign w12751 = ~w15030 & ~w11032;
assign w12752 = ~pi1769 & pi3157;
assign w12753 = w934 & pi0418;
assign w12754 = ~pi2557 & pi2920;
assign w12755 = w14138 & w3556;
assign w12756 = ~w2725 & pi0800;
assign w12757 = ~w5845 & ~w1877;
assign w12758 = ~pi0714 & w3106;
assign w12759 = ~w5285 & ~w5608;
assign w12760 = w17419 & w13002;
assign w12761 = w10818 & ~w6828;
assign w12762 = w9946 & w1100;
assign w12763 = ~pi0553 & w11739;
assign w12764 = ~pi1966 & ~w1097;
assign w12765 = pi2934 & ~pi3208;
assign w12766 = ~pi0795 & w543;
assign w12767 = pi0255 & w5113;
assign w12768 = pi1541 & ~w17935;
assign w12769 = ~pi3295 & w18259;
assign w12770 = w9440 & pi0187;
assign w12771 = ~w3059 & ~w18545;
assign w12772 = ~w7715 & ~w12972;
assign w12773 = ~pi0960 & w12197;
assign w12774 = ~w5029 & ~w3837;
assign w12775 = ~pi1161 & w1054;
assign w12776 = ~w5739 & ~w6839;
assign w12777 = ~w17854 & ~w17037;
assign w12778 = ~w11263 & ~w8834;
assign w12779 = pi0178 & w5274;
assign w12780 = pi2937 & ~w3987;
assign w12781 = ~w6785 & pi1050;
assign w12782 = w9440 & pi0199;
assign w12783 = pi3074 & ~w16502;
assign w12784 = ~pi2967 & ~pi3113;
assign w12785 = (pi0904 & ~w13509) | (pi0904 & w11527) | (~w13509 & w11527);
assign w12786 = w2742 & ~w2779;
assign w12787 = ~pi3131 & w3805;
assign w12788 = pi2499 & ~w5274;
assign w12789 = pi2310 & ~w9414;
assign w12790 = ~w11290 & ~w10790;
assign w12791 = ~w6574 & w11585;
assign w12792 = w5437 & w12087;
assign w12793 = (pi0659 & ~w13509) | (pi0659 & w15085) | (~w13509 & w15085);
assign w12794 = ~w14544 & ~w14564;
assign w12795 = ~pi2324 & w8617;
assign w12796 = ~pi3159 & w17993;
assign w12797 = ~w15954 & ~w7805;
assign w12798 = ~pi3147 & w15839;
assign w12799 = ~pi2175 & w5384;
assign w12800 = ~w15744 & ~w11295;
assign w12801 = ~w4794 & ~w12016;
assign w12802 = w5437 & w6549;
assign w12803 = (pi0641 & ~w13509) | (pi0641 & w7544) | (~w13509 & w7544);
assign w12804 = pi1861 & ~w15036;
assign w12805 = w2248 & w17796;
assign w12806 = ~pi0904 & w795;
assign w12807 = ~w2193 & ~w13977;
assign w12808 = w11031 & w8070;
assign w12809 = ~w709 & pi1295;
assign w12810 = w6649 & ~w830;
assign w12811 = w15808 & ~w1340;
assign w12812 = w13509 & w5040;
assign w12813 = ~w3000 & ~pi2773;
assign w12814 = w1509 & w15723;
assign w12815 = ~w7611 & ~w8183;
assign w12816 = w14524 & w2753;
assign w12817 = w8098 & w12535;
assign w12818 = ~w11169 & ~w1115;
assign w12819 = ~pi3350 & w18259;
assign w12820 = ~w18492 & ~w14778;
assign w12821 = ~pi2684 & w13343;
assign w12822 = w13592 & w13566;
assign w12823 = w4476 & w16232;
assign w12824 = ~w5453 & ~pi1767;
assign w12825 = ~w10087 & ~w10724;
assign w12826 = pi1402 & ~w13786;
assign w12827 = w3203 & ~w7020;
assign w12828 = (pi0567 & ~w13509) | (pi0567 & w1293) | (~w13509 & w1293);
assign w12829 = w16575 & w6293;
assign w12830 = w16575 & w6294;
assign w12831 = pi1892 & ~w15036;
assign w12832 = ~w15400 & ~w16446;
assign w12833 = ~pi2763 & w13343;
assign w12834 = ~pi1130 & pi1131;
assign w12835 = pi2937 & w13560;
assign w12836 = (pi0674 & ~w13509) | (pi0674 & w14789) | (~w13509 & w14789);
assign w12837 = (w15450 & w14073) | (w15450 & w10846) | (w14073 & w10846);
assign w12838 = w7201 & w6093;
assign w12839 = ~w2882 & ~w6075;
assign w12840 = ~pi2997 & pi2995;
assign w12841 = ~w1368 & ~pi0463;
assign w12842 = w3203 & ~w6922;
assign w12843 = ~pi3084 & w9504;
assign w12844 = ~pi0105 & w9284;
assign w12845 = pi0106 & w9284;
assign w12846 = ~pi1220 & pi3373;
assign w12847 = ~pi3132 & ~pi3160;
assign w12848 = w16067 & w4746;
assign w12849 = ~w1224 & ~w10126;
assign w12850 = w12832 & w4521;
assign w12851 = ~w8019 & ~w5499;
assign w12852 = ~pi3147 & w1843;
assign w12853 = (pi1092 & ~w13509) | (pi1092 & w430) | (~w13509 & w430);
assign w12854 = ~pi1698 & ~w11760;
assign w12855 = pi2792 & ~w11406;
assign w12856 = w4508 & w3515;
assign w12857 = pi0323 & pi3235;
assign w12858 = pi1965 & w15106;
assign w12859 = ~w15519 & ~w323;
assign w12860 = w1747 & w164;
assign w12861 = ~w6663 & ~w8945;
assign w12862 = w1368 & pi0393;
assign w12863 = ~w5805 & ~w10168;
assign w12864 = ~w6576 & ~w1783;
assign w12865 = ~w17833 & ~w4245;
assign w12866 = ~w15520 & ~w14888;
assign w12867 = w13509 & w11287;
assign w12868 = ~pi2967 & pi3125;
assign w12869 = ~w158 & w6897;
assign w12870 = (pi1060 & ~w13509) | (pi1060 & w12082) | (~w13509 & w12082);
assign w12871 = ~w7907 & ~w11150;
assign w12872 = pi2372 & ~w17683;
assign w12873 = ~pi2399 & w5384;
assign w12874 = ~w8105 & ~w8161;
assign w12875 = pi1592 & ~w16922;
assign w12876 = w17646 & w2753;
assign w12877 = pi1316 & pi1301;
assign w12878 = pi1559 & ~w13753;
assign w12879 = ~w2444 & ~w13367;
assign w12880 = ~pi1309 & ~w14094;
assign w12881 = pi2957 & w4492;
assign w12882 = w4508 & w17115;
assign w12883 = ~w8185 & ~w17352;
assign w12884 = pi3013 & ~w16502;
assign w12885 = ~w5912 & ~w12143;
assign w12886 = ~pi0919 & w17490;
assign w12887 = w1127 & ~w6012;
assign w12888 = w6785 & ~w12800;
assign w12889 = ~pi3114 & pi3164;
assign w12890 = pi1635 & ~w13753;
assign w12891 = w13509 & w12888;
assign w12892 = ~w6195 & w6479;
assign w12893 = ~w5668 & ~w4133;
assign w12894 = ~w16575 & w18452;
assign w12895 = w16575 & w18105;
assign w12896 = w13509 & w7270;
assign w12897 = pi2127 & ~w18123;
assign w12898 = ~pi3090 & w11406;
assign w12899 = ~w373 & ~w18439;
assign w12900 = pi2569 & ~w5274;
assign w12901 = ~pi3101 & w9504;
assign w12902 = w968 & ~pi0333;
assign w12903 = ~w13231 & pi0560;
assign w12904 = ~w6322 & ~w3385;
assign w12905 = ~w5981 & ~w8767;
assign w12906 = (w5517 & w2087) | (w5517 & w11319) | (w2087 & w11319);
assign w12907 = ~pi3055 & w6463;
assign w12908 = ~pi1022 & w9110;
assign w12909 = ~pi1188 & w9110;
assign w12910 = ~pi3134 & pi3207;
assign w12911 = ~w9142 & w12097;
assign w12912 = ~w13788 & ~w3518;
assign w12913 = w5867 & w55;
assign w12914 = pi1393 & ~w14918;
assign w12915 = pi0487 & pi0488;
assign w12916 = ~w9618 & ~w9765;
assign w12917 = w7703 & w3042;
assign w12918 = ~pi3428 & w15036;
assign w12919 = w5517 & w13078;
assign w12920 = w15122 & ~pi2631;
assign w12921 = w6857 & w5638;
assign w12922 = ~w1019 & w6434;
assign w12923 = ~w11863 & ~w14281;
assign w12924 = ~pi2946 & w6463;
assign w12925 = ~pi2994 & w7090;
assign w12926 = ~pi0886 & w1126;
assign w12927 = ~pi0786 & w543;
assign w12928 = pi3190 & w4899;
assign w12929 = ~w12002 & ~w11054;
assign w12930 = w13840 & pi0002;
assign w12931 = ~w17248 & ~pi0981;
assign w12932 = w11735 & w3515;
assign w12933 = w11383 & w3639;
assign w12934 = w9440 & pi0160;
assign w12935 = pi2075 & ~w17683;
assign w12936 = pi2191 & ~w11735;
assign w12937 = ~w17577 & w15877;
assign w12938 = pi1388 & ~w17935;
assign w12939 = pi0042 & ~w14148;
assign w12940 = ~pi2167 & w11313;
assign w12941 = w13807 & w2246;
assign w12942 = ~pi1234 & ~pi1258;
assign w12943 = ~w6195 & w13965;
assign w12944 = ~pi3058 & w9504;
assign w12945 = (pi1011 & ~w13509) | (pi1011 & w8699) | (~w13509 & w8699);
assign w12946 = ~pi1153 & ~w13509;
assign w12947 = pi1154 & ~w13509;
assign w12948 = ~w304 & ~w13926;
assign w12949 = ~w17835 & ~w4202;
assign w12950 = w6134 & w16784;
assign w12951 = ~w7844 & pi0593;
assign w12952 = pi1544 & ~w17935;
assign w12953 = w8658 & pi1783;
assign w12954 = ~pi3048 & w16815;
assign w12955 = w2742 & ~w7448;
assign w12956 = w14560 & pi0369;
assign w12957 = ~w9379 & ~w6709;
assign w12958 = ~w7772 & w5435;
assign w12959 = ~w13306 & ~w17224;
assign w12960 = ~w14954 & ~w8870;
assign w12961 = ~w12040 & pi0682;
assign w12962 = ~w374 & ~w13390;
assign w12963 = (pi1133 & ~w5437) | (pi1133 & w520) | (~w5437 & w520);
assign w12964 = ~pi3145 & w11132;
assign w12965 = w11383 & w9307;
assign w12966 = ~w5696 & ~w3887;
assign w12967 = ~w8434 & ~w9390;
assign w12968 = ~w4096 & ~w14841;
assign w12969 = pi2450 & ~w14524;
assign w12970 = pi1764 & ~w14951;
assign w12971 = ~pi3100 & w16815;
assign w12972 = pi2543 & w605;
assign w12973 = (~pi0051 & ~w5642) | (~pi0051 & w192) | (~w5642 & w192);
assign w12974 = ~w15935 & ~w4195;
assign w12975 = w7688 & w5382;
assign w12976 = pi2375 & ~w15883;
assign w12977 = ~w2014 & w10381;
assign w12978 = ~pi0998 & w795;
assign w12979 = w15122 & ~pi2653;
assign w12980 = ~pi3159 & w3982;
assign w12981 = w7703 & w12595;
assign w12982 = ~w14616 & ~w7949;
assign w12983 = w12868 & pi3034;
assign w12984 = pi1161 & ~pi0077;
assign w12985 = w8954 & w16513;
assign w12986 = ~pi3441 & w15036;
assign w12987 = pi1763 & pi3164;
assign w12988 = w13509 & w765;
assign w12989 = ~pi0288 & w4058;
assign w12990 = ~w16575 & w10652;
assign w12991 = w709 & pi1868;
assign w12992 = ~pi0176 & ~pi0201;
assign w12993 = pi1708 & ~w7946;
assign w12994 = ~w8247 & ~w7987;
assign w12995 = w11383 & w8017;
assign w12996 = pi1517 & ~w14918;
assign w12997 = ~w14228 & pi0615;
assign w12998 = ~w6782 & ~w9393;
assign w12999 = ~w6369 & ~w16675;
assign w13000 = ~w2895 & ~w3103;
assign w13001 = ~w14560 & pi0245;
assign w13002 = ~w11025 & ~w4001;
assign w13003 = (~pi0286 & ~w6857) | (~pi0286 & w5973) | (~w6857 & w5973);
assign w13004 = ~w13620 & w2613;
assign w13005 = ~w4113 & ~w5385;
assign w13006 = ~pi0661 & w12197;
assign w13007 = w14228 & ~w14465;
assign w13008 = (pi1042 & ~w13509) | (pi1042 & w9505) | (~w13509 & w9505);
assign w13009 = ~w3000 & ~pi2747;
assign w13010 = w13509 & w11908;
assign w13011 = ~pi2192 & w2151;
assign w13012 = ~pi0664 & w12197;
assign w13013 = w3223 & w3515;
assign w13014 = (pi0401 & w5560) | (pi0401 & w12072) | (w5560 & w12072);
assign w13015 = ~pi1953 & w11688;
assign w13016 = ~w1265 & ~w10897;
assign w13017 = ~pi2079 & w17439;
assign w13018 = w7799 & w7947;
assign w13019 = ~w4522 & w5944;
assign w13020 = ~w3316 & w12486;
assign w13021 = w13509 & w1947;
assign w13022 = ~w5945 & ~w1695;
assign w13023 = ~w1962 & pi0652;
assign w13024 = ~pi3086 & w6463;
assign w13025 = pi1312 & ~pi3362;
assign w13026 = ~w8652 & ~w981;
assign w13027 = pi2293 & ~w3555;
assign w13028 = ~w11670 & ~w15765;
assign w13029 = w5396 & pi0053;
assign w13030 = ~w15952 & w11810;
assign w13031 = w15808 & ~w6922;
assign w13032 = ~pi2392 & w8617;
assign w13033 = ~w3203 & pi0574;
assign w13034 = ~w15181 & ~w4419;
assign w13035 = ~w14593 & ~w2877;
assign w13036 = ~pi0142 & pi0191;
assign w13037 = ~pi3047 & w261;
assign w13038 = pi2657 & ~w15235;
assign w13039 = ~pi0677 & w12197;
assign w13040 = ~w7049 & ~w738;
assign w13041 = pi1575 & ~w13753;
assign w13042 = pi1239 & pi3223;
assign w13043 = w1962 & ~w1340;
assign w13044 = ~w5560 & w2728;
assign w13045 = ~w12993 & ~w7468;
assign w13046 = ~w10687 & ~w12124;
assign w13047 = w299 & w16299;
assign w13048 = ~w13959 & ~w1363;
assign w13049 = w13509 & w4663;
assign w13050 = ~pi2972 & pi3111;
assign w13051 = (pi1014 & ~w13509) | (pi1014 & w14866) | (~w13509 & w14866);
assign w13052 = ~w8440 & ~w2828;
assign w13053 = ~w5388 & ~w3173;
assign w13054 = ~pi3054 & w9504;
assign w13055 = w13509 & w18069;
assign w13056 = pi2660 & ~w15235;
assign w13057 = ~pi0505 & ~pi1345;
assign w13058 = ~w9924 & ~w12990;
assign w13059 = w3203 & ~w10947;
assign w13060 = pi2989 & ~w7212;
assign w13061 = ~w13304 & ~w13966;
assign w13062 = pi1819 & ~w653;
assign w13063 = ~pi1986 & ~w15450;
assign w13064 = w968 & ~pi0297;
assign w13065 = w3556 & w2246;
assign w13066 = w5189 & ~w17513;
assign w13067 = ~w7495 & ~w1642;
assign w13068 = pi1401 & ~w13786;
assign w13069 = ~w4644 & ~w14102;
assign w13070 = pi3184 & pi3239;
assign w13071 = ~pi1336 & pi1878;
assign w13072 = ~w13620 & w28;
assign w13073 = ~pi2957 & ~w4492;
assign w13074 = ~pi1714 & pi3155;
assign w13075 = pi1715 & ~pi3154;
assign w13076 = ~w14447 & ~w2416;
assign w13077 = ~w17141 & ~w17946;
assign w13078 = ~pi2967 & ~pi3076;
assign w13079 = ~pi3086 & w16815;
assign w13080 = ~pi3147 & w15048;
assign w13081 = ~w14560 & pi0233;
assign w13082 = w15907 & w4333;
assign w13083 = ~w14566 & ~w1024;
assign w13084 = ~w15505 & ~w12384;
assign w13085 = ~w484 & ~pi0491;
assign w13086 = pi2966 & pi2586;
assign w13087 = ~w16986 & ~w4871;
assign w13088 = ~w16983 & w5492;
assign w13089 = pi0495 & ~pi1142;
assign w13090 = pi1985 & w314;
assign w13091 = pi1529 & w13753;
assign w13092 = w14109 & pi0426;
assign w13093 = w13509 & w3460;
assign w13094 = ~w18347 & ~w8319;
assign w13095 = ~w5877 & ~w10685;
assign w13096 = (pi0886 & ~w13509) | (pi0886 & w12171) | (~w13509 & w12171);
assign w13097 = pi2564 & ~w5274;
assign w13098 = pi1899 & ~w15036;
assign w13099 = ~w12040 & pi0697;
assign w13100 = ~w6785 & pi0855;
assign w13101 = pi2341 & ~w18123;
assign w13102 = ~w18166 & ~w10159;
assign w13103 = ~pi3131 & w13570;
assign w13104 = ~pi3336 & w6072;
assign w13105 = w13509 & w15095;
assign w13106 = ~w8166 & ~w2559;
assign w13107 = ~w14828 & w6506;
assign w13108 = w13149 & w2531;
assign w13109 = w13509 & w8548;
assign w13110 = ~w11456 & ~w2244;
assign w13111 = ~w5560 & w14931;
assign w13112 = ~w5783 & ~w3310;
assign w13113 = ~w3544 & ~pi0511;
assign w13114 = w13509 & w2514;
assign w13115 = pi1912 & ~w10299;
assign w13116 = w14352 & w11517;
assign w13117 = ~w15204 & ~w8635;
assign w13118 = pi3146 & w18497;
assign w13119 = ~w724 & ~w570;
assign w13120 = pi1815 & ~w653;
assign w13121 = ~w7844 & pi0901;
assign w13122 = ~pi0821 & w1147;
assign w13123 = ~pi0733 & w17899;
assign w13124 = w15808 & ~w3374;
assign w13125 = pi2259 & ~w11671;
assign w13126 = pi0187 & w5274;
assign w13127 = ~w18124 & ~w10377;
assign w13128 = ~w10784 & w17286;
assign w13129 = w16278 & ~w14143;
assign w13130 = ~w15808 & pi0753;
assign w13131 = ~w13703 & w8905;
assign w13132 = ~w3203 & pi0584;
assign w13133 = ~pi2477 & w5384;
assign w13134 = ~pi3095 & w3555;
assign w13135 = w3988 & w4333;
assign w13136 = pi2590 & ~w5274;
assign w13137 = ~w9440 & ~w18338;
assign w13138 = w1391 & ~w6680;
assign w13139 = w15450 & w18490;
assign w13140 = ~w16769 & ~w1914;
assign w13141 = (pi0855 & ~w13509) | (pi0855 & w13100) | (~w13509 & w13100);
assign w13142 = w11505 & w2905;
assign w13143 = ~w5510 & ~w3968;
assign w13144 = w13509 & w1806;
assign w13145 = ~w14656 & ~w17821;
assign w13146 = ~w17769 & ~w7625;
assign w13147 = ~w10903 & ~w10323;
assign w13148 = pi0436 & w17173;
assign w13149 = w15612 & w9941;
assign w13150 = pi1670 & w4683;
assign w13151 = (~pi0332 & ~w6857) | (~pi0332 & w8438) | (~w6857 & w8438);
assign w13152 = ~w11834 & ~w5707;
assign w13153 = ~w6139 & ~w18248;
assign w13154 = pi2713 & ~w16815;
assign w13155 = w3747 & w12732;
assign w13156 = (pi0762 & ~w13509) | (pi0762 & w12402) | (~w13509 & w12402);
assign w13157 = ~pi2204 & w5075;
assign w13158 = ~w2014 & w11816;
assign w13159 = w11209 & ~w3101;
assign w13160 = w1368 & pi0385;
assign w13161 = w15359 & w14199;
assign w13162 = ~w756 & ~w16855;
assign w13163 = w5517 & w1114;
assign w13164 = ~pi0903 & w1147;
assign w13165 = ~pi0091 & w9284;
assign w13166 = pi0092 & w9284;
assign w13167 = ~w2341 & pi0846;
assign w13168 = ~w17873 & ~w10844;
assign w13169 = w1127 & ~w17022;
assign w13170 = ~w4823 & ~w12416;
assign w13171 = pi1852 & ~w2732;
assign w13172 = pi2643 & ~w3555;
assign w13173 = ~pi3155 & pi3166;
assign w13174 = (~pi2920 & ~w384) | (~pi2920 & w8216) | (~w384 & w8216);
assign w13175 = w2742 & ~w7592;
assign w13176 = pi0064 & w6393;
assign w13177 = ~w618 & ~w6260;
assign w13178 = ~w7335 & ~w8074;
assign w13179 = (pi0589 & ~w13509) | (pi0589 & w18537) | (~w13509 & w18537);
assign w13180 = w11345 & w7001;
assign w13181 = pi1625 & ~w18259;
assign w13182 = ~pi0915 & w6200;
assign w13183 = (pi0576 & ~w13509) | (pi0576 & w9301) | (~w13509 & w9301);
assign w13184 = ~w3055 & w1748;
assign w13185 = ~w3243 & pi0321;
assign w13186 = ~pi2320 & w16041;
assign w13187 = pi2227 & ~w11735;
assign w13188 = w7703 & w7797;
assign w13189 = ~w453 & w8487;
assign w13190 = ~w14824 & ~w4734;
assign w13191 = ~w17818 & ~w4473;
assign w13192 = ~w8588 & w3223;
assign w13193 = ~w9561 & ~w10653;
assign w13194 = w8337 & pi3329;
assign w13195 = ~w2510 & ~w4895;
assign w13196 = pi1780 & ~w8829;
assign w13197 = ~w15472 & ~w5598;
assign w13198 = pi0261 & w5274;
assign w13199 = (~pi0973 & ~w13509) | (~pi0973 & w7872) | (~w13509 & w7872);
assign w13200 = w16506 & ~w10947;
assign w13201 = ~w12692 & ~w3393;
assign w13202 = ~w11766 & ~w17386;
assign w13203 = ~w1892 & w5293;
assign w13204 = w2425 & w3556;
assign w13205 = w18267 & ~w1620;
assign w13206 = (pi1262 & ~w5437) | (pi1262 & w15882) | (~w5437 & w15882);
assign w13207 = ~w16632 & ~w8960;
assign w13208 = ~w4344 & ~w7559;
assign w13209 = ~w815 & ~w2817;
assign w13210 = ~pi3139 & w17669;
assign w13211 = pi0013 & ~w3748;
assign w13212 = ~pi0483 & pi3387;
assign w13213 = ~w6785 & pi0850;
assign w13214 = (pi0724 & ~w13509) | (pi0724 & w2267) | (~w13509 & w2267);
assign w13215 = ~w6697 & ~pi0960;
assign w13216 = pi2257 & ~w11671;
assign w13217 = (~w7428 & ~w1516) | (~w7428 & w16616) | (~w1516 & w16616);
assign w13218 = (pi1024 & ~w13509) | (pi1024 & w16374) | (~w13509 & w16374);
assign w13219 = (~pi3109 & w12651) | (~pi3109 & w11245) | (w12651 & w11245);
assign w13220 = ~pi3081 & pi3139;
assign w13221 = ~w2034 & ~w12795;
assign w13222 = ~pi1970 & ~w5274;
assign w13223 = ~pi3059 & w6463;
assign w13224 = pi0056 & pi0067;
assign w13225 = ~w11089 & ~w7673;
assign w13226 = w10647 & ~w11572;
assign w13227 = ~w17987 & w8410;
assign w13228 = pi3164 & w3987;
assign w13229 = ~w18053 & w10571;
assign w13230 = ~pi3135 & w17387;
assign w13231 = w6676 & w13679;
assign w13232 = w1500 & pi0262;
assign w13233 = w8337 & pi3312;
assign w13234 = ~pi1933 & w2151;
assign w13235 = pi2773 & ~w6463;
assign w13236 = ~pi2874 & w2431;
assign w13237 = ~w11219 & ~w1039;
assign w13238 = ~pi3154 & pi3207;
assign w13239 = ~w13157 & ~w1769;
assign w13240 = ~w3609 & ~w8750;
assign w13241 = ~w5031 & ~pi1233;
assign w13242 = ~w2280 & ~pi0061;
assign w13243 = ~w1013 & ~w11557;
assign w13244 = w13509 & w6951;
assign w13245 = ~w11547 & ~w1156;
assign w13246 = (pi0708 & ~w13509) | (pi0708 & w1581) | (~w13509 & w1581);
assign w13247 = ~pi3336 & w6448;
assign w13248 = ~w11655 & w6551;
assign w13249 = ~w10388 & w2568;
assign w13250 = w9440 & w12460;
assign w13251 = ~w220 & w12707;
assign w13252 = pi1496 & ~w13753;
assign w13253 = ~pi2814 & w13343;
assign w13254 = ~w5847 & w15956;
assign w13255 = w968 & ~pi0274;
assign w13256 = pi2842 & w14148;
assign w13257 = ~pi2353 & w12755;
assign w13258 = w3203 & ~w11978;
assign w13259 = ~w869 & ~w3990;
assign w13260 = pi2935 & ~pi3205;
assign w13261 = ~w14648 & ~pi2713;
assign w13262 = ~w12326 & ~w12194;
assign w13263 = ~w2341 & pi0826;
assign w13264 = ~w4903 & w4892;
assign w13265 = w11752 & w6007;
assign w13266 = pi1284 & pi1345;
assign w13267 = ~w1447 & ~w7865;
assign w13268 = w14560 & pi0347;
assign w13269 = (pi0903 & ~w13509) | (pi0903 & w17180) | (~w13509 & w17180);
assign w13270 = pi0230 & ~w15142;
assign w13271 = ~w8412 & ~w7812;
assign w13272 = ~pi2967 & pi3081;
assign w13273 = ~pi2967 & ~pi3080;
assign w13274 = w9640 & w5495;
assign w13275 = ~w131 & w12775;
assign w13276 = ~w16575 & w4277;
assign w13277 = ~pi0742 & w17490;
assign w13278 = pi2439 & ~w3223;
assign w13279 = ~w4573 & w9697;
assign w13280 = pi3169 & ~pi3171;
assign w13281 = ~w12937 & ~w18538;
assign w13282 = pi1876 & ~w15036;
assign w13283 = ~w3514 & ~w5570;
assign w13284 = w4240 & w11459;
assign w13285 = w709 & pi1894;
assign w13286 = ~w5458 & ~w9207;
assign w13287 = ~w4605 & ~w10495;
assign w13288 = pi2540 & w14148;
assign w13289 = w17619 & w5778;
assign w13290 = ~pi2975 & w4420;
assign w13291 = ~w15022 & ~w10981;
assign w13292 = w384 & w4642;
assign w13293 = ~w4580 & ~w1267;
assign w13294 = (pi0769 & ~w13509) | (pi0769 & w14488) | (~w13509 & w14488);
assign w13295 = ~pi3092 & w6463;
assign w13296 = ~w6195 & w15927;
assign w13297 = ~w2638 & ~w18393;
assign w13298 = (~pi0979 & ~w13509) | (~pi0979 & w10754) | (~w13509 & w10754);
assign w13299 = ~w12460 & w5977;
assign w13300 = (pi0605 & ~w13509) | (pi0605 & w4127) | (~w13509 & w4127);
assign w13301 = ~w1791 & w14559;
assign w13302 = w5437 & w14983;
assign w13303 = (pi0757 & ~w13509) | (pi0757 & w940) | (~w13509 & w940);
assign w13304 = pi1740 & ~w4058;
assign w13305 = pi3160 & ~pi3484;
assign w13306 = w6857 & w11218;
assign w13307 = w968 & ~pi0290;
assign w13308 = (~w13367 & w17577) | (~w13367 & w4501) | (w17577 & w4501);
assign w13309 = w13231 & w4470;
assign w13310 = ~pi2103 & w12724;
assign w13311 = ~w14988 & ~w15366;
assign w13312 = ~pi3227 & ~pi3371;
assign w13313 = w15808 & ~w16498;
assign w13314 = w17646 & w6320;
assign w13315 = (pi0314 & w3055) | (pi0314 & w10710) | (w3055 & w10710);
assign w13316 = ~pi0314 & pi3229;
assign w13317 = ~pi3350 & w7090;
assign w13318 = pi0063 & pi0068;
assign w13319 = ~w8106 & ~w12257;
assign w13320 = ~w15534 & ~w3664;
assign w13321 = ~w9810 & w13756;
assign w13322 = (pi0734 & ~w13509) | (pi0734 & w2712) | (~w13509 & w2712);
assign w13323 = ~w18495 & ~w12135;
assign w13324 = w13509 & w18089;
assign w13325 = pi2539 & w15191;
assign w13326 = ~w17654 & ~w12248;
assign w13327 = w7307 & w4710;
assign w13328 = ~w5216 & ~w18116;
assign w13329 = w16620 & w9476;
assign w13330 = ~w601 & ~w15436;
assign w13331 = ~w12763 & ~w6264;
assign w13332 = ~w4979 & ~w10788;
assign w13333 = ~pi3153 & w12427;
assign w13334 = ~pi2040 & w13204;
assign w13335 = (pi0396 & w5560) | (pi0396 & w6229) | (w5560 & w6229);
assign w13336 = ~w12040 & pi0689;
assign w13337 = ~pi3092 & w15235;
assign w13338 = ~w4061 & ~w413;
assign w13339 = w17562 & pi2565;
assign w13340 = ~w709 & pi1276;
assign w13341 = pi1419 & ~w6072;
assign w13342 = ~w10939 & ~w15735;
assign w13343 = ~w1791 & w7307;
assign w13344 = w7254 & w4470;
assign w13345 = pi0019 & ~w14148;
assign w13346 = ~w1117 & w5477;
assign w13347 = ~w12878 & w894;
assign w13348 = pi2207 & ~w3223;
assign w13349 = w14109 & pi0430;
assign w13350 = ~w5189 & pi0547;
assign w13351 = pi3363 & w13367;
assign w13352 = ~w18414 & ~w1406;
assign w13353 = w6857 & w12753;
assign w13354 = ~w1488 & w5957;
assign w13355 = pi1317 & ~w107;
assign w13356 = w1368 & pi0402;
assign w13357 = ~w11213 & ~w252;
assign w13358 = ~pi3158 & w3805;
assign w13359 = ~pi3315 & w9781;
assign w13360 = ~w11809 & ~w9141;
assign w13361 = ~pi1254 & w11655;
assign w13362 = (pi0575 & ~w13509) | (pi0575 & w7099) | (~w13509 & w7099);
assign w13363 = ~pi3049 & w261;
assign w13364 = pi1771 & ~w5457;
assign w13365 = pi1703 & w4683;
assign w13366 = (pi1794 & w7215) | (pi1794 & w14099) | (w7215 & w14099);
assign w13367 = ~pi0483 & w11345;
assign w13368 = pi2989 & pi3179;
assign w13369 = (pi1184 & ~w5437) | (pi1184 & w13648) | (~w5437 & w13648);
assign w13370 = ~w7596 & w15405;
assign w13371 = ~w12021 & ~w5940;
assign w13372 = pi0173 & ~pi0179;
assign w13373 = w11383 & w10881;
assign w13374 = ~w7033 & w9323;
assign w13375 = ~w5189 & pi0738;
assign w13376 = pi1874 & ~w15036;
assign w13377 = w10189 & ~pi0457;
assign w13378 = w13509 & w14238;
assign w13379 = pi0087 & w3748;
assign w13380 = pi0062 & w922;
assign w13381 = w16136 & w18483;
assign w13382 = ~w13329 & ~w13367;
assign w13383 = ~pi3330 & w17935;
assign w13384 = w16506 & w1217;
assign w13385 = ~w17665 & ~w11385;
assign w13386 = w15117 & w9577;
assign w13387 = (pi0626 & ~w13509) | (pi0626 & w3380) | (~w13509 & w3380);
assign w13388 = ~pi2318 & w5075;
assign w13389 = (pi0649 & ~w13509) | (pi0649 & w1384) | (~w13509 & w1384);
assign w13390 = ~pi1690 & w17213;
assign w13391 = w9440 & pi0148;
assign w13392 = ~pi3172 & w12427;
assign w13393 = w13509 & w7613;
assign w13394 = ~pi2252 & w18209;
assign w13395 = ~w8066 & w10008;
assign w13396 = w13509 & w8460;
assign w13397 = ~pi3152 & pi2950;
assign w13398 = w7077 & ~w7449;
assign w13399 = w9501 & w1239;
assign w13400 = pi1337 & ~pi0250;
assign w13401 = pi1337 & pi0251;
assign w13402 = ~pi3200 & w3522;
assign w13403 = w14833 & w14078;
assign w13404 = w934 & pi0413;
assign w13405 = w13509 & w415;
assign w13406 = pi2322 & ~w15883;
assign w13407 = pi2398 & ~w3223;
assign w13408 = pi3028 & ~pi3157;
assign w13409 = ~w12573 & ~w11629;
assign w13410 = w7844 & ~w17210;
assign w13411 = ~w15122 & ~pi2679;
assign w13412 = w11416 & w11024;
assign w13413 = ~w6765 & ~w14461;
assign w13414 = ~w1641 & w7025;
assign w13415 = ~w8625 & ~w10358;
assign w13416 = ~pi3099 & w16815;
assign w13417 = w1127 & ~w11533;
assign w13418 = pi3111 & ~w16502;
assign w13419 = ~pi3085 & w16815;
assign w13420 = ~w4948 & ~w8691;
assign w13421 = ~w3239 & ~w2291;
assign w13422 = pi2421 & ~w3223;
assign w13423 = ~w9653 & w10314;
assign w13424 = (pi0366 & w6195) | (pi0366 & w16036) | (w6195 & w16036);
assign w13425 = ~w1791 & w11918;
assign w13426 = w13454 & w4881;
assign w13427 = pi0085 & pi3254;
assign w13428 = w6926 & w11697;
assign w13429 = w13509 & w4456;
assign w13430 = w17286 & ~w5855;
assign w13431 = ~w9677 & ~w7050;
assign w13432 = ~pi2179 & w2151;
assign w13433 = pi1781 & ~w8829;
assign w13434 = ~w168 & w8828;
assign w13435 = w6649 & ~w16303;
assign w13436 = w13862 & w6044;
assign w13437 = ~w9791 & ~w3880;
assign w13438 = pi1618 & w13753;
assign w13439 = ~w14648 & ~pi2886;
assign w13440 = ~pi3333 & w14918;
assign w13441 = ~w14648 & ~pi2622;
assign w13442 = pi2086 & ~w17683;
assign w13443 = w3987 & w16680;
assign w13444 = w3223 & w9407;
assign w13445 = ~w18208 & ~w9156;
assign w13446 = ~w3463 & ~w436;
assign w13447 = ~w6785 & pi1205;
assign w13448 = ~w4812 & ~w12031;
assign w13449 = ~pi3133 & w8515;
assign w13450 = w10158 & w14078;
assign w13451 = ~pi1263 & pi2958;
assign w13452 = pi2870 & w15191;
assign w13453 = ~w9774 & ~w10543;
assign w13454 = ~w16561 & ~w911;
assign w13455 = w18258 & w17824;
assign w13456 = ~pi1840 & w13065;
assign w13457 = ~pi1068 & w93;
assign w13458 = (~pi0512 & w17577) | (~pi0512 & w3775) | (w17577 & w3775);
assign w13459 = w13509 & w17834;
assign w13460 = ~pi3169 & w15839;
assign w13461 = w15008 & w5574;
assign w13462 = w13509 & w6751;
assign w13463 = pi0258 & w5274;
assign w13464 = w14648 & ~pi2618;
assign w13465 = pi1520 & ~w14918;
assign w13466 = ~pi3315 & w18259;
assign w13467 = ~w6216 & ~w14410;
assign w13468 = (pi0614 & ~w13509) | (pi0614 & w15061) | (~w13509 & w15061);
assign w13469 = pi2468 & ~w17646;
assign w13470 = w6857 & w18588;
assign w13471 = ~w13414 & ~w3593;
assign w13472 = pi1224 & pi1211;
assign w13473 = ~pi0859 & w15707;
assign w13474 = ~pi3290 & w7090;
assign w13475 = ~w17189 & w11479;
assign w13476 = w13321 & ~w1749;
assign w13477 = w9028 & w16244;
assign w13478 = ~pi3093 & w16815;
assign w13479 = pi3160 & ~w3384;
assign w13480 = w6857 & w14191;
assign w13481 = ~w625 & ~w13367;
assign w13482 = ~w13612 & ~w2082;
assign w13483 = ~w9728 & ~w1622;
assign w13484 = ~w1136 & ~w7260;
assign w13485 = w16575 & w11855;
assign w13486 = pi0490 & pi1137;
assign w13487 = ~pi0489 & ~pi1136;
assign w13488 = w384 & w9076;
assign w13489 = pi2756 & ~w11406;
assign w13490 = pi2055 & ~w10158;
assign w13491 = ~pi3169 & w3805;
assign w13492 = ~w12660 & w6064;
assign w13493 = ~pi3315 & w6072;
assign w13494 = ~pi0801 & w543;
assign w13495 = ~w3942 & ~w15624;
assign w13496 = w18123 & w614;
assign w13497 = (w15842 & ~w16893) | (w15842 & w5544) | (~w16893 & w5544);
assign w13498 = w4420 & w14078;
assign w13499 = ~pi0719 & w17899;
assign w13500 = w11345 & w13212;
assign w13501 = ~pi3147 & w17993;
assign w13502 = w14648 & ~pi2735;
assign w13503 = w13509 & w3921;
assign w13504 = pi1873 & ~w15036;
assign w13505 = pi1920 & ~w15271;
assign w13506 = w15883 & w2753;
assign w13507 = ~pi2661 & w17213;
assign w13508 = ~w17603 & ~w4518;
assign w13509 = w18200 & ~w1313;
assign w13510 = ~w7825 & ~w7273;
assign w13511 = w16506 & ~w7199;
assign w13512 = ~w18392 & ~w13877;
assign w13513 = pi1548 & w13753;
assign w13514 = ~pi1129 & ~w14073;
assign w13515 = (pi0861 & ~w13509) | (pi0861 & w11792) | (~w13509 & w11792);
assign w13516 = ~w11127 & ~w866;
assign w13517 = pi3160 & ~pi3483;
assign w13518 = pi0108 & w9284;
assign w13519 = ~pi1139 & w9420;
assign w13520 = w2041 & w8585;
assign w13521 = w13509 & w16716;
assign w13522 = pi2749 & ~w5274;
assign w13523 = ~pi3157 & ~pi3160;
assign w13524 = w6785 & ~w6033;
assign w13525 = ~pi0280 & w2196;
assign w13526 = w13509 & w82;
assign w13527 = ~w1153 & ~w5254;
assign w13528 = w7844 & ~w6647;
assign w13529 = (~pi1238 & ~w11505) | (~pi1238 & w3720) | (~w11505 & w3720);
assign w13530 = ~w15808 & pi0740;
assign w13531 = ~w1962 & pi0944;
assign w13532 = w13509 & w11123;
assign w13533 = ~w9202 & ~w16282;
assign w13534 = w13509 & w11124;
assign w13535 = pi2171 & ~w15271;
assign w13536 = ~w4669 & ~w1490;
assign w13537 = w13509 & w1935;
assign w13538 = w14560 & pi0365;
assign w13539 = ~w13487 & ~w427;
assign w13540 = ~w17734 & ~w14749;
assign w13541 = w7000 & w3280;
assign w13542 = ~w17363 & ~w13288;
assign w13543 = pi0020 & ~w14148;
assign w13544 = pi1820 & ~w653;
assign w13545 = ~w15045 & w3656;
assign w13546 = pi0082 & w12161;
assign w13547 = ~w4554 & ~pi2969;
assign w13548 = ~w4091 & ~w12303;
assign w13549 = ~w6651 & ~w15399;
assign w13550 = w17562 & pi2749;
assign w13551 = ~w7109 & w442;
assign w13552 = pi1193 & ~w12581;
assign w13553 = ~w10764 & ~w3848;
assign w13554 = w384 & w5488;
assign w13555 = ~w17534 & pi0138;
assign w13556 = pi3149 & w12583;
assign w13557 = w13509 & w8263;
assign w13558 = ~pi3049 & w16815;
assign w13559 = ~w13761 & ~w9137;
assign w13560 = (w14137 & w13116) | (w14137 & w12518) | (w13116 & w12518);
assign w13561 = w15341 & w9821;
assign w13562 = pi1611 & ~w7090;
assign w13563 = (~pi0325 & ~w325) | (~pi0325 & w319) | (~w325 & w319);
assign w13564 = (pi0326 & ~w325) | (pi0326 & w320) | (~w325 & w320);
assign w13565 = ~w10501 & ~w10769;
assign w13566 = w9694 & w16527;
assign w13567 = ~w16506 & pi1142;
assign w13568 = pi0483 & ~pi2960;
assign w13569 = pi2969 & ~w8789;
assign w13570 = ~w4020 & w17683;
assign w13571 = ~pi3049 & w6463;
assign w13572 = ~pi0827 & w93;
assign w13573 = ~w10260 & ~w14452;
assign w13574 = (pi0393 & w5560) | (pi0393 & w12862) | (w5560 & w12862);
assign w13575 = (pi0657 & ~w13509) | (pi0657 & w18221) | (~w13509 & w18221);
assign w13576 = ~pi1948 & w11688;
assign w13577 = (pi0628 & ~w13509) | (pi0628 & w9763) | (~w13509 & w9763);
assign w13578 = ~w17992 & ~w8601;
assign w13579 = ~pi3133 & pi0197;
assign w13580 = (pi0679 & ~w13509) | (pi0679 & w7524) | (~w13509 & w7524);
assign w13581 = ~w11003 & ~w10982;
assign w13582 = pi2806 & ~w6463;
assign w13583 = ~pi3171 & w4310;
assign w13584 = ~pi2982 & pi2995;
assign w13585 = ~pi1244 & w11655;
assign w13586 = w3987 & w637;
assign w13587 = ~w11161 & ~pi0514;
assign w13588 = ~w7077 & pi0803;
assign w13589 = ~w4549 & ~w8744;
assign w13590 = ~pi0323 & ~pi3235;
assign w13591 = ~w5966 & ~w16178;
assign w13592 = ~w16544 & w13112;
assign w13593 = pi2595 & ~w9504;
assign w13594 = ~w7814 & w7305;
assign w13595 = w10647 & ~w17777;
assign w13596 = pi2148 & ~w11671;
assign w13597 = ~w5583 & ~w17258;
assign w13598 = pi2053 & ~w10158;
assign w13599 = ~w8215 & ~w8545;
assign w13600 = ~pi3095 & w16815;
assign w13601 = ~w6288 & w12433;
assign w13602 = ~pi0223 & pi0224;
assign w13603 = (pi0736 & ~w13509) | (pi0736 & w2824) | (~w13509 & w2824);
assign w13604 = (pi0545 & ~w13509) | (pi0545 & w15575) | (~w13509 & w15575);
assign w13605 = ~pi1985 & w314;
assign w13606 = w5647 & w3629;
assign w13607 = pi2492 & ~w15235;
assign w13608 = (~pi0295 & ~w6857) | (~pi0295 & w14625) | (~w6857 & w14625);
assign w13609 = pi1544 & w13753;
assign w13610 = w14524 & w3515;
assign w13611 = ~pi0574 & w795;
assign w13612 = pi2733 & ~w5274;
assign w13613 = (pi0354 & w6195) | (pi0354 & w9525) | (w6195 & w9525);
assign w13614 = w13509 & w13043;
assign w13615 = ~w5532 & ~w13422;
assign w13616 = pi2509 & ~w15235;
assign w13617 = pi2465 & ~w13367;
assign w13618 = ~pi2162 & w13065;
assign w13619 = ~pi3288 & w6072;
assign w13620 = w15037 & w7651;
assign w13621 = ~pi3418 & w15036;
assign w13622 = w6982 & w10186;
assign w13623 = pi2651 & ~w16815;
assign w13624 = ~w266 & w332;
assign w13625 = pi1676 & ~w16237;
assign w13626 = ~w16833 & w10084;
assign w13627 = pi3171 & w653;
assign w13628 = pi1230 & ~w8011;
assign w13629 = w7703 & w14817;
assign w13630 = w13509 & w17314;
assign w13631 = ~w10345 & ~w7663;
assign w13632 = ~pi0654 & w3791;
assign w13633 = ~pi3298 & w16922;
assign w13634 = ~w13582 & ~w16196;
assign w13635 = ~w15497 & ~w2002;
assign w13636 = pi2812 & ~w15235;
assign w13637 = w13509 & w4205;
assign w13638 = ~pi2059 & w8617;
assign w13639 = w9440 & pi0192;
assign w13640 = w13509 & w17700;
assign w13641 = ~w9687 & ~w4134;
assign w13642 = w1391 & ~w6647;
assign w13643 = ~w12013 & ~w6167;
assign w13644 = ~pi0865 & w15707;
assign w13645 = (pi0690 & ~w13509) | (pi0690 & w2760) | (~w13509 & w2760);
assign w13646 = ~w13218 & ~w14333;
assign w13647 = ~w2775 & ~w12989;
assign w13648 = ~w16506 & pi1184;
assign w13649 = ~w6781 & ~w3363;
assign w13650 = ~w13767 & ~w9114;
assign w13651 = ~w6399 & ~w7473;
assign w13652 = ~w15986 & ~w8775;
assign w13653 = ~w3000 & ~pi2805;
assign w13654 = (pi1266 & ~w14094) | (pi1266 & w5404) | (~w14094 & w5404);
assign w13655 = pi1763 & ~w14951;
assign w13656 = ~w16278 & pi1106;
assign w13657 = pi1807 & ~w9520;
assign w13658 = pi2600 & ~w9504;
assign w13659 = ~w8087 & w14234;
assign w13660 = ~pi3298 & w14918;
assign w13661 = w9440 & pi0165;
assign w13662 = ~w15146 & ~pi0513;
assign w13663 = (pi0894 & ~w13509) | (pi0894 & w16584) | (~w13509 & w16584);
assign w13664 = (pi0943 & ~w13509) | (pi0943 & w8861) | (~w13509 & w8861);
assign w13665 = w539 & ~w1331;
assign w13666 = ~w2014 & w14195;
assign w13667 = (pi0590 & ~w13509) | (pi0590 & w2072) | (~w13509 & w2072);
assign w13668 = ~pi2055 & w13204;
assign w13669 = ~pi2014 & w11688;
assign w13670 = w16965 & ~pi2971;
assign w13671 = ~w1814 & ~w17727;
assign w13672 = w3203 & ~w1236;
assign w13673 = ~pi3349 & w14918;
assign w13674 = ~w12144 & ~w18226;
assign w13675 = ~w13759 & ~w933;
assign w13676 = w15706 & w4065;
assign w13677 = w13509 & w3800;
assign w13678 = ~pi1101 & w17899;
assign w13679 = pi1167 & ~pi1176;
assign w13680 = ~w12454 & ~w13055;
assign w13681 = ~w5453 & ~pi1764;
assign w13682 = ~pi0730 & w17899;
assign w13683 = ~w652 & ~w763;
assign w13684 = pi1957 & ~w15883;
assign w13685 = ~w15353 & ~w15911;
assign w13686 = ~w10729 & ~w1283;
assign w13687 = ~pi3103 & w226;
assign w13688 = w5453 & pi2577;
assign w13689 = ~pi3150 & w12427;
assign w13690 = ~w16920 & w4635;
assign w13691 = w6523 & ~w10026;
assign w13692 = pi2764 & ~w226;
assign w13693 = pi1607 & w13753;
assign w13694 = ~w17867 & ~w9758;
assign w13695 = ~w13758 & ~w3856;
assign w13696 = (pi0571 & ~w13509) | (pi0571 & w3913) | (~w13509 & w3913);
assign w13697 = ~w5982 & ~w2304;
assign w13698 = ~w17522 & ~w2576;
assign w13699 = ~w18165 & ~w6067;
assign w13700 = ~w14842 & ~w18114;
assign w13701 = ~w3054 & w5273;
assign w13702 = (pi0848 & ~w13509) | (pi0848 & w11941) | (~w13509 & w11941);
assign w13703 = w12447 & w11949;
assign w13704 = ~w5692 & ~w17138;
assign w13705 = w6649 & ~w3154;
assign w13706 = w2725 & ~w4043;
assign w13707 = ~w10646 & w1867;
assign w13708 = pi0440 & w17173;
assign w13709 = ~pi0439 & w17173;
assign w13710 = ~w14605 & ~w1686;
assign w13711 = ~w17587 & ~w14715;
assign w13712 = ~pi0287 & w2196;
assign w13713 = ~w4502 & ~w2800;
assign w13714 = pi1767 & ~w14951;
assign w13715 = w9440 & pi0204;
assign w13716 = ~w9348 & w10366;
assign w13717 = (pi0835 & ~w13509) | (pi0835 & w17977) | (~w13509 & w17977);
assign w13718 = ~pi3150 & w17669;
assign w13719 = ~pi3054 & w16815;
assign w13720 = ~w9976 & ~w16400;
assign w13721 = ~pi1311 & w882;
assign w13722 = ~w2989 & ~w7080;
assign w13723 = ~w8824 & ~w6613;
assign w13724 = (pi0871 & ~w13509) | (pi0871 & w3497) | (~w13509 & w3497);
assign w13725 = (pi0902 & ~w13509) | (pi0902 & w12218) | (~w13509 & w12218);
assign w13726 = pi2622 & ~w16815;
assign w13727 = (~pi0962 & ~w13509) | (~pi0962 & w10042) | (~w13509 & w10042);
assign w13728 = ~w14633 & w13226;
assign w13729 = ~pi1923 & ~pi1967;
assign w13730 = ~w4020 & w11671;
assign w13731 = ~pi2756 & w13343;
assign w13732 = pi1895 & ~w15036;
assign w13733 = pi2926 & ~w11406;
assign w13734 = ~w12200 & ~w2146;
assign w13735 = ~w15925 & ~w6616;
assign w13736 = w14384 & w18512;
assign w13737 = w6697 & ~w12800;
assign w13738 = ~pi2691 & w17213;
assign w13739 = pi2200 & ~w10299;
assign w13740 = pi3160 & ~pi3493;
assign w13741 = pi2683 & ~w11406;
assign w13742 = pi0418 & w17173;
assign w13743 = w11232 & w1908;
assign w13744 = (pi2958 & w2014) | (pi2958 & w6603) | (w2014 & w6603);
assign w13745 = ~w3794 & ~w15435;
assign w13746 = ~pi2681 & w13343;
assign w13747 = w5567 & w16132;
assign w13748 = pi1616 & ~w7090;
assign w13749 = w5189 & ~w3430;
assign w13750 = w3594 & w12778;
assign w13751 = pi1310 & ~w4232;
assign w13752 = pi2407 & ~w10158;
assign w13753 = ~w10458 & ~w15815;
assign w13754 = ~w18375 & ~w7326;
assign w13755 = w13509 & w2583;
assign w13756 = (w2460 & ~w11232) | (w2460 & w6879) | (~w11232 & w6879);
assign w13757 = w13509 & w18217;
assign w13758 = (~w3351 & w3055) | (~w3351 & w6476) | (w3055 & w6476);
assign w13759 = w11383 & w11009;
assign w13760 = w11232 & w11316;
assign w13761 = pi2626 & ~w16815;
assign w13762 = ~w4946 & w15136;
assign w13763 = w2570 & pi0041;
assign w13764 = ~w18466 & ~w16387;
assign w13765 = w11383 & w10799;
assign w13766 = ~w2272 & ~w18181;
assign w13767 = ~pi3159 & w11701;
assign w13768 = pi3166 & w2848;
assign w13769 = ~pi3295 & w14918;
assign w13770 = ~pi1006 & w14641;
assign w13771 = ~pi1138 & w9420;
assign w13772 = w412 & w6320;
assign w13773 = ~w17133 & ~w17416;
assign w13774 = w10299 & w2753;
assign w13775 = ~w15959 & ~w6150;
assign w13776 = ~w3104 & ~w1187;
assign w13777 = pi1751 & ~w8113;
assign w13778 = w1391 & w1217;
assign w13779 = pi1461 & ~w7090;
assign w13780 = w9102 & ~w17871;
assign w13781 = ~w13032 & ~w1672;
assign w13782 = ~pi0802 & w543;
assign w13783 = ~w5453 & ~pi1803;
assign w13784 = ~w5280 & ~w87;
assign w13785 = ~w3859 & ~w14700;
assign w13786 = w10249 & w876;
assign w13787 = ~w11267 & ~w7665;
assign w13788 = pi1658 & ~w6072;
assign w13789 = w7703 & w18564;
assign w13790 = (pi0493 & ~w11345) | (pi0493 & w9169) | (~w11345 & w9169);
assign w13791 = pi2884 & ~w5274;
assign w13792 = ~pi2449 & w9340;
assign w13793 = ~w10942 & ~w16566;
assign w13794 = pi3131 & pi3207;
assign w13795 = ~w6785 & pi1049;
assign w13796 = w17220 & w15365;
assign w13797 = ~w1897 & ~w1049;
assign w13798 = ~w7844 & ~pi0955;
assign w13799 = ~w4668 & ~w18551;
assign w13800 = ~w1891 & ~w15732;
assign w13801 = w14345 & w15806;
assign w13802 = w5453 & pi2589;
assign w13803 = ~pi2236 & w2151;
assign w13804 = ~pi1082 & w543;
assign w13805 = ~pi0328 & w4058;
assign w13806 = (~w7580 & ~w1206) | (~w7580 & w6977) | (~w1206 & w6977);
assign w13807 = w16650 & ~w1929;
assign w13808 = w10494 & w14056;
assign w13809 = w10818 & ~w11413;
assign w13810 = (pi0773 & ~w13509) | (pi0773 & w16599) | (~w13509 & w16599);
assign w13811 = w8337 & pi3273;
assign w13812 = pi0435 & ~pi2486;
assign w13813 = ~w12234 & ~w676;
assign w13814 = ~w14560 & pi0240;
assign w13815 = pi2229 & ~w15271;
assign w13816 = ~pi2073 & w17439;
assign w13817 = ~w6679 & ~w4378;
assign w13818 = pi3365 & w137;
assign w13819 = ~w3267 & ~w2564;
assign w13820 = ~w2341 & pi0845;
assign w13821 = pi2678 & ~w226;
assign w13822 = w6857 & w7669;
assign w13823 = ~w5289 & ~w8010;
assign w13824 = ~w17044 & ~w15533;
assign w13825 = ~w14666 & ~w16484;
assign w13826 = pi3169 & w13786;
assign w13827 = w7703 & w1819;
assign w13828 = ~w184 & ~w12342;
assign w13829 = ~pi3169 & w11132;
assign w13830 = w10189 & pi0401;
assign w13831 = ~w8704 & ~w6015;
assign w13832 = ~pi1061 & w14641;
assign w13833 = w17248 & ~w13195;
assign w13834 = w14158 & w17495;
assign w13835 = ~w13171 & ~w3677;
assign w13836 = w15271 & w17115;
assign w13837 = ~w2890 & w2385;
assign w13838 = (pi1873 & w2014) | (pi1873 & w4141) | (w2014 & w4141);
assign w13839 = pi2350 & ~w4508;
assign w13840 = ~pi2981 & ~pi2982;
assign w13841 = ~w6257 & ~w2169;
assign w13842 = ~w2603 & ~w5958;
assign w13843 = ~w17577 & w11343;
assign w13844 = ~pi1996 & w3019;
assign w13845 = ~w5463 & ~w460;
assign w13846 = (~w11020 & ~w9420) | (~w11020 & w12372) | (~w9420 & w12372);
assign w13847 = w13509 & w4861;
assign w13848 = ~w1231 & ~w12477;
assign w13849 = ~pi2967 & pi3074;
assign w13850 = ~pi2967 & ~pi3073;
assign w13851 = ~w12040 & pi0926;
assign w13852 = ~w9070 & ~w707;
assign w13853 = ~pi0513 & ~pi1345;
assign w13854 = w10634 & w7931;
assign w13855 = ~w17916 & ~w1704;
assign w13856 = ~w12717 & ~w2487;
assign w13857 = pi2556 & ~w5274;
assign w13858 = (w3050 & ~w1516) | (w3050 & w10147) | (~w1516 & w10147);
assign w13859 = ~w15016 & ~w18363;
assign w13860 = (pi0816 & ~w13509) | (pi0816 & w15645) | (~w13509 & w15645);
assign w13861 = ~pi2998 & ~w6263;
assign w13862 = ~w5233 & ~w1942;
assign w13863 = pi2454 & ~w10299;
assign w13864 = ~pi3287 & w6072;
assign w13865 = ~w12216 & ~w7520;
assign w13866 = w8337 & pi3334;
assign w13867 = ~pi1167 & pi1176;
assign w13868 = ~pi1827 & w3567;
assign w13869 = ~w11924 & ~w721;
assign w13870 = ~w12766 & ~w1094;
assign w13871 = ~w11387 & ~w5330;
assign w13872 = w13509 & w12714;
assign w13873 = pi1712 & w4683;
assign w13874 = ~pi0792 & w543;
assign w13875 = w12040 & ~w1236;
assign w13876 = w2363 & pi1351;
assign w13877 = pi0252 & w5274;
assign w13878 = w4039 & w3598;
assign w13879 = ~pi3000 & ~w3987;
assign w13880 = pi3001 & ~w3987;
assign w13881 = pi2550 & w14148;
assign w13882 = (pi0693 & ~w13509) | (pi0693 & w18251) | (~w13509 & w18251);
assign w13883 = (pi0760 & ~w13509) | (pi0760 & w6170) | (~w13509 & w6170);
assign w13884 = pi1599 & ~w9781;
assign w13885 = ~w3849 & ~w9617;
assign w13886 = w7621 & ~w7079;
assign w13887 = ~pi1342 & pi3001;
assign w13888 = w7077 & ~w7707;
assign w13889 = w14838 & w10196;
assign w13890 = ~w1391 & pi1035;
assign w13891 = ~w6731 & ~w8143;
assign w13892 = pi2355 & ~w17683;
assign w13893 = ~w12053 & ~w3731;
assign w13894 = w16506 & ~w7449;
assign w13895 = pi1863 & ~w458;
assign w13896 = ~pi3128 & w11406;
assign w13897 = ~pi2640 & w15122;
assign w13898 = ~pi3153 & pi3159;
assign w13899 = ~w3359 & ~w17304;
assign w13900 = pi2612 & ~w261;
assign w13901 = ~w5223 & pi1297;
assign w13902 = pi1856 & ~w3555;
assign w13903 = w6649 & ~w449;
assign w13904 = ~w2725 & pi0791;
assign w13905 = w12460 & w14745;
assign w13906 = ~pi0172 & pi0192;
assign w13907 = pi1870 & ~w15036;
assign w13908 = ~w15887 & ~w537;
assign w13909 = ~w15122 & ~pi2875;
assign w13910 = ~pi0962 & w9110;
assign w13911 = ~w16756 & ~w16315;
assign w13912 = ~pi2157 & w15122;
assign w13913 = ~w14955 & w6718;
assign w13914 = ~pi3150 & w3805;
assign w13915 = ~w3657 & ~w13858;
assign w13916 = ~pi2987 & w261;
assign w13917 = ~w4487 & ~w15243;
assign w13918 = pi1857 & ~w9504;
assign w13919 = pi1972 & ~w10694;
assign w13920 = (pi0995 & ~w13509) | (pi0995 & w4728) | (~w13509 & w4728);
assign w13921 = (pi0406 & w5560) | (pi0406 & w8051) | (w5560 & w8051);
assign w13922 = pi2297 & ~w15883;
assign w13923 = pi3042 & ~pi3160;
assign w13924 = pi1610 & ~w9781;
assign w13925 = ~pi2239 & w2151;
assign w13926 = pi2094 & ~w4420;
assign w13927 = w14560 & pi0343;
assign w13928 = ~w4810 & ~w3520;
assign w13929 = ~w3474 & ~w166;
assign w13930 = ~pi0487 & ~pi1135;
assign w13931 = pi2838 & w14148;
assign w13932 = (pi0924 & ~w13509) | (pi0924 & w11141) | (~w13509 & w11141);
assign w13933 = ~pi1400 & ~pi1709;
assign w13934 = ~w1172 & ~w9780;
assign w13935 = ~w10826 & ~w9466;
assign w13936 = ~w6674 & ~w13238;
assign w13937 = w5437 & w1714;
assign w13938 = w13509 & w1166;
assign w13939 = ~w2195 & ~w14539;
assign w13940 = ~pi3103 & w15235;
assign w13941 = ~w16919 & ~w4367;
assign w13942 = pi1413 & ~w13753;
assign w13943 = ~w7221 & ~w3234;
assign w13944 = pi0189 & w5274;
assign w13945 = ~w9039 & w17724;
assign w13946 = ~pi0426 & w17173;
assign w13947 = ~w2725 & pi0802;
assign w13948 = ~w18287 & ~w11358;
assign w13949 = w10367 & w5515;
assign w13950 = ~w14228 & pi1004;
assign w13951 = ~pi3353 & w7090;
assign w13952 = ~w5432 & ~w6632;
assign w13953 = w15122 & ~pi2601;
assign w13954 = ~pi0263 & ~w18374;
assign w13955 = pi1369 & ~w5043;
assign w13956 = w12460 & w327;
assign w13957 = ~w11807 & w8808;
assign w13958 = w10189 & pi0390;
assign w13959 = (pi0623 & ~w13509) | (pi0623 & w17693) | (~w13509 & w17693);
assign w13960 = w16088 & w7157;
assign w13961 = ~w17540 & w18332;
assign w13962 = ~pi2091 & w12724;
assign w13963 = w1127 & ~w10461;
assign w13964 = pi2915 & ~w2423;
assign w13965 = ~w14560 & pi0228;
assign w13966 = ~pi0290 & w4058;
assign w13967 = ~w362 & ~w16551;
assign w13968 = ~w5622 & ~w3347;
assign w13969 = ~w6049 & w18214;
assign w13970 = pi3032 & ~w16502;
assign w13971 = ~w5415 & w13321;
assign w13972 = ~w877 & ~w1525;
assign w13973 = ~pi3425 & w15036;
assign w13974 = pi3157 & w3987;
assign w13975 = ~w11140 & ~w2827;
assign w13976 = ~w2317 & ~w1255;
assign w13977 = pi2914 & ~pi3205;
assign w13978 = ~w5189 & pi1099;
assign w13979 = pi2040 & ~w10158;
assign w13980 = ~w6091 & ~w2399;
assign w13981 = ~pi1131 & pi1181;
assign w13982 = w14228 & ~w14597;
assign w13983 = ~pi0043 & w922;
assign w13984 = pi0044 & w922;
assign w13985 = ~pi3189 & ~w11966;
assign w13986 = ~pi2306 & w12724;
assign w13987 = w6857 & w729;
assign w13988 = ~pi2166 & w11313;
assign w13989 = ~pi3054 & w6463;
assign w13990 = ~w3243 & pi0319;
assign w13991 = w13509 & w11717;
assign w13992 = pi1995 & ~w9414;
assign w13993 = ~w1118 & ~w9928;
assign w13994 = w11383 & w4480;
assign w13995 = pi1474 & w13753;
assign w13996 = (pi0506 & ~w9282) | (pi0506 & ~w17577) | (~w9282 & ~w17577);
assign w13997 = ~w8868 & ~w16157;
assign w13998 = ~w9051 & ~w2894;
assign w13999 = ~w14648 & ~pi2702;
assign w14000 = w10642 & w5343;
assign w14001 = ~w5968 & ~pi1337;
assign w14002 = ~w18110 & ~w4777;
assign w14003 = ~w720 & w10522;
assign w14004 = w16378 & w6041;
assign w14005 = ~w7623 & ~w1979;
assign w14006 = w5437 & w2884;
assign w14007 = w5189 & ~w1236;
assign w14008 = pi1337 & pi0253;
assign w14009 = ~w9263 & ~w10418;
assign w14010 = pi3077 & w16502;
assign w14011 = ~w18163 & ~pi0489;
assign w14012 = pi0314 & ~pi3229;
assign w14013 = ~w15633 & ~w5862;
assign w14014 = w8658 & pi1784;
assign w14015 = ~w88 & w10572;
assign w14016 = ~w14381 & ~w8448;
assign w14017 = pi3160 & ~pi3489;
assign w14018 = ~w12677 & ~w10929;
assign w14019 = (pi1138 & ~w5437) | (pi1138 & w18147) | (~w5437 & w18147);
assign w14020 = w2742 & ~w5205;
assign w14021 = ~w1952 & ~w9461;
assign w14022 = ~w12831 & ~w3508;
assign w14023 = pi2941 & ~w13367;
assign w14024 = ~w15808 & pi0923;
assign w14025 = ~pi2466 & w5384;
assign w14026 = ~w9177 & ~w3260;
assign w14027 = ~pi0042 & w922;
assign w14028 = pi3131 & w13786;
assign w14029 = w14228 & ~w6922;
assign w14030 = ~w10424 & ~w17767;
assign w14031 = ~w952 & ~w11149;
assign w14032 = pi3133 & w2732;
assign w14033 = ~w3846 & ~w17737;
assign w14034 = ~w13741 & ~w6732;
assign w14035 = (pi0731 & ~w13509) | (pi0731 & w7813) | (~w13509 & w7813);
assign w14036 = ~w3054 & w4552;
assign w14037 = ~pi3169 & w11701;
assign w14038 = ~w17665 & ~w9716;
assign w14039 = pi1670 & ~w18497;
assign w14040 = pi2596 & ~w9504;
assign w14041 = pi3165 & w15767;
assign w14042 = w6340 & w16341;
assign w14043 = ~w2542 & ~w1050;
assign w14044 = (pi0552 & ~w13509) | (pi0552 & w15823) | (~w13509 & w15823);
assign w14045 = pi1721 & ~w8113;
assign w14046 = ~pi3142 & w4310;
assign w14047 = ~w12514 & ~w11609;
assign w14048 = ~w6251 & ~w10709;
assign w14049 = w3203 & ~w15173;
assign w14050 = ~pi3097 & w9504;
assign w14051 = ~pi3172 & w17387;
assign w14052 = w9440 & pi0153;
assign w14053 = ~w7171 & ~w7247;
assign w14054 = ~w13762 & w3836;
assign w14055 = pi3134 & w14951;
assign w14056 = ~w14909 & ~w7600;
assign w14057 = w9857 & w16439;
assign w14058 = pi2026 & ~w17646;
assign w14059 = ~pi3049 & w15235;
assign w14060 = ~w13192 & ~w4545;
assign w14061 = ~w13249 & ~w2715;
assign w14062 = w8337 & pi3300;
assign w14063 = pi3057 & pi3160;
assign w14064 = w12460 & w8610;
assign w14065 = (pi1075 & ~w13509) | (pi1075 & w2652) | (~w13509 & w2652);
assign w14066 = ~w11252 & ~w9069;
assign w14067 = ~pi2983 & ~w14742;
assign w14068 = w10290 & pi1179;
assign w14069 = ~w16892 & ~w9747;
assign w14070 = ~w9238 & ~w12943;
assign w14071 = ~pi1209 & w11010;
assign w14072 = ~w14930 & ~w9067;
assign w14073 = ~w860 & ~w17924;
assign w14074 = w3121 & w11354;
assign w14075 = ~w10997 & ~w2375;
assign w14076 = ~w12478 & ~w16504;
assign w14077 = ~w15718 & ~w14533;
assign w14078 = ~pi3141 & ~w4020;
assign w14079 = ~w15492 & ~w12696;
assign w14080 = (pi1030 & ~w13509) | (pi1030 & w3300) | (~w13509 & w3300);
assign w14081 = w14228 & ~w2776;
assign w14082 = w11356 & w8679;
assign w14083 = ~w12534 & ~w7815;
assign w14084 = ~w7077 & ~pi0964;
assign w14085 = ~w2014 & w2052;
assign w14086 = ~pi1012 & w12197;
assign w14087 = ~pi3150 & w15839;
assign w14088 = ~w11519 & ~w2520;
assign w14089 = ~w3203 & pi0905;
assign w14090 = ~pi3054 & w226;
assign w14091 = w14560 & pi0361;
assign w14092 = w16810 & w1020;
assign w14093 = ~w10958 & ~w18578;
assign w14094 = (~pi0444 & w8562) | (~pi0444 & w882) | (w8562 & w882);
assign w14095 = ~pi2067 & w8617;
assign w14096 = (pi0890 & ~w13509) | (pi0890 & w14346) | (~w13509 & w14346);
assign w14097 = ~w554 & w1253;
assign w14098 = w12040 & ~w6647;
assign w14099 = w8658 & pi1794;
assign w14100 = pi1348 & w4140;
assign w14101 = w12258 & w16000;
assign w14102 = w13509 & w16846;
assign w14103 = ~w15301 & ~w13486;
assign w14104 = w539 & ~w16528;
assign w14105 = ~pi0358 & ~pi0359;
assign w14106 = w11247 & w12230;
assign w14107 = ~w3883 & ~w8386;
assign w14108 = ~w6066 & ~w13295;
assign w14109 = ~w5855 & w1093;
assign w14110 = ~w15146 & ~w13367;
assign w14111 = (pi0810 & ~w13509) | (pi0810 & w7671) | (~w13509 & w7671);
assign w14112 = ~w1791 & w1173;
assign w14113 = w1127 & ~w8820;
assign w14114 = ~pi0512 & ~pi1345;
assign w14115 = ~w12897 & ~w6258;
assign w14116 = ~w6553 & w1834;
assign w14117 = w13509 & w3379;
assign w14118 = ~pi0601 & w12825;
assign w14119 = ~pi2497 & w17213;
assign w14120 = w6857 & w14592;
assign w14121 = w501 & w4372;
assign w14122 = ~pi1021 & w9110;
assign w14123 = ~w10369 & w9098;
assign w14124 = pi1573 & ~w13753;
assign w14125 = ~pi0502 & pi1377;
assign w14126 = ~w17248 & pi0881;
assign w14127 = ~w12400 & w4922;
assign w14128 = (pi0749 & ~w13509) | (pi0749 & w6793) | (~w13509 & w6793);
assign w14129 = ~pi1946 & w7455;
assign w14130 = ~w15463 & ~w13337;
assign w14131 = ~pi1345 & ~pi2938;
assign w14132 = pi1403 & ~w7946;
assign w14133 = ~w176 & ~w3549;
assign w14134 = w6857 & w16915;
assign w14135 = ~pi3337 & w18259;
assign w14136 = ~pi3142 & w11132;
assign w14137 = ~pi3120 & pi3207;
assign w14138 = ~w7681 & w8067;
assign w14139 = (pi1040 & ~w13509) | (pi1040 & w1079) | (~w13509 & w1079);
assign w14140 = w5642 & w12371;
assign w14141 = (pi0915 & ~w13509) | (pi0915 & w12304) | (~w13509 & w12304);
assign w14142 = ~w11581 & w7284;
assign w14143 = ~w8065 & ~w13057;
assign w14144 = w6697 & ~w6647;
assign w14145 = ~pi2435 & w5075;
assign w14146 = (pi1070 & ~w13509) | (pi1070 & w1055) | (~w13509 & w1055);
assign w14147 = w1391 & w15609;
assign w14148 = ~w11059 & ~w1975;
assign w14149 = w539 & ~w1244;
assign w14150 = ~pi0984 & w15707;
assign w14151 = (pi1111 & ~w13509) | (pi1111 & w15373) | (~w13509 & w15373);
assign w14152 = pi1799 & pi3170;
assign w14153 = w6649 & ~w17762;
assign w14154 = ~w11840 & ~w954;
assign w14155 = pi2253 & ~w15883;
assign w14156 = pi2335 & ~w4508;
assign w14157 = ~pi3314 & w18259;
assign w14158 = w17477 & w2258;
assign w14159 = w539 & ~w15632;
assign w14160 = ~pi3050 & w261;
assign w14161 = ~w9023 & w6530;
assign w14162 = ~w5485 & ~w10654;
assign w14163 = w7 & w4013;
assign w14164 = (pi1062 & ~w13509) | (pi1062 & w8627) | (~w13509 & w8627);
assign w14165 = pi3169 & w3987;
assign w14166 = ~w9440 & ~pi0896;
assign w14167 = (pi0634 & ~w13509) | (pi0634 & w57) | (~w13509 & w57);
assign w14168 = ~pi2988 & w261;
assign w14169 = ~pi0602 & w12825;
assign w14170 = ~pi3147 & w8515;
assign w14171 = ~w15138 & w2781;
assign w14172 = ~w5861 & ~w17445;
assign w14173 = w17828 & w4995;
assign w14174 = ~pi3165 & w3805;
assign w14175 = w10189 & pi0379;
assign w14176 = (~pi0954 & ~w13509) | (~pi0954 & w15299) | (~w13509 & w15299);
assign w14177 = ~w581 & ~w17958;
assign w14178 = pi1580 & ~w14918;
assign w14179 = ~w2802 & ~w3476;
assign w14180 = ~w14228 & pi0631;
assign w14181 = ~w5961 & ~w17494;
assign w14182 = ~w17996 & ~w12020;
assign w14183 = pi1382 & w13753;
assign w14184 = ~w14648 & ~pi2651;
assign w14185 = w7703 & w8505;
assign w14186 = w9364 & w14787;
assign w14187 = pi1417 & ~w6072;
assign w14188 = pi0269 & w5274;
assign w14189 = w17758 & w2118;
assign w14190 = pi0098 & w3748;
assign w14191 = w8337 & pi3278;
assign w14192 = ~w10029 & ~w4721;
assign w14193 = w14186 & w306;
assign w14194 = ~w18465 & ~w13757;
assign w14195 = ~w709 & pi1272;
assign w14196 = ~w18163 & ~w13367;
assign w14197 = ~pi3047 & w226;
assign w14198 = ~w9893 & ~w4402;
assign w14199 = ~w12596 & ~w7831;
assign w14200 = ~w1368 & ~pi0477;
assign w14201 = pi2928 & ~w3555;
assign w14202 = ~w9411 & w4674;
assign w14203 = ~w10238 & ~w5836;
assign w14204 = ~w7814 & w4224;
assign w14205 = ~pi3299 & w7090;
assign w14206 = w13509 & w2694;
assign w14207 = pi1997 & ~w9414;
assign w14208 = pi1771 & ~pi3150;
assign w14209 = pi1919 & ~w11735;
assign w14210 = w9227 & w17562;
assign w14211 = ~w5445 & ~w1268;
assign w14212 = pi2264 & ~w11671;
assign w14213 = w6857 & w4874;
assign w14214 = w934 & pi0427;
assign w14215 = w6857 & w3939;
assign w14216 = w6584 & w15612;
assign w14217 = w13412 & w13889;
assign w14218 = ~w2413 & ~w16814;
assign w14219 = ~w12690 & ~w11369;
assign w14220 = ~w10991 & ~w14884;
assign w14221 = pi2618 & ~w261;
assign w14222 = w15118 & ~w4896;
assign w14223 = pi2863 & w14148;
assign w14224 = ~w18329 & ~w12235;
assign w14225 = pi2814 & ~w11406;
assign w14226 = w16278 & ~w6680;
assign w14227 = w16278 & w15609;
assign w14228 = w28 & w13867;
assign w14229 = pi2913 & ~w13753;
assign w14230 = ~pi3106 & w16502;
assign w14231 = ~w11515 & w9261;
assign w14232 = ~w17577 & w9488;
assign w14233 = w2363 & pi1364;
assign w14234 = w2206 & ~w14158;
assign w14235 = w12460 & w2936;
assign w14236 = (pi1155 & ~w5437) | (pi1155 & w3610) | (~w5437 & w3610);
assign w14237 = pi0483 & ~pi0502;
assign w14238 = w3203 & ~w4179;
assign w14239 = w13509 & w6969;
assign w14240 = ~w709 & pi1286;
assign w14241 = ~w16624 & w14364;
assign w14242 = ~w107 & w15876;
assign w14243 = ~pi3094 & w11406;
assign w14244 = ~pi1984 & w3981;
assign w14245 = pi1985 & w3981;
assign w14246 = ~w14560 & pi0216;
assign w14247 = pi2875 & ~w226;
assign w14248 = pi0896 & ~w7219;
assign w14249 = w15122 & ~pi2511;
assign w14250 = ~pi2089 & w12724;
assign w14251 = ~pi1337 & ~pi2911;
assign w14252 = ~w12485 & ~w6519;
assign w14253 = ~w11881 & ~w10210;
assign w14254 = w1127 & ~w8600;
assign w14255 = ~w18179 & ~w4550;
assign w14256 = ~w17248 & pi1174;
assign w14257 = w4470 & w12040;
assign w14258 = pi2795 & w14148;
assign w14259 = pi1554 & ~w18259;
assign w14260 = ~pi3085 & w226;
assign w14261 = ~w9102 & w17871;
assign w14262 = pi1479 & ~w9781;
assign w14263 = ~w15875 & ~w16522;
assign w14264 = w14788 & w13841;
assign w14265 = w10647 & ~w9260;
assign w14266 = ~w990 & ~w2020;
assign w14267 = ~pi1685 & ~w7300;
assign w14268 = ~w15531 & ~w6736;
assign w14269 = pi0483 & pi2465;
assign w14270 = ~pi1834 & w13204;
assign w14271 = pi1601 & w13753;
assign w14272 = w13509 & w7953;
assign w14273 = ~w15517 & ~w17078;
assign w14274 = ~w16506 & pi1158;
assign w14275 = ~w1643 & ~w16296;
assign w14276 = ~pi3166 & w4310;
assign w14277 = ~pi2656 & w17213;
assign w14278 = ~w4284 & ~w13503;
assign w14279 = w8961 & w1985;
assign w14280 = w13243 & w13929;
assign w14281 = w13509 & w5389;
assign w14282 = ~w12821 & ~w14912;
assign w14283 = (pi1083 & ~w13509) | (pi1083 & w5602) | (~w13509 & w5602);
assign w14284 = ~w1452 & ~w117;
assign w14285 = ~w12391 & ~w3118;
assign w14286 = w12471 & ~w14750;
assign w14287 = pi3154 & ~pi3172;
assign w14288 = pi1582 & w13753;
assign w14289 = ~w18164 & ~w2749;
assign w14290 = pi0487 & pi1135;
assign w14291 = ~pi0488 & ~pi1193;
assign w14292 = ~w6697 & pi0677;
assign w14293 = ~w12337 & ~w10437;
assign w14294 = w7799 & w10347;
assign w14295 = w13509 & w3392;
assign w14296 = ~w8803 & ~w11573;
assign w14297 = ~w17396 & ~w15419;
assign w14298 = ~w15687 & ~w13050;
assign w14299 = w2725 & ~w14143;
assign w14300 = ~pi3059 & w9504;
assign w14301 = ~w1315 & ~w5659;
assign w14302 = w13509 & w4842;
assign w14303 = ~w8132 & ~w4928;
assign w14304 = w13381 & w6495;
assign w14305 = w2341 & ~w7707;
assign w14306 = ~pi3003 & ~w3987;
assign w14307 = pi3004 & ~w3987;
assign w14308 = ~pi2057 & w13204;
assign w14309 = w13509 & w15549;
assign w14310 = pi2772 & ~w11406;
assign w14311 = (pi1899 & w2014) | (pi1899 & w4571) | (w2014 & w4571);
assign w14312 = w6697 & w15609;
assign w14313 = pi2188 & ~w11735;
assign w14314 = ~w1221 & ~w10052;
assign w14315 = ~w11424 & ~w14929;
assign w14316 = w2636 & w10067;
assign w14317 = ~w6931 & ~w5779;
assign w14318 = ~w15808 & pi1097;
assign w14319 = w13509 & w16829;
assign w14320 = ~w18395 & ~w4672;
assign w14321 = pi2149 & ~w11671;
assign w14322 = ~w7486 & w443;
assign w14323 = ~w7423 & ~w4198;
assign w14324 = ~w15331 & ~w18131;
assign w14325 = ~w15122 & w7703;
assign w14326 = pi2261 & ~w11671;
assign w14327 = pi2514 & ~w226;
assign w14328 = ~w10884 & w9153;
assign w14329 = ~w12970 & ~w7457;
assign w14330 = ~pi0937 & w9110;
assign w14331 = w6785 & ~w3430;
assign w14332 = w384 & w8194;
assign w14333 = w13509 & w5586;
assign w14334 = pi3018 & pi3020;
assign w14335 = (pi0680 & ~w13509) | (pi0680 & w15566) | (~w13509 & w15566);
assign w14336 = w7077 & ~w14978;
assign w14337 = ~w15847 & ~w16501;
assign w14338 = ~w12828 & ~w5706;
assign w14339 = ~w6529 & ~w13557;
assign w14340 = ~w7142 & ~w17467;
assign w14341 = ~pi1983 & pi1985;
assign w14342 = ~pi1983 & ~pi1984;
assign w14343 = pi1704 & w4667;
assign w14344 = ~pi1032 & w17490;
assign w14345 = ~w17751 & ~w17001;
assign w14346 = ~w17248 & pi0890;
assign w14347 = ~pi1692 & ~pi1805;
assign w14348 = pi2093 & ~w4420;
assign w14349 = ~pi0850 & w15707;
assign w14350 = ~pi0483 & pi3400;
assign w14351 = pi3069 & ~w16502;
assign w14352 = ~pi1159 & ~pi1160;
assign w14353 = ~w16278 & pi0711;
assign w14354 = pi1805 & w13430;
assign w14355 = ~w5453 & ~pi1759;
assign w14356 = ~pi0691 & w9110;
assign w14357 = w934 & pi0447;
assign w14358 = ~w5636 & ~w10880;
assign w14359 = ~w9417 & ~w18485;
assign w14360 = ~pi0485 & ~pi1134;
assign w14361 = ~w14111 & ~w1071;
assign w14362 = ~w7844 & pi0611;
assign w14363 = ~w865 & ~w12625;
assign w14364 = ~w17665 & ~w3553;
assign w14365 = ~w4547 & ~w12627;
assign w14366 = ~w11368 & ~w7405;
assign w14367 = w12040 & ~w3374;
assign w14368 = ~w5048 & ~w1181;
assign w14369 = pi1364 & ~w13108;
assign w14370 = pi1686 & w6960;
assign w14371 = ~pi1856 & w15122;
assign w14372 = pi3146 & w12558;
assign w14373 = pi0054 & w14782;
assign w14374 = pi0304 & pi0325;
assign w14375 = w360 & w18411;
assign w14376 = w11383 & w16024;
assign w14377 = pi1568 & ~w13753;
assign w14378 = ~pi3130 & ~pi1260;
assign w14379 = pi3246 & w3163;
assign w14380 = ~w9487 & ~w4301;
assign w14381 = ~pi0818 & w1147;
assign w14382 = ~w10714 & ~w12736;
assign w14383 = ~w3054 & w4038;
assign w14384 = w11733 & w2006;
assign w14385 = w12975 & w13060;
assign w14386 = pi0151 & w5274;
assign w14387 = (pi0987 & ~w13509) | (pi0987 & w2858) | (~w13509 & w2858);
assign w14388 = ~pi0283 & w2196;
assign w14389 = w13509 & w14147;
assign w14390 = ~w1962 & pi1118;
assign w14391 = ~w3217 & ~w17562;
assign w14392 = w968 & ~pi0331;
assign w14393 = ~w6297 & ~w7585;
assign w14394 = w15271 & w9407;
assign w14395 = pi1130 & w14073;
assign w14396 = ~w16517 & ~w1105;
assign w14397 = ~pi3158 & w4310;
assign w14398 = ~w14435 & ~w2927;
assign w14399 = w16278 & w11302;
assign w14400 = ~pi3138 & w8515;
assign w14401 = pi1566 & ~w13753;
assign w14402 = ~pi0499 & ~pi1345;
assign w14403 = w11800 & w16507;
assign w14404 = ~w17274 & ~w11282;
assign w14405 = pi1784 & ~w17817;
assign w14406 = ~pi3164 & w17993;
assign w14407 = ~pi2016 & w11688;
assign w14408 = ~pi1072 & w1147;
assign w14409 = ~pi2219 & w2151;
assign w14410 = ~pi1075 & w6200;
assign w14411 = ~pi0906 & w795;
assign w14412 = ~w12462 & ~w2976;
assign w14413 = w2725 & ~w13028;
assign w14414 = ~pi3201 & ~w2752;
assign w14415 = w13509 & w7975;
assign w14416 = ~w10263 & w16305;
assign w14417 = pi2974 & w12881;
assign w14418 = ~pi3287 & w16922;
assign w14419 = ~w10094 & ~w7667;
assign w14420 = w17998 & w9334;
assign w14421 = ~w16506 & ~pi1235;
assign w14422 = ~w15157 & ~w445;
assign w14423 = pi2886 & ~w16815;
assign w14424 = ~w18009 & ~w1311;
assign w14425 = ~w36 & ~w2709;
assign w14426 = w14228 & ~w4043;
assign w14427 = pi1727 & ~w4058;
assign w14428 = (pi0798 & ~w13509) | (pi0798 & w3401) | (~w13509 & w3401);
assign w14429 = ~w5189 & pi1028;
assign w14430 = ~w17173 & ~w4066;
assign w14431 = ~pi2356 & w3019;
assign w14432 = ~w1391 & pi0766;
assign w14433 = pi2081 & ~w17683;
assign w14434 = w13840 & w735;
assign w14435 = pi2352 & ~w4420;
assign w14436 = ~pi1036 & w6200;
assign w14437 = w1368 & pi0386;
assign w14438 = pi1325 & w458;
assign w14439 = w11671 & w14078;
assign w14440 = ~w15868 & ~w6654;
assign w14441 = ~w2341 & pi0844;
assign w14442 = ~w14576 & ~w8964;
assign w14443 = ~pi1837 & w12724;
assign w14444 = w13509 & w12123;
assign w14445 = ~w3569 & ~w18252;
assign w14446 = ~pi3102 & ~pi3112;
assign w14447 = pi2789 & ~w11406;
assign w14448 = pi1528 & ~w14918;
assign w14449 = ~w4587 & ~w2677;
assign w14450 = ~w5702 & w16641;
assign w14451 = pi1504 & ~w16922;
assign w14452 = pi2068 & ~w4508;
assign w14453 = ~pi2499 & w17562;
assign w14454 = ~w8286 & ~w16605;
assign w14455 = ~pi3159 & w4310;
assign w14456 = pi3163 & pi3207;
assign w14457 = ~pi3162 & pi3207;
assign w14458 = pi0144 & w5274;
assign w14459 = ~w10374 & ~w18341;
assign w14460 = w16534 & w6569;
assign w14461 = ~pi3349 & w6072;
assign w14462 = pi1337 & ~w6659;
assign w14463 = pi2199 & ~w10299;
assign w14464 = ~w17434 & ~w8270;
assign w14465 = ~w4496 & ~w10493;
assign w14466 = w16506 & ~w15296;
assign w14467 = ~w16240 & ~w3489;
assign w14468 = pi2009 & ~w14833;
assign w14469 = ~w3313 & ~w4011;
assign w14470 = ~w14406 & ~w17184;
assign w14471 = ~pi3350 & w9781;
assign w14472 = pi1742 & w1924;
assign w14473 = pi2240 & ~w11735;
assign w14474 = pi1737 & ~w4058;
assign w14475 = w1155 & w12657;
assign w14476 = pi1585 & w13753;
assign w14477 = ~w2838 & ~w12935;
assign w14478 = pi2883 & ~w226;
assign w14479 = ~w16029 & ~w15219;
assign w14480 = ~w1962 & pi0638;
assign w14481 = pi2901 & ~w5274;
assign w14482 = ~w1307 & w12242;
assign w14483 = w539 & ~w9486;
assign w14484 = w7307 & w17713;
assign w14485 = pi0306 & w5274;
assign w14486 = ~w10479 & ~w6417;
assign w14487 = ~w3943 & ~w17950;
assign w14488 = ~w1391 & pi0769;
assign w14489 = ~w18144 & w13809;
assign w14490 = w14109 & pi0410;
assign w14491 = (pi0648 & ~w13509) | (pi0648 & w16123) | (~w13509 & w16123);
assign w14492 = ~w7814 & w12308;
assign w14493 = ~w12113 & ~w16358;
assign w14494 = pi1900 & ~w15036;
assign w14495 = w968 & ~pi0279;
assign w14496 = ~pi0916 & w11739;
assign w14497 = (pi0867 & ~w13509) | (pi0867 & w10532) | (~w13509 & w10532);
assign w14498 = ~w2014 & w5229;
assign w14499 = ~pi3090 & w6463;
assign w14500 = w17248 & ~w10947;
assign w14501 = ~w2122 & ~w16688;
assign w14502 = w2725 & ~w4179;
assign w14503 = ~w5197 & w10246;
assign w14504 = w14228 & ~w1236;
assign w14505 = ~w428 & ~w11917;
assign w14506 = ~w7005 & ~w9918;
assign w14507 = pi0049 & ~w14148;
assign w14508 = (pi0808 & ~w13509) | (pi0808 & w8503) | (~w13509 & w8503);
assign w14509 = ~w7011 & ~w14807;
assign w14510 = ~pi3053 & w9504;
assign w14511 = ~w14648 & ~pi2931;
assign w14512 = ~w13932 & ~w17460;
assign w14513 = w2613 & ~pi1176;
assign w14514 = ~w15057 & ~w17172;
assign w14515 = ~pi2967 & ~pi3005;
assign w14516 = ~pi2967 & pi3006;
assign w14517 = (pi1785 & w7215) | (pi1785 & w15080) | (w7215 & w15080);
assign w14518 = pi1673 & w1924;
assign w14519 = w13509 & w14029;
assign w14520 = ~w14385 & ~w15242;
assign w14521 = ~pi2349 & w3019;
assign w14522 = ~pi1202 & w1147;
assign w14523 = pi0033 & ~w3748;
assign w14524 = pi1985 & w8370;
assign w14525 = ~w9011 & ~w15607;
assign w14526 = ~w5453 & ~pi1800;
assign w14527 = ~w13322 & ~w1799;
assign w14528 = pi2346 & ~w412;
assign w14529 = w9440 & pi0185;
assign w14530 = (~pi0288 & ~w6857) | (~pi0288 & w4403) | (~w6857 & w4403);
assign w14531 = ~w6697 & pi0662;
assign w14532 = pi2409 & ~w17646;
assign w14533 = ~pi3047 & w11406;
assign w14534 = ~w9764 & ~w17107;
assign w14535 = ~w880 & w6477;
assign w14536 = w7630 & w4340;
assign w14537 = ~w17421 & w18206;
assign w14538 = w13231 & ~w14465;
assign w14539 = ~pi3055 & w11406;
assign w14540 = pi2135 & ~w15883;
assign w14541 = pi1564 & ~w13753;
assign w14542 = w16965 & ~w9991;
assign w14543 = w11209 & ~w2307;
assign w14544 = (pi0825 & ~w13509) | (pi0825 & w8927) | (~w13509 & w8927);
assign w14545 = ~w3000 & ~pi2751;
assign w14546 = w10818 & ~w15039;
assign w14547 = ~w9818 & ~w7464;
assign w14548 = w16278 & ~w7020;
assign w14549 = ~w14660 & ~w5800;
assign w14550 = ~w16017 & ~w13030;
assign w14551 = pi1390 & w13753;
assign w14552 = ~w16506 & pi1137;
assign w14553 = pi1444 & ~w13753;
assign w14554 = ~pi3346 & w16922;
assign w14555 = pi3160 & ~pi3486;
assign w14556 = ~w7694 & ~w5234;
assign w14557 = w7656 & pi2913;
assign w14558 = ~w9849 & ~w13396;
assign w14559 = ~pi2714 & w15122;
assign w14560 = ~pi2960 & w1638;
assign w14561 = ~pi1000 & w12825;
assign w14562 = (~w14583 & ~w5566) | (~w14583 & w1879) | (~w5566 & w1879);
assign w14563 = ~pi0510 & ~pi1345;
assign w14564 = w13509 & w13888;
assign w14565 = pi1333 & ~w9699;
assign w14566 = pi1879 & ~w16815;
assign w14567 = ~w1962 & pi1008;
assign w14568 = ~w14648 & ~pi2605;
assign w14569 = ~pi2995 & w2460;
assign w14570 = ~w11285 & ~w5933;
assign w14571 = ~w10620 & ~w4268;
assign w14572 = w8337 & pi3305;
assign w14573 = ~w13358 & ~w12112;
assign w14574 = pi1691 & ~w11406;
assign w14575 = ~pi2359 & w8617;
assign w14576 = ~pi0568 & w11739;
assign w14577 = ~w7077 & pi0824;
assign w14578 = ~pi1836 & ~w17683;
assign w14579 = ~w6815 & ~w8498;
assign w14580 = ~w13504 & ~w2058;
assign w14581 = ~w11190 & ~w3096;
assign w14582 = ~w9351 & ~w11626;
assign w14583 = pi1375 & ~pi2913;
assign w14584 = w3223 & w17115;
assign w14585 = ~w1368 & ~pi0480;
assign w14586 = (pi1897 & w2014) | (pi1897 & w17657) | (w2014 & w17657);
assign w14587 = ~w15421 & w13967;
assign w14588 = ~pi3162 & w13730;
assign w14589 = ~w18112 & ~w2517;
assign w14590 = ~w17463 & ~w5354;
assign w14591 = ~w1791 & w8724;
assign w14592 = w8337 & pi3283;
assign w14593 = ~pi0973 & w1126;
assign w14594 = ~w10689 & w12775;
assign w14595 = ~w2667 & ~w2995;
assign w14596 = pi2449 & ~w10299;
assign w14597 = ~w1632 & ~w3786;
assign w14598 = pi1352 & ~w13786;
assign w14599 = pi1579 & ~w14918;
assign w14600 = ~w3787 & ~w11890;
assign w14601 = pi1535 & ~w17935;
assign w14602 = ~w8517 & w9400;
assign w14603 = ~w3203 & pi0581;
assign w14604 = ~w1905 & w8186;
assign w14605 = ~pi1999 & w3019;
assign w14606 = ~w9847 & w9145;
assign w14607 = ~pi3135 & w11701;
assign w14608 = ~w7995 & ~w11857;
assign w14609 = ~w1377 & ~w7435;
assign w14610 = ~w13545 & ~w8456;
assign w14611 = (pi0516 & ~w13509) | (pi0516 & w1574) | (~w13509 & w1574);
assign w14612 = ~w10341 & w2111;
assign w14613 = ~w10581 & ~w4752;
assign w14614 = ~w3243 & pi0267;
assign w14615 = w13509 & w1607;
assign w14616 = ~pi3159 & w11132;
assign w14617 = ~w5173 & ~w8807;
assign w14618 = w15842 & pi2554;
assign w14619 = ~w6088 & ~w558;
assign w14620 = (~pi1301 & ~w2325) | (~pi1301 & w215) | (~w2325 & w215);
assign w14621 = ~pi3141 & pi3207;
assign w14622 = pi3142 & pi3207;
assign w14623 = ~w3034 & ~w8654;
assign w14624 = w5383 & pi2535;
assign w14625 = w968 & ~pi0295;
assign w14626 = ~pi1973 & ~pi3370;
assign w14627 = w12460 & w5482;
assign w14628 = pi2568 & w7935;
assign w14629 = ~pi0483 & pi3390;
assign w14630 = w12040 & ~w14597;
assign w14631 = w2725 & ~w16498;
assign w14632 = ~pi3086 & w3555;
assign w14633 = pi1441 & ~w13753;
assign w14634 = ~w3210 & ~w16408;
assign w14635 = ~w2341 & pi1203;
assign w14636 = pi1151 & w9420;
assign w14637 = ~pi1150 & w9420;
assign w14638 = ~pi1046 & w93;
assign w14639 = w15808 & ~w1236;
assign w14640 = pi0068 & ~w14148;
assign w14641 = w12543 & w17490;
assign w14642 = ~w6623 & ~w11650;
assign w14643 = w14746 & w3207;
assign w14644 = pi3170 & w8829;
assign w14645 = ~w16062 & ~w395;
assign w14646 = ~w5848 & ~w4780;
assign w14647 = ~pi3018 & pi3207;
assign w14648 = ~w13184 & ~w6868;
assign w14649 = w1368 & pi0403;
assign w14650 = ~w12205 & w9385;
assign w14651 = pi1983 & ~pi1984;
assign w14652 = (pi0268 & ~w325) | (pi0268 & w9733) | (~w325 & w9733);
assign w14653 = pi1687 & w9205;
assign w14654 = pi2797 & ~w15235;
assign w14655 = ~w16312 & w13131;
assign w14656 = (pi0722 & ~w13509) | (pi0722 & w2178) | (~w13509 & w2178);
assign w14657 = (~pi0963 & ~w13509) | (~pi0963 & w3090) | (~w13509 & w3090);
assign w14658 = w706 & w10354;
assign w14659 = pi3022 & w16502;
assign w14660 = pi2493 & ~w261;
assign w14661 = w13509 & w16718;
assign w14662 = ~w14178 & ~w9813;
assign w14663 = w9653 & w16318;
assign w14664 = ~w16495 & ~w13402;
assign w14665 = pi2699 & ~w16815;
assign w14666 = ~pi2325 & w16041;
assign w14667 = w16630 & w17029;
assign w14668 = ~w13468 & ~w14519;
assign w14669 = ~w2797 & ~w7633;
assign w14670 = w13509 & w16278;
assign w14671 = ~w3128 & ~w8251;
assign w14672 = w13509 & w9833;
assign w14673 = w12460 & w1579;
assign w14674 = ~pi1064 & w93;
assign w14675 = w13509 & w12449;
assign w14676 = pi1515 & w13753;
assign w14677 = ~pi3031 & pi3154;
assign w14678 = ~pi0761 & w6200;
assign w14679 = w8710 & w5360;
assign w14680 = ~w7306 & ~w10081;
assign w14681 = ~w17310 & ~w2333;
assign w14682 = w7307 & w8271;
assign w14683 = pi2258 & ~w11671;
assign w14684 = ~pi2248 & w12941;
assign w14685 = pi2260 & ~w11671;
assign w14686 = ~pi2269 & w13065;
assign w14687 = pi1571 & ~w18259;
assign w14688 = w7703 & w1271;
assign w14689 = ~w7688 & ~w15600;
assign w14690 = pi0144 & pi0150;
assign w14691 = ~w18422 & ~w18587;
assign w14692 = pi1743 & ~w4058;
assign w14693 = ~w18340 & ~w16007;
assign w14694 = w7844 & ~w4179;
assign w14695 = ~pi1239 & ~w14094;
assign w14696 = ~pi3153 & w3982;
assign w14697 = w13509 & w7549;
assign w14698 = ~pi2358 & ~w15450;
assign w14699 = ~pi3146 & w13570;
assign w14700 = ~w649 & w209;
assign w14701 = w3203 & ~w17513;
assign w14702 = pi1348 & ~w7363;
assign w14703 = w7656 & ~pi1224;
assign w14704 = pi2860 & ~w3555;
assign w14705 = ~w6607 & ~w3002;
assign w14706 = pi1567 & ~w13753;
assign w14707 = pi2890 & ~w226;
assign w14708 = ~pi2796 & w17213;
assign w14709 = ~w11242 & ~w9770;
assign w14710 = w16506 & ~w12800;
assign w14711 = ~pi3343 & w18259;
assign w14712 = w13651 & w9926;
assign w14713 = pi1935 & ~w412;
assign w14714 = pi0086 & w3748;
assign w14715 = ~pi0613 & w12825;
assign w14716 = pi1472 & ~w7090;
assign w14717 = ~pi3126 & pi3160;
assign w14718 = ~w4489 & ~w12758;
assign w14719 = ~w1375 & ~w11372;
assign w14720 = pi0148 & w5274;
assign w14721 = w1127 & ~w15451;
assign w14722 = (~pi0982 & ~w13509) | (~pi0982 & w4625) | (~w13509 & w4625);
assign w14723 = w13509 & w5773;
assign w14724 = w13509 & w1652;
assign w14725 = (pi1110 & ~w13509) | (pi1110 & w12328) | (~w13509 & w12328);
assign w14726 = ~pi3047 & w6463;
assign w14727 = pi3074 & ~pi3133;
assign w14728 = pi0006 & ~w14148;
assign w14729 = w14648 & ~pi2731;
assign w14730 = pi2639 & ~w3555;
assign w14731 = pi1484 & ~w9781;
assign w14732 = ~w716 & w17615;
assign w14733 = pi2441 & ~w4508;
assign w14734 = ~w11593 & ~w12048;
assign w14735 = ~w1711 & ~w11397;
assign w14736 = ~w10300 & ~w3501;
assign w14737 = ~w18222 & ~w14702;
assign w14738 = pi0263 & pi0303;
assign w14739 = w17665 & w12680;
assign w14740 = ~w4144 & ~w7739;
assign w14741 = (~pi1260 & ~w545) | (~pi1260 & w14378) | (~w545 & w14378);
assign w14742 = pi2998 & w6263;
assign w14743 = ~pi3159 & w13730;
assign w14744 = ~w15808 & pi0743;
assign w14745 = w9440 & pi0158;
assign w14746 = ~w5267 & ~w14984;
assign w14747 = ~pi3293 & w18259;
assign w14748 = w5453 & pi2578;
assign w14749 = ~pi0331 & w4058;
assign w14750 = ~pi0045 & ~w9240;
assign w14751 = pi2137 & ~w15883;
assign w14752 = ~w7790 & ~w4631;
assign w14753 = ~w4020 & w18123;
assign w14754 = w13509 & w10497;
assign w14755 = (~pi0247 & ~w325) | (~pi0247 & w15493) | (~w325 & w15493);
assign w14756 = pi1621 & ~w7090;
assign w14757 = ~pi1190 & w543;
assign w14758 = ~w1391 & pi1038;
assign w14759 = ~w9988 & ~w9737;
assign w14760 = pi1634 & ~w18259;
assign w14761 = pi2647 & ~w3555;
assign w14762 = pi2642 & ~w261;
assign w14763 = pi3153 & w8829;
assign w14764 = ~pi2987 & w9504;
assign w14765 = ~w14019 & ~w9088;
assign w14766 = (pi0839 & ~w13509) | (pi0839 & w7190) | (~w13509 & w7190);
assign w14767 = pi1678 & ~w6499;
assign w14768 = ~w97 & ~w915;
assign w14769 = w16278 & ~w6033;
assign w14770 = w5189 & ~w2741;
assign w14771 = ~w14451 & ~w498;
assign w14772 = pi2425 & ~w15271;
assign w14773 = w13004 & w13867;
assign w14774 = ~w9233 & ~w10188;
assign w14775 = pi1772 & ~pi3133;
assign w14776 = w13509 & w16206;
assign w14777 = pi1248 & w11655;
assign w14778 = w13509 & w1613;
assign w14779 = w13509 & w4442;
assign w14780 = ~w3821 & ~w6739;
assign w14781 = pi1468 & ~w7090;
assign w14782 = w5642 & w12476;
assign w14783 = pi0339 & pi2967;
assign w14784 = ~w3203 & pi0591;
assign w14785 = ~w4527 & ~w11703;
assign w14786 = pi1923 & ~w7177;
assign w14787 = ~w289 & ~w17726;
assign w14788 = ~w13728 & ~w130;
assign w14789 = ~w6697 & pi0674;
assign w14790 = pi3082 & w9504;
assign w14791 = w14076 & w6730;
assign w14792 = w15064 & w17626;
assign w14793 = w10189 & ~pi0479;
assign w14794 = ~w18333 & ~w2126;
assign w14795 = (pi0709 & ~w13509) | (pi0709 & w9278) | (~w13509 & w9278);
assign w14796 = ~w18197 & ~w13805;
assign w14797 = ~pi0626 & w14641;
assign w14798 = ~w9573 & ~w10542;
assign w14799 = w1391 & ~w12800;
assign w14800 = ~pi2981 & pi1357;
assign w14801 = pi1497 & ~w16922;
assign w14802 = ~pi0282 & w4058;
assign w14803 = w2809 & w4840;
assign w14804 = pi2585 & ~w5274;
assign w14805 = pi2020 & ~w14833;
assign w14806 = ~pi0887 & w1126;
assign w14807 = pi0175 & w5274;
assign w14808 = ~pi0861 & w15707;
assign w14809 = ~w5189 & pi1101;
assign w14810 = w11760 & ~pi3369;
assign w14811 = w13509 & w9022;
assign w14812 = ~w18041 & w10163;
assign w14813 = pi2442 & ~w10299;
assign w14814 = pi0262 & pi0302;
assign w14815 = pi1386 & ~w17935;
assign w14816 = w934 & pi0422;
assign w14817 = ~w15122 & ~pi2775;
assign w14818 = ~w4365 & ~w10093;
assign w14819 = ~w12881 & w1326;
assign w14820 = w13509 & w9555;
assign w14821 = ~w8588 & w17646;
assign w14822 = ~w17300 & ~w464;
assign w14823 = pi3138 & w2732;
assign w14824 = w13509 & w16668;
assign w14825 = ~w1083 & w7356;
assign w14826 = w16278 & ~w1340;
assign w14827 = pi2465 & pi3125;
assign w14828 = pi1363 & w6297;
assign w14829 = w11671 & w3515;
assign w14830 = ~w35 & ~w14496;
assign w14831 = w3203 & ~w3374;
assign w14832 = w17844 & w3833;
assign w14833 = w10635 & w14244;
assign w14834 = (pi0592 & ~w13509) | (pi0592 & w17065) | (~w13509 & w17065);
assign w14835 = pi2593 & ~w7017;
assign w14836 = ~w588 & ~w16629;
assign w14837 = ~pi3314 & w7090;
assign w14838 = ~w15270 & ~w3009;
assign w14839 = (~w13165 & ~w5517) | (~w13165 & w11013) | (~w5517 & w11013);
assign w14840 = ~pi3051 & pi3158;
assign w14841 = pi3160 & ~w858;
assign w14842 = w14782 & w126;
assign w14843 = pi0435 & w17173;
assign w14844 = ~w18601 & w13913;
assign w14845 = w17665 & ~w17967;
assign w14846 = ~pi2125 & w16041;
assign w14847 = ~pi0428 & w6928;
assign w14848 = ~pi2357 & w12755;
assign w14849 = pi2373 & ~w412;
assign w14850 = ~w11069 & ~w6232;
assign w14851 = ~w3151 & ~w68;
assign w14852 = ~pi3113 & pi3150;
assign w14853 = pi2929 & ~w226;
assign w14854 = (pi1885 & w2014) | (pi1885 & w10829) | (w2014 & w10829);
assign w14855 = w3243 & w9511;
assign w14856 = w13328 & w7183;
assign w14857 = ~pi3094 & w6463;
assign w14858 = ~w8357 & w6854;
assign w14859 = ~w18073 & ~w8916;
assign w14860 = ~w17619 & ~pi0508;
assign w14861 = ~pi2891 & w17213;
assign w14862 = ~pi0603 & w12825;
assign w14863 = pi1657 & ~w6072;
assign w14864 = ~pi3138 & w1843;
assign w14865 = ~pi0681 & w9110;
assign w14866 = ~w6697 & pi1014;
assign w14867 = w4599 & w840;
assign w14868 = ~pi0874 & w1126;
assign w14869 = ~w18042 & ~w16931;
assign w14870 = ~pi3155 & w15839;
assign w14871 = ~w7881 & ~w4730;
assign w14872 = ~w10719 & w6918;
assign w14873 = ~w18191 & w13058;
assign w14874 = ~w2086 & ~w15110;
assign w14875 = ~w10600 & ~w6391;
assign w14876 = ~w13433 & ~w1084;
assign w14877 = pi3078 & ~pi3143;
assign w14878 = ~w17665 & ~w9943;
assign w14879 = ~pi0508 & ~pi1345;
assign w14880 = ~w11491 & ~w14936;
assign w14881 = ~w12803 & ~w18171;
assign w14882 = ~w10632 & ~w15554;
assign w14883 = pi2102 & ~w4420;
assign w14884 = pi1931 & ~w15271;
assign w14885 = (pi0681 & ~w13509) | (pi0681 & w4882) | (~w13509 & w4882);
assign w14886 = w13509 & w14513;
assign w14887 = ~w12460 & w7013;
assign w14888 = ~pi2049 & w13204;
assign w14889 = pi3136 & w7946;
assign w14890 = ~w16280 & ~w9054;
assign w14891 = w5453 & pi2590;
assign w14892 = ~pi1025 & w3106;
assign w14893 = w14404 & w4974;
assign w14894 = (pi0913 & ~w13509) | (pi0913 & w5060) | (~w13509 & w5060);
assign w14895 = ~w3190 & ~w9262;
assign w14896 = ~w7904 & w14038;
assign w14897 = pi1490 & w13753;
assign w14898 = ~w6507 & ~w15851;
assign w14899 = w8832 & w17250;
assign w14900 = ~w17317 & ~w1779;
assign w14901 = w560 & w4276;
assign w14902 = ~w16027 & ~w333;
assign w14903 = w7742 & w6255;
assign w14904 = ~pi3157 & pi3207;
assign w14905 = ~pi3133 & w13730;
assign w14906 = ~w4436 & ~w7991;
assign w14907 = ~w7077 & pi1067;
assign w14908 = (w5435 & ~w7631) | (w5435 & w12958) | (~w7631 & w12958);
assign w14909 = w11209 & ~w410;
assign w14910 = w13509 & w1725;
assign w14911 = ~w13367 & w13996;
assign w14912 = w7307 & w11212;
assign w14913 = ~w1566 & w8648;
assign w14914 = ~w7883 & ~w13346;
assign w14915 = ~pi1938 & w11688;
assign w14916 = ~w17556 & ~w7848;
assign w14917 = ~w16214 & ~w7785;
assign w14918 = ~pi1371 & w11399;
assign w14919 = ~w5523 & ~w16102;
assign w14920 = pi1867 & ~w458;
assign w14921 = ~w8781 & ~w14889;
assign w14922 = ~w6398 & ~w9785;
assign w14923 = ~w2794 & w5187;
assign w14924 = pi0108 & w3748;
assign w14925 = ~pi2362 & w12755;
assign w14926 = ~w8588 & w4508;
assign w14927 = w6109 & ~pi1241;
assign w14928 = w7307 & w8533;
assign w14929 = pi2056 & ~w10158;
assign w14930 = (~pi0265 & ~w18262) | (~pi0265 & w16958) | (~w18262 & w16958);
assign w14931 = ~w1368 & ~pi0459;
assign w14932 = ~w11324 & ~w13234;
assign w14933 = pi1357 & ~w13786;
assign w14934 = ~w836 & ~w14439;
assign w14935 = w6605 & w7516;
assign w14936 = ~pi0500 & pi1156;
assign w14937 = ~pi1119 & w3791;
assign w14938 = ~pi3316 & w9781;
assign w14939 = w2560 & w18573;
assign w14940 = ~w3000 & ~pi2666;
assign w14941 = w13509 & w16;
assign w14942 = ~pi3341 & w7090;
assign w14943 = w5437 & w381;
assign w14944 = ~pi3048 & w6463;
assign w14945 = ~w14140 & w16732;
assign w14946 = ~w16149 & ~w13049;
assign w14947 = ~w7998 & ~w7971;
assign w14948 = ~w14648 & ~pi2652;
assign w14949 = w17248 & ~w1236;
assign w14950 = pi2796 & ~w15235;
assign w14951 = w6447 & w11545;
assign w14952 = ~pi1038 & w6200;
assign w14953 = w539 & ~w16853;
assign w14954 = ~pi3171 & w3805;
assign w14955 = pi0443 & w6090;
assign w14956 = w16844 & w16956;
assign w14957 = w11209 & ~w9027;
assign w14958 = pi2379 & ~w4508;
assign w14959 = w6857 & w1193;
assign w14960 = pi0258 & w5113;
assign w14961 = pi3167 & w15106;
assign w14962 = ~pi2657 & w17213;
assign w14963 = ~w18156 & ~w14977;
assign w14964 = ~pi2076 & w17439;
assign w14965 = pi0177 & w5274;
assign w14966 = ~pi3354 & w14918;
assign w14967 = pi0060 & ~w14148;
assign w14968 = ~w15460 & ~w16261;
assign w14969 = w9720 & pi1713;
assign w14970 = pi0429 & ~w2165;
assign w14971 = w13606 & w512;
assign w14972 = ~w5125 & ~w9365;
assign w14973 = ~pi0614 & w14641;
assign w14974 = ~w17665 & ~w17837;
assign w14975 = ~w13030 & ~w2049;
assign w14976 = pi1742 & ~w4058;
assign w14977 = w8098 & w15470;
assign w14978 = ~w3592 & ~w11448;
assign w14979 = (pi0929 & ~w13509) | (pi0929 & w11066) | (~w13509 & w11066);
assign w14980 = w9227 & w12817;
assign w14981 = ~w10856 & w528;
assign w14982 = w6649 & ~w1129;
assign w14983 = w16506 & ~w6033;
assign w14984 = ~pi0171 & pi0177;
assign w14985 = pi1656 & ~w6072;
assign w14986 = w7961 & w1209;
assign w14987 = ~pi1165 & pi3216;
assign w14988 = (pi1108 & ~w13509) | (pi1108 & w16431) | (~w13509 & w16431);
assign w14989 = ~w16764 & w17464;
assign w14990 = ~w1631 & w17771;
assign w14991 = w14782 & w13763;
assign w14992 = pi0335 & ~pi0337;
assign w14993 = ~w6104 & ~w11740;
assign w14994 = ~w6123 & ~w6496;
assign w14995 = w3203 & ~w15296;
assign w14996 = ~w3006 & ~w8079;
assign w14997 = w7703 & w6578;
assign w14998 = w16127 & w16079;
assign w14999 = (pi0399 & w5560) | (pi0399 & w1380) | (w5560 & w1380);
assign w15000 = ~w13717 & ~w17661;
assign w15001 = ~w11713 & ~w18356;
assign w15002 = w7307 & w15757;
assign w15003 = ~pi1691 & w13343;
assign w15004 = w5189 & ~w6647;
assign w15005 = ~pi0899 & w14641;
assign w15006 = w12040 & ~w14465;
assign w15007 = ~pi3169 & w17669;
assign w15008 = w11644 & w14101;
assign w15009 = pi2913 & pi1211;
assign w15010 = pi1784 & ~w15767;
assign w15011 = w17814 & w16545;
assign w15012 = w17248 & ~w6647;
assign w15013 = ~w5551 & w10105;
assign w15014 = ~w15502 & ~w7065;
assign w15015 = pi3134 & w3987;
assign w15016 = ~pi3131 & w17669;
assign w15017 = (pi1080 & ~w13509) | (pi1080 & w4423) | (~w13509 & w4423);
assign w15018 = ~w7845 & ~w15141;
assign w15019 = ~w17898 & w10951;
assign w15020 = ~pi0545 & w795;
assign w15021 = ~pi0483 & pi3380;
assign w15022 = pi3025 & ~w3987;
assign w15023 = ~w3230 & ~w17942;
assign w15024 = (pi0864 & ~w13509) | (pi0864 & w16450) | (~w13509 & w16450);
assign w15025 = ~w10167 & ~w3563;
assign w15026 = pi0057 & w922;
assign w15027 = w2494 & w2867;
assign w15028 = ~pi3086 & w9504;
assign w15029 = ~w1433 & w12571;
assign w15030 = pi2620 & ~w16815;
assign w15031 = ~pi0289 & w2196;
assign w15032 = ~w14308 & ~w16837;
assign w15033 = w12040 & ~w4179;
assign w15034 = w16506 & ~w16498;
assign w15035 = pi3035 & ~pi3145;
assign w15036 = w11345 & w9063;
assign w15037 = ~w17781 & w1816;
assign w15038 = ~w17409 & ~w11223;
assign w15039 = pi1513 & w13753;
assign w15040 = ~w6195 & w13001;
assign w15041 = ~w11336 & ~w10254;
assign w15042 = pi1456 & ~w7090;
assign w15043 = ~w14782 & w1560;
assign w15044 = ~pi3131 & w11701;
assign w15045 = pi1562 & ~w13753;
assign w15046 = ~w15728 & ~w3854;
assign w15047 = w8789 & ~pi0393;
assign w15048 = ~w4020 & w17646;
assign w15049 = pi2531 & w14148;
assign w15050 = ~w4283 & ~w16391;
assign w15051 = ~pi0507 & ~pi1345;
assign w15052 = pi2825 & ~w16815;
assign w15053 = pi2016 & ~w14833;
assign w15054 = ~w9911 & ~w4564;
assign w15055 = pi2353 & ~w412;
assign w15056 = ~w4654 & ~w12894;
assign w15057 = pi1853 & ~w2732;
assign w15058 = ~w7656 & ~pi1221;
assign w15059 = ~pi3068 & pi3159;
assign w15060 = w14899 & w13622;
assign w15061 = ~w14228 & pi0614;
assign w15062 = pi0117 & w3748;
assign w15063 = (w10183 & w4903) | (w10183 & w2902) | (w4903 & w2902);
assign w15064 = w14782 & w852;
assign w15065 = ~w9931 & ~w15049;
assign w15066 = pi1710 & ~pi3143;
assign w15067 = ~w883 & ~w7216;
assign w15068 = ~w18182 & ~w13298;
assign w15069 = pi1756 & ~w15767;
assign w15070 = ~w11681 & ~w12789;
assign w15071 = ~pi0128 & pi1220;
assign w15072 = w12423 & w16655;
assign w15073 = w8337 & pi3327;
assign w15074 = ~w3210 & ~w16190;
assign w15075 = ~w4382 & w6986;
assign w15076 = w8789 & w11653;
assign w15077 = ~w17653 & ~w423;
assign w15078 = ~w709 & pi1282;
assign w15079 = ~w7054 & ~w4718;
assign w15080 = w8658 & pi1785;
assign w15081 = w1858 & w7824;
assign w15082 = ~w18040 & ~w973;
assign w15083 = ~w2725 & pi0793;
assign w15084 = w11743 & ~w18315;
assign w15085 = ~w6697 & pi0659;
assign w15086 = w13509 & w16660;
assign w15087 = pi0247 & w5113;
assign w15088 = ~pi0139 & pi1878;
assign w15089 = pi1474 & ~w9781;
assign w15090 = ~w2875 & ~w4062;
assign w15091 = w5189 & ~w17210;
assign w15092 = ~w14122 & ~w16262;
assign w15093 = ~w10503 & ~w1707;
assign w15094 = ~pi3318 & w6448;
assign w15095 = w5189 & ~w13028;
assign w15096 = w7307 & w11727;
assign w15097 = ~w12623 & ~w832;
assign w15098 = ~w15924 & ~w16208;
assign w15099 = ~w13231 & pi0572;
assign w15100 = ~w8643 & ~w18285;
assign w15101 = ~w4059 & ~w3547;
assign w15102 = pi1172 & ~w13509;
assign w15103 = w5189 & ~w14597;
assign w15104 = pi1485 & ~w9781;
assign w15105 = ~w16020 & ~w12247;
assign w15106 = pi2943 & ~pi3123;
assign w15107 = ~w5560 & w18022;
assign w15108 = ~w2418 & ~w677;
assign w15109 = ~w3041 & ~w4907;
assign w15110 = ~pi2457 & w9340;
assign w15111 = w5437 & w13384;
assign w15112 = ~w9650 & ~w14290;
assign w15113 = ~w14376 & w3768;
assign w15114 = ~w13347 & ~w15358;
assign w15115 = w11383 & w6334;
assign w15116 = w10189 & ~pi0455;
assign w15117 = ~w13910 & ~w12506;
assign w15118 = ~w14248 & ~w16751;
assign w15119 = ~pi3020 & pi3109;
assign w15120 = ~w11078 & ~w12049;
assign w15121 = ~w3445 & ~w2711;
assign w15122 = ~w10373 & ~w7483;
assign w15123 = w17057 & w18084;
assign w15124 = ~w16678 & ~w16031;
assign w15125 = ~pi2368 & w12941;
assign w15126 = w9424 & w16582;
assign w15127 = w1962 & ~w305;
assign w15128 = w5437 & w17606;
assign w15129 = (pi1081 & ~w13509) | (pi1081 & w3869) | (~w13509 & w3869);
assign w15130 = (pi1048 & ~w13509) | (pi1048 & w6634) | (~w13509 & w6634);
assign w15131 = pi1487 & ~w9781;
assign w15132 = ~w5246 & ~w9877;
assign w15133 = w8337 & pi3310;
assign w15134 = w709 & pi1888;
assign w15135 = w2341 & ~w2776;
assign w15136 = w2591 & w2201;
assign w15137 = ~pi1910 & w5384;
assign w15138 = ~w14073 & w9303;
assign w15139 = ~w4463 & ~w1423;
assign w15140 = (pi0910 & ~w13509) | (pi0910 & w15810) | (~w13509 & w15810);
assign w15141 = ~pi3318 & w14918;
assign w15142 = (pi0197 & ~w10992) | (pi0197 & w13579) | (~w10992 & w13579);
assign w15143 = ~pi0665 & w12197;
assign w15144 = ~w17662 & ~w17855;
assign w15145 = ~pi3133 & w12427;
assign w15146 = w625 & w2547;
assign w15147 = (pi1064 & ~w13509) | (pi1064 & w10415) | (~w13509 & w10415);
assign w15148 = ~w10032 & ~w14615;
assign w15149 = ~pi0737 & w17899;
assign w15150 = (pi0793 & ~w13509) | (pi0793 & w15083) | (~w13509 & w15083);
assign w15151 = ~w6175 & ~w11000;
assign w15152 = pi2566 & ~w5274;
assign w15153 = ~w3334 & ~w1259;
assign w15154 = ~w10346 & ~w3525;
assign w15155 = ~w8709 & w16811;
assign w15156 = w11383 & w3627;
assign w15157 = (pi0883 & ~w13509) | (pi0883 & w5881) | (~w13509 & w5881);
assign w15158 = w10762 & w269;
assign w15159 = ~pi2027 & w7455;
assign w15160 = ~w2449 & w18518;
assign w15161 = ~w7277 & ~w13546;
assign w15162 = w11345 & w15841;
assign w15163 = ~pi3165 & w4310;
assign w15164 = ~w15808 & pi0919;
assign w15165 = (pi1126 & ~w13509) | (pi1126 & w10515) | (~w13509 & w10515);
assign w15166 = ~w16165 & ~w5472;
assign w15167 = ~w3039 & ~w17120;
assign w15168 = ~pi3100 & w15235;
assign w15169 = ~w11146 & ~w15989;
assign w15170 = pi1617 & ~w13753;
assign w15171 = ~w14397 & ~w2982;
assign w15172 = pi2603 & ~w16815;
assign w15173 = ~w10585 & ~w10911;
assign w15174 = ~w14542 & w7804;
assign w15175 = pi2935 & ~w6045;
assign w15176 = w7698 & w254;
assign w15177 = ~pi0788 & w543;
assign w15178 = pi2828 & ~w3555;
assign w15179 = w14648 & ~pi2614;
assign w15180 = pi0494 & pi0511;
assign w15181 = ~pi3172 & w13730;
assign w15182 = ~w6785 & pi0870;
assign w15183 = w11345 & w3307;
assign w15184 = (pi0362 & w6195) | (pi0362 & w16612) | (w6195 & w16612);
assign w15185 = w11383 & w14729;
assign w15186 = w8658 & pi1795;
assign w15187 = ~w15024 & ~w8266;
assign w15188 = w15558 & w15302;
assign w15189 = w13509 & w6157;
assign w15190 = ~pi0684 & w9110;
assign w15191 = w16893 & w8238;
assign w15192 = ~w1312 & w2460;
assign w15193 = pi2237 & ~w11735;
assign w15194 = w7844 & w11302;
assign w15195 = ~w2443 & ~w10265;
assign w15196 = pi2099 & ~w4420;
assign w15197 = w15122 & ~pi2636;
assign w15198 = pi1488 & w13753;
assign w15199 = (pi0870 & ~w13509) | (pi0870 & w15182) | (~w13509 & w15182);
assign w15200 = w13509 & w1625;
assign w15201 = pi2709 & ~w9504;
assign w15202 = pi1770 & pi1810;
assign w15203 = pi0306 & ~pi0307;
assign w15204 = (pi0797 & ~w13509) | (pi0797 & w6937) | (~w13509 & w6937);
assign w15205 = ~w7283 & ~w9170;
assign w15206 = pi3174 & pi3348;
assign w15207 = pi2744 & ~w11406;
assign w15208 = (w4836 & w9096) | (w4836 & w548) | (w9096 & w548);
assign w15209 = ~pi3298 & w6448;
assign w15210 = ~pi1993 & w3019;
assign w15211 = ~pi0491 & ~pi1345;
assign w15212 = ~w11622 & w11120;
assign w15213 = pi3001 & w18047;
assign w15214 = pi1439 & ~w6448;
assign w15215 = w13509 & w9469;
assign w15216 = w13509 & w12088;
assign w15217 = w4240 & w18012;
assign w15218 = ~pi1699 & w4667;
assign w15219 = ~pi3168 & pi3207;
assign w15220 = pi3169 & pi3207;
assign w15221 = ~w17974 & w8018;
assign w15222 = pi2680 & ~w11406;
assign w15223 = w233 & w12501;
assign w15224 = w4312 & ~w11879;
assign w15225 = ~pi2056 & w13204;
assign w15226 = ~w8203 & ~w7184;
assign w15227 = ~pi3424 & w15036;
assign w15228 = w13509 & w17248;
assign w15229 = ~pi0856 & w15707;
assign w15230 = pi3136 & w3987;
assign w15231 = ~w6195 & w17720;
assign w15232 = w17433 & w9231;
assign w15233 = pi2722 & ~w9504;
assign w15234 = w5189 & w11302;
assign w15235 = w1804 & w12686;
assign w15236 = ~pi3153 & w11132;
assign w15237 = pi0016 & ~w3748;
assign w15238 = ~w4977 & ~w4704;
assign w15239 = ~pi3000 & ~pi3207;
assign w15240 = w9440 & pi0146;
assign w15241 = ~w5590 & ~w12293;
assign w15242 = w7388 & w12854;
assign w15243 = ~pi2128 & w16041;
assign w15244 = (w2460 & ~w11232) | (w2460 & w5170) | (~w11232 & w5170);
assign w15245 = pi1337 & pi0306;
assign w15246 = ~pi2207 & w5075;
assign w15247 = ~w7378 & ~w12214;
assign w15248 = pi2555 & ~w5274;
assign w15249 = ~pi3163 & w11132;
assign w15250 = pi1778 & pi0085;
assign w15251 = ~w9144 & ~w14209;
assign w15252 = ~pi1693 & ~w8869;
assign w15253 = w6379 & w14693;
assign w15254 = ~pi2117 & w12755;
assign w15255 = ~pi1681 & ~w7177;
assign w15256 = pi1682 & ~w7177;
assign w15257 = ~w2366 & ~w6196;
assign w15258 = ~w8413 & ~w717;
assign w15259 = w17248 & ~w6033;
assign w15260 = w9720 & pi1718;
assign w15261 = ~w889 & ~w14663;
assign w15262 = pi2249 & ~w4420;
assign w15263 = ~w1368 & ~pi0462;
assign w15264 = ~pi0720 & w17899;
assign w15265 = ~w6160 & ~w15174;
assign w15266 = w4508 & w14078;
assign w15267 = w12040 & ~w13028;
assign w15268 = ~w5177 & ~w1175;
assign w15269 = w6697 & ~w6680;
assign w15270 = pi1132 & pi2938;
assign w15271 = w10635 & w7140;
assign w15272 = w10818 & ~w6153;
assign w15273 = w13509 & w2430;
assign w15274 = pi1223 & ~w5768;
assign w15275 = ~w5577 & w12580;
assign w15276 = (pi1259 & w302) | (pi1259 & w8733) | (w302 & w8733);
assign w15277 = ~w11760 & ~w14385;
assign w15278 = w11046 & w1789;
assign w15279 = ~w18309 & ~w10422;
assign w15280 = ~pi0701 & w3106;
assign w15281 = ~w3355 & w4590;
assign w15282 = ~pi0589 & w795;
assign w15283 = ~w7844 & pi0604;
assign w15284 = pi2457 & ~w10299;
assign w15285 = ~pi3133 & w11132;
assign w15286 = ~w13080 & ~w17325;
assign w15287 = pi2807 & ~w11406;
assign w15288 = ~pi1205 & w15707;
assign w15289 = ~w3941 & ~w17702;
assign w15290 = pi1379 & pi3160;
assign w15291 = ~w13250 & ~w1322;
assign w15292 = pi1242 & pi1229;
assign w15293 = pi2544 & w605;
assign w15294 = ~w9009 & ~w7141;
assign w15295 = ~w1962 & pi0643;
assign w15296 = ~w17344 & ~w14114;
assign w15297 = ~w5453 & ~pi1797;
assign w15298 = ~pi0921 & w17490;
assign w15299 = ~w3203 & ~pi0954;
assign w15300 = ~w16859 & ~w13248;
assign w15301 = ~pi0497 & ~pi1191;
assign w15302 = w9722 & w17995;
assign w15303 = ~pi3093 & w9504;
assign w15304 = ~w18509 & ~w5770;
assign w15305 = pi1722 & ~w8113;
assign w15306 = ~w5150 & ~w7886;
assign w15307 = ~w4409 & w17264;
assign w15308 = pi3162 & w619;
assign w15309 = pi1212 & ~pi1221;
assign w15310 = ~w18599 & ~w7355;
assign w15311 = ~pi3295 & w9781;
assign w15312 = pi0107 & w9284;
assign w15313 = ~w5052 & ~w10885;
assign w15314 = pi2024 & ~w17646;
assign w15315 = ~w7948 & ~w6821;
assign w15316 = ~pi3164 & w13570;
assign w15317 = ~w1791 & w3206;
assign w15318 = w13509 & w906;
assign w15319 = w15450 & ~w12297;
assign w15320 = ~pi0796 & w543;
assign w15321 = pi2654 & ~w15235;
assign w15322 = ~pi3036 & w16502;
assign w15323 = ~w18342 & w801;
assign w15324 = ~w16978 & ~w9419;
assign w15325 = w13509 & w11725;
assign w15326 = ~w12040 & pi1022;
assign w15327 = w1946 & pi0249;
assign w15328 = ~w13280 & ~w6863;
assign w15329 = w14537 & w3985;
assign w15330 = ~pi0997 & w795;
assign w15331 = (pi0707 & ~w13509) | (pi0707 & w12444) | (~w13509 & w12444);
assign w15332 = ~w2341 & pi1047;
assign w15333 = ~pi1236 & ~pi1237;
assign w15334 = ~w2185 & ~w16989;
assign w15335 = w15717 & ~w1575;
assign w15336 = ~pi3153 & w8515;
assign w15337 = ~w16920 & ~w13560;
assign w15338 = pi1396 & w12285;
assign w15339 = ~w14228 & pi0619;
assign w15340 = ~w3000 & ~pi2753;
assign w15341 = w6639 & w10421;
assign w15342 = ~pi3170 & ~w1793;
assign w15343 = pi0095 & w3748;
assign w15344 = w8692 & w5133;
assign w15345 = ~w8670 & ~w12553;
assign w15346 = ~pi0878 & w1126;
assign w15347 = (pi1202 & w4470) | (pi1202 & w8555) | (w4470 & w8555);
assign w15348 = pi1960 & ~w14833;
assign w15349 = ~pi1265 & w10552;
assign w15350 = ~pi1677 & w17562;
assign w15351 = w1381 & w12950;
assign w15352 = ~w3431 & ~w18071;
assign w15353 = ~pi1170 & ~pi3192;
assign w15354 = pi1135 & w9420;
assign w15355 = pi1523 & w13753;
assign w15356 = ~pi3164 & w15839;
assign w15357 = w7799 & w3278;
assign w15358 = ~w1273 & w14153;
assign w15359 = ~w7775 & ~w1703;
assign w15360 = ~pi2045 & w13204;
assign w15361 = ~pi3337 & w7090;
assign w15362 = ~w6759 & ~w679;
assign w15363 = w16861 & w7293;
assign w15364 = ~pi3150 & w11132;
assign w15365 = ~w11002 & ~w14095;
assign w15366 = w13509 & w6779;
assign w15367 = pi3168 & w18497;
assign w15368 = ~w14864 & ~w11558;
assign w15369 = ~pi2705 & ~pi2966;
assign w15370 = w15808 & ~w17210;
assign w15371 = ~pi1080 & w795;
assign w15372 = ~w5936 & ~w15308;
assign w15373 = ~w6697 & pi1111;
assign w15374 = ~w14728 & ~w16168;
assign w15375 = pi1571 & ~w13753;
assign w15376 = pi2173 & ~w15271;
assign w15377 = ~w6351 & ~w6089;
assign w15378 = pi3143 & w2253;
assign w15379 = ~w4667 & ~w302;
assign w15380 = ~w2435 & ~w6400;
assign w15381 = (pi1173 & ~w13509) | (pi1173 & w1167) | (~w13509 & w1167);
assign w15382 = ~pi0443 & w17173;
assign w15383 = w7799 & w11721;
assign w15384 = w12040 & ~w4043;
assign w15385 = ~w6291 & ~w17009;
assign w15386 = w11383 & w4504;
assign w15387 = ~w5937 & ~w4008;
assign w15388 = ~pi3145 & w13730;
assign w15389 = ~w16161 & pi0000;
assign w15390 = w17969 & w8922;
assign w15391 = ~w14723 & ~w2419;
assign w15392 = ~pi1353 & ~w8804;
assign w15393 = ~w7932 & ~w11596;
assign w15394 = ~pi3139 & w3805;
assign w15395 = w6785 & w15609;
assign w15396 = w11010 & w1864;
assign w15397 = ~w1124 & ~w12243;
assign w15398 = w551 & ~pi1219;
assign w15399 = ~pi1117 & w3791;
assign w15400 = ~w1798 & w4380;
assign w15401 = w14103 & w13865;
assign w15402 = (pi0556 & ~w13509) | (pi0556 & w10205) | (~w13509 & w10205);
assign w15403 = ~w12441 & ~w2164;
assign w15404 = pi1245 & ~w11655;
assign w15405 = w10818 & ~w8700;
assign w15406 = ~pi3104 & w16502;
assign w15407 = ~w8530 & ~w10233;
assign w15408 = pi2194 & ~w10299;
assign w15409 = ~w9391 & ~w10770;
assign w15410 = ~w14141 & ~w1241;
assign w15411 = ~w14073 & w10290;
assign w15412 = w9440 & pi0190;
assign w15413 = ~w8050 & ~w17385;
assign w15414 = ~w2819 & ~w9735;
assign w15415 = ~w1368 & ~pi0468;
assign w15416 = ~w15222 & ~w11428;
assign w15417 = pi0975 & pi0076;
assign w15418 = ~w8090 & ~w13991;
assign w15419 = ~pi1152 & pi1176;
assign w15420 = w6649 & ~w4785;
assign w15421 = ~w16281 & ~w1774;
assign w15422 = ~pi0920 & w12197;
assign w15423 = ~pi3133 & w1843;
assign w15424 = ~w7608 & w12885;
assign w15425 = ~w5568 & ~w2411;
assign w15426 = ~pi3090 & w16815;
assign w15427 = pi1179 & ~w14073;
assign w15428 = ~w2148 & ~w2693;
assign w15429 = (pi0002 & ~w10992) | (pi0002 & w6460) | (~w10992 & w6460);
assign w15430 = ~w2292 & ~w10251;
assign w15431 = pi2837 & ~w11406;
assign w15432 = ~w14757 & ~w14522;
assign w15433 = ~w14283 & ~w3964;
assign w15434 = w14109 & pi0421;
assign w15435 = ~pi3337 & w17935;
assign w15436 = ~pi3104 & ~w3987;
assign w15437 = w13509 & w13066;
assign w15438 = ~pi2987 & w3555;
assign w15439 = ~w4831 & ~w15273;
assign w15440 = pi1398 & w13753;
assign w15441 = w6649 & ~w1018;
assign w15442 = pi1386 & w13753;
assign w15443 = pi2447 & ~w10299;
assign w15444 = ~w3000 & ~pi2809;
assign w15445 = (pi1008 & ~w13509) | (pi1008 & w14567) | (~w13509 & w14567);
assign w15446 = pi0029 & ~w3748;
assign w15447 = pi2296 & ~w3223;
assign w15448 = ~w3395 & ~w4760;
assign w15449 = ~pi2077 & w17439;
assign w15450 = pi0134 & ~pi3206;
assign w15451 = pi1392 & w13753;
assign w15452 = w3988 & w13344;
assign w15453 = ~w4997 & ~w12005;
assign w15454 = w7703 & w12979;
assign w15455 = pi2012 & ~w14833;
assign w15456 = ~w2014 & w4581;
assign w15457 = w13509 & w14500;
assign w15458 = w934 & pi0417;
assign w15459 = ~pi3151 & ~pi3160;
assign w15460 = ~pi1175 & ~pi3209;
assign w15461 = pi2028 & ~w17646;
assign w15462 = (~pi0960 & ~w13509) | (~pi0960 & w13215) | (~w13509 & w13215);
assign w15463 = pi2661 & ~w15235;
assign w15464 = pi3162 & w15767;
assign w15465 = ~w17552 & w14018;
assign w15466 = w1820 & w11885;
assign w15467 = pi1438 & ~w13753;
assign w15468 = ~pi1231 & pi1267;
assign w15469 = ~pi3142 & w15048;
assign w15470 = w5383 & pi1396;
assign w15471 = (pi0675 & ~w13509) | (pi0675 & w17393) | (~w13509 & w17393);
assign w15472 = pi1866 & ~w15036;
assign w15473 = w16893 & w8091;
assign w15474 = w9903 & w9559;
assign w15475 = ~w469 & ~w450;
assign w15476 = w6385 & w14791;
assign w15477 = pi1557 & ~w13753;
assign w15478 = ~w3133 & ~w1035;
assign w15479 = ~w2645 & ~w5021;
assign w15480 = ~w8813 & ~w15930;
assign w15481 = ~pi3055 & w16815;
assign w15482 = w384 & w17634;
assign w15483 = pi1148 & w9420;
assign w15484 = w412 & w614;
assign w15485 = w384 & w10535;
assign w15486 = ~w6785 & pi0985;
assign w15487 = ~w16382 & ~w16273;
assign w15488 = w1962 & ~w2741;
assign w15489 = w10158 & w9407;
assign w15490 = w13509 & w18372;
assign w15491 = pi3006 & ~w16502;
assign w15492 = (pi1031 & ~w13509) | (pi1031 & w584) | (~w13509 & w584);
assign w15493 = pi1337 & ~pi0247;
assign w15494 = ~w2483 & ~w12729;
assign w15495 = pi1872 & ~w458;
assign w15496 = w13509 & w18460;
assign w15497 = pi2476 & ~w14524;
assign w15498 = ~pi3313 & w14918;
assign w15499 = pi3116 & ~pi3132;
assign w15500 = pi0066 & ~w14148;
assign w15501 = ~pi1113 & w3791;
assign w15502 = ~pi3163 & w13730;
assign w15503 = ~pi1754 & pi3162;
assign w15504 = w11232 & w17545;
assign w15505 = (pi0748 & ~w13509) | (pi0748 & w18087) | (~w13509 & w18087);
assign w15506 = w3409 & w2158;
assign w15507 = ~w4262 & ~w6899;
assign w15508 = w13509 & w12000;
assign w15509 = ~w5189 & pi0719;
assign w15510 = ~pi0940 & w9110;
assign w15511 = ~w14065 & ~w12649;
assign w15512 = w13509 & w15259;
assign w15513 = pi1370 & ~w480;
assign w15514 = ~pi0277 & w2196;
assign w15515 = ~pi0698 & w3106;
assign w15516 = ~w7058 & ~w14438;
assign w15517 = ~pi2131 & w16041;
assign w15518 = w9242 & w4793;
assign w15519 = pi2739 & ~w15235;
assign w15520 = ~pi1921 & w11313;
assign w15521 = pi1471 & w13753;
assign w15522 = ~w5808 & ~w9237;
assign w15523 = w16278 & ~w6647;
assign w15524 = (pi0373 & w6195) | (pi0373 & w1967) | (w6195 & w1967);
assign w15525 = w11209 & ~w9565;
assign w15526 = ~w14275 & w15689;
assign w15527 = ~pi1220 & ~pi3375;
assign w15528 = ~w16181 & ~w13359;
assign w15529 = ~w14411 & ~w243;
assign w15530 = pi2679 & ~w226;
assign w15531 = ~pi3154 & w17993;
assign w15532 = ~w9072 & ~w15976;
assign w15533 = pi2036 & ~w17646;
assign w15534 = pi1567 & ~w18259;
assign w15535 = ~pi3165 & pi3207;
assign w15536 = pi3166 & pi3207;
assign w15537 = ~pi1799 & ~pi3170;
assign w15538 = ~w4326 & ~w3010;
assign w15539 = (~w13518 & ~w5517) | (~w13518 & w10579) | (~w5517 & w10579);
assign w15540 = w12489 & w16617;
assign w15541 = pi2905 & ~w9504;
assign w15542 = w5453 & pi2884;
assign w15543 = ~w14080 & ~w9628;
assign w15544 = w13509 & w3659;
assign w15545 = pi2256 & ~w11671;
assign w15546 = (pi0790 & ~w13509) | (pi0790 & w9218) | (~w13509 & w9218);
assign w15547 = pi0126 & pi1220;
assign w15548 = ~w9440 & w18583;
assign w15549 = w12040 & ~w2741;
assign w15550 = ~w9858 & ~w844;
assign w15551 = ~pi3172 & w1843;
assign w15552 = ~pi3055 & w261;
assign w15553 = (pi0205 & w2726) | (pi0205 & w11408) | (w2726 & w11408);
assign w15554 = ~w14373 & w15212;
assign w15555 = (pi0905 & ~w13509) | (pi0905 & w14089) | (~w13509 & w14089);
assign w15556 = ~w3829 & ~w16924;
assign w15557 = w13509 & w7339;
assign w15558 = ~w8243 & w16743;
assign w15559 = ~w14051 & ~w5307;
assign w15560 = ~pi3157 & w8515;
assign w15561 = pi3364 & ~pi3365;
assign w15562 = ~w18541 & ~w10088;
assign w15563 = pi1470 & w13753;
assign w15564 = ~pi1972 & ~pi2252;
assign w15565 = ~w18212 & ~w16170;
assign w15566 = ~w12040 & pi0680;
assign w15567 = w14228 & ~w17513;
assign w15568 = ~pi3153 & w13730;
assign w15569 = (pi0703 & ~w13509) | (pi0703 & w10538) | (~w13509 & w10538);
assign w15570 = ~w3700 & w16372;
assign w15571 = ~w17208 & ~w3825;
assign w15572 = ~w3000 & ~pi2668;
assign w15573 = pi0024 & ~w3748;
assign w15574 = ~w6370 & ~w14059;
assign w15575 = ~w3203 & pi0545;
assign w15576 = ~pi1108 & w9110;
assign w15577 = ~pi0648 & w3791;
assign w15578 = ~pi0334 & w4058;
assign w15579 = ~pi3142 & w13730;
assign w15580 = ~w3646 & w11939;
assign w15581 = w1368 & pi0360;
assign w15582 = w17793 & w1427;
assign w15583 = w539 & ~w5913;
assign w15584 = w13509 & w4101;
assign w15585 = ~pi1772 & pi3133;
assign w15586 = ~w12036 & ~w11761;
assign w15587 = w17286 & w489;
assign w15588 = ~w14455 & ~w14528;
assign w15589 = ~pi3053 & w11406;
assign w15590 = (w2460 & ~w384) | (w2460 & w6180) | (~w384 & w6180);
assign w15591 = ~w2830 & ~w17742;
assign w15592 = ~w9435 & w4789;
assign w15593 = w7346 & w16881;
assign w15594 = ~w2725 & pi1085;
assign w15595 = ~w8878 & ~w15231;
assign w15596 = w9720 & pi1723;
assign w15597 = ~w1130 & ~w1964;
assign w15598 = ~w5189 & pi0721;
assign w15599 = ~w10174 & ~w13974;
assign w15600 = ~w4077 & w3279;
assign w15601 = ~w7844 & pi0598;
assign w15602 = (~w17562 & ~w384) | (~w17562 & w14391) | (~w384 & w14391);
assign w15603 = pi3136 & w4324;
assign w15604 = w9897 & w7763;
assign w15605 = (pi1001 & ~w13509) | (pi1001 & w103) | (~w13509 & w103);
assign w15606 = ~pi3150 & w8515;
assign w15607 = ~pi3086 & w15235;
assign w15608 = ~pi0868 & w15707;
assign w15609 = ~w18311 & ~w10584;
assign w15610 = ~pi2428 & w5075;
assign w15611 = ~pi2975 & w14524;
assign w15612 = ~pi2997 & w9474;
assign w15613 = ~pi3165 & w11701;
assign w15614 = pi3006 & ~pi3162;
assign w15615 = ~w12207 & ~w8951;
assign w15616 = ~w2311 & w16276;
assign w15617 = ~w16506 & pi1132;
assign w15618 = ~pi2061 & w8617;
assign w15619 = w12030 & w15684;
assign w15620 = ~w6195 & w16186;
assign w15621 = w14971 & w11321;
assign w15622 = w8383 & w6111;
assign w15623 = w13509 & w18303;
assign w15624 = w9414 & w6320;
assign w15625 = ~w14373 & w14839;
assign w15626 = w11936 & w9092;
assign w15627 = pi1651 & ~w6072;
assign w15628 = ~pi3147 & w11132;
assign w15629 = ~pi2262 & w13065;
assign w15630 = pi0298 & w5274;
assign w15631 = w13509 & w4383;
assign w15632 = w7481 & w14284;
assign w15633 = (pi0384 & w5560) | (pi0384 & w3721) | (w5560 & w3721);
assign w15634 = w9720 & pi1755;
assign w15635 = ~pi3133 & pi3207;
assign w15636 = ~w444 & ~w17643;
assign w15637 = ~pi3096 & w3555;
assign w15638 = ~w5163 & w3807;
assign w15639 = ~w7807 & ~w18425;
assign w15640 = pi1427 & ~w13753;
assign w15641 = pi3160 & ~pi3482;
assign w15642 = pi1606 & w13753;
assign w15643 = pi1785 & ~w8073;
assign w15644 = w6162 & w3157;
assign w15645 = ~w7077 & pi0816;
assign w15646 = w3252 & w7786;
assign w15647 = w8789 & pi0360;
assign w15648 = ~w11625 & ~w9927;
assign w15649 = w11383 & w10176;
assign w15650 = ~pi1104 & w17899;
assign w15651 = (pi0697 & ~w13509) | (pi0697 & w13099) | (~w13509 & w13099);
assign w15652 = ~w17299 & ~w6083;
assign w15653 = ~w4332 & ~w13063;
assign w15654 = pi1498 & ~w16922;
assign w15655 = ~w4138 & ~w63;
assign w15656 = (pi0637 & ~w13509) | (pi0637 & w10596) | (~w13509 & w10596);
assign w15657 = ~w13544 & ~w17682;
assign w15658 = ~pi2370 & w16041;
assign w15659 = ~w7574 & ~w14992;
assign w15660 = w15122 & ~pi2600;
assign w15661 = ~w13303 & ~w6026;
assign w15662 = pi2775 & ~w226;
assign w15663 = ~w7614 & ~w9766;
assign w15664 = ~pi3146 & w11132;
assign w15665 = ~w10402 & ~w9005;
assign w15666 = ~pi3089 & w9504;
assign w15667 = pi2385 & ~w18123;
assign w15668 = w10818 & ~w6309;
assign w15669 = pi0147 & w5274;
assign w15670 = pi0146 & ~w9966;
assign w15671 = ~pi3157 & w11132;
assign w15672 = w13509 & w15809;
assign w15673 = ~w4853 & ~w8094;
assign w15674 = ~w11600 & w6077;
assign w15675 = ~w2909 & w2960;
assign w15676 = w13509 & w4632;
assign w15677 = ~pi1920 & w11313;
assign w15678 = ~w8591 & ~w14223;
assign w15679 = w7844 & ~w6033;
assign w15680 = ~w5189 & pi0723;
assign w15681 = ~w8928 & ~w4139;
assign w15682 = pi0174 & pi0175;
assign w15683 = ~pi3097 & w6463;
assign w15684 = w425 & w3644;
assign w15685 = (pi0386 & w5560) | (pi0386 & w14437) | (w5560 & w14437);
assign w15686 = ~w12040 & pi0695;
assign w15687 = pi3105 & ~pi3169;
assign w15688 = ~pi3133 & ~pi3160;
assign w15689 = ~w7420 & ~w14587;
assign w15690 = ~pi2100 & w12724;
assign w15691 = ~w10413 & ~w3818;
assign w15692 = ~pi3150 & w3982;
assign w15693 = ~w5189 & pi1103;
assign w15694 = ~w485 & pi1299;
assign w15695 = (pi1781 & w7215) | (pi1781 & w2682) | (w7215 & w2682);
assign w15696 = pi1780 & ~w13787;
assign w15697 = ~pi2095 & w12724;
assign w15698 = w17562 & pi2571;
assign w15699 = pi2867 & w15191;
assign w15700 = (pi0581 & ~w13509) | (pi0581 & w14603) | (~w13509 & w14603);
assign w15701 = w1391 & ~w11978;
assign w15702 = ~w13546 & ~w13374;
assign w15703 = w8741 & w8798;
assign w15704 = (pi0677 & ~w13509) | (pi0677 & w14292) | (~w13509 & w14292);
assign w15705 = w4959 & w696;
assign w15706 = ~w11537 & ~w5226;
assign w15707 = w12543 & w93;
assign w15708 = ~w11111 & ~w12537;
assign w15709 = ~w10298 & ~w17170;
assign w15710 = w14109 & pi0425;
assign w15711 = ~pi3145 & w17387;
assign w15712 = w9335 & w16075;
assign w15713 = w16575 & w10120;
assign w15714 = pi1777 & ~w14951;
assign w15715 = ~pi1220 & pi3374;
assign w15716 = w8789 & pi0476;
assign w15717 = ~w5560 & w14557;
assign w15718 = pi2681 & ~w11406;
assign w15719 = pi2201 & ~w10299;
assign w15720 = pi0045 & ~w14148;
assign w15721 = ~pi3058 & w226;
assign w15722 = ~w1791 & w10425;
assign w15723 = w12607 & w16169;
assign w15724 = w13509 & w7635;
assign w15725 = ~w11884 & ~w6436;
assign w15726 = ~w12750 & w4499;
assign w15727 = ~w1132 & ~w11993;
assign w15728 = pi2741 & ~w15235;
assign w15729 = ~w5500 & ~w4722;
assign w15730 = (pi1029 & ~w13509) | (pi1029 & w1409) | (~w13509 & w1409);
assign w15731 = ~w10863 & ~w9581;
assign w15732 = ~pi3341 & w18259;
assign w15733 = pi1406 & ~pi2910;
assign w15734 = ~pi1042 & w1147;
assign w15735 = ~pi3328 & w17935;
assign w15736 = ~w15346 & ~w11465;
assign w15737 = (~pi0278 & ~w6857) | (~pi0278 & w1896) | (~w6857 & w1896);
assign w15738 = ~w13630 & ~w14722;
assign w15739 = w18295 & w1044;
assign w15740 = ~w7403 & ~w2369;
assign w15741 = ~pi0695 & w9110;
assign w15742 = w13509 & w13138;
assign w15743 = ~w180 & w4454;
assign w15744 = pi1292 & pi1345;
assign w15745 = ~w11508 & ~w18158;
assign w15746 = (pi0599 & ~w13509) | (pi0599 & w4432) | (~w13509 & w4432);
assign w15747 = ~w2342 & ~w3294;
assign w15748 = w6857 & w11865;
assign w15749 = ~w1794 & ~w17333;
assign w15750 = ~w1576 & ~w2945;
assign w15751 = pi1263 & ~pi2958;
assign w15752 = ~pi0847 & w93;
assign w15753 = ~w105 & ~w6832;
assign w15754 = pi3068 & ~w16502;
assign w15755 = ~w10438 & ~w10850;
assign w15756 = ~w9462 & w4219;
assign w15757 = ~w3000 & ~pi2770;
assign w15758 = ~w7776 & ~w18369;
assign w15759 = ~w4929 & ~w2958;
assign w15760 = w8337 & pi3332;
assign w15761 = ~w11795 & w11804;
assign w15762 = w13509 & w14769;
assign w15763 = w13509 & w14770;
assign w15764 = ~w14387 & ~w743;
assign w15765 = ~pi0498 & ~pi1345;
assign w15766 = ~w3988 & ~w15907;
assign w15767 = w2531 & w3550;
assign w15768 = pi1902 & w10959;
assign w15769 = ~w17248 & pi0949;
assign w15770 = ~w476 & ~w6372;
assign w15771 = ~w5189 & pi0725;
assign w15772 = w1368 & pi0387;
assign w15773 = w657 & w5218;
assign w15774 = w5712 & w13710;
assign w15775 = ~w8277 & ~w4701;
assign w15776 = ~pi0651 & w3791;
assign w15777 = pi1719 & ~pi3151;
assign w15778 = ~w3538 & ~w14006;
assign w15779 = w16506 & ~w11978;
assign w15780 = ~w11691 & ~w8395;
assign w15781 = pi1433 & ~w6448;
assign w15782 = ~w10379 & ~w15002;
assign w15783 = w1962 & ~w4179;
assign w15784 = ~w2662 & w14546;
assign w15785 = (pi0612 & ~w13509) | (pi0612 & w3245) | (~w13509 & w3245);
assign w15786 = ~w11556 & ~w3815;
assign w15787 = ~w6316 & ~w15028;
assign w15788 = pi1914 & ~w10299;
assign w15789 = ~w12908 & ~w7445;
assign w15790 = ~w9378 & ~w1524;
assign w15791 = ~pi3034 & ~w16502;
assign w15792 = pi3035 & ~w16502;
assign w15793 = ~w2341 & pi1046;
assign w15794 = ~w14560 & pi0241;
assign w15795 = (pi0617 & ~w13509) | (pi0617 & w789) | (~w13509 & w789);
assign w15796 = ~w4057 & ~w912;
assign w15797 = ~w10266 & ~w17206;
assign w15798 = (~w13367 & w17577) | (~w13367 & w14196) | (w17577 & w14196);
assign w15799 = ~w6148 & ~w5992;
assign w15800 = ~w1876 & ~w4859;
assign w15801 = w5639 & w16313;
assign w15802 = pi1533 & w13753;
assign w15803 = ~pi3062 & w226;
assign w15804 = w7200 & w2180;
assign w15805 = ~w7814 & w2511;
assign w15806 = ~w13494 & ~w4511;
assign w15807 = (pi0602 & ~w13509) | (pi0602 & w294) | (~w13509 & w294);
assign w15808 = w7254 & w13867;
assign w15809 = w6785 & ~w10235;
assign w15810 = ~w1391 & pi0910;
assign w15811 = ~w15122 & ~pi2432;
assign w15812 = pi2893 & ~w226;
assign w15813 = ~pi2206 & w5075;
assign w15814 = ~w13231 & pi0573;
assign w15815 = ~w5560 & w14703;
assign w15816 = ~pi2412 & w13204;
assign w15817 = pi0113 & ~w16965;
assign w15818 = ~w1572 & ~w12323;
assign w15819 = ~w13780 & ~w14261;
assign w15820 = ~w14648 & ~pi2725;
assign w15821 = w10299 & w614;
assign w15822 = pi2703 & ~w3555;
assign w15823 = ~w13231 & pi0552;
assign w15824 = ~pi1839 & ~w15883;
assign w15825 = ~w17621 & ~w9094;
assign w15826 = ~pi0697 & w9110;
assign w15827 = ~w6733 & ~w7597;
assign w15828 = w16679 & w13472;
assign w15829 = w2725 & w15609;
assign w15830 = ~w11764 & ~w13832;
assign w15831 = pi1434 & ~w6448;
assign w15832 = w12460 & w6834;
assign w15833 = ~w7009 & ~w4050;
assign w15834 = pi1323 & w458;
assign w15835 = ~pi2118 & w12755;
assign w15836 = w2341 & ~w1236;
assign w15837 = ~w11386 & ~w1248;
assign w15838 = ~w17248 & pi1056;
assign w15839 = ~w4020 & w10158;
assign w15840 = ~w8239 & ~w17580;
assign w15841 = ~pi0483 & pi3403;
assign w15842 = pi2920 & ~pi2966;
assign w15843 = pi1622 & ~w16922;
assign w15844 = ~pi3088 & w226;
assign w15845 = ~w9734 & ~w18036;
assign w15846 = ~w15214 & ~w8164;
assign w15847 = pi1869 & ~w15036;
assign w15848 = ~w5189 & pi0727;
assign w15849 = ~pi1009 & w3791;
assign w15850 = w13679 & w17130;
assign w15851 = pi2303 & ~w3223;
assign w15852 = pi1566 & ~w18259;
assign w15853 = ~w3884 & ~w1123;
assign w15854 = ~w5548 & ~w154;
assign w15855 = ~w9578 & w1649;
assign w15856 = ~pi3165 & w12427;
assign w15857 = w2725 & ~w14978;
assign w15858 = w1127 & ~w2550;
assign w15859 = ~w16172 & ~w4637;
assign w15860 = ~w9206 & ~w2942;
assign w15861 = pi1498 & ~w13753;
assign w15862 = pi2763 & ~w11406;
assign w15863 = w5453 & pi2579;
assign w15864 = ~pi0622 & w14641;
assign w15865 = ~pi1707 & pi3147;
assign w15866 = ~w16189 & ~w5401;
assign w15867 = w659 & ~w16543;
assign w15868 = (pi1103 & ~w13509) | (pi1103 & w15693) | (~w13509 & w15693);
assign w15869 = (pi0569 & ~w13509) | (pi0569 & w2606) | (~w13509 & w2606);
assign w15870 = ~w5087 & ~w9449;
assign w15871 = ~pi0994 & w795;
assign w15872 = ~w10689 & ~w17786;
assign w15873 = w13509 & w6734;
assign w15874 = w11383 & w13261;
assign w15875 = (pi1039 & ~w13509) | (pi1039 & w8818) | (~w13509 & w8818);
assign w15876 = w62 & ~w242;
assign w15877 = w9488 & pi0493;
assign w15878 = ~pi0512 & ~pi1150;
assign w15879 = ~w18066 & ~w49;
assign w15880 = w11383 & w3874;
assign w15881 = ~w9203 & ~w8193;
assign w15882 = ~w16506 & pi1262;
assign w15883 = w14651 & w13605;
assign w15884 = w13509 & w1667;
assign w15885 = ~w10499 & ~w3623;
assign w15886 = pi2916 & ~w6045;
assign w15887 = (pi0704 & ~w13509) | (pi0704 & w18378) | (~w13509 & w18378);
assign w15888 = ~w1352 & ~w4723;
assign w15889 = (~pi0046 & ~w14782) | (~pi0046 & w9837) | (~w14782 & w9837);
assign w15890 = w11232 & w3026;
assign w15891 = ~pi2474 & w11688;
assign w15892 = ~pi2434 & w13343;
assign w15893 = ~w18100 & ~w17076;
assign w15894 = ~w11075 & ~w7059;
assign w15895 = ~w9158 & pi0484;
assign w15896 = w9396 & w791;
assign w15897 = w7703 & w18205;
assign w15898 = w6785 & ~w4043;
assign w15899 = ~pi3047 & w15235;
assign w15900 = ~w7844 & pi1003;
assign w15901 = ~pi2643 & w15122;
assign w15902 = ~w10502 & ~w9397;
assign w15903 = w12040 & ~w7020;
assign w15904 = ~w5079 & w6081;
assign w15905 = w5341 & w18241;
assign w15906 = (~pi0281 & ~w6857) | (~pi0281 & w4714) | (~w6857 & w4714);
assign w15907 = ~pi1167 & ~pi1176;
assign w15908 = w10647 & ~w13995;
assign w15909 = w1803 & w13239;
assign w15910 = ~pi2257 & w13065;
assign w15911 = pi1170 & pi3192;
assign w15912 = ~w13206 & ~w18575;
assign w15913 = ~w14385 & ~w8350;
assign w15914 = ~pi3171 & w17669;
assign w15915 = pi3073 & ~pi3153;
assign w15916 = pi0056 & w6288;
assign w15917 = pi1662 & w1924;
assign w15918 = pi1744 & w1924;
assign w15919 = w15883 & w3515;
assign w15920 = w18244 & w1066;
assign w15921 = (~pi0969 & ~w13509) | (~pi0969 & w2011) | (~w13509 & w2011);
assign w15922 = ~w2993 & w11512;
assign w15923 = pi1688 & ~w261;
assign w15924 = pi2788 & ~w6463;
assign w15925 = w5189 & w11010;
assign w15926 = pi2154 & ~w11671;
assign w15927 = ~w14560 & pi0229;
assign w15928 = (w4503 & ~w914) | (w4503 & w16461) | (~w914 & w16461);
assign w15929 = pi1253 & w11655;
assign w15930 = ~pi3299 & w17935;
assign w15931 = w9440 & pi0151;
assign w15932 = ~pi3061 & w6463;
assign w15933 = ~w16969 & ~w16016;
assign w15934 = ~w14073 & w14068;
assign w15935 = pi2581 & ~w5274;
assign w15936 = ~w16077 & ~w11108;
assign w15937 = ~w4527 & ~w4720;
assign w15938 = ~pi0486 & ~pi1133;
assign w15939 = ~pi0506 & ~pi1345;
assign w15940 = ~w7634 & ~w17895;
assign w15941 = pi1751 & ~pi3158;
assign w15942 = pi2774 & ~w11406;
assign w15943 = ~w8847 & w5680;
assign w15944 = (pi1188 & w4470) | (pi1188 & w17207) | (w4470 & w17207);
assign w15945 = w7703 & w15197;
assign w15946 = ~w18180 & w9863;
assign w15947 = ~w12040 & pi0687;
assign w15948 = w13509 & w5011;
assign w15949 = pi1710 & ~w2253;
assign w15950 = ~w12964 & ~w1031;
assign w15951 = w10990 & pi0251;
assign w15952 = w12722 & w1379;
assign w15953 = w10867 & w11041;
assign w15954 = pi0017 & ~w14148;
assign w15955 = ~w13374 & w3119;
assign w15956 = w6649 & ~w15563;
assign w15957 = pi1768 & ~w5457;
assign w15958 = w14109 & pi0429;
assign w15959 = (pi0756 & ~w13509) | (pi0756 & w3926) | (~w13509 & w3926);
assign w15960 = ~w5291 & ~w14672;
assign w15961 = pi2017 & ~w14833;
assign w15962 = pi3014 & w16502;
assign w15963 = w13509 & w6456;
assign w15964 = ~w6960 & ~w14653;
assign w15965 = ~w9403 & ~w2955;
assign w15966 = ~pi2992 & ~pi3207;
assign w15967 = ~pi2177 & w5384;
assign w15968 = ~pi2018 & w11688;
assign w15969 = ~w9031 & ~w2585;
assign w15970 = pi1129 & pi1177;
assign w15971 = ~w15069 & ~w16569;
assign w15972 = ~pi2704 & w15122;
assign w15973 = ~w14044 & ~w13677;
assign w15974 = w16721 & w3229;
assign w15975 = ~w9131 & ~w16361;
assign w15976 = w13509 & w7605;
assign w15977 = ~w13367 & ~pi0501;
assign w15978 = w1368 & pi0404;
assign w15979 = pi2697 & ~w16815;
assign w15980 = w15808 & ~w15173;
assign w15981 = ~w12460 & w18525;
assign w15982 = ~w12556 & ~w15816;
assign w15983 = ~w12040 & pi0941;
assign w15984 = ~pi1232 & pi1973;
assign w15985 = ~w6195 & w4528;
assign w15986 = w914 & w1500;
assign w15987 = w13231 & ~w16498;
assign w15988 = w7307 & w1602;
assign w15989 = ~pi0958 & w3791;
assign w15990 = pi1337 & pi0308;
assign w15991 = ~w10018 & ~w9775;
assign w15992 = w18449 & w11175;
assign w15993 = ~pi3346 & w18259;
assign w15994 = (pi0811 & ~w13509) | (pi0811 & w12451) | (~w13509 & w12451);
assign w15995 = ~w10743 & ~w14197;
assign w15996 = w18558 & w5014;
assign w15997 = ~w5695 & ~w5591;
assign w15998 = pi1337 & ~pi0270;
assign w15999 = pi1328 & w458;
assign w16000 = ~w401 & ~w4651;
assign w16001 = ~pi0881 & w1126;
assign w16002 = pi1704 & w4683;
assign w16003 = ~w9056 & ~w11224;
assign w16004 = ~w16220 & ~w9951;
assign w16005 = ~pi2023 & w7455;
assign w16006 = ~w15606 & ~w12544;
assign w16007 = ~pi1074 & w1147;
assign w16008 = w16506 & w17718;
assign w16009 = ~w9313 & ~w6395;
assign w16010 = ~pi0430 & w13806;
assign w16011 = ~pi2227 & w2151;
assign w16012 = ~w4936 & ~pi0487;
assign w16013 = ~pi0817 & w1147;
assign w16014 = w11383 & w1260;
assign w16015 = pi2533 & w14148;
assign w16016 = ~w11655 & w14927;
assign w16017 = w12460 & w462;
assign w16018 = ~w3386 & w2460;
assign w16019 = pi1388 & w13753;
assign w16020 = pi2855 & ~w226;
assign w16021 = w18557 & w922;
assign w16022 = ~w12641 & ~w9710;
assign w16023 = ~pi2342 & w12724;
assign w16024 = w14648 & ~pi2727;
assign w16025 = ~pi3108 & ~pi3207;
assign w16026 = ~w2340 & w2497;
assign w16027 = pi1664 & w1924;
assign w16028 = w12040 & ~w15173;
assign w16029 = ~pi3004 & ~pi3207;
assign w16030 = (pi1376 & ~w8966) | (pi1376 & w17902) | (~w8966 & w17902);
assign w16031 = pi0255 & w5274;
assign w16032 = pi1454 & w13753;
assign w16033 = ~pi0259 & w5082;
assign w16034 = pi2869 & w15191;
assign w16035 = w17248 & ~w6922;
assign w16036 = w14560 & pi0366;
assign w16037 = pi1781 & ~w16886;
assign w16038 = ~w4203 & ~w6415;
assign w16039 = ~w16647 & ~w10172;
assign w16040 = pi1131 & ~pi1181;
assign w16041 = w14138 & w17559;
assign w16042 = ~w13123 & ~w9914;
assign w16043 = ~pi0507 & ~pi1151;
assign w16044 = ~w16724 & ~w2928;
assign w16045 = w8789 & ~pi0449;
assign w16046 = w5459 & w1036;
assign w16047 = ~w12362 & ~w4170;
assign w16048 = ~w15994 & ~w5474;
assign w16049 = ~w1742 & ~w17390;
assign w16050 = ~w709 & ~pi1291;
assign w16051 = ~w709 & pi1292;
assign w16052 = w14228 & ~w9852;
assign w16053 = ~w12301 & ~w6274;
assign w16054 = ~w16082 & ~w15177;
assign w16055 = ~pi3024 & ~pi3025;
assign w16056 = ~pi0397 & w871;
assign w16057 = ~w11104 & ~w2364;
assign w16058 = ~w13525 & ~w10655;
assign w16059 = ~pi1051 & w15707;
assign w16060 = pi1327 & w458;
assign w16061 = pi3009 & w16502;
assign w16062 = ~w3369 & ~w15342;
assign w16063 = pi1867 & ~w15036;
assign w16064 = ~pi0747 & w17490;
assign w16065 = ~w12417 & ~w16158;
assign w16066 = ~w669 & ~w12017;
assign w16067 = w4297 & w17127;
assign w16068 = ~pi0483 & pi3393;
assign w16069 = ~pi3311 & w6072;
assign w16070 = ~w14087 & ~w13752;
assign w16071 = w3223 & w614;
assign w16072 = w17248 & ~w2587;
assign w16073 = ~pi3354 & w6072;
assign w16074 = pi3154 & w619;
assign w16075 = ~w4960 & ~w8154;
assign w16076 = ~w17773 & ~w12022;
assign w16077 = (pi0780 & ~w13509) | (pi0780 & w5793) | (~w13509 & w5793);
assign w16078 = w13546 & w7060;
assign w16079 = w2742 & ~w13365;
assign w16080 = ~w11612 & ~w1940;
assign w16081 = ~pi1913 & w11313;
assign w16082 = ~pi0942 & w12197;
assign w16083 = ~w1082 & ~w9629;
assign w16084 = ~w188 & ~w7708;
assign w16085 = w13509 & w2658;
assign w16086 = pi2134 & ~w15883;
assign w16087 = ~pi3139 & ~pi3160;
assign w16088 = ~w12739 & w7233;
assign w16089 = ~w1285 & ~w3650;
assign w16090 = ~w11826 & ~w16100;
assign w16091 = w9908 & w6537;
assign w16092 = ~pi2021 & w11688;
assign w16093 = ~pi3163 & w12427;
assign w16094 = pi1156 & w9420;
assign w16095 = ~w9550 & ~w16346;
assign w16096 = pi2980 & ~w3987;
assign w16097 = ~w234 & ~pi0499;
assign w16098 = ~pi3036 & ~pi3207;
assign w16099 = ~w3054 & w15260;
assign w16100 = ~pi3287 & w9781;
assign w16101 = ~pi2181 & w5384;
assign w16102 = ~w4032 & ~w18305;
assign w16103 = w8869 & ~w1341;
assign w16104 = ~w14039 & ~w13118;
assign w16105 = pi3012 & w16502;
assign w16106 = w539 & ~w7528;
assign w16107 = ~w13388 & ~w17952;
assign w16108 = w5437 & w13511;
assign w16109 = w14524 & w14078;
assign w16110 = w6941 & w17523;
assign w16111 = w15122 & ~pi2719;
assign w16112 = w7703 & w6810;
assign w16113 = ~w5475 & ~w11085;
assign w16114 = pi0139 & w5274;
assign w16115 = ~w6697 & ~pi0961;
assign w16116 = w7307 & w10135;
assign w16117 = w574 & w16565;
assign w16118 = ~pi1128 & w14073;
assign w16119 = pi1129 & w14073;
assign w16120 = ~pi3020 & ~w3384;
assign w16121 = ~w5376 & ~w301;
assign w16122 = ~w923 & ~w3697;
assign w16123 = ~w1962 & pi0648;
assign w16124 = ~w7149 & ~w1548;
assign w16125 = ~w13821 & ~w3056;
assign w16126 = w968 & ~pi0277;
assign w16127 = ~w12319 & w2207;
assign w16128 = pi2959 & ~w13367;
assign w16129 = pi1953 & ~w14833;
assign w16130 = w7498 & w14233;
assign w16131 = pi1887 & ~w15036;
assign w16132 = ~w17907 & ~w10039;
assign w16133 = ~w14648 & ~pi1749;
assign w16134 = w8658 & pi1786;
assign w16135 = ~w8231 & ~w10677;
assign w16136 = ~w2675 & ~w10315;
assign w16137 = ~w5650 & pi1162;
assign w16138 = w7299 & w15401;
assign w16139 = w16713 & w2420;
assign w16140 = w6697 & ~w7020;
assign w16141 = ~w8588 & w10299;
assign w16142 = ~pi2240 & w2151;
assign w16143 = pi1473 & w13753;
assign w16144 = pi1753 & ~w8113;
assign w16145 = pi1510 & ~w13753;
assign w16146 = ~w7844 & pi1073;
assign w16147 = ~w14096 & ~w3621;
assign w16148 = ~w16023 & ~w4858;
assign w16149 = (pi0866 & ~w13509) | (pi0866 & w3540) | (~w13509 & w3540);
assign w16150 = w13509 & w2332;
assign w16151 = ~w17248 & pi0876;
assign w16152 = w13509 & w3172;
assign w16153 = ~pi3349 & w9781;
assign w16154 = ~pi2084 & w17439;
assign w16155 = pi2448 & ~w10299;
assign w16156 = ~w16506 & pi1148;
assign w16157 = pi1752 & pi3157;
assign w16158 = ~pi2384 & ~w15450;
assign w16159 = ~w2321 & ~w411;
assign w16160 = ~w10477 & ~w13324;
assign w16161 = w1498 & ~w13869;
assign w16162 = ~w15122 & ~pi2693;
assign w16163 = pi0206 & pi0207;
assign w16164 = w14228 & ~w4179;
assign w16165 = pi1786 & ~w15767;
assign w16166 = w15122 & ~pi2696;
assign w16167 = ~w17371 & ~w7765;
assign w16168 = ~pi2873 & w14148;
assign w16169 = ~w6036 & ~w14231;
assign w16170 = ~pi1934 & w12724;
assign w16171 = ~w3000 & ~pi2670;
assign w16172 = ~w9440 & ~w9949;
assign w16173 = (~w16820 & ~w5517) | (~w16820 & w18260) | (~w5517 & w18260);
assign w16174 = pi0274 & w14001;
assign w16175 = (~pi1760 & ~w7799) | (~pi1760 & w5070) | (~w7799 & w5070);
assign w16176 = w8939 & w18136;
assign w16177 = w5453 & pi2483;
assign w16178 = ~pi3333 & w18259;
assign w16179 = pi1657 & ~w13753;
assign w16180 = ~w16254 & ~w1297;
assign w16181 = pi1478 & ~w9781;
assign w16182 = w3779 & w6693;
assign w16183 = ~pi0820 & w1147;
assign w16184 = ~w3484 & ~w8346;
assign w16185 = ~pi3164 & w17387;
assign w16186 = ~w14560 & pi0217;
assign w16187 = ~pi1939 & w11688;
assign w16188 = pi3075 & ~pi3170;
assign w16189 = ~pi2305 & w12941;
assign w16190 = ~w16119 & w12837;
assign w16191 = ~w256 & w7777;
assign w16192 = pi2139 & ~w15883;
assign w16193 = w3203 & w11302;
assign w16194 = pi2140 & ~w15883;
assign w16195 = w15883 & w614;
assign w16196 = ~pi3098 & w6463;
assign w16197 = pi2636 & ~w9504;
assign w16198 = w8789 & pi0404;
assign w16199 = w14648 & ~pi2515;
assign w16200 = pi2387 & ~w412;
assign w16201 = pi1683 & w5274;
assign w16202 = ~w12783 & ~w9226;
assign w16203 = ~w2341 & pi1045;
assign w16204 = pi1391 & ~w17935;
assign w16205 = pi0222 & w7536;
assign w16206 = w3203 & ~w6033;
assign w16207 = ~w4328 & w15379;
assign w16208 = ~pi3100 & w6463;
assign w16209 = ~w6697 & pi1114;
assign w16210 = w14782 & w2570;
assign w16211 = ~w2326 & ~w12554;
assign w16212 = pi0492 & pi0493;
assign w16213 = ~w2930 & ~w1202;
assign w16214 = w7799 & w5051;
assign w16215 = ~w7454 & ~w13992;
assign w16216 = ~pi2988 & w226;
assign w16217 = ~w17964 & ~w5700;
assign w16218 = ~pi0152 & ~pi0203;
assign w16219 = w458 & w9579;
assign w16220 = ~w9812 & w13275;
assign w16221 = w968 & ~pi0293;
assign w16222 = ~pi2109 & w12755;
assign w16223 = ~pi2367 & w17439;
assign w16224 = ~w1289 & ~w1812;
assign w16225 = w10818 & ~w6864;
assign w16226 = (pi0862 & ~w13509) | (pi0862 & w10603) | (~w13509 & w10603);
assign w16227 = ~w11704 & ~w5600;
assign w16228 = ~pi1299 & ~pi1317;
assign w16229 = ~w3384 & w8607;
assign w16230 = w11077 & w13547;
assign w16231 = w14228 & ~w305;
assign w16232 = ~w18265 & ~w7911;
assign w16233 = w13509 & w17402;
assign w16234 = ~w17893 & ~w8436;
assign w16235 = w3402 & w18501;
assign w16236 = w384 & w10207;
assign w16237 = ~w9960 & w9569;
assign w16238 = ~pi3074 & pi3133;
assign w16239 = (~w17562 & ~w384) | (~w17562 & w718) | (~w384 & w718);
assign w16240 = (pi0806 & ~w13509) | (pi0806 & w17570) | (~w13509 & w17570);
assign w16241 = pi1326 & w458;
assign w16242 = ~w4709 & ~w16015;
assign w16243 = ~w17819 & ~w14945;
assign w16244 = ~w7689 & ~w2762;
assign w16245 = ~w9368 & ~w17186;
assign w16246 = pi2367 & ~w17683;
assign w16247 = ~w14228 & pi0630;
assign w16248 = ~w15808 & pi0752;
assign w16249 = (pi1205 & ~w13509) | (pi1205 & w13447) | (~w13509 & w13447);
assign w16250 = pi2760 & w7965;
assign w16251 = ~w14706 & w12283;
assign w16252 = ~w12617 & ~w14772;
assign w16253 = ~w1887 & ~w2730;
assign w16254 = pi0009 & ~w14148;
assign w16255 = ~w17017 & ~w7430;
assign w16256 = ~w1353 & ~w13463;
assign w16257 = ~pi1369 & pi3233;
assign w16258 = pi2538 & w15191;
assign w16259 = pi1146 & ~w3771;
assign w16260 = ~w7844 & pi0597;
assign w16261 = pi1175 & pi3209;
assign w16262 = ~pi1105 & w3106;
assign w16263 = (~pi0968 & ~w13509) | (~pi0968 & w10624) | (~w13509 & w10624);
assign w16264 = pi0207 & w10959;
assign w16265 = ~w2725 & pi0795;
assign w16266 = w10602 & w10272;
assign w16267 = ~pi3131 & w12427;
assign w16268 = ~w18481 & ~w1840;
assign w16269 = pi1319 & pi1345;
assign w16270 = ~pi3133 & w3982;
assign w16271 = w5517 & w16556;
assign w16272 = ~pi3159 & w14753;
assign w16273 = ~pi3429 & w15036;
assign w16274 = w12460 & w15240;
assign w16275 = w13509 & w7407;
assign w16276 = w10647 & ~w18355;
assign w16277 = pi3133 & ~pi3165;
assign w16278 = w28 & w15907;
assign w16279 = ~pi1356 & pi2995;
assign w16280 = pi2598 & ~w9504;
assign w16281 = w312 & w7312;
assign w16282 = w13509 & w16472;
assign w16283 = ~pi3131 & w17993;
assign w16284 = ~pi1945 & w7455;
assign w16285 = w5517 & w17750;
assign w16286 = w3243 & ~pi0322;
assign w16287 = ~pi0837 & w93;
assign w16288 = (pi0584 & ~w13509) | (pi0584 & w13132) | (~w13509 & w13132);
assign w16289 = ~pi3117 & ~pi3160;
assign w16290 = pi3118 & ~pi3160;
assign w16291 = ~w6186 & ~w10821;
assign w16292 = pi2223 & ~w11735;
assign w16293 = ~w13230 & ~w16292;
assign w16294 = ~w9304 & ~w17228;
assign w16295 = ~w12784 & ~w12844;
assign w16296 = ~w14285 & ~w1615;
assign w16297 = w1127 & ~w4017;
assign w16298 = w13509 & w10837;
assign w16299 = ~w16116 & ~w16872;
assign w16300 = w6697 & ~w4179;
assign w16301 = pi0303 & pi1858;
assign w16302 = ~w8447 & w6192;
assign w16303 = pi1464 & w13753;
assign w16304 = w9440 & pi0195;
assign w16305 = ~w15483 & ~w13946;
assign w16306 = w10818 & ~w18362;
assign w16307 = ~w1368 & ~pi0450;
assign w16308 = ~w3724 & w16239;
assign w16309 = ~pi2088 & w12724;
assign w16310 = ~w2725 & pi0784;
assign w16311 = ~pi2254 & w12941;
assign w16312 = w15307 & w8035;
assign w16313 = ~w9869 & ~w4958;
assign w16314 = pi2993 & w16502;
assign w16315 = ~pi2992 & w16502;
assign w16316 = ~w9782 & ~w17681;
assign w16317 = w12460 & w17102;
assign w16318 = pi3170 & w4304;
assign w16319 = w16506 & ~w15173;
assign w16320 = ~pi3286 & w9781;
assign w16321 = ~w953 & ~w5907;
assign w16322 = ~w16278 & pi0715;
assign w16323 = ~pi3355 & w6072;
assign w16324 = pi1497 & ~w13753;
assign w16325 = (pi0389 & w5560) | (pi0389 & w7802) | (w5560 & w7802);
assign w16326 = ~pi3147 & pi3207;
assign w16327 = ~pi0770 & w6200;
assign w16328 = w3203 & w15609;
assign w16329 = ~w12598 & ~w7045;
assign w16330 = ~w10964 & ~w9673;
assign w16331 = pi1911 & ~w14524;
assign w16332 = ~w3333 & ~w13367;
assign w16333 = w4251 & w3803;
assign w16334 = w3402 & w6981;
assign w16335 = ~w7571 & ~w16666;
assign w16336 = ~w5719 & ~w17664;
assign w16337 = (pi1119 & ~w13509) | (pi1119 & w211) | (~w13509 & w211);
assign w16338 = ~w17248 & pi0885;
assign w16339 = w9440 & pi0183;
assign w16340 = ~pi2939 & w1326;
assign w16341 = w18257 & w5518;
assign w16342 = ~w9383 & w348;
assign w16343 = ~pi2129 & w11313;
assign w16344 = w6546 & w8000;
assign w16345 = w9720 & ~w3054;
assign w16346 = ~w5560 & w2071;
assign w16347 = w709 & pi1861;
assign w16348 = ~w15988 & w12962;
assign w16349 = ~w4290 & ~w15641;
assign w16350 = w934 & pi0431;
assign w16351 = w7864 & w833;
assign w16352 = w11209 & ~w18308;
assign w16353 = pi2508 & ~w5274;
assign w16354 = ~pi3045 & w6463;
assign w16355 = (pi0006 & ~w1766) | (pi0006 & w8513) | (~w1766 & w8513);
assign w16356 = ~w3000 & ~pi2811;
assign w16357 = ~w11439 & ~w8944;
assign w16358 = ~pi2044 & w13204;
assign w16359 = pi1454 & ~w7090;
assign w16360 = w4020 & ~w3094;
assign w16361 = w412 & w3515;
assign w16362 = pi3029 & ~w16502;
assign w16363 = ~w6253 & ~w10195;
assign w16364 = w15808 & w1217;
assign w16365 = ~pi3035 & pi3145;
assign w16366 = pi0028 & ~w3748;
assign w16367 = ~pi0749 & w17490;
assign w16368 = ~pi2946 & w226;
assign w16369 = pi2674 & ~w226;
assign w16370 = (~pi0202 & ~w15290) | (~pi0202 & w10110) | (~w15290 & w10110);
assign w16371 = w7703 & w2335;
assign w16372 = (~w4232 & ~w9420) | (~w4232 & w13751) | (~w9420 & w13751);
assign w16373 = pi0172 & w5274;
assign w16374 = ~w16278 & pi1024;
assign w16375 = ~w9820 & ~w634;
assign w16376 = w1391 & ~w4179;
assign w16377 = (w17562 & ~w7799) | (w17562 & w11198) | (~w7799 & w11198);
assign w16378 = ~w15576 & ~w5117;
assign w16379 = w709 & pi1898;
assign w16380 = ~pi3131 & w14753;
assign w16381 = w13509 & w4093;
assign w16382 = pi1862 & ~w15036;
assign w16383 = ~pi3157 & w4310;
assign w16384 = ~w11220 & ~w6526;
assign w16385 = ~pi2498 & w17213;
assign w16386 = ~pi2921 & ~w6045;
assign w16387 = ~pi2739 & w17213;
assign w16388 = pi0491 & w7098;
assign w16389 = pi2624 & ~w16815;
assign w16390 = ~w2014 & w5353;
assign w16391 = ~w5560 & w9916;
assign w16392 = ~w1791 & w15972;
assign w16393 = ~w88 & w2139;
assign w16394 = pi0438 & w17173;
assign w16395 = ~w3055 & w6219;
assign w16396 = ~w3055 & w6220;
assign w16397 = ~pi2286 & w5075;
assign w16398 = w6649 & ~w4285;
assign w16399 = pi2856 & ~w5274;
assign w16400 = ~pi2431 & w7455;
assign w16401 = ~w1480 & ~w6357;
assign w16402 = ~w9440 & ~w1322;
assign w16403 = ~w6785 & pi0869;
assign w16404 = ~pi2826 & w13343;
assign w16405 = w8658 & pi1756;
assign w16406 = pi0504 & pi1186;
assign w16407 = ~w6465 & ~w10994;
assign w16408 = w16650 & w15450;
assign w16409 = ~pi0743 & w17490;
assign w16410 = w13509 & w8053;
assign w16411 = w7077 & ~w6647;
assign w16412 = w16278 & ~w7707;
assign w16413 = ~pi2361 & w17439;
assign w16414 = w8882 & w8062;
assign w16415 = ~pi3135 & w4310;
assign w16416 = w7703 & w10858;
assign w16417 = pi2675 & ~w226;
assign w16418 = ~w8178 & ~w16153;
assign w16419 = w14648 & ~pi2690;
assign w16420 = w766 & w14005;
assign w16421 = ~w16478 & ~w15438;
assign w16422 = ~w4072 & ~w4174;
assign w16423 = ~pi0499 & ~pi1183;
assign w16424 = ~pi3335 & w6072;
assign w16425 = w10189 & ~pi0482;
assign w16426 = w14560 & pi0344;
assign w16427 = ~w16324 & w13963;
assign w16428 = ~w3134 & ~w17005;
assign w16429 = ~w11436 & ~w16726;
assign w16430 = ~w15808 & pi1032;
assign w16431 = ~w12040 & pi1108;
assign w16432 = w17741 & w9371;
assign w16433 = ~pi3091 & w226;
assign w16434 = ~w3055 & w2205;
assign w16435 = ~w15165 & ~w5530;
assign w16436 = ~w11311 & ~w10435;
assign w16437 = w539 & ~w8728;
assign w16438 = ~pi1755 & ~pi3165;
assign w16439 = ~w8637 & ~w471;
assign w16440 = ~w5784 & w6587;
assign w16441 = ~w5683 & ~w16766;
assign w16442 = ~w11454 & ~w16840;
assign w16443 = pi1506 & ~w13753;
assign w16444 = ~pi2976 & w15235;
assign w16445 = pi1590 & ~w13753;
assign w16446 = ~w16445 & w6959;
assign w16447 = w9794 & w16794;
assign w16448 = ~w2725 & pi1041;
assign w16449 = ~w15122 & ~pi2821;
assign w16450 = ~w6785 & pi0864;
assign w16451 = ~w15897 & ~w5854;
assign w16452 = w14105 & ~w9462;
assign w16453 = pi2972 & ~w13207;
assign w16454 = (pi0344 & w6195) | (pi0344 & w16426) | (w6195 & w16426);
assign w16455 = ~pi2302 & w12941;
assign w16456 = pi3160 & ~pi3477;
assign w16457 = pi1298 & pi1270;
assign w16458 = pi3028 & ~w16502;
assign w16459 = pi2944 & ~w4868;
assign w16460 = ~w8003 & w1326;
assign w16461 = ~w1500 & w4503;
assign w16462 = w14228 & ~w7707;
assign w16463 = ~pi2226 & w2151;
assign w16464 = ~w5041 & ~w16775;
assign w16465 = pi2842 & w605;
assign w16466 = pi1573 & ~w18259;
assign w16467 = ~pi2111 & w12755;
assign w16468 = ~pi3131 & w15839;
assign w16469 = ~w5217 & ~w15155;
assign w16470 = ~pi1047 & w93;
assign w16471 = ~w16278 & pi0700;
assign w16472 = w7077 & w11302;
assign w16473 = pi1374 & ~w5724;
assign w16474 = pi2311 & ~w4508;
assign w16475 = w5189 & ~w7707;
assign w16476 = pi2294 & w15974;
assign w16477 = ~w509 & w15056;
assign w16478 = pi1975 & ~w3555;
assign w16479 = ~w2230 & w5352;
assign w16480 = pi1359 & ~w4324;
assign w16481 = ~w5369 & w11595;
assign w16482 = w6857 & w13811;
assign w16483 = ~w18381 & ~w14823;
assign w16484 = ~pi1942 & w17439;
assign w16485 = ~pi1044 & w1147;
assign w16486 = w13509 & w169;
assign w16487 = ~w17968 & ~w6764;
assign w16488 = ~w7110 & ~w3152;
assign w16489 = ~w7077 & pi0814;
assign w16490 = ~w13231 & pi0553;
assign w16491 = ~w12062 & ~w2167;
assign w16492 = w9905 & w4197;
assign w16493 = ~w2782 & ~w17633;
assign w16494 = ~w5542 & ~w3535;
assign w16495 = pi1750 & ~w3522;
assign w16496 = ~w7769 & ~w13956;
assign w16497 = (pi0789 & ~w13509) | (pi0789 & w4553) | (~w13509 & w4553);
assign w16498 = ~w9451 & ~w3516;
assign w16499 = pi1371 & w10455;
assign w16500 = ~w5564 & ~w12347;
assign w16501 = ~pi3412 & w15036;
assign w16502 = w12524 & w6801;
assign w16503 = ~pi2330 & w7455;
assign w16504 = pi1375 & ~pi3224;
assign w16505 = ~w6095 & ~pi0505;
assign w16506 = ~w14705 & w16782;
assign w16507 = pi1811 & pi1969;
assign w16508 = pi1243 & ~pi1267;
assign w16509 = ~pi0660 & w12197;
assign w16510 = ~w17282 & ~w17918;
assign w16511 = ~w16606 & ~w9356;
assign w16512 = ~w11815 & ~w4024;
assign w16513 = ~w9020 & ~w7686;
assign w16514 = w8337 & pi3303;
assign w16515 = pi2378 & ~w412;
assign w16516 = ~pi3154 & w17387;
assign w16517 = ~pi2916 & pi3205;
assign w16518 = w15450 & ~w11628;
assign w16519 = ~pi3088 & w6463;
assign w16520 = pi3079 & w16502;
assign w16521 = w16268 & w12807;
assign w16522 = w13509 & w16669;
assign w16523 = ~w10577 & ~w18498;
assign w16524 = ~w2754 & ~w6254;
assign w16525 = ~w1057 & ~w5069;
assign w16526 = pi2548 & w14148;
assign w16527 = ~w13629 & ~w17461;
assign w16528 = w15789 & w4126;
assign w16529 = pi1798 & ~w7177;
assign w16530 = pi2095 & ~w4420;
assign w16531 = ~w702 & w12187;
assign w16532 = ~w13489 & ~w8159;
assign w16533 = w5523 & w16102;
assign w16534 = pi0039 & pi0050;
assign w16535 = w11209 & ~w14658;
assign w16536 = ~w9753 & ~w17276;
assign w16537 = ~w8182 & w1314;
assign w16538 = pi2220 & ~w11735;
assign w16539 = pi2416 & ~w10158;
assign w16540 = ~w13664 & ~w10514;
assign w16541 = ~w2128 & w13366;
assign w16542 = ~pi2637 & w15122;
assign w16543 = (pi2950 & ~w545) | (pi2950 & w13397) | (~w545 & w13397);
assign w16544 = ~pi2682 & w13343;
assign w16545 = ~w8213 & ~w15031;
assign w16546 = w3889 & w6860;
assign w16547 = ~w2519 & ~w9223;
assign w16548 = ~w10466 & ~w4659;
assign w16549 = pi3014 & ~w3987;
assign w16550 = (pi1232 & w302) | (pi1232 & w7359) | (w302 & w7359);
assign w16551 = ~w4584 & w8810;
assign w16552 = w539 & ~w14004;
assign w16553 = w14228 & ~w11978;
assign w16554 = pi2794 & ~w11406;
assign w16555 = (pi1134 & ~w5437) | (pi1134 & w3952) | (~w5437 & w3952);
assign w16556 = ~pi2967 & pi3026;
assign w16557 = w15883 & w14078;
assign w16558 = w10647 & ~w3539;
assign w16559 = pi1602 & ~w9781;
assign w16560 = w5383 & pi2540;
assign w16561 = ~pi0917 & w17490;
assign w16562 = ~pi3341 & w9781;
assign w16563 = ~w13376 & ~w13621;
assign w16564 = ~w14045 & ~w17457;
assign w16565 = w2742 & ~w6337;
assign w16566 = pi1959 & ~w14833;
assign w16567 = ~w17420 & ~w2509;
assign w16568 = ~w6785 & pi0984;
assign w16569 = pi3134 & w15767;
assign w16570 = ~w1191 & ~w2773;
assign w16571 = ~pi2242 & w12941;
assign w16572 = ~w1929 & w15450;
assign w16573 = ~pi3427 & w15036;
assign w16574 = ~w7259 & ~w13290;
assign w16575 = (w14137 & ~w15136) | (w14137 & w17610) | (~w15136 & w17610);
assign w16576 = ~w6958 & ~w5465;
assign w16577 = (pi2955 & w2014) | (pi2955 & w17775) | (w2014 & w17775);
assign w16578 = pi2085 & ~w18123;
assign w16579 = pi1731 & w1924;
assign w16580 = w7703 & w7118;
assign w16581 = pi1405 & ~w12497;
assign w16582 = ~w14489 & ~w10622;
assign w16583 = w13509 & w16035;
assign w16584 = ~w17248 & pi0894;
assign w16585 = ~w6270 & ~w11528;
assign w16586 = pi2003 & ~w9414;
assign w16587 = ~w13136 & ~w13198;
assign w16588 = ~w18250 & w5460;
assign w16589 = ~pi2987 & w15235;
assign w16590 = pi3040 & ~w3987;
assign w16591 = ~w10220 & ~w10578;
assign w16592 = pi2482 & ~w5274;
assign w16593 = w12911 & w12223;
assign w16594 = ~w3011 & ~w10892;
assign w16595 = w13509 & w1878;
assign w16596 = ~w5131 & ~w15776;
assign w16597 = (pi0683 & ~w13509) | (pi0683 & w2376) | (~w13509 & w2376);
assign w16598 = ~w5366 & w6523;
assign w16599 = ~w1391 & pi0773;
assign w16600 = ~pi3115 & pi3136;
assign w16601 = ~pi3006 & pi3162;
assign w16602 = (pi1053 & ~w13509) | (pi1053 & w8974) | (~w13509 & w8974);
assign w16603 = pi3158 & w8001;
assign w16604 = w9440 & pi0156;
assign w16605 = ~w10469 & w15602;
assign w16606 = ~pi0292 & w2196;
assign w16607 = pi3160 & ~pi3498;
assign w16608 = w384 & w13550;
assign w16609 = w5453 & pi2894;
assign w16610 = w7077 & ~w7020;
assign w16611 = ~pi1971 & w10539;
assign w16612 = w14560 & pi0362;
assign w16613 = ~w1368 & ~pi0453;
assign w16614 = ~w14542 & ~w12166;
assign w16615 = w17248 & ~w17210;
assign w16616 = ~pi0250 & ~w7428;
assign w16617 = ~w13804 & ~w887;
assign w16618 = ~w15547 & ~w15527;
assign w16619 = ~pi2462 & w5384;
assign w16620 = pi0515 & w4787;
assign w16621 = ~w7688 & ~w10199;
assign w16622 = ~pi0307 & ~w8801;
assign w16623 = pi3143 & w18497;
assign w16624 = pi0271 & w5113;
assign w16625 = pi1250 & pi3226;
assign w16626 = ~pi0638 & w3791;
assign w16627 = w13509 & w14331;
assign w16628 = w13509 & w10736;
assign w16629 = pi2360 & ~w412;
assign w16630 = w17960 & w2767;
assign w16631 = ~w7868 & ~w7988;
assign w16632 = ~pi1878 & ~pi3510;
assign w16633 = (w6688 & w5901) | (w6688 & w1040) | (w5901 & w1040);
assign w16634 = ~w3469 & ~w14686;
assign w16635 = pi1337 & ~pi0272;
assign w16636 = ~w4220 & ~w16623;
assign w16637 = ~w7482 & ~w11117;
assign w16638 = ~w6981 & ~w6111;
assign w16639 = w5437 & w9295;
assign w16640 = pi1499 & ~w16922;
assign w16641 = w62 & ~w7664;
assign w16642 = ~pi3346 & w6448;
assign w16643 = w6697 & w1217;
assign w16644 = ~w8110 & w7773;
assign w16645 = ~w709 & pi1273;
assign w16646 = w12209 & w354;
assign w16647 = pi1809 & ~w8829;
assign w16648 = ~w3297 & ~w10882;
assign w16649 = ~pi2484 & w17213;
assign w16650 = ~w13514 & ~w16118;
assign w16651 = ~w7844 & pi0548;
assign w16652 = w4927 & w1706;
assign w16653 = pi1809 & ~w3795;
assign w16654 = ~pi2994 & w14918;
assign w16655 = ~w17392 & ~w6932;
assign w16656 = ~w593 & ~w7894;
assign w16657 = ~w10334 & ~w7188;
assign w16658 = ~w10750 & ~w4209;
assign w16659 = ~w2513 & ~w8689;
assign w16660 = w7077 & ~w15173;
assign w16661 = ~w6641 & ~w8450;
assign w16662 = w9674 & w11687;
assign w16663 = w6785 & ~w13195;
assign w16664 = w10189 & ~pi0458;
assign w16665 = (pi0882 & ~w13509) | (pi0882 & w9975) | (~w13509 & w9975);
assign w16666 = w13509 & w5849;
assign w16667 = pi1453 & ~w7090;
assign w16668 = w1391 & ~w7020;
assign w16669 = w1391 & ~w17513;
assign w16670 = (pi0942 & ~w13509) | (pi0942 & w6023) | (~w13509 & w6023);
assign w16671 = pi0148 & ~pi0187;
assign w16672 = ~w8442 & ~w11762;
assign w16673 = w13509 & w10828;
assign w16674 = ~w230 & ~w17111;
assign w16675 = ~pi3290 & w16922;
assign w16676 = pi0500 & ~pi1156;
assign w16677 = ~pi3153 & w15048;
assign w16678 = pi2584 & ~w5274;
assign w16679 = ~w5560 & w18464;
assign w16680 = w15106 & ~pi1858;
assign w16681 = pi1733 & w1924;
assign w16682 = ~w14601 & ~w2473;
assign w16683 = ~pi3018 & ~pi3020;
assign w16684 = w10728 & w15982;
assign w16685 = w14121 & w8787;
assign w16686 = (pi1898 & w2014) | (pi1898 & w16379) | (w2014 & w16379);
assign w16687 = ~w17935 & ~w1832;
assign w16688 = pi0100 & w3748;
assign w16689 = w11209 & ~w1724;
assign w16690 = w5189 & ~w7020;
assign w16691 = pi3005 & ~w16502;
assign w16692 = ~pi1311 & ~pi0444;
assign w16693 = pi1416 & ~w6072;
assign w16694 = pi3160 & ~w13207;
assign w16695 = pi1358 & ~w4324;
assign w16696 = pi0122 & w3748;
assign w16697 = pi0301 & w5113;
assign w16698 = (pi0706 & ~w13509) | (pi0706 & w4682) | (~w13509 & w4682);
assign w16699 = w16893 & w11776;
assign w16700 = ~w10864 & w17838;
assign w16701 = ~w3499 & ~w7208;
assign w16702 = ~pi0959 & w3791;
assign w16703 = pi0054 & pi0050;
assign w16704 = ~w6501 & ~w7762;
assign w16705 = ~w17692 & ~w3608;
assign w16706 = ~w16480 & ~w10122;
assign w16707 = ~w6357 & w16502;
assign w16708 = ~w3021 & w5652;
assign w16709 = w11383 & w13441;
assign w16710 = (pi1789 & w7215) | (pi1789 & w691) | (w7215 & w691);
assign w16711 = ~w7177 & ~w11056;
assign w16712 = w4535 & w6006;
assign w16713 = w15604 & w7521;
assign w16714 = pi1337 & ~pi0263;
assign w16715 = w41 & w2144;
assign w16716 = w7077 & ~w6680;
assign w16717 = ~w7364 & ~w14433;
assign w16718 = w13231 & w1217;
assign w16719 = ~w12493 & ~w9915;
assign w16720 = ~w18469 & ~w14825;
assign w16721 = ~pi2757 & w10862;
assign w16722 = pi1540 & ~w17935;
assign w16723 = pi1586 & ~w14918;
assign w16724 = (pi1090 & ~w13509) | (pi1090 & w6124) | (~w13509 & w6124);
assign w16725 = ~pi1383 & ~pi2913;
assign w16726 = ~pi0702 & w3106;
assign w16727 = ~w6235 & ~w3811;
assign w16728 = ~pi0130 & pi0153;
assign w16729 = ~pi1798 & ~pi1806;
assign w16730 = ~pi1400 & w8341;
assign w16731 = ~w8511 & ~w9843;
assign w16732 = ~w11576 & w11194;
assign w16733 = w11383 & w12504;
assign w16734 = ~w18218 & ~w16595;
assign w16735 = ~w6560 & ~w8519;
assign w16736 = w914 & w13232;
assign w16737 = w7353 & w9562;
assign w16738 = ~pi3165 & w15048;
assign w16739 = pi2424 & ~w10158;
assign w16740 = ~w4114 & ~w9472;
assign w16741 = ~w5189 & ~pi1199;
assign w16742 = pi1725 & ~pi1796;
assign w16743 = w18077 & w18210;
assign w16744 = w13840 & pi1700;
assign w16745 = ~w4619 & ~w3637;
assign w16746 = pi2588 & ~w5274;
assign w16747 = pi2693 & ~w226;
assign w16748 = ~pi0700 & w3106;
assign w16749 = w16778 & ~w11291;
assign w16750 = ~pi3162 & w12427;
assign w16751 = w17665 & ~w15208;
assign w16752 = ~pi2108 & w12755;
assign w16753 = w12460 & w1141;
assign w16754 = ~w4451 & ~w8048;
assign w16755 = ~pi3353 & w9781;
assign w16756 = pi3076 & ~w16502;
assign w16757 = ~w12080 & ~w16314;
assign w16758 = ~pi3048 & w261;
assign w16759 = ~pi1228 & w2235;
assign w16760 = ~pi2222 & w2151;
assign w16761 = ~w16059 & ~w1571;
assign w16762 = ~pi1039 & w6200;
assign w16763 = ~w11059 & ~w10643;
assign w16764 = w5517 & w5504;
assign w16765 = ~pi2050 & w13204;
assign w16766 = pi1329 & w458;
assign w16767 = ~w16144 & ~w11659;
assign w16768 = ~w3000 & ~pi2672;
assign w16769 = w6857 & w13233;
assign w16770 = ~w18416 & w3201;
assign w16771 = pi3125 & w7177;
assign w16772 = pi3158 & w2732;
assign w16773 = (pi1145 & ~w5437) | (pi1145 & w5470) | (~w5437 & w5470);
assign w16774 = ~w783 & ~w1434;
assign w16775 = w7703 & w17051;
assign w16776 = pi1503 & ~w16922;
assign w16777 = ~pi3097 & w261;
assign w16778 = ~w16920 & ~w14420;
assign w16779 = ~w10540 & ~pi0083;
assign w16780 = ~pi0424 & w17173;
assign w16781 = ~w16857 & w10284;
assign w16782 = pi1679 & w3163;
assign w16783 = pi1254 & pi3232;
assign w16784 = ~w12608 & ~w8197;
assign w16785 = ~w12764 & ~w11950;
assign w16786 = ~w667 & w4796;
assign w16787 = ~w9920 & ~w17301;
assign w16788 = ~w8483 & ~w12294;
assign w16789 = w1127 & ~w17411;
assign w16790 = ~pi1676 & w7388;
assign w16791 = pi2474 & ~w14833;
assign w16792 = ~w15664 & ~w2119;
assign w16793 = ~pi0885 & w1126;
assign w16794 = ~w13789 & ~w6390;
assign w16795 = (pi1010 & ~w13509) | (pi1010 & w4428) | (~w13509 & w4428);
assign w16796 = w9414 & w614;
assign w16797 = w16278 & ~w10235;
assign w16798 = (pi0672 & ~w13509) | (pi0672 & w17881) | (~w13509 & w17881);
assign w16799 = w7077 & ~w6033;
assign w16800 = ~pi2813 & w13343;
assign w16801 = (pi1376 & w13142) | (pi1376 & w1997) | (w13142 & w1997);
assign w16802 = ~w15949 & ~w15378;
assign w16803 = pi2371 & ~w4508;
assign w16804 = ~w6195 & w1959;
assign w16805 = (pi0554 & ~w13509) | (pi0554 & w17139) | (~w13509 & w17139);
assign w16806 = pi1848 & ~w12558;
assign w16807 = pi3516 & w3919;
assign w16808 = w8789 & w16442;
assign w16809 = ~w5507 & ~w5257;
assign w16810 = w12277 & w6185;
assign w16811 = (~pi0077 & w13707) | (~pi0077 & w8859) | (w13707 & w8859);
assign w16812 = ~w6570 & ~w2212;
assign w16813 = pi1667 & w1924;
assign w16814 = ~pi3432 & w15036;
assign w16815 = pi2949 & w7912;
assign w16816 = ~w13501 & ~w12594;
assign w16817 = ~pi3147 & w3982;
assign w16818 = ~w15530 & ~w3936;
assign w16819 = ~w13960 & ~w12546;
assign w16820 = ~pi0096 & w9284;
assign w16821 = pi0097 & w9284;
assign w16822 = ~w9240 & w17306;
assign w16823 = w3046 & w16054;
assign w16824 = ~w16222 & ~w2331;
assign w16825 = (pi0714 & ~w13509) | (pi0714 & w8518) | (~w13509 & w8518);
assign w16826 = ~w1325 & w6241;
assign w16827 = ~w12511 & ~w2057;
assign w16828 = pi3025 & w16502;
assign w16829 = w15808 & ~w13028;
assign w16830 = ~w8046 & w917;
assign w16831 = w13509 & w17903;
assign w16832 = ~pi3142 & w17993;
assign w16833 = w6857 & w9065;
assign w16834 = (~pi0331 & ~w6857) | (~pi0331 & w14392) | (~w6857 & w14392);
assign w16835 = w1962 & ~w6647;
assign w16836 = w14460 & w4200;
assign w16837 = ~pi2155 & w13065;
assign w16838 = (pi1037 & ~w13509) | (pi1037 & w2035) | (~w13509 & w2035);
assign w16839 = ~w4819 & ~w10976;
assign w16840 = w16575 & w10218;
assign w16841 = ~w7912 & ~w2640;
assign w16842 = pi1555 & ~w13753;
assign w16843 = ~w1368 & ~pi0482;
assign w16844 = ~w8572 & ~w2198;
assign w16845 = w15122 & ~pi2635;
assign w16846 = w16278 & ~w1236;
assign w16847 = pi0269 & w5113;
assign w16848 = ~w14307 & ~w2337;
assign w16849 = w16363 & w13319;
assign w16850 = w17683 & w14078;
assign w16851 = w3243 & pi0312;
assign w16852 = ~w1687 & ~w12910;
assign w16853 = w15393 & w13819;
assign w16854 = ~w1145 & ~w5735;
assign w16855 = w13509 & w16462;
assign w16856 = ~pi3135 & w13730;
assign w16857 = ~w17577 & w1827;
assign w16858 = ~w8013 & ~w2798;
assign w16859 = ~pi1251 & w11655;
assign w16860 = pi1252 & w11655;
assign w16861 = ~w7685 & ~w15941;
assign w16862 = ~w17947 & w15556;
assign w16863 = ~w8358 & ~w12262;
assign w16864 = pi1503 & ~w13753;
assign w16865 = pi2060 & ~w4508;
assign w16866 = w3384 & ~w8607;
assign w16867 = ~w6568 & ~w13296;
assign w16868 = ~w7534 & ~w17415;
assign w16869 = ~w7039 & w12136;
assign w16870 = w7318 & w799;
assign w16871 = ~pi3146 & w3982;
assign w16872 = w11383 & w14184;
assign w16873 = ~w11742 & w8499;
assign w16874 = w10818 & ~w6130;
assign w16875 = ~w3203 & pi0582;
assign w16876 = ~pi3154 & w8515;
assign w16877 = ~w1829 & ~w2440;
assign w16878 = w17351 & w10216;
assign w16879 = ~w8382 & ~w3271;
assign w16880 = pi1481 & w13753;
assign w16881 = ~w6029 & ~w7193;
assign w16882 = ~w5183 & ~w3548;
assign w16883 = (~pi0961 & ~w13509) | (~pi0961 & w16115) | (~w13509 & w16115);
assign w16884 = w3585 & w6599;
assign w16885 = ~pi2137 & w12941;
assign w16886 = ~w15 & ~w673;
assign w16887 = ~w10332 & ~w7091;
assign w16888 = ~w15918 & w4099;
assign w16889 = ~w14704 & ~w17074;
assign w16890 = ~w16108 & ~w18447;
assign w16891 = ~w13341 & ~w11730;
assign w16892 = ~pi1725 & ~w487;
assign w16893 = w12689 & w3481;
assign w16894 = ~pi0946 & w14641;
assign w16895 = pi2682 & ~w11406;
assign w16896 = ~w8948 & ~w13944;
assign w16897 = (w13368 & w5855) | (w13368 & w349) | (w5855 & w349);
assign w16898 = w13436 & w2661;
assign w16899 = w384 & w5832;
assign w16900 = w13509 & w5826;
assign w16901 = pi3186 & pi3248;
assign w16902 = ~pi2336 & w12755;
assign w16903 = w6857 & w8008;
assign w16904 = ~pi3165 & w17387;
assign w16905 = pi2834 & w15191;
assign w16906 = pi2033 & ~w17646;
assign w16907 = ~w11684 & ~w15408;
assign w16908 = pi1775 & pi3143;
assign w16909 = ~w571 & ~w3390;
assign w16910 = pi3153 & w3987;
assign w16911 = ~pi0583 & w795;
assign w16912 = ~pi3019 & ~pi3207;
assign w16913 = w14648 & ~pi2610;
assign w16914 = w5453 & pi2580;
assign w16915 = w934 & pi0426;
assign w16916 = w5453 & pi2885;
assign w16917 = ~w18278 & ~w10028;
assign w16918 = ~pi2038 & w7455;
assign w16919 = pi2822 & ~w11406;
assign w16920 = (w12775 & ~w9636) | (w12775 & w14594) | (~w9636 & w14594);
assign w16921 = ~pi0483 & pi3389;
assign w16922 = w5043 & w16499;
assign w16923 = ~w2194 & w9840;
assign w16924 = (~pi0333 & ~w6857) | (~pi0333 & w12902) | (~w6857 & w12902);
assign w16925 = ~pi1832 & w5384;
assign w16926 = ~w7996 & w10009;
assign w16927 = pi0086 & w9284;
assign w16928 = ~w14377 & w16306;
assign w16929 = (~pi0964 & ~w13509) | (~pi0964 & w14084) | (~w13509 & w14084);
assign w16930 = (pi1148 & ~w5437) | (pi1148 & w16156) | (~w5437 & w16156);
assign w16931 = pi2096 & ~w4420;
assign w16932 = w5189 & ~w3374;
assign w16933 = ~w4543 & ~w1205;
assign w16934 = ~w1957 & ~w8372;
assign w16935 = ~w3211 & ~w11482;
assign w16936 = pi3133 & w8113;
assign w16937 = ~w15805 & w12008;
assign w16938 = ~w16925 & ~w8327;
assign w16939 = (~w11159 & ~w8324) | (~w11159 & w18555) | (~w8324 & w18555);
assign w16940 = ~pi1214 & pi3193;
assign w16941 = ~w7638 & ~w2372;
assign w16942 = ~pi3330 & w18259;
assign w16943 = w2653 & w21;
assign w16944 = ~pi0565 & w11739;
assign w16945 = w13509 & w9528;
assign w16946 = w6359 & ~w13641;
assign w16947 = (~w15312 & ~w5517) | (~w15312 & w615) | (~w5517 & w615);
assign w16948 = w17248 & ~w16498;
assign w16949 = ~pi2915 & ~pi2953;
assign w16950 = ~w9280 & w11156;
assign w16951 = (pi1861 & w2014) | (pi1861 & w16347) | (w2014 & w16347);
assign w16952 = pi1990 & ~w9414;
assign w16953 = pi2826 & ~w11406;
assign w16954 = ~w4254 & ~w10109;
assign w16955 = pi0142 & ~pi0191;
assign w16956 = ~w9401 & ~w5024;
assign w16957 = w13509 & w14630;
assign w16958 = pi0309 & ~pi0265;
assign w16959 = ~w18062 & ~w10403;
assign w16960 = pi1623 & ~w7090;
assign w16961 = ~w17077 & ~w14763;
assign w16962 = ~pi2345 & w17439;
assign w16963 = ~w6195 & w7035;
assign w16964 = w13509 & w11927;
assign w16965 = (~pi0975 & ~w1475) | (~pi0975 & w10841) | (~w1475 & w10841);
assign w16966 = pi3138 & w9520;
assign w16967 = w11383 & w8935;
assign w16968 = w10554 & w13915;
assign w16969 = (pi1241 & w11655) | (pi1241 & w7783) | (w11655 & w7783);
assign w16970 = ~w11957 & w6133;
assign w16971 = ~w4239 & ~w71;
assign w16972 = ~pi3058 & w15235;
assign w16973 = ~w1962 & pi0653;
assign w16974 = pi1755 & pi3165;
assign w16975 = w412 & w9407;
assign w16976 = ~w7878 & ~w8943;
assign w16977 = pi2162 & ~w11671;
assign w16978 = pi1726 & w1924;
assign w16979 = w12610 & w698;
assign w16980 = w968 & ~pi0352;
assign w16981 = ~w17804 & ~w2526;
assign w16982 = pi0089 & w3748;
assign w16983 = (~pi0514 & w17577) | (~pi0514 & w13587) | (w17577 & w13587);
assign w16984 = ~w15685 & ~w7871;
assign w16985 = ~w3975 & ~w8720;
assign w16986 = pi2546 & w605;
assign w16987 = w11247 & w17295;
assign w16988 = ~w9286 & ~w9814;
assign w16989 = pi2013 & ~w14833;
assign w16990 = pi2666 & ~w6463;
assign w16991 = pi1765 & ~w14951;
assign w16992 = pi2239 & ~w11735;
assign w16993 = ~w5186 & ~w14372;
assign w16994 = ~w16592 & ~w16114;
assign w16995 = ~pi1775 & ~pi3143;
assign w16996 = ~w10738 & ~w4677;
assign w16997 = ~pi2903 & w15122;
assign w16998 = pi1511 & ~w13753;
assign w16999 = (pi0588 & ~w13509) | (pi0588 & w5729) | (~w13509 & w5729);
assign w17000 = ~pi3337 & w6448;
assign w17001 = ~pi0895 & w1126;
assign w17002 = ~w15812 & ~w2840;
assign w17003 = ~w6195 & w3838;
assign w17004 = ~w4074 & ~w3438;
assign w17005 = ~pi2277 & w3019;
assign w17006 = ~w1180 & ~w5689;
assign w17007 = pi0257 & w5113;
assign w17008 = ~pi0611 & w12825;
assign w17009 = ~pi3060 & w15235;
assign w17010 = pi1746 & ~w226;
assign w17011 = ~pi3346 & w9781;
assign w17012 = ~w10962 & ~w2031;
assign w17013 = ~w14170 & ~w14540;
assign w17014 = ~pi2837 & w13343;
assign w17015 = w1368 & pi0388;
assign w17016 = w14647 & w2878;
assign w17017 = pi2575 & ~w5274;
assign w17018 = w17277 & w14902;
assign w17019 = (pi0725 & ~w13509) | (pi0725 & w15771) | (~w13509 & w15771);
assign w17020 = ~w9584 & ~w5942;
assign w17021 = ~w13327 & w3790;
assign w17022 = pi1538 & w13753;
assign w17023 = pi2559 & ~w5274;
assign w17024 = pi1372 & w9653;
assign w17025 = ~w7319 & ~w4379;
assign w17026 = ~pi0334 & w2196;
assign w17027 = w16506 & ~w6922;
assign w17028 = ~w9680 & w5738;
assign w17029 = ~w8031 & ~w14149;
assign w17030 = ~w2923 & ~w12918;
assign w17031 = pi2735 & ~w261;
assign w17032 = ~w15651 & ~w5417;
assign w17033 = ~pi2451 & w9340;
assign w17034 = w16506 & pi2958;
assign w17035 = pi0033 & ~w14148;
assign w17036 = pi0486 & pi1133;
assign w17037 = pi3154 & w3987;
assign w17038 = w712 & w9762;
assign w17039 = w11383 & w7709;
assign w17040 = ~w10833 & ~w9529;
assign w17041 = ~w16549 & ~w12697;
assign w17042 = pi2761 & w605;
assign w17043 = ~w579 & ~w9513;
assign w17044 = ~pi3169 & w15048;
assign w17045 = ~w165 & ~w11919;
assign w17046 = ~w17332 & ~w15803;
assign w17047 = ~w18283 & ~w14530;
assign w17048 = ~w13837 & ~w9510;
assign w17049 = ~w17499 & ~w11757;
assign w17050 = ~w1142 & w10115;
assign w17051 = ~w15122 & ~pi2675;
assign w17052 = w10189 & pi0402;
assign w17053 = ~w9133 & ~w5318;
assign w17054 = ~pi3108 & w16502;
assign w17055 = ~pi3111 & pi3112;
assign w17056 = ~pi3346 & w14918;
assign w17057 = ~w5776 & w16464;
assign w17058 = ~w1113 & w13077;
assign w17059 = pi1288 & pi1345;
assign w17060 = pi1541 & w13753;
assign w17061 = ~pi2414 & w5075;
assign w17062 = pi1337 & w1341;
assign w17063 = pi0014 & ~w14148;
assign w17064 = w12460 & w18122;
assign w17065 = ~w3203 & pi0592;
assign w17066 = ~w2883 & ~w6005;
assign w17067 = w14109 & pi0440;
assign w17068 = ~pi3090 & w15235;
assign w17069 = ~pi0295 & w2196;
assign w17070 = w18123 & w2753;
assign w17071 = ~pi2407 & w13204;
assign w17072 = w6697 & ~w9852;
assign w17073 = ~w8676 & ~w925;
assign w17074 = ~pi3085 & w3555;
assign w17075 = w11383 & w5920;
assign w17076 = ~w1064 & w13903;
assign w17077 = pi1757 & ~w8829;
assign w17078 = ~pi2259 & w13065;
assign w17079 = ~w9190 & ~w4815;
assign w17080 = w8256 & ~w3047;
assign w17081 = w16278 & ~w14597;
assign w17082 = pi1697 & ~w11760;
assign w17083 = pi2921 & w6045;
assign w17084 = pi0049 & pi0058;
assign w17085 = ~w9593 & ~w7781;
assign w17086 = ~w14139 & ~w17362;
assign w17087 = ~pi3055 & w226;
assign w17088 = pi1603 & w13753;
assign w17089 = (pi0759 & ~w13509) | (pi0759 & w4166) | (~w13509 & w4166);
assign w17090 = pi1755 & ~w619;
assign w17091 = pi2333 & ~w11671;
assign w17092 = pi2966 & ~w3987;
assign w17093 = w18220 & w11005;
assign w17094 = ~w10749 & ~w13393;
assign w17095 = (~pi1152 & ~w13509) | (~pi1152 & w1847) | (~w13509 & w1847);
assign w17096 = w1463 & ~w994;
assign w17097 = ~w2286 & ~w12536;
assign w17098 = ~pi3415 & w15036;
assign w17099 = ~w964 & ~w4158;
assign w17100 = ~pi1828 & ~w9165;
assign w17101 = ~w10474 & ~w17674;
assign w17102 = w9440 & pi0144;
assign w17103 = w6111 & w2441;
assign w17104 = ~w458 & w17456;
assign w17105 = ~w1154 & ~w12181;
assign w17106 = pi3015 & w16502;
assign w17107 = (~pi0290 & ~w6857) | (~pi0290 & w13307) | (~w6857 & w13307);
assign w17108 = w2341 & ~w7449;
assign w17109 = ~w15914 & ~w17126;
assign w17110 = ~w17422 & ~w4243;
assign w17111 = w13509 & w8677;
assign w17112 = ~w18135 & ~w12743;
assign w17113 = ~w6919 & ~w12267;
assign w17114 = pi2006 & ~w14833;
assign w17115 = ~pi3151 & ~w4020;
assign w17116 = pi2743 & ~w6463;
assign w17117 = ~w2907 & w901;
assign w17118 = ~w11999 & ~w12167;
assign w17119 = pi1673 & ~w4058;
assign w17120 = pi2920 & ~w3987;
assign w17121 = ~pi3157 & w15839;
assign w17122 = ~pi2967 & pi3075;
assign w17123 = ~pi2897 & w15122;
assign w17124 = (w229 & ~w11247) | (w229 & w3289) | (~w11247 & w3289);
assign w17125 = ~w8588 & w18123;
assign w17126 = pi2011 & ~w14833;
assign w17127 = ~w8049 & ~w6102;
assign w17128 = ~w3198 & ~w10282;
assign w17129 = ~w12638 & w16479;
assign w17130 = ~w458 & w13004;
assign w17131 = w7307 & w16768;
assign w17132 = ~w12023 & w89;
assign w17133 = ~pi3135 & w13570;
assign w17134 = ~w16506 & pi1143;
assign w17135 = (pi1149 & ~w5437) | (pi1149 & w1075) | (~w5437 & w1075);
assign w17136 = ~pi0891 & w1126;
assign w17137 = ~w5560 & w8902;
assign w17138 = ~w10580 & w13169;
assign w17139 = ~w13231 & pi0554;
assign w17140 = ~pi0282 & w2196;
assign w17141 = w6857 & w7092;
assign w17142 = ~w17381 & ~w14498;
assign w17143 = w7307 & w12682;
assign w17144 = pi2082 & ~w17683;
assign w17145 = pi1332 & ~w12166;
assign w17146 = ~w14560 & pi0212;
assign w17147 = ~w3676 & ~w2001;
assign w17148 = ~w5569 & ~w3744;
assign w17149 = w13509 & w4799;
assign w17150 = ~w4286 & ~w12925;
assign w17151 = (pi0570 & ~w13509) | (pi0570 & w3244) | (~w13509 & w3244);
assign w17152 = ~w14247 & ~w6543;
assign w17153 = w11383 & w7147;
assign w17154 = ~w2846 & w1605;
assign w17155 = pi2567 & ~w5274;
assign w17156 = ~w11380 & ~w7974;
assign w17157 = ~pi3163 & w4310;
assign w17158 = pi1407 & ~pi2913;
assign w17159 = w10189 & pi0391;
assign w17160 = ~w14844 & w6114;
assign w17161 = ~w835 & ~w10483;
assign w17162 = ~w9948 & ~w8086;
assign w17163 = ~pi1164 & pi3222;
assign w17164 = ~pi0995 & w795;
assign w17165 = ~w3669 & ~w9620;
assign w17166 = ~w6835 & ~w16975;
assign w17167 = (pi1791 & w7215) | (pi1791 & w10943) | (w7215 & w10943);
assign w17168 = ~w17665 & ~w8628;
assign w17169 = ~w8167 & ~w8930;
assign w17170 = pi3170 & w18497;
assign w17171 = pi1337 & pi0303;
assign w17172 = pi3151 & w2732;
assign w17173 = w8616 & w8949;
assign w17174 = w13509 & w6403;
assign w17175 = ~w2485 & ~w11035;
assign w17176 = ~pi3290 & w18259;
assign w17177 = w9440 & pi0188;
assign w17178 = ~w10742 & w16030;
assign w17179 = ~w16409 & ~w5195;
assign w17180 = ~w7077 & pi0903;
assign w17181 = ~w8815 & ~w11391;
assign w17182 = ~pi3096 & w16815;
assign w17183 = w1127 & ~w4500;
assign w17184 = pi2359 & ~w4508;
assign w17185 = pi1716 & pi3164;
assign w17186 = ~pi2377 & w17439;
assign w17187 = pi1550 & ~w17935;
assign w17188 = ~pi1310 & ~w8804;
assign w17189 = ~pi2967 & w236;
assign w17190 = ~w14648 & ~pi2624;
assign w17191 = ~w9002 & ~w2457;
assign w17192 = pi2000 & ~w9414;
assign w17193 = ~w11674 & ~w34;
assign w17194 = ~w14174 & ~w1025;
assign w17195 = w539 & ~w5258;
assign w17196 = ~w5560 & w12415;
assign w17197 = w12515 & w9984;
assign w17198 = ~w12202 & ~w2864;
assign w17199 = ~w7137 & ~w237;
assign w17200 = pi2044 & ~w10158;
assign w17201 = pi2423 & ~w10158;
assign w17202 = ~w1653 & ~w11769;
assign w17203 = pi0511 & pi1157;
assign w17204 = ~pi1030 & w17490;
assign w17205 = pi1266 & ~pi1311;
assign w17206 = w13509 & w3879;
assign w17207 = ~w10108 & pi1188;
assign w17208 = (pi0815 & ~w13509) | (pi0815 & w10795) | (~w13509 & w10795);
assign w17209 = ~w12100 & ~w4449;
assign w17210 = ~w148 & ~w14563;
assign w17211 = w8658 & pi1787;
assign w17212 = ~pi3155 & w17387;
assign w17213 = ~w3000 & w13695;
assign w17214 = w13509 & w14226;
assign w17215 = w13509 & w14227;
assign w17216 = ~pi2946 & w3555;
assign w17217 = ~pi2151 & w13065;
assign w17218 = ~pi1838 & w5075;
assign w17219 = pi2126 & ~w18123;
assign w17220 = ~w15677 & ~w7712;
assign w17221 = ~w2353 & ~w7133;
assign w17222 = ~pi2333 & w13065;
assign w17223 = ~w16773 & ~w9841;
assign w17224 = (~pi0275 & ~w6857) | (~pi0275 & w17746) | (~w6857 & w17746);
assign w17225 = pi1810 & ~w9520;
assign w17226 = ~pi1834 & ~w10158;
assign w17227 = ~w13214 & ~w13537;
assign w17228 = ~pi3318 & w16922;
assign w17229 = ~w5306 & ~w5022;
assign w17230 = pi0109 & w9284;
assign w17231 = ~pi0612 & w12825;
assign w17232 = ~w15317 & ~w3004;
assign w17233 = w13509 & w14297;
assign w17234 = ~pi0634 & w14641;
assign w17235 = ~w13353 & w13483;
assign w17236 = ~w12040 & pi1020;
assign w17237 = (pi0885 & ~w13509) | (pi0885 & w16338) | (~w13509 & w16338);
assign w17238 = pi2380 & ~w412;
assign w17239 = ~pi2956 & pi3205;
assign w17240 = w17955 & w4828;
assign w17241 = pi2520 & w4140;
assign w17242 = (~pi2920 & ~w384) | (~pi2920 & w8568) | (~w384 & w8568);
assign w17243 = w6857 & w586;
assign w17244 = ~w9216 & ~w8629;
assign w17245 = ~w8622 & ~w6516;
assign w17246 = ~w6667 & ~w10010;
assign w17247 = w13509 & w324;
assign w17248 = w2613 & w13867;
assign w17249 = pi1144 & w9420;
assign w17250 = ~w12331 & ~w15891;
assign w17251 = ~w11133 & ~w6356;
assign w17252 = pi0315 & ~pi3235;
assign w17253 = ~w6968 & ~w1845;
assign w17254 = w1368 & pi0405;
assign w17255 = w13509 & w399;
assign w17256 = pi3155 & w3987;
assign w17257 = ~w6785 & ~pi0966;
assign w17258 = pi2534 & w14148;
assign w17259 = pi2960 & ~w13367;
assign w17260 = ~w17063 & ~w5655;
assign w17261 = ~w11307 & ~w6757;
assign w17262 = ~w10127 & ~w4484;
assign w17263 = pi2170 & ~w15271;
assign w17264 = ~w17665 & ~w597;
assign w17265 = ~w5628 & ~w5337;
assign w17266 = w12670 & w4342;
assign w17267 = ~pi3050 & w226;
assign w17268 = ~w16506 & pi1185;
assign w17269 = w2991 & w2127;
assign w17270 = pi3160 & ~pi3475;
assign w17271 = ~pi2662 & w17213;
assign w17272 = ~w112 & ~w15125;
assign w17273 = ~w18242 & ~w17858;
assign w17274 = ~pi2032 & w7455;
assign w17275 = ~w16516 & ~w9535;
assign w17276 = pi2065 & ~w4508;
assign w17277 = ~w9875 & w4037;
assign w17278 = w1516 & w10990;
assign w17279 = w3831 & w1618;
assign w17280 = w2725 & ~w6033;
assign w17281 = pi1441 & ~w6448;
assign w17282 = pi1636 & ~w18259;
assign w17283 = ~w9783 & ~w4225;
assign w17284 = w2341 & ~w6922;
assign w17285 = ~w7150 & ~w15721;
assign w17286 = ~w15715 & ~w5424;
assign w17287 = ~w13292 & ~w463;
assign w17288 = ~pi0543 & w9110;
assign w17289 = pi1217 & ~w16725;
assign w17290 = ~w6697 & pi1012;
assign w17291 = w709 & pi1871;
assign w17292 = ~w733 & ~w3967;
assign w17293 = w9440 & pi0176;
assign w17294 = ~w17103 & ~w4331;
assign w17295 = w5874 & pi0256;
assign w17296 = ~pi1935 & w12755;
assign w17297 = pi2664 & ~w15235;
assign w17298 = pi3147 & w2253;
assign w17299 = (pi0782 & ~w13509) | (pi0782 & w6952) | (~w13509 & w6952);
assign w17300 = pi2659 & ~w15235;
assign w17301 = ~pi3321 & w17935;
assign w17302 = ~pi1353 & w7177;
assign w17303 = pi3021 & w16502;
assign w17304 = ~pi3020 & w16502;
assign w17305 = ~w17860 & w13178;
assign w17306 = (~w12844 & ~w5517) | (~w12844 & w16295) | (~w5517 & w16295);
assign w17307 = w11383 & w90;
assign w17308 = ~w5106 & ~w8567;
assign w17309 = ~pi1701 & w4667;
assign w17310 = pi2307 & ~w18123;
assign w17311 = w1391 & ~w7449;
assign w17312 = pi1428 & ~w6072;
assign w17313 = ~w546 & ~w13173;
assign w17314 = w14228 & ~w7020;
assign w17315 = pi1712 & ~w7946;
assign w17316 = ~w8708 & ~w2575;
assign w17317 = (pi0875 & ~w13509) | (pi0875 & w1627) | (~w13509 & w1627);
assign w17318 = ~w16458 & ~w6962;
assign w17319 = ~w2341 & pi0836;
assign w17320 = pi3176 & w4140;
assign w17321 = (pi0667 & ~w13509) | (pi0667 & w2765) | (~w13509 & w2765);
assign w17322 = ~w11197 & ~w7604;
assign w17323 = w11405 & w15964;
assign w17324 = w13509 & w11753;
assign w17325 = pi2025 & ~w17646;
assign w17326 = w4936 & pi0487;
assign w17327 = pi2989 & ~w5366;
assign w17328 = pi0105 & w3748;
assign w17329 = ~w11474 & ~w8763;
assign w17330 = ~pi2458 & w5384;
assign w17331 = ~pi0633 & w14641;
assign w17332 = pi2646 & ~w226;
assign w17333 = ~pi2332 & w16041;
assign w17334 = ~w11268 & ~w13276;
assign w17335 = ~w14229 & ~w10737;
assign w17336 = ~w8139 & w7735;
assign w17337 = pi2462 & ~w14524;
assign w17338 = pi2769 & ~w6463;
assign w17339 = ~w2725 & pi1087;
assign w17340 = ~pi3328 & w7090;
assign w17341 = ~w5560 & w12841;
assign w17342 = ~w578 & ~w3269;
assign w17343 = ~w3544 & ~w13367;
assign w17344 = pi1294 & pi1345;
assign w17345 = ~w5456 & ~w2737;
assign w17346 = pi1439 & ~w13753;
assign w17347 = w12354 & w7508;
assign w17348 = ~w913 & ~w9416;
assign w17349 = w12436 & ~w10784;
assign w17350 = ~w4888 & ~w8594;
assign w17351 = ~w8706 & ~w7288;
assign w17352 = pi2541 & w14148;
assign w17353 = ~pi3318 & w6072;
assign w17354 = pi2824 & ~w226;
assign w17355 = w13509 & w14538;
assign w17356 = ~w9059 & ~w14751;
assign w17357 = ~w5691 & ~w1386;
assign w17358 = w1127 & ~w13513;
assign w17359 = ~w1085 & ~w9591;
assign w17360 = ~w12460 & w1689;
assign w17361 = ~w11854 & ~w13257;
assign w17362 = w13509 & w17943;
assign w17363 = pi0063 & ~w14148;
assign w17364 = ~pi3101 & w226;
assign w17365 = ~pi3410 & w15036;
assign w17366 = w2725 & ~w15173;
assign w17367 = ~pi1408 & ~pi2913;
assign w17368 = ~w11154 & ~w5857;
assign w17369 = ~w14497 & ~w2215;
assign w17370 = pi0988 & ~pi3362;
assign w17371 = pi2334 & ~w4508;
assign w17372 = w6857 & w12701;
assign w17373 = pi1871 & ~w15036;
assign w17374 = w7703 & w5956;
assign w17375 = ~w15349 & ~w8326;
assign w17376 = w14738 & w14374;
assign w17377 = pi0268 & w5113;
assign w17378 = pi0253 & pi0254;
assign w17379 = w13423 & ~w17945;
assign w17380 = (~w11235 & ~w5517) | (~w11235 & w3746) | (~w5517 & w3746);
assign w17381 = (pi1886 & w2014) | (pi1886 & w9492) | (w2014 & w9492);
assign w17382 = w7177 & w14565;
assign w17383 = w11735 & w9407;
assign w17384 = pi3071 & ~w15513;
assign w17385 = w13509 & w11191;
assign w17386 = ~w7311 & ~w6424;
assign w17387 = ~w4020 & w11735;
assign w17388 = w798 & w16301;
assign w17389 = ~pi3169 & w4310;
assign w17390 = pi3150 & w9520;
assign w17391 = (pi0308 & ~w325) | (pi0308 & w15990) | (~w325 & w15990);
assign w17392 = ~pi0981 & w1126;
assign w17393 = ~w6697 & pi0675;
assign w17394 = ~pi1828 & ~w15450;
assign w17395 = pi1268 & ~pi2959;
assign w17396 = pi1152 & ~pi1176;
assign w17397 = w968 & ~pi0282;
assign w17398 = ~pi2268 & w3019;
assign w17399 = ~w10250 & ~w7465;
assign w17400 = ~pi2272 & w17439;
assign w17401 = ~w14228 & pi0618;
assign w17402 = w12040 & ~w9852;
assign w17403 = (~w13367 & w2605) | (~w13367 & w11985) | (w2605 & w11985);
assign w17404 = pi2670 & ~w6463;
assign w17405 = ~pi3328 & w14918;
assign w17406 = w13509 & w8889;
assign w17407 = pi1213 & ~w5769;
assign w17408 = ~pi3171 & w12427;
assign w17409 = w11209 & ~w15390;
assign w17410 = ~pi3166 & w12427;
assign w17411 = pi1553 & w13753;
assign w17412 = (pi1065 & ~w13509) | (pi1065 & w5755) | (~w13509 & w5755);
assign w17413 = w7498 & w18213;
assign w17414 = (w10571 & ~w3114) | (w10571 & w13229) | (~w3114 & w13229);
assign w17415 = (~pi0330 & ~w6857) | (~pi0330 & w9855) | (~w6857 & w9855);
assign w17416 = pi2080 & ~w17683;
assign w17417 = pi2966 & pi2556;
assign w17418 = pi2729 & ~w261;
assign w17419 = ~w14960 & w3382;
assign w17420 = pi2354 & ~w4420;
assign w17421 = ~pi2774 & w13343;
assign w17422 = w12460 & w2724;
assign w17423 = w8658 & pi1757;
assign w17424 = ~w4506 & ~w3261;
assign w17425 = ~w3100 & ~w1828;
assign w17426 = ~w15184 & ~w3015;
assign w17427 = w12460 & w11561;
assign w17428 = w15518 & w7240;
assign w17429 = ~pi0556 & w11739;
assign w17430 = w8337 & pi3291;
assign w17431 = w968 & ~pi0334;
assign w17432 = ~w6655 & ~w17329;
assign w17433 = w2439 & w17272;
assign w17434 = (pi1141 & ~w5437) | (pi1141 & w9990) | (~w5437 & w9990);
assign w17435 = ~pi3162 & w15048;
assign w17436 = ~w6265 & ~w7682;
assign w17437 = ~w15754 & ~w10004;
assign w17438 = ~pi1212 & pi1213;
assign w17439 = w2425 & w5410;
assign w17440 = w9720 & pi1711;
assign w17441 = ~w2492 & ~w12769;
assign w17442 = pi2835 & ~w11406;
assign w17443 = ~w7286 & ~w11790;
assign w17444 = ~pi3067 & pi3147;
assign w17445 = pi1334 & ~w3358;
assign w17446 = ~pi0640 & w3791;
assign w17447 = pi1875 & ~w458;
assign w17448 = ~w8957 & ~w16796;
assign w17449 = ~w2860 & ~w11905;
assign w17450 = w2742 & ~w15293;
assign w17451 = ~w2725 & pi0786;
assign w17452 = ~w5757 & ~w385;
assign w17453 = pi1913 & ~w15271;
assign w17454 = w1962 & ~w10235;
assign w17455 = ~w8435 & ~w9408;
assign w17456 = w13072 & w13679;
assign w17457 = pi3135 & w8113;
assign w17458 = pi1526 & ~w14918;
assign w17459 = w15808 & ~w15296;
assign w17460 = w13509 & w14639;
assign w17461 = w7703 & w15660;
assign w17462 = w10988 & w14074;
assign w17463 = pi1774 & ~w10389;
assign w17464 = ~w12180 & ~w11236;
assign w17465 = (pi0610 & ~w13509) | (pi0610 & w6855) | (~w13509 & w6855);
assign w17466 = pi1654 & ~w13753;
assign w17467 = pi2124 & ~w412;
assign w17468 = ~w15375 & w18385;
assign w17469 = pi0003 & ~w14148;
assign w17470 = pi1258 & w5031;
assign w17471 = ~w6697 & pi0912;
assign w17472 = ~w16204 & ~w51;
assign w17473 = pi2215 & ~w15271;
assign w17474 = ~pi2991 & ~w8571;
assign w17475 = w9074 & w11173;
assign w17476 = ~pi0352 & w4058;
assign w17477 = w11356 & w7250;
assign w17478 = ~w10460 & ~w2881;
assign w17479 = ~w16742 & w11388;
assign w17480 = pi2698 & ~w9504;
assign w17481 = pi3170 & w3987;
assign w17482 = (pi0651 & ~w13509) | (pi0651 & w9104) | (~w13509 & w9104);
assign w17483 = (pi0985 & ~w13509) | (pi0985 & w15486) | (~w13509 & w15486);
assign w17484 = ~w5904 & ~w7660;
assign w17485 = w5517 & w13272;
assign w17486 = ~w2725 & pi0801;
assign w17487 = ~pi3135 & w3982;
assign w17488 = ~w4767 & ~w7175;
assign w17489 = ~w12450 & ~w6520;
assign w17490 = w3381 & w10724;
assign w17491 = ~w3773 & ~w11076;
assign w17492 = w15271 & w614;
assign w17493 = ~w6055 & ~w5538;
assign w17494 = ~pi3315 & w14918;
assign w17495 = ~pi1298 & ~pi1270;
assign w17496 = pi1941 & ~w17646;
assign w17497 = ~w8150 & ~w14328;
assign w17498 = ~pi3145 & w17669;
assign w17499 = pi2392 & ~w4508;
assign w17500 = w16506 & ~w2741;
assign w17501 = ~w680 & ~w2899;
assign w17502 = ~w709 & pi1283;
assign w17503 = pi1425 & ~w13753;
assign w17504 = ~w3048 & ~w10727;
assign w17505 = ~w12256 & ~w244;
assign w17506 = ~w9171 & ~w5059;
assign w17507 = ~pi0649 & w3791;
assign w17508 = ~w12460 & w6825;
assign w17509 = ~pi3047 & w3555;
assign w17510 = ~w4916 & ~w13440;
assign w17511 = ~w14334 & w2069;
assign w17512 = w12040 & ~w10947;
assign w17513 = ~w776 & ~w10227;
assign w17514 = ~w10722 & ~w11690;
assign w17515 = pi1925 & ~w15271;
assign w17516 = w17941 & w9361;
assign w17517 = w2742 & ~w16034;
assign w17518 = ~w10675 & ~w1577;
assign w17519 = ~w13294 & ~w3285;
assign w17520 = ~pi3153 & pi3207;
assign w17521 = ~w8911 & ~w15999;
assign w17522 = pi2748 & ~w261;
assign w17523 = ~w12609 & ~w8269;
assign w17524 = ~w7672 & w2346;
assign w17525 = ~pi2279 & w12941;
assign w17526 = w2725 & ~w17210;
assign w17527 = pi2649 & ~w3555;
assign w17528 = ~w2943 & w6132;
assign w17529 = ~pi0722 & w17899;
assign w17530 = pi3132 & w15767;
assign w17531 = w1962 & ~w2587;
assign w17532 = w17248 & ~w3430;
assign w17533 = ~w13616 & ~w6541;
assign w17534 = w6188 & w8642;
assign w17535 = w13509 & w3523;
assign w17536 = w5533 & w4116;
assign w17537 = pi0082 & pi1811;
assign w17538 = pi2736 & ~w5274;
assign w17539 = pi1937 & ~w18123;
assign w17540 = pi2564 & w384;
assign w17541 = ~w5430 & ~w14820;
assign w17542 = ~w1374 & ~w1185;
assign w17543 = ~w12376 & w1059;
assign w17544 = ~w16311 & ~w7401;
assign w17545 = pi2995 & pi1352;
assign w17546 = w3203 & ~w7449;
assign w17547 = ~w12070 & ~w1899;
assign w17548 = ~pi3159 & w12427;
assign w17549 = ~pi0745 & w17490;
assign w17550 = ~w1320 & w6001;
assign w17551 = w2341 & ~w6033;
assign w17552 = w384 & w3122;
assign w17553 = w1766 & w922;
assign w17554 = ~w1534 & ~w2486;
assign w17555 = ~pi0988 & ~pi1210;
assign w17556 = ~pi3166 & w17387;
assign w17557 = ~w2197 & ~w4757;
assign w17558 = pi2471 & ~w14524;
assign w17559 = w16650 & w1929;
assign w17560 = ~w18348 & w7365;
assign w17561 = pi1979 & ~w226;
assign w17562 = pi2920 & pi2966;
assign w17563 = pi2067 & ~w4508;
assign w17564 = w12040 & ~w12800;
assign w17565 = ~pi1777 & ~pi3134;
assign w17566 = pi1897 & ~w15036;
assign w17567 = ~w6697 & pi1109;
assign w17568 = w14524 & w17115;
assign w17569 = ~pi3138 & w12427;
assign w17570 = ~w7077 & pi0806;
assign w17571 = ~pi3139 & w1843;
assign w17572 = ~w6344 & ~w13905;
assign w17573 = ~w9574 & ~w10411;
assign w17574 = w13509 & w16835;
assign w17575 = ~pi3430 & w15036;
assign w17576 = ~pi0709 & w3106;
assign w17577 = ~w6195 & w15456;
assign w17578 = (pi1082 & ~w13509) | (pi1082 & w8838) | (~w13509 & w8838);
assign w17579 = ~w17429 & ~w12352;
assign w17580 = pi3031 & ~pi3154;
assign w17581 = ~w10057 & ~w14845;
assign w17582 = ~w2569 & ~w536;
assign w17583 = w12838 & w3519;
assign w17584 = ~w12603 & w3421;
assign w17585 = w13509 & w9184;
assign w17586 = w1913 & w609;
assign w17587 = ~pi0739 & w17899;
assign w17588 = ~w14886 & ~w10505;
assign w17589 = ~w12804 & ~w16573;
assign w17590 = ~w13210 & ~w12559;
assign w17591 = w735 & pi3178;
assign w17592 = ~w4945 & ~w4405;
assign w17593 = pi1718 & ~pi3171;
assign w17594 = pi1620 & ~w7090;
assign w17595 = pi0014 & ~w3748;
assign w17596 = ~w5560 & w3905;
assign w17597 = w2350 & w8896;
assign w17598 = ~w9342 & ~w16654;
assign w17599 = ~pi3142 & w11701;
assign w17600 = ~w3270 & ~w17249;
assign w17601 = pi2861 & w14148;
assign w17602 = pi2195 & ~w10299;
assign w17603 = pi0207 & w9021;
assign w17604 = pi2281 & ~w11671;
assign w17605 = ~w14654 & ~w862;
assign w17606 = w16506 & ~w14143;
assign w17607 = w13509 & w1318;
assign w17608 = ~w3350 & ~w4089;
assign w17609 = ~w7607 & ~w2277;
assign w17610 = w4946 & w14137;
assign w17611 = pi1165 & ~pi3216;
assign w17612 = w6857 & w16514;
assign w17613 = ~w857 & ~w12856;
assign w17614 = ~w16092 & ~w2314;
assign w17615 = (w13367 & ~w10745) | (w13367 & ~w17577) | (~w10745 & ~w17577);
assign w17616 = ~w5122 & w14914;
assign w17617 = ~pi2250 & w3019;
assign w17618 = w8730 & w2683;
assign w17619 = w625 & w1637;
assign w17620 = ~pi3153 & w17993;
assign w17621 = pi0034 & ~w3748;
assign w17622 = ~w5827 & w2666;
assign w17623 = (pi1874 & w2014) | (pi1874 & w11067) | (w2014 & w11067);
assign w17624 = w10647 & ~w7470;
assign w17625 = ~pi3092 & w11406;
assign w17626 = w10473 & w6984;
assign w17627 = w10189 & ~pi0450;
assign w17628 = w14560 & pi0376;
assign w17629 = pi0332 & ~pi1337;
assign w17630 = pi2204 & ~w3223;
assign w17631 = pi2838 & w15191;
assign w17632 = w7536 & w5841;
assign w17633 = ~w2014 & w4446;
assign w17634 = w17562 & pi2567;
assign w17635 = ~w16575 & w3149;
assign w17636 = w12775 & ~pi2969;
assign w17637 = ~pi1720 & pi3172;
assign w17638 = pi2245 & ~w18123;
assign w17639 = ~w11747 & ~w8474;
assign w17640 = ~w4667 & ~w12212;
assign w17641 = pi2832 & ~w11406;
assign w17642 = ~w6785 & pi0863;
assign w17643 = ~pi0552 & w11739;
assign w17644 = pi2327 & ~w4508;
assign w17645 = ~pi3133 & w15048;
assign w17646 = w14651 & w13090;
assign w17647 = pi2935 & w6045;
assign w17648 = ~w2947 & ~w13600;
assign w17649 = ~pi2785 & w15122;
assign w17650 = ~w5037 & w12887;
assign w17651 = w539 & ~w3572;
assign w17652 = ~w15381 & ~w17104;
assign w17653 = ~pi3160 & ~pi3162;
assign w17654 = (pi1002 & ~w13509) | (pi1002 & w7950) | (~w13509 & w7950);
assign w17655 = ~pi3316 & w18259;
assign w17656 = pi1440 & ~w13753;
assign w17657 = w709 & pi1897;
assign w17658 = ~w5874 & w3770;
assign w17659 = ~w2598 & ~w9987;
assign w17660 = (pi0775 & ~w13509) | (pi0775 & w4148) | (~w13509 & w4148);
assign w17661 = w13509 & w2557;
assign w17662 = ~w6013 & w17722;
assign w17663 = w709 & pi1860;
assign w17664 = pi1723 & ~pi3150;
assign w17665 = (~pi0896 & ~w12460) | (~pi0896 & w14166) | (~w12460 & w14166);
assign w17666 = pi1229 & ~w11655;
assign w17667 = w5189 & ~w2776;
assign w17668 = pi1894 & ~w15036;
assign w17669 = ~w4020 & w14833;
assign w17670 = pi0153 & w5274;
assign w17671 = pi0055 & ~w14148;
assign w17672 = (pi0920 & ~w13509) | (pi0920 & w7165) | (~w13509 & w7165);
assign w17673 = (~pi1258 & ~w13142) | (~pi1258 & w12942) | (~w13142 & w12942);
assign w17674 = pi2181 & ~w14524;
assign w17675 = (pi0786 & ~w13509) | (pi0786 & w17451) | (~w13509 & w17451);
assign w17676 = (pi1051 & ~w13509) | (pi1051 & w1370) | (~w13509 & w1370);
assign w17677 = pi2390 & ~w17683;
assign w17678 = ~w15122 & ~pi2510;
assign w17679 = ~w12651 & ~w9674;
assign w17680 = pi1915 & ~w15271;
assign w17681 = ~pi0548 & w12825;
assign w17682 = pi3162 & w653;
assign w17683 = w7996 & w9166;
assign w17684 = ~pi2220 & w2151;
assign w17685 = w3203 & ~w13195;
assign w17686 = ~pi3098 & w3555;
assign w17687 = ~pi3335 & w6448;
assign w17688 = pi0065 & w922;
assign w17689 = ~w701 & w1152;
assign w17690 = ~w15249 & ~w16530;
assign w17691 = ~w12482 & ~w4601;
assign w17692 = w13509 & w14426;
assign w17693 = ~w14228 & pi0623;
assign w17694 = pi1569 & ~w18259;
assign w17695 = pi2356 & ~w9414;
assign w17696 = ~pi3165 & w1843;
assign w17697 = ~w14287 & ~w3473;
assign w17698 = (~w9232 & ~w5517) | (~w9232 & w1429) | (~w5517 & w1429);
assign w17699 = ~w7017 & ~w7767;
assign w17700 = w13231 & ~w2776;
assign w17701 = ~pi0729 & w17899;
assign w17702 = ~pi0610 & w12825;
assign w17703 = ~pi1093 & w6200;
assign w17704 = (pi0788 & ~w13509) | (pi0788 & w8107) | (~w13509 & w8107);
assign w17705 = pi1945 & ~w17646;
assign w17706 = ~w4838 & ~w8252;
assign w17707 = ~w114 & ~w15376;
assign w17708 = ~w6244 & ~w17238;
assign w17709 = w7853 & w7272;
assign w17710 = ~w2866 & ~w5154;
assign w17711 = ~w3188 & ~w17568;
assign w17712 = pi0038 & ~w3748;
assign w17713 = ~w3000 & ~pi2759;
assign w17714 = pi1337 & ~w3262;
assign w17715 = ~pi2976 & w3555;
assign w17716 = ~pi3047 & w16815;
assign w17717 = w14782 & w6873;
assign w17718 = w5196 & w6214;
assign w17719 = pi3029 & ~pi3151;
assign w17720 = ~w14560 & pi0242;
assign w17721 = w9720 & pi1716;
assign w17722 = w10818 & ~w14676;
assign w17723 = pi1785 & ~w15767;
assign w17724 = ~w5535 & w6579;
assign w17725 = w14109 & pi0448;
assign w17726 = ~pi2011 & w11688;
assign w17727 = pi1745 & w1924;
assign w17728 = ~w3203 & pi1084;
assign w17729 = ~w16679 & ~w11163;
assign w17730 = pi2610 & ~w261;
assign w17731 = ~w14106 & w5613;
assign w17732 = ~w6785 & pi0858;
assign w17733 = w14923 & w12805;
assign w17734 = pi1675 & ~w4058;
assign w17735 = pi2574 & ~w5274;
assign w17736 = w6785 & w11302;
assign w17737 = pi2470 & ~w10299;
assign w17738 = ~w608 & ~w10656;
assign w17739 = ~w13278 & ~w47;
assign w17740 = pi1707 & ~w2253;
assign w17741 = w12689 & w18271;
assign w17742 = ~pi3437 & w15036;
assign w17743 = ~pi2300 & w16041;
assign w17744 = w3131 & w15801;
assign w17745 = (pi1144 & ~w5437) | (pi1144 & w1984) | (~w5437 & w1984);
assign w17746 = w968 & ~pi0275;
assign w17747 = ~w12050 & ~w6900;
assign w17748 = ~w11866 & ~w17507;
assign w17749 = ~w11045 & ~w5202;
assign w17750 = ~pi2967 & pi3068;
assign w17751 = ~pi0825 & w1147;
assign w17752 = w13509 & w12582;
assign w17753 = (pi1758 & w7215) | (pi1758 & w18479) | (w7215 & w18479);
assign w17754 = w9440 & pi0149;
assign w17755 = ~w18440 & ~w5487;
assign w17756 = ~w18169 & ~w1986;
assign w17757 = w18075 & w15739;
assign w17758 = ~w10198 & ~w465;
assign w17759 = ~w1962 & pi0945;
assign w17760 = (pi0379 & w5560) | (pi0379 & w7915) | (w5560 & w7915);
assign w17761 = pi1721 & ~pi3135;
assign w17762 = pi1458 & w13753;
assign w17763 = ~w5045 & ~w12867;
assign w17764 = w15122 & ~pi2695;
assign w17765 = w5453 & pi2904;
assign w17766 = w1962 & ~w3430;
assign w17767 = pi2752 & w605;
assign w17768 = ~w14990 & ~w13434;
assign w17769 = w12460 & w13391;
assign w17770 = pi1965 & ~w3836;
assign w17771 = w10647 & ~w10398;
assign w17772 = ~w15720 & ~w3117;
assign w17773 = ~pi3171 & w17387;
assign w17774 = ~w16723 & ~w17405;
assign w17775 = w709 & pi2955;
assign w17776 = ~w5153 & ~w12393;
assign w17777 = pi1475 & w13753;
assign w17778 = ~w14979 & ~w17215;
assign w17779 = ~pi0285 & w4058;
assign w17780 = ~w15207 & ~w2083;
assign w17781 = ~w1752 & ~w3949;
assign w17782 = ~w17622 & w16576;
assign w17783 = pi0500 & ~w1648;
assign w17784 = ~w11477 & ~w12562;
assign w17785 = ~w15043 & w15625;
assign w17786 = pi3057 & w3987;
assign w17787 = w12040 & ~w7449;
assign w17788 = pi1233 & pi1234;
assign w17789 = ~w16709 & ~w2910;
assign w17790 = ~pi3091 & w15235;
assign w17791 = pi3075 & ~w16502;
assign w17792 = ~pi1001 & w12825;
assign w17793 = w11251 & w15644;
assign w17794 = pi2125 & ~w18123;
assign w17795 = pi1605 & ~w13753;
assign w17796 = ~w14484 & ~w15649;
assign w17797 = ~w8796 & ~w6830;
assign w17798 = ~pi0845 & w93;
assign w17799 = w13509 & w1133;
assign w17800 = ~w1603 & ~w9406;
assign w17801 = pi1973 & pi3227;
assign w17802 = ~w16805 & ~w15873;
assign w17803 = ~w1232 & ~w5381;
assign w17804 = pi1398 & ~w14918;
assign w17805 = ~w18428 & ~w16216;
assign w17806 = ~pi3131 & w3982;
assign w17807 = ~w13231 & pi0555;
assign w17808 = ~w13196 & ~w2807;
assign w17809 = ~w3908 & w10180;
assign w17810 = ~pi3154 & ~pi3160;
assign w17811 = ~w149 & ~w16071;
assign w17812 = w12460 & w4713;
assign w17813 = w13509 & w16193;
assign w17814 = ~w17007 & w18029;
assign w17815 = ~w1818 & w5347;
assign w17816 = pi1338 & w8928;
assign w17817 = ~pi1763 & ~pi3164;
assign w17818 = pi1543 & ~w17935;
assign w17819 = w5642 & w5396;
assign w17820 = ~w2405 & ~w16681;
assign w17821 = w13509 & w13749;
assign w17822 = pi1817 & ~w653;
assign w17823 = pi2906 & w18405;
assign w17824 = ~w70 & ~w2074;
assign w17825 = ~pi0991 & w11739;
assign w17826 = w13509 & w9433;
assign w17827 = pi1436 & ~w13753;
assign w17828 = ~w6653 & ~w11475;
assign w17829 = ~w6125 & ~w13144;
assign w17830 = ~w17665 & ~w12420;
assign w17831 = (~pi0296 & ~w6857) | (~pi0296 & w496) | (~w6857 & w496);
assign w17832 = ~w12440 & ~w7023;
assign w17833 = ~pi2114 & w12755;
assign w17834 = w3203 & w1217;
assign w17835 = (pi0838 & ~w13509) | (pi0838 & w7828) | (~w13509 & w7828);
assign w17836 = w930 & w4735;
assign w17837 = ~w12460 & w15434;
assign w17838 = ~w13425 & ~w6701;
assign w17839 = ~w80 & w5102;
assign w17840 = w11351 & w8883;
assign w17841 = ~w16399 & ~w14188;
assign w17842 = ~w9412 & ~w9426;
assign w17843 = w16575 & w11524;
assign w17844 = ~w4121 & ~w7851;
assign w17845 = ~w15869 & ~w14661;
assign w17846 = ~pi3087 & w11406;
assign w17847 = w11209 & ~w8131;
assign w17848 = w2725 & w11302;
assign w17849 = w5345 & w12637;
assign w17850 = ~pi1321 & w458;
assign w17851 = pi1322 & w458;
assign w17852 = ~w6583 & ~w4329;
assign w17853 = ~w10027 & ~w899;
assign w17854 = pi3010 & ~w3987;
assign w17855 = ~w16179 & w439;
assign w17856 = ~w2455 & ~w12119;
assign w17857 = ~pi1312 & w17555;
assign w17858 = pi0095 & w9284;
assign w17859 = pi1967 & ~w7177;
assign w17860 = w6857 & w5407;
assign w17861 = ~w15808 & pi0742;
assign w17862 = ~pi3155 & w15048;
assign w17863 = (~pi0284 & ~w6857) | (~pi0284 & w7618) | (~w6857 & w7618);
assign w17864 = pi1791 & ~w15767;
assign w17865 = ~w2014 & w15078;
assign w17866 = ~w16185 & ~w9495;
assign w17867 = pi2349 & ~w9414;
assign w17868 = w15808 & ~w3430;
assign w17869 = pi2579 & ~w5274;
assign w17870 = ~pi3101 & w6463;
assign w17871 = ~w16277 & ~w6642;
assign w17872 = ~w14622 & ~w15966;
assign w17873 = pi1533 & ~w17935;
assign w17874 = pi2981 & w4084;
assign w17875 = ~w6637 & ~w9308;
assign w17876 = ~pi1976 & w17213;
assign w17877 = ~w1450 & ~w9026;
assign w17878 = ~w2669 & ~w14277;
assign w17879 = ~w9243 & w10604;
assign w17880 = pi2129 & ~w15271;
assign w17881 = ~w6697 & pi0672;
assign w17882 = (~pi1803 & ~w7799) | (~pi1803 & w13783) | (~w7799 & w13783);
assign w17883 = pi2868 & w14148;
assign w17884 = ~w2066 & ~w14578;
assign w17885 = w708 & w12436;
assign w17886 = w15808 & w15609;
assign w17887 = ~w12545 & ~w15053;
assign w17888 = ~pi0758 & w17490;
assign w17889 = ~pi3007 & ~pi3111;
assign w17890 = ~pi3138 & w15048;
assign w17891 = (pi2980 & w15119) | (pi2980 & w3410) | (w15119 & w3410);
assign w17892 = ~w11624 & ~w9689;
assign w17893 = w12460 & w18453;
assign w17894 = ~pi3158 & w8515;
assign w17895 = (~pi0977 & ~w13509) | (~pi0977 & w18289) | (~w13509 & w18289);
assign w17896 = ~pi0862 & w15707;
assign w17897 = ~w18298 & ~w11275;
assign w17898 = (~pi1799 & ~w7799) | (~pi1799 & w5033) | (~w7799 & w5033);
assign w17899 = w10087 & ~w10724;
assign w17900 = ~w5813 & ~w9625;
assign w17901 = ~w6195 & w7626;
assign w17902 = ~pi1236 & pi1376;
assign w17903 = w1391 & w11302;
assign w17904 = ~w5439 & ~w4520;
assign w17905 = ~pi3131 & pi3136;
assign w17906 = ~w5855 & w1500;
assign w17907 = ~pi0721 & w17899;
assign w17908 = ~w8192 & ~w3040;
assign w17909 = (pi1012 & ~w13509) | (pi1012 & w17290) | (~w13509 & w17290);
assign w17910 = (~w16821 & ~w5517) | (~w16821 & w3840) | (~w5517 & w3840);
assign w17911 = ~w3054 & w9626;
assign w17912 = pi1956 & ~w14833;
assign w17913 = pi2635 & ~w9504;
assign w17914 = (w7069 & w6837) | (w7069 & w11662) | (w6837 & w11662);
assign w17915 = ~w10878 & ~w4255;
assign w17916 = ~pi3170 & w3982;
assign w17917 = ~w8470 & ~w7787;
assign w17918 = ~pi3288 & w18259;
assign w17919 = ~pi1928 & w11313;
assign w17920 = w5587 & w6451;
assign w17921 = pi1741 & w1924;
assign w17922 = pi0299 & w5274;
assign w17923 = ~pi3054 & w3555;
assign w17924 = w8087 & ~w9462;
assign w17925 = pi1624 & ~w13753;
assign w17926 = w15808 & ~w10235;
assign w17927 = w1326 & w18461;
assign w17928 = ~pi2389 & w12755;
assign w17929 = ~pi0443 & ~pi2486;
assign w17930 = ~w3197 & ~w15669;
assign w17931 = pi0029 & ~w14148;
assign w17932 = (pi0633 & ~w13509) | (pi0633 & w10119) | (~w13509 & w10119);
assign w17933 = w934 & pi0440;
assign w17934 = pi0103 & w3748;
assign w17935 = pi1371 & w11399;
assign w17936 = ~w15017 & ~w17813;
assign w17937 = ~w17125 & ~w10546;
assign w17938 = w3756 & w3984;
assign w17939 = w3203 & ~w6647;
assign w17940 = w17240 & w18368;
assign w17941 = ~w4703 & ~w3699;
assign w17942 = (pi0549 & ~w13509) | (pi0549 & w6866) | (~w13509 & w6866);
assign w17943 = w2725 & ~w305;
assign w17944 = w4747 & w3480;
assign w17945 = pi2779 & w605;
assign w17946 = (~pi0276 & ~w6857) | (~pi0276 & w11663) | (~w6857 & w11663);
assign w17947 = w6857 & w6554;
assign w17948 = ~pi3076 & pi3142;
assign w17949 = ~w16290 & ~w7083;
assign w17950 = w13509 & w6894;
assign w17951 = pi0502 & ~pi1148;
assign w17952 = ~pi1950 & w11688;
assign w17953 = ~w216 & ~w6240;
assign w17954 = ~w2166 & ~w15734;
assign w17955 = w2742 & ~w10249;
assign w17956 = ~w13603 & ~w5467;
assign w17957 = ~w6595 & ~w4509;
assign w17958 = w5437 & w3861;
assign w17959 = pi0434 & ~pi2486;
assign w17960 = w13331 & w6666;
assign w17961 = w7077 & ~w1236;
assign w17962 = ~w17487 & ~w13535;
assign w17963 = ~pi0411 & pi1346;
assign w17964 = (pi1086 & ~w13509) | (pi1086 & w8577) | (~w13509 & w8577);
assign w17965 = pi1976 & ~w15235;
assign w17966 = ~w18394 & ~w12891;
assign w17967 = (w11653 & w1951) | (w11653 & w15076) | (w1951 & w15076);
assign w17968 = ~pi0685 & w9110;
assign w17969 = ~w3202 & ~w9509;
assign w17970 = ~pi3150 & w13570;
assign w17971 = pi0041 & pi0046;
assign w17972 = w15867 & w11731;
assign w17973 = w8988 & w8431;
assign w17974 = pi1433 & ~w13753;
assign w17975 = ~w5374 & ~w11836;
assign w17976 = ~w16575 & w14175;
assign w17977 = ~w2341 & pi0835;
assign w17978 = ~w5633 & ~w9831;
assign w17979 = w10158 & w17115;
assign w17980 = pi1674 & ~w4058;
assign w17981 = ~pi3138 & pi3145;
assign w17982 = pi1823 & ~w2732;
assign w17983 = ~pi1266 & pi1311;
assign w17984 = ~w12597 & ~w14155;
assign w17985 = ~w1391 & pi0551;
assign w17986 = ~w13250 & ~w17160;
assign w17987 = pi1761 & w3689;
assign w17988 = ~w13732 & ~w2094;
assign w17989 = ~w10902 & ~w4117;
assign w17990 = ~w16939 & pi0003;
assign w17991 = ~w2245 & ~w129;
assign w17992 = pi2007 & ~w14833;
assign w17993 = ~w4020 & w4508;
assign w17994 = w14648 & ~pi2611;
assign w17995 = ~w5428 & ~w7900;
assign w17996 = ~w3054 & w17721;
assign w17997 = w11671 & w6320;
assign w17998 = ~w17891 & w10642;
assign w17999 = pi0437 & w17173;
assign w18000 = ~w1582 & ~w17174;
assign w18001 = ~w7262 & ~w16246;
assign w18002 = pi1696 & ~pi1697;
assign w18003 = ~w4412 & w10610;
assign w18004 = ~w2761 & ~w3164;
assign w18005 = w160 & w11510;
assign w18006 = (pi1185 & ~w5437) | (pi1185 & w17268) | (~w5437 & w17268);
assign w18007 = ~pi0727 & w17899;
assign w18008 = w11345 & w18102;
assign w18009 = pi2196 & ~w10299;
assign w18010 = ~pi0313 & pi3225;
assign w18011 = ~w14863 & ~w6818;
assign w18012 = ~pi1762 & ~w18345;
assign w18013 = ~pi3337 & w6072;
assign w18014 = w13509 & w12026;
assign w18015 = ~w15467 & w8665;
assign w18016 = pi3138 & ~pi3145;
assign w18017 = ~w10351 & w17914;
assign w18018 = w13509 & w1477;
assign w18019 = ~w7992 & ~w6668;
assign w18020 = pi1366 & ~w5737;
assign w18021 = ~pi0120 & pi0126;
assign w18022 = ~w1368 & ~pi0473;
assign w18023 = ~pi3095 & w9504;
assign w18024 = ~w4337 & ~w15501;
assign w18025 = pi1738 & w1924;
assign w18026 = ~w12723 & ~w3424;
assign w18027 = ~w8573 & ~w15062;
assign w18028 = pi1659 & ~w6072;
assign w18029 = ~w17665 & ~w18574;
assign w18030 = w14109 & pi0420;
assign w18031 = ~w13725 & ~w4215;
assign w18032 = ~pi3340 & w6072;
assign w18033 = (~pi2920 & ~w2971) | (~pi2920 & w7493) | (~w2971 & w7493);
assign w18034 = ~w5560 & w8272;
assign w18035 = (~pi0959 & ~w13509) | (~pi0959 & w6100) | (~w13509 & w6100);
assign w18036 = ~pi1706 & w17562;
assign w18037 = (pi0717 & ~w13509) | (pi0717 & w2696) | (~w13509 & w2696);
assign w18038 = ~w405 & ~w12664;
assign w18039 = ~w18263 & ~w5335;
assign w18040 = pi1508 & ~w16922;
assign w18041 = ~pi2926 & w13343;
assign w18042 = ~pi3162 & w11132;
assign w18043 = w7533 & w6618;
assign w18044 = (pi1136 & ~w5437) | (pi1136 & w11047) | (~w5437 & w11047);
assign w18045 = pi2008 & ~w14833;
assign w18046 = ~w13924 & ~w2535;
assign w18047 = pi2996 & ~pi2997;
assign w18048 = pi1800 & pi3146;
assign w18049 = ~w8087 & w5411;
assign w18050 = w7703 & w133;
assign w18051 = w5437 & w5277;
assign w18052 = ~w8604 & ~w10733;
assign w18053 = ~w15890 & w1135;
assign w18054 = w13509 & w6281;
assign w18055 = ~pi3058 & w261;
assign w18056 = ~w12125 & ~w11178;
assign w18057 = ~w16580 & ~w2889;
assign w18058 = w13509 & w12555;
assign w18059 = w9440 & pi0193;
assign w18060 = ~w4185 & ~w6271;
assign w18061 = w10647 & ~w2120;
assign w18062 = pi1494 & ~w9781;
assign w18063 = w14366 & w1479;
assign w18064 = ~pi0757 & w17490;
assign w18065 = w10518 & w15893;
assign w18066 = pi3142 & w3987;
assign w18067 = w11383 & w9546;
assign w18068 = ~pi0699 & w3106;
assign w18069 = w6697 & ~w6033;
assign w18070 = ~w18590 & ~w10838;
assign w18071 = (w8562 & w16692) | (w8562 & w13721) | (w16692 & w13721);
assign w18072 = ~w1870 & ~w11869;
assign w18073 = ~w26 & w8614;
assign w18074 = ~w3626 & ~w7477;
assign w18075 = w16656 & w7053;
assign w18076 = ~w5484 & ~w10684;
assign w18077 = pi1360 & pi1793;
assign w18078 = pi3160 & ~pi3492;
assign w18079 = ~pi0285 & w2196;
assign w18080 = w5437 & w14710;
assign w18081 = ~pi2907 & ~w8304;
assign w18082 = pi1558 & ~w13753;
assign w18083 = (pi0560 & ~w13509) | (pi0560 & w12903) | (~w13509 & w12903);
assign w18084 = w16923 & w2408;
assign w18085 = w13231 & ~w9852;
assign w18086 = ~w14835 & ~w17823;
assign w18087 = ~w15808 & pi0748;
assign w18088 = w12460 & w13715;
assign w18089 = w15808 & w11302;
assign w18090 = ~pi1831 & ~w17646;
assign w18091 = ~w1569 & ~w11801;
assign w18092 = ~w3082 & w5437;
assign w18093 = ~w4231 & ~w13768;
assign w18094 = ~w752 & w5443;
assign w18095 = w13509 & w16690;
assign w18096 = w3567 & w13443;
assign w18097 = pi1252 & ~w11655;
assign w18098 = w7758 & w13736;
assign w18099 = pi2230 & ~w11735;
assign w18100 = ~w5666 & w5444;
assign w18101 = pi2601 & ~w9504;
assign w18102 = ~pi0483 & pi3402;
assign w18103 = pi3051 & ~w16502;
assign w18104 = pi0321 & pi3225;
assign w18105 = w10189 & ~pi0480;
assign w18106 = (pi0395 & w5560) | (pi0395 & w4914) | (w5560 & w4914);
assign w18107 = w14269 & w17537;
assign w18108 = w16348 & w3219;
assign w18109 = ~pi2969 & ~pi2984;
assign w18110 = pi2689 & ~w16815;
assign w18111 = ~w11262 & ~w4790;
assign w18112 = pi1542 & ~w17935;
assign w18113 = ~w15808 & pi0918;
assign w18114 = ~w6567 & w6080;
assign w18115 = (~pi1800 & ~w7799) | (~pi1800 & w14526) | (~w7799 & w14526);
assign w18116 = ~pi1087 & w543;
assign w18117 = ~w3000 & ~pi2791;
assign w18118 = w5437 & w15034;
assign w18119 = w14116 & w15290;
assign w18120 = ~w4563 & ~w6802;
assign w18121 = ~w2692 & ~w17383;
assign w18122 = w9440 & pi0181;
assign w18123 = w14245 & w14342;
assign w18124 = (w4903 & w7382) | (w4903 & w17586) | (w7382 & w17586);
assign w18125 = ~pi1010 & w3791;
assign w18126 = pi2724 & ~w16815;
assign w18127 = ~w7186 & ~w14806;
assign w18128 = w6649 & ~w358;
assign w18129 = w17302 & w10780;
assign w18130 = ~pi2964 & ~pi3160;
assign w18131 = w13509 & w2271;
assign w18132 = ~w16736 & ~w7575;
assign w18133 = ~pi3135 & w3805;
assign w18134 = ~w17571 & ~w17630;
assign w18135 = pi2676 & ~w226;
assign w18136 = w201 & w15909;
assign w18137 = ~pi0143 & pi0198;
assign w18138 = (pi0821 & ~w13509) | (pi0821 & w10569) | (~w13509 & w10569);
assign w18139 = w14301 & w8425;
assign w18140 = ~w4210 & w1838;
assign w18141 = ~w8225 & ~w15107;
assign w18142 = pi1243 & w11655;
assign w18143 = w12460 & w11048;
assign w18144 = pi1637 & ~w13753;
assign w18145 = pi1437 & ~w6448;
assign w18146 = ~w4753 & ~w5941;
assign w18147 = ~w16506 & pi1138;
assign w18148 = pi2891 & ~w15235;
assign w18149 = w10647 & ~w14271;
assign w18150 = ~w18540 & ~w3326;
assign w18151 = ~w8919 & ~w11225;
assign w18152 = ~w3049 & ~w2618;
assign w18153 = (w3987 & w12762) | (w3987 & w8788) | (w12762 & w8788);
assign w18154 = ~pi0275 & w4058;
assign w18155 = ~pi1878 & ~pi3513;
assign w18156 = w17741 & w11723;
assign w18157 = ~w12040 & pi0678;
assign w18158 = ~pi0833 & w93;
assign w18159 = w16278 & ~w3374;
assign w18160 = pi1337 & ~pi0258;
assign w18161 = pi1337 & pi0259;
assign w18162 = w5121 & w12179;
assign w18163 = w4936 & w12915;
assign w18164 = pi1493 & ~w9781;
assign w18165 = (pi0694 & ~w13509) | (pi0694 & w7619) | (~w13509 & w7619);
assign w18166 = ~pi3159 & ~pi3160;
assign w18167 = ~w18396 & ~w7800;
assign w18168 = ~w10097 & ~w1668;
assign w18169 = pi1664 & ~w4058;
assign w18170 = ~w4362 & ~w3979;
assign w18171 = w13509 & w8682;
assign w18172 = w1962 & w11302;
assign w18173 = ~w5560 & w6427;
assign w18174 = w15448 & w12584;
assign w18175 = pi2475 & ~w18123;
assign w18176 = ~w16578 & ~w6831;
assign w18177 = ~pi0288 & w2196;
assign w18178 = ~pi0993 & w11739;
assign w18179 = pi0022 & ~w3748;
assign w18180 = pi0251 & w5113;
assign w18181 = w13509 & w11686;
assign w18182 = w13509 & w15903;
assign w18183 = ~w18107 & ~w701;
assign w18184 = w4420 & w9407;
assign w18185 = w10647 & ~w16880;
assign w18186 = ~pi1246 & w11655;
assign w18187 = pi1247 & w11655;
assign w18188 = ~w14604 & w437;
assign w18189 = ~pi2047 & w13204;
assign w18190 = ~w16697 & ~w14472;
assign w18191 = w2065 & w1956;
assign w18192 = ~w10210 & ~w11323;
assign w18193 = w2341 & ~w10947;
assign w18194 = pi1209 & ~w11010;
assign w18195 = ~w15122 & ~pi2890;
assign w18196 = ~pi0870 & w15707;
assign w18197 = pi1744 & ~w4058;
assign w18198 = pi2150 & ~w11671;
assign w18199 = pi2224 & ~w11735;
assign w18200 = ~w13620 & ~w7060;
assign w18201 = ~pi0911 & w6200;
assign w18202 = ~w7488 & ~w6312;
assign w18203 = w6785 & ~w7707;
assign w18204 = ~w2016 & ~w12882;
assign w18205 = w15122 & ~pi2163;
assign w18206 = ~w7358 & ~w12405;
assign w18207 = ~w3035 & ~w16258;
assign w18208 = pi0036 & ~w14148;
assign w18209 = ~pi1972 & w10694;
assign w18210 = w16683 & w14063;
assign w18211 = ~pi3335 & w18259;
assign w18212 = ~pi1919 & w2151;
assign w18213 = w2363 & w15842;
assign w18214 = ~w4667 & ~w920;
assign w18215 = ~w929 & ~w11346;
assign w18216 = w10189 & ~pi0461;
assign w18217 = w13231 & ~w7707;
assign w18218 = (pi0630 & ~w13509) | (pi0630 & w16247) | (~w13509 & w16247);
assign w18219 = ~pi2976 & w261;
assign w18220 = ~w13925 & ~w13962;
assign w18221 = ~w6697 & pi0657;
assign w18222 = pi3136 & w7363;
assign w18223 = ~w14165 & ~w13880;
assign w18224 = w11383 & w15179;
assign w18225 = w16278 & ~w4043;
assign w18226 = ~pi3316 & w6448;
assign w18227 = w384 & w13802;
assign w18228 = w7077 & ~w1340;
assign w18229 = ~pi3350 & w6072;
assign w18230 = ~pi1040 & w543;
assign w18231 = ~w7738 & ~w11501;
assign w18232 = pi3081 & ~pi3139;
assign w18233 = ~w4738 & ~w12775;
assign w18234 = w13509 & w17667;
assign w18235 = ~w5560 & w9387;
assign w18236 = ~pi3346 & w17935;
assign w18237 = ~w17539 & ~w18488;
assign w18238 = w5874 & w5082;
assign w18239 = ~w14760 & ~w8527;
assign w18240 = pi2778 & ~w3555;
assign w18241 = ~w136 & ~w14953;
assign w18242 = pi0070 & w922;
assign w18243 = ~pi3092 & w9504;
assign w18244 = w17544 & w9228;
assign w18245 = (pi1016 & ~w13509) | (pi1016 & w2344) | (~w13509 & w2344);
assign w18246 = ~w15662 & ~w5062;
assign w18247 = pi2190 & ~w11735;
assign w18248 = pi2383 & ~w14524;
assign w18249 = pi1522 & ~w14918;
assign w18250 = w11247 & w8356;
assign w18251 = ~w12040 & pi0693;
assign w18252 = pi3013 & ~pi3134;
assign w18253 = w13509 & w10875;
assign w18254 = w13509 & w12634;
assign w18255 = ~w2795 & ~w2305;
assign w18256 = ~w12765 & ~w6343;
assign w18257 = ~w11858 & w2681;
assign w18258 = ~w10809 & ~w16702;
assign w18259 = w6097 & w10455;
assign w18260 = ~w8363 & ~w16820;
assign w18261 = ~w10022 & ~w371;
assign w18262 = ~w3055 & w5188;
assign w18263 = (pi0705 & ~w13509) | (pi0705 & w7440) | (~w13509 & w7440);
assign w18264 = w7522 & w15745;
assign w18265 = ~pi0925 & w17899;
assign w18266 = ~w5722 & ~w4986;
assign w18267 = w5517 & w12868;
assign w18268 = ~w16317 & ~w814;
assign w18269 = ~w17354 & ~w13687;
assign w18270 = ~w2281 & ~w6222;
assign w18271 = ~pi3001 & ~pi2995;
assign w18272 = ~w4475 & w14913;
assign w18273 = pi1417 & ~w13753;
assign w18274 = ~w9787 & ~w4490;
assign w18275 = (~pi0488 & w17577) | (~pi0488 & w2978) | (w17577 & w2978);
assign w18276 = pi1683 & pi0305;
assign w18277 = ~w5480 & ~w8253;
assign w18278 = pi1505 & ~w16922;
assign w18279 = w14109 & pi0424;
assign w18280 = ~w9259 & ~w7653;
assign w18281 = w3138 & w6626;
assign w18282 = pi1916 & ~w10299;
assign w18283 = w6857 & w14062;
assign w18284 = w12040 & ~w305;
assign w18285 = w12460 & w16339;
assign w18286 = w62 & w10848;
assign w18287 = pi1354 & ~w11272;
assign w18288 = ~w10145 & ~w2590;
assign w18289 = ~w7077 & ~pi0977;
assign w18290 = w8658 & pi1788;
assign w18291 = ~pi3151 & pi3207;
assign w18292 = ~w17164 & ~w5635;
assign w18293 = ~w11948 & ~w1610;
assign w18294 = ~pi2703 & w15122;
assign w18295 = ~w16406 & ~w6304;
assign w18296 = pi2949 & ~w5675;
assign w18297 = pi1457 & ~w7090;
assign w18298 = pi1901 & ~w11406;
assign w18299 = w11209 & ~w12374;
assign w18300 = ~w12875 & ~w7417;
assign w18301 = ~w17296 & ~w12481;
assign w18302 = ~pi0676 & w12197;
assign w18303 = w7077 & ~w13028;
assign w18304 = ~w4962 & ~w11850;
assign w18305 = ~w1329 & w7760;
assign w18306 = ~w9311 & ~w3467;
assign w18307 = ~w9917 & ~w9865;
assign w18308 = w18024 & w9582;
assign w18309 = pi1574 & ~w16922;
assign w18310 = ~pi1753 & pi3138;
assign w18311 = ~pi0500 & ~pi1345;
assign w18312 = ~pi3341 & w17935;
assign w18313 = ~pi3162 & w8515;
assign w18314 = ~pi2999 & ~pi3002;
assign w18315 = w12126 & w14414;
assign w18316 = ~w141 & ~w11207;
assign w18317 = ~pi2852 & w14148;
assign w18318 = pi2853 & w14148;
assign w18319 = ~pi3315 & w16922;
assign w18320 = w17562 & pi2496;
assign w18321 = w621 & ~w11215;
assign w18322 = ~w7545 & ~w17563;
assign w18323 = ~w11195 & ~w6803;
assign w18324 = w13679 & w13344;
assign w18325 = ~pi0111 & w3748;
assign w18326 = ~w14591 & ~w14962;
assign w18327 = w15920 & w11496;
assign w18328 = ~pi2972 & pi3018;
assign w18329 = pi1553 & ~w17935;
assign w18330 = ~w17243 & w18543;
assign w18331 = ~w779 & ~w17576;
assign w18332 = w17562 & ~w10211;
assign w18333 = ~w8354 & w11202;
assign w18334 = ~w7222 & ~w859;
assign w18335 = (pi0398 & w5560) | (pi0398 & w8774) | (w5560 & w8774);
assign w18336 = w17251 & w4355;
assign w18337 = ~w17248 & pi0880;
assign w18338 = (w12633 & ~w3613) | (w12633 & w3970) | (~w3613 & w3970);
assign w18339 = pi2819 & w14148;
assign w18340 = ~pi1081 & w543;
assign w18341 = ~pi1842 & ~w412;
assign w18342 = pi1672 & w1924;
assign w18343 = ~w7345 & ~w8089;
assign w18344 = ~w11059 & w12631;
assign w18345 = pi1682 & pi1684;
assign w18346 = pi2758 & ~w14123;
assign w18347 = pi1418 & ~w6072;
assign w18348 = (~pi0497 & w17577) | (~pi0497 & w3275) | (w17577 & w3275);
assign w18349 = (pi0730 & ~w13509) | (pi0730 & w2543) | (~w13509 & w2543);
assign w18350 = w13509 & w16553;
assign w18351 = w1540 & w14217;
assign w18352 = ~w1388 & w16460;
assign w18353 = pi3150 & pi3162;
assign w18354 = ~pi2136 & w12941;
assign w18355 = pi1602 & w13753;
assign w18356 = pi3170 & w12558;
assign w18357 = pi1389 & w13753;
assign w18358 = w1127 & ~w4150;
assign w18359 = w5437 & w2329;
assign w18360 = w2725 & ~w2587;
assign w18361 = ~w709 & pi1279;
assign w18362 = pi1528 & w13753;
assign w18363 = pi2021 & ~w14833;
assign w18364 = ~pi2924 & ~w2536;
assign w18365 = ~pi0483 & pi3392;
assign w18366 = w422 & w17361;
assign w18367 = ~pi2946 & w11406;
assign w18368 = ~w2987 & w11925;
assign w18369 = ~pi1107 & w3106;
assign w18370 = w11383 & w875;
assign w18371 = ~w3317 & w5310;
assign w18372 = w14228 & ~w6647;
assign w18373 = ~w9382 & ~w27;
assign w18374 = (pi0303 & ~w325) | (pi0303 & w17171) | (~w325 & w17171);
assign w18375 = (pi1263 & ~w5437) | (pi1263 & w896) | (~w5437 & w896);
assign w18376 = ~w6538 & ~w14326;
assign w18377 = ~w3963 & ~w10230;
assign w18378 = ~w16278 & pi0704;
assign w18379 = (w758 & w3631) | (w758 & w4435) | (w3631 & w4435);
assign w18380 = w1127 & ~w18387;
assign w18381 = pi1821 & ~w2732;
assign w18382 = ~w2387 & w214;
assign w18383 = ~w3203 & pi0579;
assign w18384 = w13509 & w6585;
assign w18385 = w10818 & ~w806;
assign w18386 = pi2655 & ~w15235;
assign w18387 = pi1648 & w13753;
assign w18388 = ~w9025 & ~w13429;
assign w18389 = ~w16575 & w12620;
assign w18390 = w3243 & ~pi0321;
assign w18391 = ~pi3147 & w13570;
assign w18392 = pi2582 & ~w5274;
assign w18393 = pi0090 & w3748;
assign w18394 = (pi0869 & ~w13509) | (pi0869 & w16403) | (~w13509 & w16403);
assign w18395 = pi2583 & ~w5274;
assign w18396 = pi1775 & ~w10389;
assign w18397 = ~pi3085 & w261;
assign w18398 = ~w12975 & w4756;
assign w18399 = ~pi3150 & ~pi3162;
assign w18400 = (~pi0981 & ~w13509) | (~pi0981 & w12931) | (~w13509 & w12931);
assign w18401 = ~w13235 & ~w13223;
assign w18402 = ~w4607 & ~w1808;
assign w18403 = ~pi1696 & pi1697;
assign w18404 = ~pi2978 & ~w9545;
assign w18405 = ~pi2593 & w8304;
assign w18406 = w15064 & w10473;
assign w18407 = w7703 & w16162;
assign w18408 = ~w6195 & w4461;
assign w18409 = pi3509 & w13367;
assign w18410 = ~pi0693 & w9110;
assign w18411 = ~w13370 & ~w6212;
assign w18412 = ~w6961 & ~w479;
assign w18413 = pi2122 & ~w412;
assign w18414 = ~w1791 & w5954;
assign w18415 = ~pi0864 & w15707;
assign w18416 = pi1432 & ~w13753;
assign w18417 = w7703 & w10128;
assign w18418 = pi2565 & ~w5274;
assign w18419 = ~w6697 & pi0669;
assign w18420 = w8230 & w12505;
assign w18421 = (pi0698 & ~w13509) | (pi0698 & w11400) | (~w13509 & w11400);
assign w18422 = ~pi1268 & w4880;
assign w18423 = (pi0695 & ~w13509) | (pi0695 & w15686) | (~w13509 & w15686);
assign w18424 = ~pi3150 & w17993;
assign w18425 = ~w14637 & w12178;
assign w18426 = ~pi2070 & w8617;
assign w18427 = ~pi2097 & w12724;
assign w18428 = pi2432 & ~w226;
assign w18429 = w12460 & w14052;
assign w18430 = ~w2080 & w3931;
assign w18431 = ~w12073 & ~w14408;
assign w18432 = pi2362 & ~w412;
assign w18433 = w17840 & w635;
assign w18434 = w8337 & pi3301;
assign w18435 = ~pi3516 & w12206;
assign w18436 = ~w12475 & w10222;
assign w18437 = (w5855 & w17629) | (w5855 & w8655) | (w17629 & w8655);
assign w18438 = pi0304 & w5274;
assign w18439 = ~pi3060 & w226;
assign w18440 = pi1539 & ~w17935;
assign w18441 = pi2529 & w14148;
assign w18442 = ~pi2975 & w11735;
assign w18443 = ~w3224 & ~w1727;
assign w18444 = pi2027 & ~w17646;
assign w18445 = ~w3597 & ~w4732;
assign w18446 = ~w18523 & ~w1198;
assign w18447 = (pi1230 & ~w5437) | (pi1230 & w11331) | (~w5437 & w11331);
assign w18448 = ~pi3431 & w15036;
assign w18449 = ~w6348 & ~w6716;
assign w18450 = ~w3158 & ~w10906;
assign w18451 = pi1640 & ~w6448;
assign w18452 = w10189 & pi0405;
assign w18453 = w9440 & pi0154;
assign w18454 = w9323 & w12678;
assign w18455 = ~w9683 & ~w9971;
assign w18456 = (pi0631 & ~w13509) | (pi0631 & w14180) | (~w13509 & w14180);
assign w18457 = ~w1962 & pi0639;
assign w18458 = ~w1391 & pi0914;
assign w18459 = pi1596 & ~w16922;
assign w18460 = w16278 & ~w13195;
assign w18461 = ~w8571 & ~w18314;
assign w18462 = pi1421 & ~w13753;
assign w18463 = w13431 & w4700;
assign w18464 = w7656 & ~pi1180;
assign w18465 = (pi0573 & ~w13509) | (pi0573 & w15814) | (~w13509 & w15814);
assign w18466 = ~w1791 & w207;
assign w18467 = pi1356 & ~w13786;
assign w18468 = ~w821 & w15441;
assign w18469 = ~w238 & w11028;
assign w18470 = ~w7077 & pi0804;
assign w18471 = w12040 & ~w17513;
assign w18472 = ~pi2972 & pi3207;
assign w18473 = ~pi3170 & w15048;
assign w18474 = w12040 & w1217;
assign w18475 = ~pi2823 & w17213;
assign w18476 = ~w14503 & w5274;
assign w18477 = ~w16825 & ~w2707;
assign w18478 = ~pi0278 & w4058;
assign w18479 = w8658 & pi1758;
assign w18480 = ~pi3087 & w15235;
assign w18481 = pi2940 & ~pi3208;
assign w18482 = ~pi0486 & ~pi1345;
assign w18483 = ~w16760 & ~w495;
assign w18484 = w7703 & w11824;
assign w18485 = ~pi3089 & w6463;
assign w18486 = w384 & w8556;
assign w18487 = ~pi2452 & w9340;
assign w18488 = ~pi3154 & w14753;
assign w18489 = w13509 & w10307;
assign w18490 = (pi1179 & ~w773) | (pi1179 & ~w14073) | (~w773 & ~w14073);
assign w18491 = w1962 & ~w14978;
assign w18492 = (pi0676 & ~w13509) | (pi0676 & w11709) | (~w13509 & w11709);
assign w18493 = ~w12460 & w15958;
assign w18494 = w1962 & ~w11978;
assign w18495 = (pi0796 & ~w13509) | (pi0796 & w2256) | (~w13509 & w2256);
assign w18496 = w7077 & ~w11978;
assign w18497 = w4683 & w4304;
assign w18498 = w13509 & w5821;
assign w18499 = (pi0645 & ~w13509) | (pi0645 & w4393) | (~w13509 & w4393);
assign w18500 = ~w5943 & ~w17256;
assign w18501 = w137 & w1278;
assign w18502 = ~w5083 & ~w15892;
assign w18503 = ~pi1796 & w11388;
assign w18504 = ~w12561 & ~w7456;
assign w18505 = ~pi3153 & w14753;
assign w18506 = ~w14968 & w2036;
assign w18507 = pi0325 & w5113;
assign w18508 = w7766 & w1817;
assign w18509 = w17786 & w16662;
assign w18510 = pi2866 & w14148;
assign w18511 = ~w709 & pi1293;
assign w18512 = w5104 & w4656;
assign w18513 = ~w14707 & ~w17267;
assign w18514 = ~w9856 & ~w8043;
assign w18515 = ~pi0293 & w2196;
assign w18516 = pi1333 & pi2966;
assign w18517 = w10189 & pi0394;
assign w18518 = (w15842 & ~w384) | (w15842 & w10520) | (~w384 & w10520);
assign w18519 = ~pi1118 & w3791;
assign w18520 = (~w16725 & ~w15717) | (~w16725 & w17289) | (~w15717 & w17289);
assign w18521 = ~w11513 & ~w838;
assign w18522 = ~w12040 & pi0685;
assign w18523 = pi1733 & ~w4058;
assign w18524 = ~pi0315 & pi3235;
assign w18525 = w14109 & pi0428;
assign w18526 = w62 & w7926;
assign w18527 = w14105 & pi1318;
assign w18528 = ~w6747 & ~w457;
assign w18529 = w6697 & ~w3374;
assign w18530 = w10206 & w6117;
assign w18531 = w15122 & ~pi2634;
assign w18532 = w14269 & ~w9516;
assign w18533 = pi2059 & ~w4508;
assign w18534 = ~pi3162 & w17993;
assign w18535 = ~pi1345 & ~pi2941;
assign w18536 = ~w17599 & ~w6943;
assign w18537 = ~w3203 & pi0589;
assign w18538 = (w8541 & w17577) | (w8541 & w2992) | (w17577 & w2992);
assign w18539 = ~w17248 & pi0889;
assign w18540 = pi2437 & ~w3223;
assign w18541 = ~pi0954 & w795;
assign w18542 = pi1499 & ~w13753;
assign w18543 = ~w6378 & ~w7505;
assign w18544 = pi2785 & ~w3555;
assign w18545 = ~pi1116 & w3791;
assign w18546 = (~w8629 & ~w1007) | (~w8629 & w17244) | (~w1007 & w17244);
assign w18547 = ~pi1722 & pi3133;
assign w18548 = ~pi1930 & w2151;
assign w18549 = w539 & ~w10824;
assign w18550 = ~w13914 & ~w2966;
assign w18551 = pi2543 & w14148;
assign w18552 = ~pi3160 & ~pi3163;
assign w18553 = w15842 & w10676;
assign w18554 = pi1591 & ~w16922;
assign w18555 = ~w13475 & ~w11159;
assign w18556 = (pi0671 & ~w13509) | (pi0671 & w4791) | (~w13509 & w4791);
assign w18557 = (~pi0061 & ~w17103) | (~pi0061 & w13242) | (~w17103 & w13242);
assign w18558 = w6675 & w1529;
assign w18559 = pi1220 & ~pi3120;
assign w18560 = ~w6933 & ~w1885;
assign w18561 = (~w13367 & w17577) | (~w13367 & w10595) | (w17577 & w10595);
assign w18562 = ~w161 & ~w15468;
assign w18563 = ~pi1878 & ~pi3511;
assign w18564 = ~w15122 & ~pi2674;
assign w18565 = pi3136 & w11608;
assign w18566 = pi1482 & ~w9781;
assign w18567 = pi2847 & w605;
assign w18568 = ~w18423 & ~w7746;
assign w18569 = (~pi0255 & ~w325) | (~pi0255 & w1523) | (~w325 & w1523);
assign w18570 = ~pi1125 & w1126;
assign w18571 = w3203 & ~w2741;
assign w18572 = ~w10644 & ~w13847;
assign w18573 = ~w9532 & w11068;
assign w18574 = ~w12460 & w2108;
assign w18575 = w5437 & w5290;
assign w18576 = ~w14560 & pi0237;
assign w18577 = ~pi0738 & w17899;
assign w18578 = ~pi0561 & w11739;
assign w18579 = ~w15923 & ~w7757;
assign w18580 = w7348 & w3641;
assign w18581 = pi3072 & ~pi3171;
assign w18582 = ~w13073 & w14819;
assign w18583 = ~pi1676 & pi1698;
assign w18584 = ~w9961 & ~w7903;
assign w18585 = pi1410 & ~pi3240;
assign w18586 = ~pi0425 & w1599;
assign w18587 = pi0436 & ~pi2486;
assign w18588 = w934 & pi0415;
assign w18589 = pi1545 & ~w17935;
assign w18590 = pi3067 & ~w16502;
assign w18591 = w7807 & w15327;
assign w18592 = ~w7078 & ~w1222;
assign w18593 = (pi0989 & ~w13509) | (pi0989 & w8871) | (~w13509 & w8871);
assign w18594 = w7688 & w3111;
assign w18595 = ~w17435 & ~w4942;
assign w18596 = ~pi3135 & w17993;
assign w18597 = pi0274 & ~pi1337;
assign w18598 = pi0263 & w5274;
assign w18599 = w11383 & w13502;
assign w18600 = ~w14846 & ~w7292;
assign w18601 = pi1693 & w293;
assign w18602 = ~w1619 & ~w6355;
assign one = 1;
assign po0000 = ~w8579;// level 1
assign po0001 = pi0988;// level 0
assign po0002 = pi1312;// level 0
assign po0003 = pi1210;// level 0
assign po0004 = ~pi0339;// level 0
assign po0005 = pi0340;// level 0
assign po0006 = pi0336;// level 0
assign po0007 = one;// level 0
assign po0008 = pi2964;// level 0
assign po0009 = pi3127;// level 0
assign po0010 = pi3183;// level 0
assign po0011 = pi1259;// level 0
assign po0012 = pi1859;// level 0
assign po0013 = pi3195;// level 0
assign po0014 = pi1227;// level 0
assign po0015 = pi1225;// level 0
assign po0016 = pi1226;// level 0
assign po0017 = pi3119;// level 0
assign po0018 = pi0127;// level 0
assign po0019 = pi0121;// level 0
assign po0020 = pi0125;// level 0
assign po0021 = pi1347;// level 0
assign po0022 = pi0445;// level 0
assign po0023 = pi0219;// level 0
assign po0024 = pi0132;// level 0
assign po0025 = pi0221;// level 0
assign po0026 = pi0220;// level 0
assign po0027 = pi0231;// level 0
assign po0028 = pi0213;// level 0
assign po0029 = pi0229;// level 0
assign po0030 = pi0242;// level 0
assign po0031 = pi0243;// level 0
assign po0032 = pi0217;// level 0
assign po0033 = pi0218;// level 0
assign po0034 = pi0244;// level 0
assign po0035 = pi0245;// level 0
assign po0036 = pi0246;// level 0
assign po0037 = pi0208;// level 0
assign po0038 = pi0209;// level 0
assign po0039 = pi0232;// level 0
assign po0040 = pi0233;// level 0
assign po0041 = pi0234;// level 0
assign po0042 = pi0225;// level 0
assign po0043 = pi0210;// level 0
assign po0044 = pi0235;// level 0
assign po0045 = pi0211;// level 0
assign po0046 = pi0212;// level 0
assign po0047 = pi0236;// level 0
assign po0048 = pi0214;// level 0
assign po0049 = pi0215;// level 0
assign po0050 = pi0237;// level 0
assign po0051 = pi0226;// level 0
assign po0052 = pi0227;// level 0
assign po0053 = pi0238;// level 0
assign po0054 = pi0228;// level 0
assign po0055 = pi0239;// level 0
assign po0056 = pi0240;// level 0
assign po0057 = pi0216;// level 0
assign po0058 = pi0241;// level 0
assign po0059 = pi0069;// level 0
assign po0060 = pi0070;// level 0
assign po0061 = pi0065;// level 0
assign po0062 = pi0059;// level 0
assign po0063 = pi0060;// level 0
assign po0064 = pi0061;// level 0
assign po0065 = pi0062;// level 0
assign po0066 = pi0068;// level 0
assign po0067 = pi0063;// level 0
assign po0068 = pi0064;// level 0
assign po0069 = pi0051;// level 0
assign po0070 = pi0052;// level 0
assign po0071 = pi0053;// level 0
assign po0072 = pi0056;// level 0
assign po0073 = pi0055;// level 0
assign po0074 = pi0067;// level 0
assign po0075 = pi0054;// level 0
assign po0076 = pi0050;// level 0
assign po0077 = pi0066;// level 0
assign po0078 = pi0039;// level 0
assign po0079 = pi0042;// level 0
assign po0080 = pi0044;// level 0
assign po0081 = pi0040;// level 0
assign po0082 = pi0057;// level 0
assign po0083 = pi0041;// level 0
assign po0084 = pi0046;// level 0
assign po0085 = pi0058;// level 0
assign po0086 = pi0043;// level 0
assign po0087 = pi0047;// level 0
assign po0088 = pi0049;// level 0
assign po0089 = pi0045;// level 0
assign po0090 = pi0048;// level 0
assign po0091 = pi0007;// level 0
assign po0092 = pi0015;// level 0
assign po0093 = pi0026;// level 0
assign po0094 = pi0028;// level 0
assign po0095 = pi0029;// level 0
assign po0096 = pi0030;// level 0
assign po0097 = pi0031;// level 0
assign po0098 = pi0037;// level 0
assign po0099 = pi0032;// level 0
assign po0100 = pi0033;// level 0
assign po0101 = pi0008;// level 0
assign po0102 = pi0009;// level 0
assign po0103 = pi0010;// level 0
assign po0104 = pi0011;// level 0
assign po0105 = pi0035;// level 0
assign po0106 = pi0038;// level 0
assign po0107 = pi0012;// level 0
assign po0108 = pi0013;// level 0
assign po0109 = pi0036;// level 0
assign po0110 = pi0014;// level 0
assign po0111 = pi0016;// level 0
assign po0112 = pi0017;// level 0
assign po0113 = pi0018;// level 0
assign po0114 = pi0019;// level 0
assign po0115 = pi0020;// level 0
assign po0116 = pi0021;// level 0
assign po0117 = pi0022;// level 0
assign po0118 = pi0023;// level 0
assign po0119 = pi0024;// level 0
assign po0120 = pi0025;// level 0
assign po0121 = pi0034;// level 0
assign po0122 = pi0027;// level 0
assign po0123 = pi0930;// level 0
assign po0124 = pi0536;// level 0
assign po0125 = pi0537;// level 0
assign po0126 = pi0534;// level 0
assign po0127 = pi0535;// level 0
assign po0128 = pi0533;// level 0
assign po0129 = pi0931;// level 0
assign po0130 = pi0531;// level 0
assign po0131 = pi0530;// level 0
assign po0132 = pi0532;// level 0
assign po0133 = pi0934;// level 0
assign po0134 = pi0528;// level 0
assign po0135 = pi0933;// level 0
assign po0136 = pi0527;// level 0
assign po0137 = pi0526;// level 0
assign po0138 = pi0525;// level 0
assign po0139 = pi0935;// level 0
assign po0140 = pi0523;// level 0
assign po0141 = pi0524;// level 0
assign po0142 = pi0522;// level 0
assign po0143 = pi0938;// level 0
assign po0144 = pi0521;// level 0
assign po0145 = pi0520;// level 0
assign po0146 = pi0519;// level 0
assign po0147 = pi0939;// level 0
assign po0148 = pi0529;// level 0
assign po0149 = pi0538;// level 0
assign po0150 = pi0542;// level 0
assign po0151 = pi0541;// level 0
assign po0152 = pi0540;// level 0
assign po0153 = pi0928;// level 0
assign po0154 = pi0539;// level 0
assign po0155 = pi0200;// level 0
assign po0156 = pi0193;// level 0
assign po0157 = pi0163;// level 0
assign po0158 = pi0170;// level 0
assign po0159 = pi0164;// level 0
assign po0160 = pi0165;// level 0
assign po0161 = pi0166;// level 0
assign po0162 = pi0167;// level 0
assign po0163 = pi0169;// level 0
assign po0164 = pi0188;// level 0
assign po0165 = pi0180;// level 0
assign po0166 = pi0154;// level 0
assign po0167 = pi0155;// level 0
assign po0168 = pi0156;// level 0
assign po0169 = pi0157;// level 0
assign po0170 = pi0158;// level 0
assign po0171 = pi0181;// level 0
assign po0172 = pi0182;// level 0
assign po0173 = pi0183;// level 0
assign po0174 = pi0184;// level 0
assign po0175 = pi0186;// level 0
assign po0176 = pi0196;// level 0
assign po0177 = pi0185;// level 0
assign po0178 = pi0168;// level 0
assign po0179 = pi0159;// level 0
assign po0180 = pi0204;// level 0
assign po0181 = pi0199;// level 0
assign po0182 = pi0160;// level 0
assign po0183 = pi0162;// level 0
assign po0184 = pi0161;// level 0
assign po0185 = pi0194;// level 0
assign po0186 = pi0131;// level 0
assign po0187 = pi0003;// level 0
assign po0188 = pi0004;// level 0
assign po0189 = pi0005;// level 0
assign po0190 = pi0006;// level 0
assign po0191 = pi2405;// level 0
assign po0192 = pi2404;// level 0
assign po0193 = pi1982;// level 0
assign po0194 = pi1981;// level 0
assign po0195 = pi0137;// level 0
assign po0196 = pi1343;// level 0
assign po0197 = pi0138;// level 0
assign po0198 = pi0140;// level 0
assign po0199 = pi0000;// level 0
assign po0200 = pi0080;// level 0
assign po0201 = pi0001;// level 0
assign po0202 = pi3368;// level 0
assign po0203 = one;// level 0
assign po0204 = pi3359;// level 0
assign po0205 = ~w9147;// level 11
assign po0206 = ~w3008;// level 11
assign po0207 = pi3367;// level 0
assign po0208 = ~w3618;// level 6
assign po0209 = ~w7497;// level 11
assign po0210 = ~w6503;// level 11
assign po0211 = ~w737;// level 11
assign po0212 = ~w17028;// level 11
assign po0213 = ~w1383;// level 11
assign po0214 = ~w10928;// level 11
assign po0215 = ~w8492;// level 11
assign po0216 = ~w2131;// level 11
assign po0217 = ~w13297;// level 11
assign po0218 = ~w12287;// level 11
assign po0219 = ~w3213;// level 11
assign po0220 = ~w8454;// level 11
assign po0221 = ~w12728;// level 11
assign po0222 = ~w7711;// level 11
assign po0223 = ~w11340;// level 11
assign po0224 = ~w1279;// level 11
assign po0225 = ~w11835;// level 11
assign po0226 = ~w14501;// level 11
assign po0227 = ~w10509;// level 11
assign po0228 = ~w14255;// level 11
assign po0229 = ~w12496;// level 11
assign po0230 = ~w5438;// level 11
assign po0231 = ~w8641;// level 11
assign po0232 = ~w290;// level 11
assign po0233 = ~w5400;// level 11
assign po0234 = ~w10507;// level 11
assign po0235 = ~w5420;// level 11
assign po0236 = ~w10111;// level 11
assign po0237 = ~w18027;// level 11
assign po0238 = ~w10966;// level 11
assign po0239 = ~w3922;// level 11
assign po0240 = ~w15825;// level 11
assign po0241 = ~w2625;// level 11
assign po0242 = ~w6218;// level 11
assign po0243 = ~w18304;// level 11
assign po0244 = ~w3240;// level 11
assign po0245 = w16053;// level 10
assign po0246 = w9213;// level 10
assign po0247 = w10521;// level 10
assign po0248 = w757;// level 9
assign po0249 = w10915;// level 10
assign po0250 = w13700;// level 10
assign po0251 = ~w8794;// level 10
assign po0252 = ~w9533;// level 9
assign po0253 = w9713;// level 10
assign po0254 = ~w12791;// level 9
assign po0255 = w4925;// level 9
assign po0256 = w14882;// level 10
assign po0257 = ~w2904;// level 8
assign po0258 = w16243;// level 10
assign po0259 = w808;// level 10
assign po0260 = w17785;// level 9
assign po0261 = w3718;// level 10
assign po0262 = w8580;// level 10
assign po0263 = ~w6754;// level 10
assign po0264 = w2022;// level 10
assign po0265 = w15281;// level 8
assign po0266 = w6557;// level 9
assign po0267 = w9646;// level 8
assign po0268 = w11027;// level 9
assign po0269 = w12138;// level 9
assign po0270 = w9321;// level 8
assign po0271 = w17294;// level 9
assign po0272 = w6339;// level 9
assign po0273 = w3918;// level 9
assign po0274 = w13624;// level 8
assign po0275 = ~w14989;// level 9
assign po0276 = ~w2268;// level 9
assign po0277 = w12064;// level 3
assign po0278 = ~w16735;// level 8
assign po0279 = ~w5946;// level 8
assign po0280 = ~w8836;// level 8
assign po0281 = ~w4424;// level 8
assign po0282 = w12957;// level 4
assign po0283 = w16469;// level 12
assign po0284 = w9700;// level 9
assign po0285 = ~w12344;// level 9
assign po0286 = ~w12173;// level 11
assign po0287 = w1330;// level 9
assign po0288 = ~w3579;// level 9
assign po0289 = ~w12655;// level 15
assign po0290 = ~w3199;// level 15
assign po0291 = ~w924;// level 15
assign po0292 = ~w14475;// level 15
assign po0293 = ~w15344;// level 15
assign po0294 = ~w16593;// level 15
assign po0295 = ~w10429;// level 15
assign po0296 = ~w2214;// level 15
assign po0297 = ~w7253;// level 15
assign po0298 = ~w1045;// level 15
assign po0299 = ~w7476;// level 15
assign po0300 = ~w12688;// level 15
assign po0301 = ~w9719;// level 15
assign po0302 = ~w9730;// level 15
assign po0303 = ~w6869;// level 15
assign po0304 = ~w9681;// level 15
assign po0305 = ~w12296;// level 15
assign po0306 = ~w12822;// level 15
assign po0307 = ~w7127;// level 15
assign po0308 = ~w17269;// level 15
assign po0309 = ~w15619;// level 15
assign po0310 = ~w9292;// level 15
assign po0311 = ~w8528;// level 15
assign po0312 = ~w8561;// level 15
assign po0313 = ~w10253;// level 15
assign po0314 = ~w6687;// level 15
assign po0315 = ~w10061;// level 15
assign po0316 = ~w5803;// level 15
assign po0317 = ~w17733;// level 15
assign po0318 = ~w5979;// level 15
assign po0319 = ~w1029;// level 15
assign po0320 = ~w5116;// level 15
assign po0321 = ~w12266;// level 15
assign po0322 = ~w16344;// level 15
assign po0323 = ~w14042;// level 15
assign po0324 = ~w1161;// level 15
assign po0325 = ~w15123;// level 15
assign po0326 = w16004;// level 11
assign po0327 = ~w15804;// level 15
assign po0328 = ~w1777;// level 15
assign po0329 = ~w4817;// level 15
assign po0330 = w1718;// level 11
assign po0331 = w8276;// level 12
assign po0332 = ~w4544;// level 14
assign po0333 = ~w10416;// level 12
assign po0334 = ~w14222;// level 12
assign po0335 = w4544;// level 14
assign po0336 = ~w8200;// level 6
assign po0337 = w2607;// level 8
assign po0338 = ~w2856;// level 8
assign po0339 = ~w2525;// level 8
assign po0340 = ~w5852;// level 8
assign po0341 = ~w11128;// level 8
assign po0342 = ~w12330;// level 8
assign po0343 = ~w15859;// level 8
assign po0344 = ~w2504;// level 11
assign po0345 = ~w17432;// level 11
assign po0346 = ~w7071;// level 11
assign po0347 = ~w18268;// level 11
assign po0348 = ~w17110;// level 11
assign po0349 = ~w7294;// level 11
assign po0350 = ~w340;// level 11
assign po0351 = ~w13146;// level 11
assign po0352 = ~w18072;// level 11
assign po0353 = ~w150;// level 11
assign po0354 = ~w4349;// level 11
assign po0355 = ~w9823;// level 11
assign po0356 = ~w5304;// level 11
assign po0357 = ~w16234;// level 11
assign po0358 = ~w5599;// level 11
assign po0359 = ~w17609;// level 11
assign po0360 = ~w2589;// level 11
assign po0361 = ~w17572;// level 11
assign po0362 = ~w11521;// level 11
assign po0363 = ~w8714;// level 11
assign po0364 = ~w4505;// level 11
assign po0365 = ~w6774;// level 11
assign po0366 = ~w6851;// level 11
assign po0367 = ~w1170;// level 11
assign po0368 = ~w6841;// level 11
assign po0369 = ~w3927;// level 11
assign po0370 = ~w15120;// level 11
assign po0371 = ~w2546;// level 11
assign po0372 = ~w1165;// level 11
assign po0373 = ~w10995;// level 11
assign po0374 = ~w10614;// level 11
assign po0375 = ~w10768;// level 11
assign po0376 = ~w3161;// level 11
assign po0377 = ~w14550;// level 11
assign po0378 = ~w4238;// level 11
assign po0379 = ~w6548;// level 11
assign po0380 = ~w4299;// level 11
assign po0381 = ~w3925;// level 11
assign po0382 = ~w8306;// level 11
assign po0383 = ~w12056;// level 11
assign po0384 = ~w1871;// level 11
assign po0385 = ~w14975;// level 11
assign po0386 = ~w15100;// level 11
assign po0387 = ~w6467;// level 11
assign po0388 = ~w2783;// level 11
assign po0389 = ~w16496;// level 11
assign po0390 = ~w16909;// level 11
assign po0391 = ~w11972;// level 11
assign po0392 = ~w6504;// level 11
assign po0393 = ~w13471;// level 11
assign po0394 = ~w10699;// level 11
assign po0395 = ~w14253;// level 12
assign po0396 = ~w705;// level 11
assign po0397 = ~w18192;// level 12
assign po0398 = ~w2512;// level 11
assign po0399 = ~w14608;// level 11
assign po0400 = ~w13270;// level 6
assign po0401 = ~w6016;// level 12
assign po0402 = ~w10015;// level 12
assign po0403 = ~w13886;// level 12
assign po0404 = ~w847;// level 12
assign po0405 = w9954;// level 13
assign po0406 = ~w7859;// level 12
assign po0407 = ~w6877;// level 12
assign po0408 = ~w17616;// level 7
assign po0409 = ~w14858;// level 7
assign po0410 = ~w3478;// level 7
assign po0411 = ~w7282;// level 9
assign po0412 = ~w2857;// level 9
assign po0413 = ~w9921;// level 9
assign po0414 = ~w3907;// level 9
assign po0415 = ~w12264;// level 9
assign po0416 = ~w1988;// level 9
assign po0417 = ~w13734;// level 9
assign po0418 = ~w14021;// level 9
assign po0419 = ~w9644;// level 9
assign po0420 = ~w710;// level 9
assign po0421 = ~w11951;// level 9
assign po0422 = ~w2839;// level 13
assign po0423 = ~w17972;// level 14
assign po0424 = ~w15867;// level 13
assign po0425 = ~w9534;// level 3
assign po0426 = ~w9859;// level 9
assign po0427 = ~w6710;// level 9
assign po0428 = ~w12103;// level 9
assign po0429 = ~w14070;// level 9
assign po0430 = ~w16867;// level 9
assign po0431 = w17972;// level 14
assign po0432 = ~w6721;// level 9
assign po0433 = ~w17426;// level 9
assign po0434 = ~w407;// level 9
assign po0435 = ~w668;// level 9
assign po0436 = ~w3696;// level 9
assign po0437 = ~w986;// level 9
assign po0438 = ~w3142;// level 9
assign po0439 = ~w13208;// level 9
assign po0440 = ~w17452;// level 9
assign po0441 = ~w10968;// level 9
assign po0442 = ~w3066;// level 9
assign po0443 = ~w15595;// level 9
assign po0444 = ~w8114;// level 9
assign po0445 = ~w15648;// level 9
assign po0446 = ~w10162;// level 9
assign po0447 = ~w11627;// level 9
assign po0448 = w16531;// level 10
assign po0449 = w11597;// level 9
assign po0450 = w2722;// level 10
assign po0451 = w12446;// level 9
assign po0452 = ~w4633;// level 9
assign po0453 = w4524;// level 10
assign po0454 = w13106;// level 10
assign po0455 = w5486;// level 10
assign po0456 = w1717;// level 10
assign po0457 = w12286;// level 10
assign po0458 = w5676;// level 10
assign po0459 = w4681;// level 10
assign po0460 = w151;// level 10
assign po0461 = w3860;// level 9
assign po0462 = w13652;// level 9
assign po0463 = w2371;// level 9
assign po0464 = w17516;// level 9
assign po0465 = ~w18330;// level 8
assign po0466 = ~w14072;// level 10
assign po0467 = ~w10896;// level 11
assign po0468 = w3912;// level 9
assign po0469 = w10921;// level 9
assign po0470 = w3989;// level 10
assign po0471 = w12412;// level 10
assign po0472 = w4952;// level 10
assign po0473 = w16968;// level 9
assign po0474 = ~w811;// level 7
assign po0475 = ~w18026;// level 7
assign po0476 = ~w5268;// level 8
assign po0477 = ~w17058;// level 8
assign po0478 = ~w18140;// level 8
assign po0479 = ~w12869;// level 8
assign po0480 = ~w4010;// level 8
assign po0481 = ~w15904;// level 8
assign po0482 = ~w9336;// level 8
assign po0483 = ~w955;// level 8
assign po0484 = ~w7908;// level 8
assign po0485 = ~w1776;// level 8
assign po0486 = ~w17235;// level 8
assign po0487 = ~w5332;// level 8
assign po0488 = ~w17524;// level 8
assign po0489 = ~w12547;// level 8
assign po0490 = ~w10751;// level 8
assign po0491 = ~w10091;// level 8
assign po0492 = ~w13626;// level 8
assign po0493 = ~w5750;// level 8
assign po0494 = ~w1782;// level 8
assign po0495 = ~w12539;// level 8
assign po0496 = ~w9645;// level 8
assign po0497 = ~w4773;// level 8
assign po0498 = ~w17305;// level 8
assign po0499 = w284;// level 10
assign po0500 = w9384;// level 10
assign po0501 = w10925;// level 10
assign po0502 = w6307;// level 9
assign po0503 = w15639;// level 10
assign po0504 = ~w8076;// level 9
assign po0505 = w1440;// level 10
assign po0506 = ~w5887;// level 8
assign po0507 = ~w9500;// level 8
assign po0508 = ~w15570;// level 8
assign po0509 = ~w10278;// level 8
assign po0510 = w10591;// level 10
assign po0511 = ~w7706;// level 10
assign po0512 = w9888;// level 10
assign po0513 = ~w14993;// level 10
assign po0514 = ~w2868;// level 9
assign po0515 = ~w7940;// level 9
assign po0516 = ~w4031;// level 9
assign po0517 = w9392;// level 9
assign po0518 = w2796;// level 9
assign po0519 = w4983;// level 9
assign po0520 = w5110;// level 9
assign po0521 = w14609;// level 9
assign po0522 = w10690;// level 9
assign po0523 = ~w8052;// level 9
assign po0524 = w17053;// level 9
assign po0525 = w14154;// level 9
assign po0526 = w13716;// level 10
assign po0527 = ~w18430;// level 8
assign po0528 = ~w11848;// level 8
assign po0529 = ~w8004;// level 8
assign po0530 = ~w3670;// level 8
assign po0531 = ~w5923;// level 8
assign po0532 = ~w1086;// level 8
assign po0533 = ~w9327;// level 7
assign po0534 = ~w16862;// level 8
assign po0535 = ~w16869;// level 8
assign po0536 = ~w14648;// level 9
assign po0537 = w598;// level 10
assign po0538 = w3000;// level 9
assign po0539 = w15122;// level 9
assign po0540 = w17553;// level 9
assign po0541 = ~w16176;// level 16
assign po0542 = ~w8663;// level 16
assign po0543 = ~w17347;// level 16
assign po0544 = ~w11177;// level 16
assign po0545 = ~w3287;// level 16
assign po0546 = ~w17973;// level 16
assign po0547 = ~w2544;// level 16
assign po0548 = ~w9538;// level 16
assign po0549 = ~w404;// level 16
assign po0550 = ~w1367;// level 16
assign po0551 = ~w10293;// level 16
assign po0552 = ~w12437;// level 8
assign po0553 = ~w10256;// level 16
assign po0554 = ~w2697;// level 16
assign po0555 = ~w3268;// level 16
assign po0556 = ~w4843;// level 16
assign po0557 = ~w17462;// level 16
assign po0558 = ~w8650;// level 16
assign po0559 = ~w10871;// level 16
assign po0560 = ~w15268;// level 8
assign po0561 = ~w15582;// level 16
assign po0562 = ~w17583;// level 16
assign po0563 = ~w12626;// level 16
assign po0564 = ~w12386;// level 16
assign po0565 = ~w9208;// level 16
assign po0566 = ~w8153;// level 16
assign po0567 = ~w16646;// level 16
assign po0568 = ~w1909;// level 16
assign po0569 = ~w16139;// level 16
assign po0570 = ~w5972;// level 16
assign po0571 = ~w3573;// level 16
assign po0572 = ~w10439;// level 16
assign po0573 = ~w1983;// level 16
assign po0574 = ~w18327;// level 16
assign po0575 = ~w6792;// level 16
assign po0576 = ~w3415;// level 16
assign po0577 = w4292;// level 8
assign po0578 = w15050;// level 8
assign po0579 = w6321;// level 8
assign po0580 = ~pi0411;// level 0
assign po0581 = w8862;// level 8
assign po0582 = w15827;// level 8
assign po0583 = w10419;// level 8
assign po0584 = w14013;// level 8
assign po0585 = w10060;// level 8
assign po0586 = w16984;// level 8
assign po0587 = w9643;// level 8
assign po0588 = w11233;// level 8
assign po0589 = w2338;// level 8
assign po0590 = w10071;// level 8
assign po0591 = w17246;// level 8
assign po0592 = w3365;// level 8
assign po0593 = w2502;// level 8
assign po0594 = w16727;// level 8
assign po0595 = w5605;// level 8
assign po0596 = w2922;// level 8
assign po0597 = w14323;// level 8
assign po0598 = w10598;// level 8
assign po0599 = w8464;// level 8
assign po0600 = w18141;// level 8
assign po0601 = w9448;// level 8
assign po0602 = w4468;// level 8
assign po0603 = w13332;// level 8
assign po0604 = w7874;// level 8
assign po0605 = w5365;// level 8
assign po0606 = w9358;// level 8
assign po0607 = w14780;// level 8
assign po0608 = w6285;// level 8
assign po0609 = w4081;// level 8
assign po0610 = ~w16685;// level 16
assign po0611 = ~w9129;// level 1
assign po0612 = ~w16492;// level 16
assign po0613 = ~w16333;// level 16
assign po0614 = ~w10712;// level 16
assign po0615 = ~w8865;// level 16
assign po0616 = ~w13461;// level 16
assign po0617 = ~w14092;// level 16
assign po0618 = ~w5685;// level 16
assign po0619 = ~w15593;// level 16
assign po0620 = ~w121;// level 16
assign po0621 = ~w13808;// level 16
assign po0622 = ~w10165;// level 16
assign po0623 = ~w2622;// level 16
assign po0624 = ~w135;// level 16
assign po0625 = ~w6371;// level 16
assign po0626 = ~w10774;// level 16
assign po0627 = ~w16715;// level 16
assign po0628 = ~w16546;// level 16
assign po0629 = ~w12552;// level 16
assign po0630 = ~w17920;// level 16
assign po0631 = ~w14536;// level 16
assign po0632 = ~w6004;// level 16
assign po0633 = ~w9272;// level 16
assign po0634 = ~w14901;// level 16
assign po0635 = ~w18043;// level 16
assign po0636 = ~w6461;// level 16
assign po0637 = ~w12090;// level 16
assign po0638 = ~w14667;// level 16
assign po0639 = ~w1939;// level 16
assign po0640 = ~w2695;// level 16
assign po0641 = ~w18433;// level 16
assign po0642 = ~w15621;// level 16
assign po0643 = ~w15905;// level 16
assign po0644 = ~w9515;// level 16
assign po0645 = w9129;// level 1
assign po0646 = ~w6269;// level 16
assign po0647 = ~w3994;// level 16
assign po0648 = ~w10200;// level 16
assign po0649 = ~w9878;// level 13
assign po0650 = ~w5265;// level 13
assign po0651 = ~w3877;// level 13
assign po0652 = ~w10843;// level 7
assign po0653 = ~w10672;// level 13
assign po0654 = ~w15126;// level 13
assign po0655 = ~w16870;// level 13
assign po0656 = ~w5284;// level 13
assign po0657 = ~w9220;// level 13
assign po0658 = ~w14375;// level 13
assign po0659 = ~w4854;// level 13
assign po0660 = ~w8377;// level 13
assign po0661 = ~w14264;// level 13
assign po0662 = ~w1635;// level 13
assign po0663 = ~w9369;// level 13
assign po0664 = ~w14280;// level 13
assign po0665 = ~w592;// level 13
assign po0666 = ~w14712;// level 13
assign po0667 = ~w8856;// level 13
assign po0668 = ~w18065;// level 13
assign po0669 = ~w7989;// level 13
assign po0670 = ~w12850;// level 13
assign po0671 = ~w14935;// level 13
assign po0672 = ~w104;// level 13
assign po0673 = ~w118;// level 13
assign po0674 = ~w11429;// level 13
assign po0675 = ~w13750;// level 13
assign po0676 = ~w10568;// level 13
assign po0677 = ~w8422;// level 13
assign po0678 = ~w10760;// level 13
assign po0679 = ~w7237;// level 13
assign po0680 = ~w1301;// level 13
assign po0681 = ~w12628;// level 13
assign po0682 = ~w11616;// level 13
assign po0683 = w3453;// level 12
assign po0684 = ~w2019;// level 9
assign po0685 = ~w2935;// level 11
assign po0686 = ~w15205;// level 11
assign po0687 = ~w13776;// level 11
assign po0688 = ~w15090;// level 11
assign po0689 = ~w4494;// level 12
assign po0690 = ~w1317;// level 11
assign po0691 = ~w9200;// level 11
assign po0692 = w14142;// level 11
assign po0693 = w13281;// level 10
assign po0694 = w2833;// level 11
assign po0695 = ~w15414;// level 11
assign po0696 = ~w10523;// level 12
assign po0697 = ~w8353;// level 11
assign po0698 = ~w8792;// level 12
assign po0699 = ~w10573;// level 12
assign po0700 = ~w4212;// level 12
assign po0701 = w13020;// level 11
assign po0702 = ~w6976;// level 11
assign po0703 = ~w10394;// level 12
assign po0704 = ~w788;// level 12
assign po0705 = ~w17497;// level 11
assign po0706 = ~w8459;// level 12
assign po0707 = ~w10805;// level 12
assign po0708 = ~w5656;// level 12
assign po0709 = w9790;// level 9
assign po0710 = ~w4319;// level 12
assign po0711 = ~w12122;// level 11
assign po0712 = ~w10583;// level 11
assign po0713 = ~w15597;// level 12
assign po0714 = ~w4699;// level 11
assign po0715 = ~w6156;// level 11
assign po0716 = w11441;// level 8
assign po0717 = w6820;// level 8
assign po0718 = w16488;// level 8
assign po0719 = w14875;// level 13
assign po0720 = w14875;// level 13
assign po0721 = w14875;// level 13
assign po0722 = w14875;// level 13
assign po0723 = w14875;// level 13
assign po0724 = w14875;// level 13
assign po0725 = w14875;// level 13
assign po0726 = w14875;// level 13
assign po0727 = w14875;// level 13
assign po0728 = w14875;// level 13
assign po0729 = w14875;// level 13
assign po0730 = w14875;// level 13
assign po0731 = w8390;// level 8
assign po0732 = w10170;// level 8
assign po0733 = w2104;// level 8
assign po0734 = w14595;// level 8
assign po0735 = w140;// level 8
assign po0736 = w14469;// level 8
assign po0737 = w15023;// level 8
assign po0738 = w16858;// level 8
assign po0739 = w8233;// level 8
assign po0740 = w15973;// level 8
assign po0741 = w14547;// level 8
assign po0742 = w17802;// level 8
assign po0743 = w13371;// level 8
assign po0744 = w804;// level 8
assign po0745 = w14048;// level 8
assign po0746 = w12612;// level 8
assign po0747 = w16523;// level 8
assign po0748 = w11964;// level 8
assign po0749 = w17541;// level 8
assign po0750 = w3804;// level 8
assign po0751 = w4792;// level 8
assign po0752 = w5123;// level 8
assign po0753 = w13536;// level 8
assign po0754 = w3413;// level 8
assign po0755 = w14338;// level 8
assign po0756 = w6678;// level 8
assign po0757 = w17845;// level 8
assign po0758 = w4748;// level 8
assign po0759 = w2518;// level 8
assign po0760 = w2030;// level 8
assign po0761 = w14194;// level 8
assign po0762 = w18170;// level 8
assign po0763 = w617;// level 8
assign po0764 = w10289;// level 8
assign po0765 = w2209;// level 8
assign po0766 = w5270;// level 8
assign po0767 = w17491;// level 8
assign po0768 = w573;// level 8
assign po0769 = w8296;// level 8
assign po0770 = w5786;// level 8
assign po0771 = w14642;// level 8
assign po0772 = w1157;// level 8
assign po0773 = w13267;// level 8
assign po0774 = w15902;// level 8
assign po0775 = w4467;// level 8
assign po0776 = w7588;// level 8
assign po0777 = w8621;// level 8
assign po0778 = w9862;// level 8
assign po0779 = w17484;// level 8
assign po0780 = w3328;// level 8
assign po0781 = w3526;// level 8
assign po0782 = w16335;// level 8
assign po0783 = w10504;// level 8
assign po0784 = w16863;// level 8
assign po0785 = w9471;// level 8
assign po0786 = w6590;// level 8
assign po0787 = w1628;// level 8
assign po0788 = w6621;// level 8
assign po0789 = w2396;// level 8
assign po0790 = w6366;// level 8
assign po0791 = w7275;// level 8
assign po0792 = w9183;// level 8
assign po0793 = w12389;// level 8
assign po0794 = w17261;// level 8
assign po0795 = w5970;// level 8
assign po0796 = w12730;// level 8
assign po0797 = w15418;// level 8
assign po0798 = w7913;// level 8
assign po0799 = w17175;// level 8
assign po0800 = w1107;// level 8
assign po0801 = w14752;// level 8
assign po0802 = w14668;// level 8
assign po0803 = w2612;// level 8
assign po0804 = w17829;// level 8
assign po0805 = w4971;// level 8
assign po0806 = w11107;// level 8
assign po0807 = w8592;// level 8
assign po0808 = w12510;// level 8
assign po0809 = w15731;// level 8
assign po0810 = w13697;// level 8
assign po0811 = w13048;// level 8
assign po0812 = w5804;// level 8
assign po0813 = w15079;// level 8
assign po0814 = w12574;// level 8
assign po0815 = w9983;// level 8
assign po0816 = w9195;// level 8
assign po0817 = w6845;// level 8
assign po0818 = w16734;// level 8
assign po0819 = w246;// level 8
assign po0820 = w9219;// level 8
assign po0821 = w7809;// level 8
assign po0822 = w10555;// level 8
assign po0823 = w5553;// level 8
assign po0824 = w7280;// level 8
assign po0825 = w2496;// level 8
assign po0826 = w6209;// level 8
assign po0827 = w11615;// level 8
assign po0828 = w17505;// level 8
assign po0829 = w14881;// level 8
assign po0830 = w16591;// level 8
assign po0831 = w8687;// level 8
assign po0832 = w138;// level 8
assign po0833 = w7510;// level 8
assign po0834 = w6861;// level 8
assign po0835 = w5084;// level 8
assign po0836 = w8797;// level 8
assign po0837 = w10365;// level 8
assign po0838 = w9811;// level 8
assign po0839 = w11174;// level 8
assign po0840 = w17020;// level 8
assign po0841 = w15615;// level 8
assign po0842 = w4377;// level 8
assign po0843 = w4726;// level 8
assign po0844 = w13823;// level 8
assign po0845 = w4160;// level 8
assign po0846 = w14582;// level 8
assign po0847 = w7641;// level 8
assign po0848 = w13680;// level 8
assign po0849 = w16089;// level 8
assign po0850 = w4300;// level 8
assign po0851 = w2062;// level 8
assign po0852 = w2438;// level 8
assign po0853 = w15067;// level 8
assign po0854 = w18231;// level 8
assign po0855 = w8488;// level 8
assign po0856 = w9124;// level 8
assign po0857 = w4316;// level 8
assign po0858 = w7466;// level 8
assign po0859 = w12748;// level 8
assign po0860 = w11791;// level 8
assign po0861 = w11543;// level 8
assign po0862 = w2644;// level 8
assign po0863 = w4865;// level 8
assign po0864 = w12820;// level 8
assign po0865 = w72;// level 8
assign po0866 = w10471;// level 8
assign po0867 = w2105;// level 8
assign po0868 = w53;// level 8
assign po0869 = w5835;// level 8
assign po0870 = w14219;// level 8
assign po0871 = w3533;// level 8
assign po0872 = w10933;// level 8
assign po0873 = w2373;// level 8
assign po0874 = w3712;// level 8
assign po0875 = w12702;// level 8
assign po0876 = w14487;// level 8
assign po0877 = w9641;// level 8
assign po0878 = w7719;// level 8
assign po0879 = w5230;// level 8
assign po0880 = w8116;// level 8
assign po0881 = w11768;// level 8
assign po0882 = w13699;// level 8
assign po0883 = w18568;// level 8
assign po0884 = w4191;// level 8
assign po0885 = w17032;// level 8
assign po0886 = w4226;// level 8
assign po0887 = w904;// level 8
assign po0888 = w7503;// level 8
assign po0889 = w6239;// level 8
assign po0890 = w4416;// level 8
assign po0891 = w4443;// level 8
assign po0892 = w13908;// level 8
assign po0893 = w18039;// level 8
assign po0894 = w3571;// level 8
assign po0895 = w14324;// level 8
assign po0896 = w1251;// level 8
assign po0897 = w7255;// level 8
assign po0898 = w15708;// level 8
assign po0899 = w2312;// level 8
assign po0900 = w7471;// level 8
assign po0901 = w10404;// level 8
assign po0902 = w18477;// level 8
assign po0903 = w8234;// level 8
assign po0904 = w4426;// level 8
assign po0905 = w7362;// level 8
assign po0906 = w3376;// level 8
assign po0907 = w4445;// level 8
assign po0908 = w3141;// level 8
assign po0909 = w15403;// level 8
assign po0910 = w13145;// level 8
assign po0911 = w13271;// level 8
assign po0912 = w17227;// level 8
assign po0913 = w10089;// level 8
assign po0914 = w17425;// level 8
assign po0915 = w12033;// level 8
assign po0916 = w10842;// level 8
assign po0917 = w3153;// level 8
assign po0918 = w6867;// level 8
assign po0919 = w4705;// level 8
assign po0920 = w2679;// level 8
assign po0921 = w8224;// level 8
assign po0922 = w14527;// level 8
assign po0923 = w9291;// level 8
assign po0924 = w17956;// level 8
assign po0925 = w17877;// level 8
assign po0926 = w12156;// level 8
assign po0927 = w195;// level 8
assign po0928 = w7075;// level 8
assign po0929 = w17803;// level 8
assign po0930 = w13225;// level 8
assign po0931 = w18266;// level 8
assign po0932 = w14736;// level 8
assign po0933 = w15860;// level 8
assign po0934 = w5915;// level 8
assign po0935 = w1403;// level 8
assign po0936 = w13084;// level 8
assign po0937 = w3135;// level 8
assign po0938 = w9185;// level 8
assign po0939 = w3966;// level 8
assign po0940 = w11293;// level 8
assign po0941 = w3896;// level 8
assign po0942 = w3789;// level 8
assign po0943 = w15770;// level 8
assign po0944 = w13775;// level 8
assign po0945 = w15661;// level 8
assign po0946 = w13201;// level 8
assign po0947 = w12204;// level 8
assign po0948 = w6247;// level 8
assign po0949 = w14179;// level 8
assign po0950 = w4673;// level 8
assign po0951 = w7298;// level 8
assign po0952 = w4267;// level 8
assign po0953 = w4479;// level 8
assign po0954 = w3881;// level 8
assign po0955 = w7615;// level 8
assign po0956 = w5885;// level 8
assign po0957 = w17519;// level 8
assign po0958 = w10002;// level 8
assign po0959 = w18000;// level 8
assign po0960 = w11326;// level 8
assign po0961 = w9221;// level 8
assign po0962 = w984;// level 8
assign po0963 = w10102;// level 8
assign po0964 = w15313;// level 8
assign po0965 = w6068;// level 8
assign po0966 = w7261;// level 8
assign po0967 = w12790;// level 8
assign po0968 = w15936;// level 8
assign po0969 = w13766;// level 8
assign po0970 = w15652;// level 8
assign po0971 = w5305;// level 8
assign po0972 = w7472;// level 8
assign po0973 = w17763;// level 8
assign po0974 = w11092;// level 8
assign po0975 = w14278;// level 8
assign po0976 = w3661;// level 8
assign po0977 = w6596;// level 8
assign po0978 = w6363;// level 8
assign po0979 = w18455;// level 8
assign po0980 = w15753;// level 8
assign po0981 = w6105;// level 8
assign po0982 = w15439;// level 8
assign po0983 = w14075;// level 8
assign po0984 = w13323;// level 8
assign po0985 = w13117;// level 8
assign po0986 = w4918;// level 8
assign po0987 = w10030;// level 8
assign po0988 = w16083;// level 8
assign po0989 = w3250;// level 8
assign po0990 = w15833;// level 8
assign po0991 = w310;// level 8
assign po0992 = w7036;// level 8
assign po0993 = w607;// level 8
assign po0994 = w14467;// level 8
assign po0995 = w15380;// level 8
assign po0996 = w9447;// level 8
assign po0997 = w18572;// level 8
assign po0998 = w14361;// level 8
assign po0999 = w16048;// level 8
assign po1000 = w4805;// level 8
assign po1001 = w5794;// level 8
assign po1002 = w6513;// level 8
assign po1003 = w15571;// level 8
assign po1004 = w8713;// level 8
assign po1005 = w6234;// level 8
assign po1006 = w16224;// level 8
assign po1007 = w14339;// level 8
assign po1008 = w813;// level 8
assign po1009 = w11832;// level 8
assign po1010 = w13713;// level 8
assign po1011 = w11184;// level 8
assign po1012 = w13934;// level 8
assign po1013 = w12794;// level 8
assign po1014 = w17957;// level 8
assign po1015 = w15747;// level 8
assign po1016 = w1228;// level 8
assign po1017 = w8998;// level 8
assign po1018 = w4386;// level 8
assign po1019 = w3440;// level 8
assign po1020 = w3917;// level 8
assign po1021 = w17245;// level 8
assign po1022 = w17900;// level 8
assign po1023 = w15000;// level 8
assign po1024 = w1669;// level 8
assign po1025 = w1761;// level 8
assign po1026 = w12949;// level 8
assign po1027 = w6907;// level 8
assign po1028 = w8910;// level 8
assign po1029 = w11538;// level 8
assign po1030 = w17489;// level 8
assign po1031 = w17105;// level 8
assign po1032 = w7778;// level 8
assign po1033 = w10617;// level 8
assign po1034 = w6096;// level 8
assign po1035 = w15413;// level 8
assign po1036 = w7243;// level 8
assign po1037 = w11276;// level 8
assign po1038 = w7185;// level 8
assign po1039 = w12199;// level 8
assign po1040 = w7642;// level 8
assign po1041 = w12361;// level 8
assign po1042 = w6614;// level 8
assign po1043 = w9526;// level 8
assign po1044 = w6159;// level 8
assign po1045 = w16003;// level 8
assign po1046 = w4567;// level 8
assign po1047 = w16934;// level 8
assign po1048 = w17253;// level 8
assign po1049 = w12270;// level 8
assign po1050 = w1111;// level 8
assign po1051 = w3304;// level 8
assign po1052 = w15187;// level 8
assign po1053 = w2844;// level 8
assign po1054 = w14946;// level 8
assign po1055 = w17369;// level 8
assign po1056 = w17691;// level 8
assign po1057 = w17966;// level 8
assign po1058 = w1713;// level 8
assign po1059 = w10112;// level 8
assign po1060 = w713;// level 8
assign po1061 = w11874;// level 8
assign po1062 = w17169;// level 8
assign po1063 = w14900;// level 8
assign po1064 = w8241;// level 8
assign po1065 = w10600;// level 6
assign po1066 = w2772;// level 8
assign po1067 = w11719;// level 8
assign po1068 = w3951;// level 8
assign po1069 = w3754;// level 8
assign po1070 = w5817;// level 8
assign po1071 = w14422;// level 8
assign po1072 = w15960;// level 8
assign po1073 = w11886;// level 8
assign po1074 = w6735;// level 8
assign po1075 = w15790;// level 8
assign po1076 = w10137;// level 8
assign po1077 = w12528;// level 8
assign po1078 = w16147;// level 8
assign po1079 = w794;// level 8
assign po1080 = w1067;// level 8
assign po1081 = w13283;// level 8
assign po1082 = w7144;// level 8
assign po1083 = w10907;// level 8
assign po1084 = w6391;// level 12
assign po1085 = w6169;// level 8
assign po1086 = w86;// level 8
assign po1087 = w9298;// level 8
assign po1088 = w6856;// level 8
assign po1089 = w3221;// level 8
assign po1090 = w18031;// level 8
assign po1091 = w3218;// level 8
assign po1092 = w11451;// level 8
assign po1093 = w827;// level 8
assign po1094 = w18323;// level 8
assign po1095 = w6772;// level 8
assign po1096 = w616;// level 8
assign po1097 = w7561;// level 8
assign po1098 = w10576;// level 8
assign po1099 = w1164;// level 8
assign po1100 = w4400;// level 8
assign po1101 = w4187;// level 8
assign po1102 = w8047;// level 8
assign po1103 = w15410;// level 8
assign po1104 = w6233;// level 8
assign po1105 = w5748;// level 8
assign po1106 = w77;// level 8
assign po1107 = w10431;// level 8
assign po1108 = w2279;// level 8
assign po1109 = w11079;// level 8
assign po1110 = w14613;// level 8
assign po1111 = w17292;// level 8
assign po1112 = w14512;// level 8
assign po1113 = w15522;// level 8
assign po1114 = w5013;// level 8
assign po1115 = w17399;// level 8
assign po1116 = w17778;// level 8
assign po1117 = w17917;// level 8
assign po1118 = w13069;// level 8
assign po1119 = w1346;// level 8
assign po1120 = w8174;// level 8
assign po1121 = w31;// level 8
assign po1122 = w11473;// level 8
assign po1123 = w16540;// level 8
assign po1124 = w15315;// level 8
assign po1125 = w1305;// level 8
assign po1126 = w13162;// level 8
assign po1127 = w1491;// level 8
assign po1128 = w15148;// level 8
assign po1129 = w5320;// level 8
assign po1130 = ~w18120;// level 8
assign po1131 = ~w8480;// level 8
assign po1132 = ~w8603;// level 8
assign po1133 = ~w15691;// level 8
assign po1134 = ~w12487;// level 8
assign po1135 = ~w15780;// level 8
assign po1136 = ~w9085;// level 8
assign po1137 = ~w16705;// level 8
assign po1138 = ~w16357;// level 8
assign po1139 = ~w1032;// level 8
assign po1140 = ~w8122;// level 8
assign po1141 = ~w9937;// level 8
assign po1142 = ~w3599;// level 8
assign po1143 = ~w2124;// level 8
assign po1144 = ~w4068;// level 8
assign po1145 = ~w8903;// level 8
assign po1146 = ~w17908;// level 8
assign po1147 = ~w7394;// level 8
assign po1148 = ~w3703;// level 8
assign po1149 = ~w2377;// level 8
assign po1150 = ~w4498;// level 8
assign po1151 = ~w10970;// level 8
assign po1152 = ~w19;// level 8
assign po1153 = ~w2038;// level 8
assign po1154 = ~w15391;// level 8
assign po1155 = w16614;// level 8
assign po1156 = ~w1884;// level 8
assign po1157 = ~w15940;// level 8
assign po1158 = ~w4645;// level 8
assign po1159 = ~w15068;// level 8
assign po1160 = ~w13190;// level 8
assign po1161 = ~w2183;// level 8
assign po1162 = ~w15738;// level 8
assign po1163 = w6542;// level 8
assign po1164 = w10150;// level 8
assign po1165 = w4844;// level 8
assign po1166 = w11523;// level 8
assign po1167 = w15764;// level 8
assign po1168 = ~w11093;// level 9
assign po1169 = w8894;// level 8
assign po1170 = w8391;// level 8
assign po1171 = w12801;// level 8
assign po1172 = w7438;// level 8
assign po1173 = w11779;// level 8
assign po1174 = w8612;// level 8
assign po1175 = w5072;// level 8
assign po1176 = w9701;// level 8
assign po1177 = w17308;// level 8
assign po1178 = w9119;// level 8
assign po1179 = w1763;// level 8
assign po1180 = w9922;// level 8
assign po1181 = w5801;// level 8
assign po1182 = w13326;// level 8
assign po1183 = w2691;// level 8
assign po1184 = w1837;// level 8
assign po1185 = w5792;// level 8
assign po1186 = w5588;// level 8
assign po1187 = w2806;// level 8
assign po1188 = w9815;// level 8
assign po1189 = w1719;// level 8
assign po1190 = w10488;// level 8
assign po1191 = w5575;// level 8
assign po1192 = w3568;// level 8
assign po1193 = w2594;// level 8
assign po1194 = w9876;// level 8
assign po1195 = w2476;// level 8
assign po1196 = w11870;// level 8
assign po1197 = w2718;// level 8
assign po1198 = w17099;// level 8
assign po1199 = w12774;// level 8
assign po1200 = w17265;// level 8
assign po1201 = w15377;// level 8
assign po1202 = w2172;// level 8
assign po1203 = w13589;// level 8
assign po1204 = w13646;// level 8
assign po1205 = w10693;// level 8
assign po1206 = w1073;// level 8
assign po1207 = w8032;// level 8
assign po1208 = w5871;// level 8
assign po1209 = w4090;// level 8
assign po1210 = w15543;// level 8
assign po1211 = w14079;// level 8
assign po1212 = w17478;// level 8
assign po1213 = w10732;// level 8
assign po1214 = w11607;// level 8
assign po1215 = w7197;// level 8
assign po1216 = w6930;// level 8
assign po1217 = w4902;// level 8
assign po1218 = w14031;// level 8
assign po1219 = w14263;// level 8
assign po1220 = w17086;// level 8
assign po1221 = w13240;// level 8
assign po1222 = w8235;// level 8
assign po1223 = w13533;// level 8
assign po1224 = w3695;// level 8
assign po1225 = w6262;// level 8
assign po1226 = w14556;// level 8
assign po1227 = w17749;// level 8
assign po1228 = w7933;// level 8
assign po1229 = w13053;// level 8
assign po1230 = w9112;// level 8
assign po1231 = w12740;// level 8
assign po1232 = w16160;// level 8
assign po1233 = w10948;// level 8
assign po1234 = w10082;// level 8
assign po1235 = w10442;// level 8
assign po1236 = w15797;// level 8
assign po1237 = w17191;// level 8
assign po1238 = w7679;// level 8
assign po1239 = w17094;// level 8
assign po1240 = w10796;// level 8
assign po1241 = w6859;// level 8
assign po1242 = w5073;// level 8
assign po1243 = w14558;// level 8
assign po1244 = w2876;// level 8
assign po1245 = w8967;// level 8
assign po1246 = w6712;// level 8
assign po1247 = w12456;// level 8
assign po1248 = w18388;// level 8
assign po1249 = w4063;// level 8
assign po1250 = w1471;// level 8
assign po1251 = w15532;// level 8
assign po1252 = w4579;// level 8
assign po1253 = w511;// level 8
assign po1254 = w828;// level 8
assign po1255 = w15511;// level 8
assign po1256 = w15108;// level 8
assign po1257 = w12718;// level 8
assign po1258 = w1654;// level 8
assign po1259 = w18052;// level 8
assign po1260 = w17936;// level 8
assign po1261 = w5115;// level 8
assign po1262 = w12413;// level 8
assign po1263 = w15433;// level 8
assign po1264 = w5172;// level 8
assign po1265 = w8061;// level 8
assign po1266 = w16217;// level 8
assign po1267 = w210;// level 8
assign po1268 = w17147;// level 8
assign po1269 = w3704;// level 8
assign po1270 = w16044;// level 8
assign po1271 = w9952;// level 8
assign po1272 = w4533;// level 8
assign po1273 = w11265;// level 8
assign po1274 = w13722;// level 8
assign po1275 = w2719;// level 8
assign po1276 = w9712;// level 8
assign po1277 = w4614;// level 8
assign po1278 = w12520;// level 8
assign po1279 = w1428;// level 8
assign po1280 = w4531;// level 8
assign po1281 = w12923;// level 8
assign po1282 = w6773;// level 8
assign po1283 = w14440;// level 8
assign po1284 = w13871;// level 8
assign po1285 = w3396;// level 8
assign po1286 = w12089;// level 8
assign po1287 = w9604;// level 8
assign po1288 = w13311;// level 8
assign po1289 = w1470;// level 8
assign po1290 = w10450;// level 8
assign po1291 = w7267;// level 8
assign po1292 = w1323;// level 8
assign po1293 = w15550;// level 8
assign po1294 = w9757;// level 8
assign po1295 = w15345;// level 8
assign po1296 = w17832;// level 8
assign po1297 = w14317;// level 8
assign po1298 = w12502;// level 8
assign po1299 = w10043;// level 8
assign po1300 = w18019;// level 8
assign po1301 = w1651;// level 8
assign po1302 = w16494;// level 8
assign po1303 = w8453;// level 8
assign po1304 = w9725;// level 8
assign po1305 = w4879;// level 8
assign po1306 = w16435;// level 8
assign po1307 = w16674;// level 8
assign po1308 = w14634;// level 11
assign po1309 = ~w15074;// level 10
assign po1310 = w3620;// level 11
assign po1311 = w17073;// level 11
assign po1312 = w3102;// level 8
assign po1313 = w9491;// level 8
assign po1314 = w7032;// level 8
assign po1315 = w5505;// level 8
assign po1316 = w11802;// level 8
assign po1317 = w13831;// level 8
assign po1318 = w14765;// level 8
assign po1319 = w686;// level 8
assign po1320 = w6452;// level 8
assign po1321 = w14464;// level 8
assign po1322 = w10649;// level 8
assign po1323 = w17322;// level 8
assign po1324 = w1310;// level 8
assign po1325 = w17223;// level 8
assign po1326 = w4814;// level 8
assign po1327 = w1376;// level 8
assign po1328 = w3233;// level 8
assign po1329 = w4309;// level 8
assign po1330 = w11710;// level 8
assign po1331 = w15478;// level 8
assign po1332 = w10475;// level 8
assign po1333 = w4953;// level 9
assign po1334 = ~w9767;// level 8
assign po1335 = w8843;// level 8
assign po1336 = w6565;// level 8
assign po1337 = w3349;// level 8
assign po1338 = w10318;// level 8
assign po1339 = w17080;// level 12
assign po1340 = w3047;// level 11
assign po1341 = ~w8256;// level 10
assign po1342 = w5780;// level 11
assign po1343 = ~w10360;// level 9
assign po1344 = ~w14171;// level 9
assign po1345 = ~w5508;// level 9
assign po1346 = w2407;// level 8
assign po1347 = ~w11472;// level 8
assign po1348 = ~w1290;// level 8
assign po1349 = ~w12818;// level 8
assign po1350 = ~w12316;// level 8
assign po1351 = ~w5534;// level 8
assign po1352 = ~w3148;// level 8
assign po1353 = w17652;// level 9
assign po1354 = w12871;// level 9
assign po1355 = ~w7239;// level 8
assign po1356 = ~w17588;// level 8
assign po1357 = ~w11460;// level 10
assign po1358 = ~w10467;// level 9
assign po1359 = w14203;// level 11
assign po1360 = w15937;// level 10
assign po1361 = w1556;// level 11
assign po1362 = ~w6625;// level 8
assign po1363 = w14177;// level 8
assign po1364 = w4252;// level 8
assign po1365 = w3857;// level 8
assign po1366 = w5493;// level 8
assign po1367 = w11534;// level 8
assign po1368 = w5883;// level 10
assign po1369 = w8361;// level 11
assign po1370 = w7086;// level 10
assign po1371 = w15778;// level 8
assign po1372 = w6862;// level 8
assign po1373 = w6806;// level 8
assign po1374 = ~w6428;// level 10
assign po1375 = w14996;// level 8
assign po1376 = w17915;// level 8
assign po1377 = w3820;// level 10
assign po1378 = w7325;// level 10
assign po1379 = ~w13735;// level 8
assign po1380 = w7835;// level 10
assign po1381 = ~w1504;// level 8
assign po1382 = w11634;// level 10
assign po1383 = w13357;// level 10
assign po1384 = w11900;// level 11
assign po1385 = w10228;// level 10
assign po1386 = w2763;// level 10
assign po1387 = w5701;// level 11
assign po1388 = w5916;// level 8
assign po1389 = w10930;// level 8
assign po1390 = w6331;// level 9
assign po1391 = w3062;// level 10
assign po1392 = w17335;// level 10
assign po1393 = w15494;// level 10
assign po1394 = ~w12632;// level 9
assign po1395 = ~w9637;// level 9
assign po1396 = ~w2789;// level 9
assign po1397 = ~w7134;// level 9
assign po1398 = ~w15965;// level 8
assign po1399 = ~w922;// level 6
assign po1400 = ~w15506;// level 11
assign po1401 = ~w14785;// level 10
assign po1402 = ~w13957;// level 9
assign po1403 = ~w12742;// level 9
assign po1404 = ~w6512;// level 10
assign po1405 = w15506;// level 11
assign po1406 = w6822;// level 5
assign po1407 = w4052;// level 9
assign po1408 = w16890;// level 8
assign po1409 = ~w10087;// level 9
assign po1410 = w14689;// level 10
assign po1411 = w2803;// level 5
assign po1412 = w6657;// level 5
assign po1413 = ~w17316;// level 8
assign po1414 = w17178;// level 3
assign po1415 = w1805;// level 4
assign po1416 = w8287;// level 4
assign po1417 = w7406;// level 11
assign po1418 = w15750;// level 9
assign po1419 = ~w15933;// level 9
assign po1420 = w5074;// level 9
assign po1421 = ~w6575;// level 9
assign po1422 = ~w11486;// level 9
assign po1423 = ~w14412;// level 9
assign po1424 = ~w11082;// level 9
assign po1425 = w9741;// level 9
assign po1426 = w10986;// level 9
assign po1427 = w4083;// level 9
assign po1428 = w12994;// level 9
assign po1429 = w15300;// level 9
assign po1430 = ~w11851;// level 9
assign po1431 = w12041;// level 9
assign po1432 = w671;// level 9
assign po1433 = ~w3492;// level 9
assign po1434 = ~w3381;// level 9
assign po1435 = w12037;// level 4
assign po1436 = w9896;// level 5
assign po1437 = w16621;// level 10
assign po1438 = ~w12360;// level 9
assign po1439 = w9086;// level 9
assign po1440 = ~w15912;// level 8
assign po1441 = ~w13754;// level 8
assign po1442 = ~w3016;// level 8
assign po1443 = w3407;// level 8
assign po1444 = w2225;// level 9
assign po1445 = ~w10724;// level 9
assign po1446 = ~w4173;// level 8
assign po1447 = w4566;// level 8
assign po1448 = w5124;// level 8
assign po1449 = ~w92;// level 9
assign po1450 = w9246;// level 8
assign po1451 = w8236;// level 8
assign po1452 = w7909;// level 8
assign po1453 = w4453;// level 8
assign po1454 = w506;// level 8
assign po1455 = w17142;// level 8
assign po1456 = w753;// level 8
assign po1457 = w12587;// level 8
assign po1458 = w8433;// level 8
assign po1459 = w16493;// level 8
assign po1460 = w8987;// level 8
assign po1461 = w856;// level 8
assign po1462 = w17784;// level 8
assign po1463 = w12381;// level 8
assign po1464 = w17710;// level 8
assign po1465 = w4041;// level 8
assign po1466 = w16839;// level 8
assign po1467 = ~w9631;// level 8
assign po1468 = ~w12602;// level 8
assign po1469 = ~w2729;// level 8
assign po1470 = w14579;// level 8
assign po1471 = w2400;// level 8
assign po1472 = w734;// level 8
assign po1473 = w17004;// level 8
assign po1474 = w8547;// level 7
assign po1475 = w6345;// level 7
assign po1476 = w14450;// level 8
assign po1477 = w14242;// level 8
assign po1478 = w18286;// level 7
assign po1479 = w18526;// level 7
assign po1480 = w3116;// level 7
assign po1481 = w15013;// level 7
assign po1482 = w5235;// level 7
assign po1483 = w17262;// level 9
assign po1484 = w6473;// level 7
assign po1485 = ~w15352;// level 9
assign po1486 = w9439;// level 8
assign po1487 = w8680;// level 9
assign po1488 = w17188;// level 8
assign po1489 = w11958;// level 9
assign po1490 = ~w10786;// level 9
assign po1491 = w11682;// level 8
assign po1492 = w2252;// level 7
assign po1493 = w10498;// level 8
assign po1494 = w9211;// level 7
assign po1495 = w8731;// level 8
assign po1496 = w8461;// level 7
assign po1497 = w10116;// level 9
assign po1498 = w6947;// level 9
assign po1499 = ~w7927;// level 9
assign po1500 = w1844;// level 9
assign po1501 = w8257;// level 9
assign po1502 = w7014;// level 9
assign po1503 = w15516;// level 9
assign po1504 = w8969;// level 9
assign po1505 = w3170;// level 9
assign po1506 = w17521;// level 9
assign po1507 = w16441;// level 9
assign po1508 = w9312;// level 8
assign po1509 = w5872;// level 9
assign po1510 = ~w8054;// level 9
assign po1511 = ~w9457;// level 7
assign po1512 = ~w14172;// level 7
assign po1513 = w15681;// level 8
assign po1514 = ~w11657;// level 10
assign po1515 = ~w9134;// level 10
assign po1516 = ~w17554;// level 7
assign po1517 = ~w18093;// level 7
assign po1518 = ~w3702;// level 7
assign po1519 = ~w3828;// level 7
assign po1520 = ~w8294;// level 7
assign po1521 = ~w16548;// level 10
assign po1522 = w12373;// level 8
assign po1523 = w15702;// level 7
assign po1524 = w9556;// level 16
assign po1525 = ~w14737;// level 6
assign po1526 = ~w2655;// level 7
assign po1527 = ~w14314;// level 7
assign po1528 = ~w4837;// level 6
assign po1529 = ~w4739;// level 7
assign po1530 = w6695;// level 9
assign po1531 = ~w13948;// level 7
assign po1532 = ~w17506;// level 7
assign po1533 = ~w6409;// level 7
assign po1534 = ~w3541;// level 7
assign po1535 = ~w7759;// level 6
assign po1536 = ~w16706;// level 6
assign po1537 = ~w12600;// level 6
assign po1538 = ~w2262;// level 6
assign po1539 = ~w4237;// level 6
assign po1540 = ~w6552;// level 7
assign po1541 = ~w7132;// level 7
assign po1542 = ~w15261;// level 6
assign po1543 = ~w4005;// level 9
assign po1544 = ~w1836;// level 7
assign po1545 = ~w3903;// level 7
assign po1546 = ~w12521;// level 9
assign po1547 = ~w17384;// level 7
assign po1548 = ~w3742;// level 7
assign po1549 = ~w5239;// level 7
assign po1550 = ~w4548;// level 10
assign po1551 = w6586;// level 13
assign po1552 = ~w8898;// level 7
assign po1553 = ~w612;// level 8
assign po1554 = ~w13026;// level 7
assign po1555 = ~w10148;// level 7
assign po1556 = ~w2043;// level 6
assign po1557 = w8457;// level 9
assign po1558 = w2162;// level 10
assign po1559 = w12232;// level 10
assign po1560 = w11945;// level 7
assign po1561 = w18521;// level 10
assign po1562 = w2578;// level 10
assign po1563 = w3343;// level 10
assign po1564 = w16787;// level 10
assign po1565 = w5798;// level 10
assign po1566 = w15151;// level 10
assign po1567 = w7857;// level 10
assign po1568 = w17472;// level 10
assign po1569 = w11522;// level 10
assign po1570 = w5876;// level 10
assign po1571 = w13975;// level 10
assign po1572 = ~w13170;// level 6
assign po1573 = ~w16022;// level 6
assign po1574 = ~w9350;// level 6
assign po1575 = w16981;// level 10
assign po1576 = ~w14211;// level 7
assign po1577 = ~w11166;// level 6
assign po1578 = ~w10036;// level 7
assign po1579 = ~w1089;// level 7
assign po1580 = ~w5787;// level 6
assign po1581 = ~w15885;// level 6
assign po1582 = w4421;// level 8
assign po1583 = w18074;// level 7
assign po1584 = ~w16687;// level 9
assign po1585 = w1833;// level 7
assign po1586 = w6289;// level 7
assign po1587 = ~w17639;// level 7
assign po1588 = w16704;// level 10
assign po1589 = w12629;// level 10
assign po1590 = w477;// level 10
assign po1591 = w12419;// level 10
assign po1592 = w3091;// level 10
assign po1593 = w6910;// level 10
assign po1594 = w4042;// level 10
assign po1595 = w13094;// level 10
assign po1596 = w16891;// level 10
assign po1597 = w18450;// level 10
assign po1598 = w17856;// level 10
assign po1599 = w13413;// level 10
assign po1600 = w5379;// level 10
assign po1601 = w8915;// level 10
assign po1602 = w12078;// level 10
assign po1603 = w2063;// level 10
assign po1604 = w16887;// level 10
assign po1605 = w11610;// level 10
assign po1606 = w5085;// level 10
assign po1607 = w12851;// level 10
assign po1608 = w4869;// level 10
assign po1609 = w12348;// level 10
assign po1610 = w3715;// level 10
assign po1611 = w7978;// level 10
assign po1612 = w4180;// level 10
assign po1613 = w13845;// level 10
assign po1614 = w14;// level 10
assign po1615 = w13674;// level 10
assign po1616 = w15846;// level 10
assign po1617 = w18270;// level 10
assign po1618 = w8258;// level 10
assign po1619 = w7801;// level 10
assign po1620 = w14709;// level 10
assign po1621 = w12673;// level 10
assign po1622 = w15894;// level 10
assign po1623 = w8342;// level 10
assign po1624 = w13980;// level 10
assign po1625 = w14380;// level 10
assign po1626 = w1758;// level 10
assign po1627 = w13046;// level 10
assign po1628 = w9389;// level 10
assign po1629 = w13885;// level 9
assign po1630 = w2820;// level 9
assign po1631 = w7115;// level 9
assign po1632 = w5938;// level 9
assign po1633 = w7067;// level 9
assign po1634 = w7226;// level 9
assign po1635 = w8857;// level 9
assign po1636 = w12272;// level 9
assign po1637 = w434;// level 9
assign po1638 = w7501;// level 9
assign po1639 = w16971;// level 9
assign po1640 = w18056;// level 9
assign po1641 = w16637;// level 9
assign po1642 = w8427;// level 9
assign po1643 = w3954;// level 9
assign po1644 = w17150;// level 9
assign po1645 = w11729;// level 9
assign po1646 = w4510;// level 9
assign po1647 = w15799;// level 9
assign po1648 = w9484;// level 9
assign po1649 = w2237;// level 9
assign po1650 = w17852;// level 9
assign po1651 = w884;// level 9
assign po1652 = w16090;// level 9
assign po1653 = w12685;// level 9
assign po1654 = w6284;// level 9
assign po1655 = w15528;// level 9
assign po1656 = w1014;// level 9
assign po1657 = w16422;// level 9
assign po1658 = w11849;// level 9
assign po1659 = w969;// level 9
assign po1660 = w2261;// level 9
assign po1661 = w2924;// level 9
assign po1662 = w3419;// level 9
assign po1663 = w861;// level 9
assign po1664 = w7048;// level 9
assign po1665 = w13040;// level 9
assign po1666 = w2489;// level 9
assign po1667 = w8102;// level 9
assign po1668 = w4754;// level 9
assign po1669 = w11289;// level 9
assign po1670 = w14289;// level 9
assign po1671 = w16959;// level 9
assign po1672 = w18592;// level 8
assign po1673 = w12999;// level 8
assign po1674 = w7414;// level 8
assign po1675 = w5286;// level 8
assign po1676 = w8852;// level 8
assign po1677 = w13415;// level 8
assign po1678 = w3916;// level 8
assign po1679 = w13852;// level 8
assign po1680 = w4358;// level 8
assign po1681 = w14771;// level 8
assign po1682 = w16917;// level 8
assign po1683 = w12055;// level 8
assign po1684 = w8516;// level 8
assign po1685 = w15082;// level 8
assign po1686 = w3336;// level 8
assign po1687 = w6000;// level 8
assign po1688 = w3798;// level 8
assign po1689 = w989;// level 8
assign po1690 = w6597;// level 10
assign po1691 = w3841;// level 10
assign po1692 = w2232;// level 10
assign po1693 = w17989;// level 10
assign po1694 = w239;// level 10
assign po1695 = w14181;// level 10
assign po1696 = w17209;// level 10
assign po1697 = w7351;// level 10
assign po1698 = w17510;// level 10
assign po1699 = w10561;// level 10
assign po1700 = w6796;// level 10
assign po1701 = w15018;// level 10
assign po1702 = w232;// level 10
assign po1703 = w1938;// level 10
assign po1704 = w17776;// level 10
assign po1705 = w1693;// level 10
assign po1706 = w5986;// level 10
assign po1707 = w942;// level 10
assign po1708 = w3530;// level 10
assign po1709 = w11023;// level 10
assign po1710 = w13168;// level 10
assign po1711 = w13342;// level 10
assign po1712 = w16682;// level 10
assign po1713 = w1590;// level 10
assign po1714 = w2224;// level 10
assign po1715 = w4715;// level 10
assign po1716 = w17755;// level 10
assign po1717 = w10683;// level 10
assign po1718 = w10537;// level 10
assign po1719 = w14589;// level 10
assign po1720 = w13191;// level 10
assign po1721 = w11144;// level 10
assign po1722 = w12527;// level 10
assign po1723 = w12563;// level 10
assign po1724 = w15480;// level 10
assign po1725 = w7204;// level 10
assign po1726 = w13797;// level 10
assign po1727 = w12425;// level 10
assign po1728 = w16525;// level 10
assign po1729 = w1076;// level 10
assign po1730 = w14224;// level 10
assign po1731 = w4930;// level 9
assign po1732 = w8014;// level 9
assign po1733 = w17079;// level 9
assign po1734 = w1675;// level 9
assign po1735 = w7577;// level 9
assign po1736 = w7203;// level 9
assign po1737 = w343;// level 9
assign po1738 = w13591;// level 9
assign po1739 = w5372;// level 9
assign po1740 = w13631;// level 9
assign po1741 = w18306;// level 9
assign po1742 = w17582;// level 9
assign po1743 = w805;// level 9
assign po1744 = w13320;// level 9
assign po1745 = w13800;// level 9
assign po1746 = w5856;// level 9
assign po1747 = w15800;// level 9
assign po1748 = w11542;// level 9
assign po1749 = w8821;// level 9
assign po1750 = w7841;// level 9
assign po1751 = w15279;// level 8
assign po1752 = w1972;// level 8
assign po1753 = w13022;// level 10
assign po1754 = w17598;// level 10
assign po1755 = w1338;// level 10
assign po1756 = w7928;// level 10
assign po1757 = w14662;// level 10
assign po1758 = w13891;// level 10
assign po1759 = w8524;// level 10
assign po1760 = w10333;// level 10
assign po1761 = w9608;// level 8
assign po1762 = w587;// level 10
assign po1763 = w17774;// level 10
assign po1764 = w16294;// level 8
assign po1765 = w6692;// level 9
assign po1766 = ~w7076;// level 6
assign po1767 = w7205;// level 8
assign po1768 = w5114;// level 8
assign po1769 = w18300;// level 8
assign po1770 = w16330;// level 8
assign po1771 = w9234;// level 8
assign po1772 = ~w10153;// level 7
assign po1773 = w627;// level 8
assign po1774 = w17443;// level 8
assign po1775 = w6708;// level 8
assign po1776 = w10886;// level 9
assign po1777 = w12513;// level 9
assign po1778 = w6592;// level 9
assign po1779 = w9850;// level 9
assign po1780 = w16418;// level 9
assign po1781 = w11221;// level 9
assign po1782 = w16827;// level 9
assign po1783 = w1810;// level 9
assign po1784 = w1990;// level 9
assign po1785 = w16080;// level 9
assign po1786 = w12849;// level 9
assign po1787 = w18046;// level 9
assign po1788 = w7609;// level 9
assign po1789 = w18151;// level 9
assign po1790 = w1390;// level 9
assign po1791 = w17608;// level 9
assign po1792 = w7044;// level 9
assign po1793 = w1773;// level 9
assign po1794 = w13287;// level 8
assign po1795 = w416;// level 9
assign po1796 = w10370;// level 8
assign po1797 = w6407;// level 9
assign po1798 = w7114;// level 9
assign po1799 = w1981;// level 8
assign po1800 = w2107;// level 9
assign po1801 = w17797;// level 10
assign po1802 = w9572;// level 9
assign po1803 = w17342;// level 10
assign po1804 = w5184;// level 9
assign po1805 = w8793;// level 9
assign po1806 = w17202;// level 9
assign po1807 = w15818;// level 9
assign po1808 = w18277;// level 10
assign po1809 = w5346;// level 10
assign po1810 = w17441;// level 9
assign po1811 = w18239;// level 9
assign po1812 = w3958;// level 10
assign po1813 = w16510;// level 9
assign po1814 = w6790;// level 9
assign po1815 = w12069;// level 10
assign po1816 = w7566;// level 9
assign po1817 = w2427;// level 10
assign po1818 = w5630;// level 10
assign po1819 = w2053;// level 9
assign po1820 = w4621;// level 9
assign po1821 = w16321;// level 10
assign po1822 = w3834;// level 10
assign po1823 = w16877;// level 10
assign po1824 = w5137;// level 10
assign po1825 = w13745;// level 10
assign po1826 = w11852;// level 10
assign po1827 = w8199;// level 10
assign po1828 = w863;// level 10
assign po1829 = w8864;// level 10
assign po1830 = w1017;// level 10
assign po1831 = w874;// level 10
assign po1832 = w15428;// level 10
assign po1833 = w1606;// level 10
assign po1834 = w18011;// level 10
assign po1835 = w12912;// level 10
assign po1836 = w5026;// level 10
assign po1837 = w17118;// level 10
assign po1838 = w459;// level 10
assign po1839 = ~w5759;// level 8
assign po1840 = ~w15729;// level 8
assign po1841 = ~w17756;// level 8
assign po1842 = ~w6346;// level 8
assign po1843 = ~w15025;// level 8
assign po1844 = ~w10516;// level 8
assign po1845 = ~w17181;// level 8
assign po1846 = ~w13647;// level 8
assign po1847 = ~w16104;// level 6
assign po1848 = ~w12233;// level 8
assign po1849 = ~w6438;// level 8
assign po1850 = ~w4474;// level 8
assign po1851 = ~w11780;// level 8
assign po1852 = ~w13540;// level 8
assign po1853 = w5527;// level 8
assign po1854 = ~w4429;// level 6
assign po1855 = ~w1750;// level 8
assign po1856 = ~w11011;// level 7
assign po1857 = ~w14266;// level 8
assign po1858 = ~w11699;// level 8
assign po1859 = ~w10454;// level 9
assign po1860 = ~w8037;// level 9
assign po1861 = ~w2580;// level 9
assign po1862 = w12338;// level 3
assign po1863 = w3113;// level 7
assign po1864 = ~w17323;// level 8
assign po1865 = w18579;// level 8
assign po1866 = w6964;// level 10
assign po1867 = w7081;// level 9
assign po1868 = w418;// level 10
assign po1869 = w664;// level 7
assign po1870 = ~w9333;// level 8
assign po1871 = ~w8237;// level 7
assign po1872 = w11998;// level 5
assign po1873 = w7830;// level 7
assign po1874 = ~w163;// level 7
assign po1875 = w14520;// level 8
assign po1876 = ~w15709;// level 6
assign po1877 = ~w13581;// level 6
assign po1878 = ~w6978;// level 6
assign po1879 = ~w12647;// level 6
assign po1880 = ~w16636;// level 6
assign po1881 = ~w4338;// level 6
assign po1882 = ~w10607;// level 6
assign po1883 = ~w14921;// level 6
assign po1884 = ~w4411;// level 8
assign po1885 = ~w13045;// level 6
assign po1886 = ~w15362;// level 6
assign po1887 = ~w16802;// level 8
assign po1888 = ~w13828;// level 8
assign po1889 = ~w9685;// level 6
assign po1890 = ~w17113;// level 8
assign po1891 = ~w11437;// level 8
assign po1892 = ~w12147;// level 8
assign po1893 = ~w18602;// level 8
assign po1894 = ~w8971;// level 8
assign po1895 = ~w7727;// level 8
assign po1896 = ~w3045;// level 8
assign po1897 = ~w11097;// level 8
assign po1898 = ~w16564;// level 8
assign po1899 = ~w8245;// level 8
assign po1900 = ~w14449;// level 8
assign po1901 = ~w2390;// level 9
assign po1902 = w855;// level 10
assign po1903 = ~w6598;// level 8
assign po1904 = ~w7387;// level 8
assign po1905 = ~w11902;// level 8
assign po1906 = ~w3739;// level 8
assign po1907 = ~w3529;// level 8
assign po1908 = ~w9979;// level 8
assign po1909 = ~w11541;// level 8
assign po1910 = ~w18446;// level 8
assign po1911 = ~w11308;// level 8
assign po1912 = ~w265;// level 8
assign po1913 = ~w6660;// level 8
assign po1914 = ~w2474;// level 8
assign po1915 = ~w10698;// level 8
assign po1916 = ~w5772;// level 8
assign po1917 = ~w13061;// level 8
assign po1918 = ~w10855;// level 8
assign po1919 = ~w6622;// level 8
assign po1920 = ~w11250;// level 8
assign po1921 = ~w14796;// level 8
assign po1922 = ~w602;// level 8
assign po1923 = w7729;// level 10
assign po1924 = w11706;// level 10
assign po1925 = w10860;// level 10
assign po1926 = w851;// level 10
assign po1927 = w2013;// level 12
assign po1928 = ~w8129;// level 8
assign po1929 = ~w10787;// level 8
assign po1930 = ~w16767;// level 8
assign po1931 = ~w15372;// level 8
assign po1932 = ~w10064;// level 8
assign po1933 = ~w15971;// level 7
assign po1934 = ~w16961;// level 7
assign po1935 = ~w8467;// level 7
assign po1936 = ~w14425;// level 6
assign po1937 = ~w12656;// level 6
assign po1938 = w9429;// level 12
assign po1939 = ~w13107;// level 9
assign po1940 = ~w8521;// level 8
assign po1941 = ~w14329;// level 8
assign po1942 = ~w8168;// level 8
assign po1943 = ~w9854;// level 8
assign po1944 = ~w1734;// level 8
assign po1945 = ~w11860;// level 6
assign po1946 = ~w7701;// level 6
assign po1947 = ~w15665;// level 6
assign po1948 = ~w3826;// level 6
assign po1949 = ~w6126;// level 6
assign po1950 = ~w12893;// level 6
assign po1951 = ~w14590;// level 6
assign po1952 = ~w18167;// level 6
assign po1953 = ~w1467;// level 6
assign po1954 = ~w11487;// level 8
assign po1955 = ~w1451;// level 8
assign po1956 = ~w10918;// level 7
assign po1957 = ~w17808;// level 7
assign po1958 = ~w14876;// level 7
assign po1959 = ~w11893;// level 7
assign po1960 = ~w15538;// level 7
assign po1961 = ~w10482;// level 7
assign po1962 = ~w3371;// level 7
assign po1963 = ~w15166;// level 7
assign po1964 = ~w11847;// level 7
assign po1965 = ~w6889;// level 7
assign po1966 = ~w14066;// level 7
assign po1967 = ~w7687;// level 7
assign po1968 = ~w12713;// level 7
assign po1969 = ~w16049;// level 7
assign po1970 = ~w12263;// level 7
assign po1971 = ~w3231;// level 7
assign po1972 = ~w17514;// level 7
assign po1973 = w167;// level 9
assign po1974 = ~w8022;// level 6
assign po1975 = ~w7792;// level 7
assign po1976 = ~w2398;// level 6
assign po1977 = ~w18255;// level 6
assign po1978 = ~w17975;// level 8
assign po1979 = ~w8636;// level 6
assign po1980 = ~w15139;// level 6
assign po1981 = ~w10916;// level 8
assign po1982 = w316;// level 9
assign po1983 = ~w14393;// level 7
assign po1984 = ~w12512;// level 7
assign po1985 = ~w6544;// level 7
assign po1986 = ~w16039;// level 7
assign po1987 = ~w4228;// level 7
assign po1988 = ~w16711;// level 6
assign po1989 = ~w12105;// level 7
assign po1990 = w11376;// level 7
assign po1991 = ~w4852;// level 7
assign po1992 = ~w4418;// level 7
assign po1993 = w9079;// level 11
assign po1994 = ~w9001;// level 7
assign po1995 = ~w3214;// level 7
assign po1996 = ~w7968;// level 7
assign po1997 = ~w15657;// level 7
assign po1998 = ~w16483;// level 7
assign po1999 = ~w16754;// level 7
assign po2000 = ~w6988;// level 7
assign po2001 = ~w5328;// level 7
assign po2002 = ~w9703;// level 7
assign po2003 = ~w10139;// level 7
assign po2004 = ~w2751;// level 9
assign po2005 = w7939;// level 11
assign po2006 = ~w11553;// level 13
assign po2007 = ~w1394;// level 13
assign po2008 = ~w2870;// level 13
assign po2009 = ~w5418;// level 14
assign po2010 = ~w6454;// level 13
assign po2011 = ~w1294;// level 13
assign po2012 = ~w455;// level 13
assign po2013 = ~w17884;// level 12
assign po2014 = ~w13;// level 13
assign po2015 = ~w14060;// level 14
assign po2016 = ~w7636;// level 13
assign po2017 = ~w12776;// level 14
assign po2018 = ~w10092;// level 13
assign po2019 = ~w14459;// level 13
assign po2020 = ~w17937;// level 13
assign po2021 = ~w2586;// level 14
assign po2022 = ~w3652;// level 7
assign po2023 = ~w17162;// level 7
assign po2024 = ~w3638;// level 7
assign po2025 = ~w4870;// level 7
assign po2026 = ~w15001;// level 7
assign po2027 = ~w16993;// level 7
assign po2028 = ~w6272;// level 7
assign po2029 = ~w13835;// level 7
assign po2030 = ~w14514;// level 7
assign po2031 = ~w17953;// level 7
assign po2032 = ~w7458;// level 7
assign po2033 = w3645;// level 10
assign po2034 = w11432;// level 10
assign po2035 = ~w14430;// level 9
assign po2036 = w15913;// level 8
assign po2037 = w15591;// level 6
assign po2038 = w17589;// level 6
assign po2039 = w15487;// level 6
assign po2040 = w1842;// level 6
assign po2041 = w14218;// level 6
assign po2042 = w767;// level 6
assign po2043 = w13197;// level 6
assign po2044 = w8465;// level 6
assign po2045 = w6636;// level 6
assign po2046 = w14337;// level 6
assign po2047 = w2698;// level 6
assign po2048 = w7246;// level 6
assign po2049 = w16038;// level 6
assign po2050 = w14580;// level 6
assign po2051 = w16563;// level 6
assign po2052 = w4368;// level 6
assign po2053 = w3531;// level 6
assign po2054 = w3583;// level 10
assign po2055 = ~w8473;// level 8
assign po2056 = w13083;// level 10
assign po2057 = w11603;// level 8
assign po2058 = w8036;// level 9
assign po2059 = w892;// level 10
assign po2060 = w1448;// level 10
assign po2061 = w12213;// level 10
assign po2062 = w4046;// level 6
assign po2063 = w2210;// level 6
assign po2064 = w4813;// level 6
assign po2065 = w4996;// level 6
assign po2066 = w14107;// level 6
assign po2067 = w5932;// level 10
assign po2068 = w938;// level 6
assign po2069 = w14022;// level 6
assign po2070 = w17030;// level 6
assign po2071 = w1987;// level 6
assign po2072 = w17988;// level 6
assign po2073 = w12619;// level 6
assign po2074 = w11526;// level 6
assign po2075 = w15870;// level 6
assign po2076 = w641;// level 6
assign po2077 = w11423;// level 6
assign po2078 = w17897;// level 10
assign po2079 = ~w6608;// level 7
assign po2080 = w15154;// level 10
assign po2081 = w16585;// level 9
assign po2082 = w79;// level 14
assign po2083 = w7506;// level 14
assign po2084 = w983;// level 14
assign po2085 = w1961;// level 15
assign po2086 = w4036;// level 15
assign po2087 = w1412;// level 15
assign po2088 = w9175;// level 14
assign po2089 = w10395;// level 15
assign po2090 = w7979;// level 14
assign po2091 = w4569;// level 15
assign po2092 = w5579;// level 14
assign po2093 = w8586;// level 14
assign po2094 = w13855;// level 14
assign po2095 = w2548;// level 14
assign po2096 = w15251;// level 14
assign po2097 = w9874;// level 14
assign po2098 = w647;// level 13
assign po2099 = w5431;// level 14
assign po2100 = w14786;// level 6
assign po2101 = w1587;// level 13
assign po2102 = w5434;// level 14
assign po2103 = w3247;// level 14
assign po2104 = w2716;// level 15
assign po2105 = w18168;// level 13
assign po2106 = w9285;// level 14
assign po2107 = w7930;// level 14
assign po2108 = w14220;// level 14
assign po2109 = w3037;// level 14
assign po2110 = w9679;// level 14
assign po2111 = w10506;// level 14
assign po2112 = w10708;// level 14
assign po2113 = w8697;// level 13
assign po2114 = w18237;// level 14
assign po2115 = w5157;// level 14
assign po2116 = w704;// level 14
assign po2117 = w12379;// level 12
assign po2118 = w6911;// level 14
assign po2119 = w14570;// level 12
assign po2120 = w16935;// level 14
assign po2121 = w4056;// level 14
assign po2122 = w4993;// level 13
assign po2123 = w9115;// level 14
assign po2124 = w1080;// level 14
assign po2125 = w5713;// level 13
assign po2126 = w7108;// level 13
assign po2127 = w15655;// level 14
assign po2128 = w985;// level 13
assign po2129 = w9778;// level 14
assign po2130 = w274;// level 14
assign po2131 = w5469;// level 13
assign po2132 = w13005;// level 14
assign po2133 = w2295;// level 14
assign po2134 = w10075;// level 14
assign po2135 = w16291;// level 14
assign po2136 = w13793;// level 14
assign po2137 = w2964;// level 14
assign po2138 = w18288;// level 14
assign po2139 = w16500;// level 14
assign po2140 = w9638;// level 14
assign po2141 = w666;// level 14
assign po2142 = w687;// level 15
assign po2143 = ~w16785;// level 9
assign po2144 = w17859;// level 6
assign po2145 = w9776;// level 6
assign po2146 = w4136;// level 6
assign po2147 = w9531;// level 9
assign po2148 = ~w5554;// level 8
assign po2149 = w14047;// level 9
assign po2150 = ~w15913;// level 8
assign po2151 = w3542;// level 10
assign po2152 = w16421;// level 10
assign po2153 = w3738;// level 9
assign po2154 = w13516;// level 10
assign po2155 = w17198;// level 10
assign po2156 = w9798;// level 10
assign po2157 = w4143;// level 10
assign po2158 = w8473;// level 8
assign po2159 = ~w6577;// level 13
assign po2160 = w4334;// level 10
assign po2161 = w8140;// level 12
assign po2162 = w7733;// level 10
assign po2163 = w17448;// level 13
assign po2164 = w9480;// level 14
assign po2165 = w16009;// level 13
assign po2166 = w2918;// level 14
assign po2167 = w17590;// level 14
assign po2168 = w13495;// level 13
assign po2169 = w13553;// level 14
assign po2170 = w9651;// level 14
assign po2171 = w16215;// level 14
assign po2172 = w7674;// level 14
assign po2173 = w1382;// level 14
assign po2174 = w8656;// level 13
assign po2175 = w11871;// level 14
assign po2176 = w10651;// level 14
assign po2177 = w18550;// level 14
assign po2178 = w1226;// level 14
assign po2179 = w6411;// level 14
assign po2180 = w11157;// level 14
assign po2181 = w6037;// level 14
assign po2182 = w9668;// level 13
assign po2183 = w13578;// level 13
assign po2184 = w157;// level 13
assign po2185 = w7539;// level 14
assign po2186 = w5795;// level 13
assign po2187 = w17109;// level 14
assign po2188 = w1889;// level 14
assign po2189 = w15334;// level 14
assign po2190 = w11409;// level 14
assign po2191 = w10808;// level 14
assign po2192 = w17887;// level 14
assign po2193 = w1405;// level 14
assign po2194 = w16745;// level 14
assign po2195 = w5464;// level 14
assign po2196 = w12704;// level 14
assign po2197 = w13859;// level 14
assign po2198 = w12007;// level 13
assign po2199 = w6752;// level 13
assign po2200 = w10443;// level 13
assign po2201 = w15286;// level 14
assign po2202 = w1404;// level 14
assign po2203 = w5311;// level 13
assign po2204 = w11256;// level 14
assign po2205 = w10146;// level 14
assign po2206 = w11878;// level 14
assign po2207 = w18595;// level 14
assign po2208 = w8510;// level 14
assign po2209 = w8685;// level 14
assign po2210 = w5282;// level 14
assign po2211 = w12517;// level 14
assign po2212 = w13824;// level 14
assign po2213 = w736;// level 14
assign po2214 = w13245;// level 14
assign po2215 = w7179;// level 13
assign po2216 = w7287;// level 13
assign po2217 = w1676;// level 13
assign po2218 = w14895;// level 14
assign po2219 = w12529;// level 13
assign po2220 = w522;// level 14
assign po2221 = w12541;// level 14
assign po2222 = w9942;// level 14
assign po2223 = w8953;// level 14
assign po2224 = w12709;// level 14
assign po2225 = w8348;// level 13
assign po2226 = w8758;// level 14
assign po2227 = w12117;// level 14
assign po2228 = w9686;// level 14
assign po2229 = w1621;// level 14
assign po2230 = w13935;// level 14
assign po2231 = w5331;// level 14
assign po2232 = w14315;// level 14
assign po2233 = w6296;// level 14
assign po2234 = w12457;// level 14
assign po2235 = w6227;// level 14
assign po2236 = w7316;// level 13
assign po2237 = w17613;// level 13
assign po2238 = w16816;// level 14
assign po2239 = w7148;// level 13
assign po2240 = w8574;// level 14
assign po2241 = w16536;// level 14
assign po2242 = w17165;// level 14
assign po2243 = w18322;// level 14
assign po2244 = w13573;// level 14
assign po2245 = w7962;// level 14
assign po2246 = w3344;// level 14
assign po2247 = w262;// level 14
assign po2248 = w5356;// level 12
assign po2249 = w15881;// level 13
assign po2250 = w15796;// level 13
assign po2251 = w14477;// level 13
assign po2252 = w9522;// level 13
assign po2253 = w13527;// level 13
assign po2254 = w9866;// level 13
assign po2255 = w9718;// level 13
assign po2256 = w13773;// level 13
assign po2257 = w16717;// level 13
assign po2258 = w9755;// level 13
assign po2259 = w9518;// level 13
assign po2260 = w2367;// level 13
assign po2261 = w18176;// level 14
assign po2262 = w10817;// level 13
assign po2263 = w6999;// level 13
assign po2264 = w8471;// level 14
assign po2265 = w695;// level 13
assign po2266 = w11587;// level 14
assign po2267 = w7751;// level 14
assign po2268 = w526;// level 13
assign po2269 = w8317;// level 14
assign po2270 = w12948;// level 14
assign po2271 = w17690;// level 14
assign po2272 = w14869;// level 14
assign po2273 = w8151;// level 14
assign po2274 = w1760;// level 14
assign po2275 = w12644;// level 13
assign po2276 = w8506;// level 14
assign po2277 = w3084;// level 14
assign po2278 = w119;// level 14
assign po2279 = w9870;// level 14
assign po2280 = w15950;// level 14
assign po2281 = w12982;// level 14
assign po2282 = w13152;// level 14
assign po2283 = w11315;// level 13
assign po2284 = w3822;// level 13
assign po2285 = w15975;// level 13
assign po2286 = w7754;// level 14
assign po2287 = w11044;// level 14
assign po2288 = w17166;// level 13
assign po2289 = w3397;// level 14
assign po2290 = w5007;// level 14
assign po2291 = w6800;// level 14
assign po2292 = w1358;// level 14
assign po2293 = w8152;// level 14
assign po2294 = w8335;// level 14
assign po2295 = w4404;// level 14
assign po2296 = w11994;// level 14
assign po2297 = w11651;// level 14
assign po2298 = w5506;// level 14
assign po2299 = w5412;// level 14
assign po2300 = w14340;// level 14
assign po2301 = w4781;// level 14
assign po2302 = w6392;// level 13
assign po2303 = w14115;// level 14
assign po2304 = w8157;// level 14
assign po2305 = w4863;// level 13
assign po2306 = w10007;// level 14
assign po2307 = w263;// level 14
assign po2308 = w3204;// level 14
assign po2309 = w9404;// level 14
assign po2310 = w5241;// level 13
assign po2311 = w17013;// level 14
assign po2312 = w4900;// level 13
assign po2313 = w17356;// level 14
assign po2314 = w15257;// level 14
assign po2315 = w4216;// level 14
assign po2316 = w12176;// level 14
assign po2317 = w5789;// level 14
assign po2318 = w2676;// level 13
assign po2319 = w16006;// level 14
assign po2320 = w12177;// level 14
assign po2321 = w9898;// level 14
assign po2322 = w3495;// level 14
assign po2323 = w12142;// level 15
assign po2324 = w10983;// level 15
assign po2325 = w4;// level 15
assign po2326 = w11880;// level 15
assign po2327 = w10234;// level 15
assign po2328 = w7461;// level 15
assign po2329 = w15247;// level 15
assign po2330 = w10326;// level 15
assign po2331 = w16384;// level 15
assign po2332 = w5709;// level 15
assign po2333 = w3112;// level 10
assign po2334 = w12725;// level 10
assign po2335 = w14083;// level 12
assign po2336 = w1395;// level 13
assign po2337 = w16996;// level 14
assign po2338 = w4184;// level 15
assign po2339 = w8522;// level 10
assign po2340 = ~w15853;// level 8
assign po2341 = w13420;// level 13
assign po2342 = w16407;// level 13
assign po2343 = w5478;// level 14
assign po2344 = w10934;// level 14
assign po2345 = w3108;// level 14
assign po2346 = w12034;// level 14
assign po2347 = w17962;// level 14
assign po2348 = w9179;// level 14
assign po2349 = w17707;// level 14
assign po2350 = w10014;// level 14
assign po2351 = w12160;// level 15
assign po2352 = w10789;// level 15
assign po2353 = w895;// level 15
assign po2354 = w16524;// level 15
assign po2355 = w11136;// level 14
assign po2356 = w3814;// level 15
assign po2357 = w17101;// level 15
assign po2358 = w13968;// level 15
assign po2359 = w13650;// level 15
assign po2360 = w22;// level 15
assign po2361 = w17547;// level 13
assign po2362 = w16076;// level 14
assign po2363 = w2102;// level 14
assign po2364 = w6338;// level 14
assign po2365 = w14916;// level 14
assign po2366 = w3934;// level 14
assign po2367 = w6975;// level 14
assign po2368 = w10049;// level 14
assign po2369 = w17012;// level 15
assign po2370 = w16907;// level 15
assign po2371 = w777;// level 15
assign po2372 = w14424;// level 14
assign po2373 = w5314;// level 15
assign po2374 = w7024;// level 14
assign po2375 = w12516;// level 15
assign po2376 = w356;// level 15
assign po2377 = w4149;// level 14
assign po2378 = w16657;// level 13
assign po2379 = w16574;// level 13
assign po2380 = w18134;// level 15
assign po2381 = w10229;// level 15
assign po2382 = w12145;// level 15
assign po2383 = w9696;// level 15
assign po2384 = w5948;// level 15
assign po2385 = w14972;// level 15
assign po2386 = w18316;// level 14
assign po2387 = w14192;// level 15
assign po2388 = w3139;// level 13
assign po2389 = w13784;// level 14
assign po2390 = w13052;// level 14
assign po2391 = w8809;// level 14
assign po2392 = w3602;// level 14
assign po2393 = w5893;// level 13
assign po2394 = w613;// level 14
assign po2395 = w9879;// level 14
assign po2396 = w7064;// level 14
assign po2397 = w8312;// level 14
assign po2398 = w15559;// level 14
assign po2399 = w16293;// level 14
assign po2400 = w12693;// level 14
assign po2401 = w16124;// level 13
assign po2402 = w10449;// level 14
assign po2403 = w4696;// level 13
assign po2404 = w6807;// level 13
assign po2405 = w2351;// level 13
assign po2406 = w11969;// level 14
assign po2407 = w17161;// level 14
assign po2408 = w17275;// level 14
assign po2409 = w16879;// level 13
assign po2410 = w14581;// level 13
assign po2411 = w18121;// level 13
assign po2412 = w17866;// level 14
assign po2413 = w1732;// level 14
assign po2414 = w13286;// level 13
assign po2415 = w2816;// level 14
assign po2416 = w10179;// level 13
assign po2417 = w7279;// level 14
assign po2418 = w1176;// level 14
assign po2419 = w2627;// level 14
assign po2420 = w10500;// level 13
assign po2421 = w2493;// level 14
assign po2422 = w14871;// level 14
assign po2423 = w17424;// level 14
assign po2424 = w8365;// level 14
assign po2425 = w7546;// level 14
assign po2426 = w1665;// level 14
assign po2427 = w8984;// level 14
assign po2428 = w9835;// level 10
assign po2429 = w17984;// level 14
assign po2430 = w4970;// level 14
assign po2431 = w13034;// level 15
assign po2432 = w9816;// level 15
assign po2433 = w5032;// level 15
assign po2434 = w8100;// level 15
assign po2435 = w2409;// level 15
assign po2436 = w5096;// level 15
assign po2437 = w18376;// level 15
assign po2438 = w15014;// level 15
assign po2439 = w17348;// level 15
assign po2440 = w3554;// level 14
assign po2441 = w10062;// level 15
assign po2442 = w13237;// level 15
assign po2443 = w14573;// level 14
assign po2444 = w8311;// level 14
assign po2445 = w3914;// level 14
assign po2446 = w17875;// level 13
assign po2447 = w10636;// level 12
assign po2448 = w12681;// level 12
assign po2449 = w9109;// level 13
assign po2450 = w9566;// level 14
assign po2451 = w4457;// level 14
assign po2452 = w17738;// level 14
assign po2453 = w11187;// level 14
assign po2454 = w18;// level 15
assign po2455 = w6329;// level 14
assign po2456 = w14363;// level 15
assign po2457 = w7135;// level 15
assign po2458 = w18504;// level 14
assign po2459 = w11303;// level 15
assign po2460 = w6955;// level 10
assign po2461 = ~w11444;// level 9
assign po2462 = w6121;// level 15
assign po2463 = w14268;// level 14
assign po2464 = w7336;// level 13
assign po2465 = w8355;// level 8
assign po2466 = w7747;// level 13
assign po2467 = w5203;// level 14
assign po2468 = w8009;// level 10
assign po2469 = w4189;// level 10
assign po2470 = w9772;// level 7
assign po2471 = w9478;// level 8
assign po2472 = w4053;// level 15
assign po2473 = w12611;// level 13
assign po2474 = w8729;// level 14
assign po2475 = w18204;// level 13
assign po2476 = w2135;// level 13
assign po2477 = w18076;// level 13
assign po2478 = w10063;// level 14
assign po2479 = w14898;// level 15
assign po2480 = w12052;// level 14
assign po2481 = w10974;// level 14
assign po2482 = w6412;// level 14
assign po2483 = w14681;// level 14
assign po2484 = w11488;// level 14
assign po2485 = w6238;// level 14
assign po2486 = w15070;// level 14
assign po2487 = w1190;// level 14
assign po2488 = w17853;// level 14
assign po2489 = w18261;// level 14
assign po2490 = w521;// level 14
assign po2491 = w6991;// level 14
assign po2492 = w17194;// level 14
assign po2493 = w1796;// level 14
assign po2494 = w3288;// level 15
assign po2495 = w12960;// level 14
assign po2496 = w2098;// level 13
assign po2497 = w9583;// level 14
assign po2498 = w1327;// level 14
assign po2499 = w8039;// level 14
assign po2500 = w7159;// level 14
assign po2501 = w6494;// level 13
assign po2502 = w5844;// level 14
assign po2503 = w420;// level 14
assign po2504 = w245;// level 14
assign po2505 = w3418;// level 14
assign po2506 = w16113;// level 14
assign po2507 = w13000;// level 14
assign po2508 = w10570;// level 14
assign po2509 = w7354;// level 15
assign po2510 = w16167;// level 13
assign po2511 = w10508;// level 14
assign po2512 = w15171;// level 14
assign po2513 = w731;// level 13
assign po2514 = w793;// level 13
assign po2515 = w1159;// level 13
assign po2516 = w3127;// level 15
assign po2517 = w1617;// level 14
assign po2518 = w17283;// level 13
assign po2519 = w16792;// level 14
assign po2520 = w7432;// level 14
assign po2521 = w2527;// level 13
assign po2522 = w15588;// level 14
assign po2523 = w8608;// level 14
assign po2524 = w6948;// level 14
assign po2525 = w13694;// level 13
assign po2526 = w7942;// level 14
assign po2527 = w2939;// level 14
assign po2528 = w14398;// level 13
assign po2529 = w29;// level 14
assign po2530 = w16567;// level 13
assign po2531 = w2308;// level 12
assign po2532 = w12010;// level 13
assign po2533 = w2012;// level 14
assign po2534 = ~w8158;// level 10
assign po2535 = w14470;// level 14
assign po2536 = w14836;// level 14
assign po2537 = w15153;// level 13
assign po2538 = w295;// level 14
assign po2539 = w4076;// level 14
assign po2540 = w4371;// level 15
assign po2541 = w12404;// level 13
assign po2542 = w12268;// level 14
assign po2543 = w18001;// level 13
assign po2544 = w8791;// level 14
assign po2545 = w6904;// level 13
assign po2546 = w12495;// level 14
assign po2547 = w6401;// level 13
assign po2548 = w11777;// level 13
assign po2549 = w2872;// level 14
assign po2550 = w6313;// level 15
assign po2551 = w10854;// level 13
assign po2552 = w3855;// level 14
assign po2553 = w7119;// level 13
assign po2554 = w2746;// level 13
assign po2555 = w5264;// level 14
assign po2556 = w17708;// level 14
assign po2557 = w663;// level 13
assign po2558 = w15755;// level 14
assign po2559 = w13153;// level 15
assign po2560 = w2897;// level 12
assign po2561 = w1102;// level 14
assign po2562 = w6122;// level 14
assign po2563 = w3014;// level 13
assign po2564 = w4047;// level 14
assign po2565 = w6707;// level 14
assign po2566 = w4917;// level 12
assign po2567 = w12904;// level 14
assign po2568 = w17049;// level 13
assign po2569 = w6705;// level 14
assign po2570 = w681;// level 15
assign po2571 = w17659;// level 14
assign po2572 = w12967;// level 14
assign po2573 = w2967;// level 15
assign po2574 = w2103;// level 15
assign po2575 = w17711;// level 14
assign po2576 = w10372;// level 13
assign po2577 = w18536;// level 15
assign po2578 = w12916;// level 14
assign po2579 = w9953;// level 13
assign po2580 = w3617;// level 15
assign po2581 = w16070;// level 14
assign po2582 = w10173;// level 14
assign po2583 = w5987;// level 14
assign po2584 = w14947;// level 15
assign po2585 = w7321;// level 14
assign po2586 = w12759;// level 14
assign po2587 = w9012;// level 15
assign po2588 = w15854;// level 15
assign po2589 = w7590;// level 14
assign po2590 = w12459;// level 14
assign po2591 = w5837;// level 14
assign po2592 = w15368;// level 15
assign po2593 = w9659;// level 13
assign po2594 = w9611;// level 14
assign po2595 = w13615;// level 15
assign po2596 = w3025;// level 15
assign po2597 = w8742;// level 14
assign po2598 = w8526;// level 13
assign po2599 = w16252;// level 14
assign po2600 = w11457;// level 14
assign po2601 = w1420;// level 14
assign po2602 = w6970;// level 15
assign po2603 = w2025;// level 14
assign po2604 = w5231;// level 14
assign po2605 = w16084;// level 14
assign po2606 = w17805;// level 10
assign po2607 = w14623;// level 14
assign po2608 = w8025;// level 10
assign po2609 = w17592;// level 15
assign po2610 = w8743;// level 9
assign po2611 = w18150;// level 14
assign po2612 = w935;// level 15
assign po2613 = w17739;// level 14
assign po2614 = w17811;// level 14
assign po2615 = w730;// level 13
assign po2616 = w12645;// level 15
assign po2617 = w1506;// level 15
assign po2618 = w7849;// level 15
assign po2619 = w10144;// level 15
assign po2620 = w13565;// level 15
assign po2621 = w655;// level 15
assign po2622 = w8553;// level 15
assign po2623 = w8726;// level 15
assign po2624 = w3028;// level 15
assign po2625 = w4551;// level 15
assign po2626 = w18146;// level 15
assign po2627 = w8581;// level 15
assign po2628 = w8981;// level 15
assign po2629 = w4296;// level 14
assign po2630 = w17518;// level 15
assign po2631 = w2948;// level 15
assign po2632 = w16253;// level 15
assign po2633 = w3324;// level 14
assign po2634 = w14934;// level 14
assign po2635 = ~w9319;// level 7
assign po2636 = w7899;// level 14
assign po2637 = w11787;// level 7
assign po2638 = w2595;// level 15
assign po2639 = ~w10562;// level 7
assign po2640 = w9773;// level 15
assign po2641 = w17193;// level 10
assign po2642 = w10965;// level 13
assign po2643 = w12228;// level 15
assign po2644 = w14033;// level 15
assign po2645 = w6742;// level 14
assign po2646 = w3414;// level 15
assign po2647 = w5980;// level 15
assign po2648 = w8325;// level 13
assign po2649 = w5537;// level 13
assign po2650 = w13635;// level 14
assign po2651 = w9861;// level 15
assign po2652 = w1679;// level 14
assign po2653 = ~w8449;// level 9
assign po2654 = ~w5999;// level 9
assign po2655 = w15574;// level 9
assign po2656 = ~w16994;// level 9
assign po2657 = ~w6099;// level 9
assign po2658 = w6967;// level 9
assign po2659 = ~w11404;// level 8
assign po2660 = ~w4392;// level 7
assign po2661 = w7761;// level 10
assign po2662 = ~w5909;// level 9
assign po2663 = ~w6949;// level 9
assign po2664 = w14525;// level 9
assign po2665 = w3892;// level 10
assign po2666 = w8077;// level 9
assign po2667 = w14549;// level 8
assign po2668 = w1096;// level 10
assign po2669 = w9270;// level 10
assign po2670 = ~w3915;// level 9
assign po2671 = w9795;// level 9
assign po2672 = w2384;// level 9
assign po2673 = ~w7737;// level 9
assign po2674 = w9372;// level 10
assign po2675 = ~w14906;// level 9
assign po2676 = ~w6909;// level 9
assign po2677 = ~w13943;// level 9
assign po2678 = w6413;// level 10
assign po2679 = ~w2186;// level 9
assign po2680 = ~w1339;// level 9
assign po2681 = w10629;// level 10
assign po2682 = ~w4275;// level 9
assign po2683 = w17533;// level 9
assign po2684 = w12899;// level 10
assign po2685 = w13643;// level 10
assign po2686 = w5619;// level 10
assign po2687 = w15995;// level 10
assign po2688 = w45;// level 10
assign po2689 = w4536;// level 8
assign po2690 = w9363;// level 10
assign po2691 = w12410;// level 10
assign po2692 = ~w3640;// level 9
assign po2693 = w1831;// level 8
assign po2694 = w16763;// level 7
assign po2695 = w5990;// level 7
assign po2696 = w11877;// level 8
assign po2697 = w3079;// level 8
assign po2698 = w15888;// level 8
assign po2699 = w3257;// level 10
assign po2700 = w8651;// level 10
assign po2701 = ~w16882;// level 8
assign po2702 = ~w8512;// level 8
assign po2703 = ~w1088;// level 8
assign po2704 = ~w12245;// level 8
assign po2705 = ~w15065;// level 8
assign po2706 = ~w8082;// level 8
assign po2707 = ~w16242;// level 8
assign po2708 = ~w13597;// level 8
assign po2709 = ~w260;// level 8
assign po2710 = ~w13095;// level 8
assign po2711 = ~w17221;// level 8
assign po2712 = ~w74;// level 8
assign po2713 = ~w15054;// level 8
assign po2714 = ~w13542;// level 8
assign po2715 = ~w12883;// level 8
assign po2716 = ~w16180;// level 8
assign po2717 = ~w13799;// level 8
assign po2718 = ~w6531;// level 8
assign po2719 = ~w15093;// level 8
assign po2720 = ~w17260;// level 8
assign po2721 = ~w12797;// level 8
assign po2722 = ~w8839;// level 8
assign po2723 = ~w5101;// level 8
assign po2724 = ~w10472;// level 8
assign po2725 = ~w6191;// level 8
assign po2726 = ~w46;// level 8
assign po2727 = ~w7357;// level 9
assign po2728 = ~w11125;// level 9
assign po2729 = ~w6353;// level 9
assign po2730 = ~w4848;// level 9
assign po2731 = ~w16896;// level 9
assign po2732 = ~w11257;// level 9
assign po2733 = ~w6384;// level 9
assign po2734 = ~w10496;// level 9
assign po2735 = ~w9727;// level 9
assign po2736 = ~w14509;// level 9
assign po2737 = ~w4538;// level 9
assign po2738 = ~w1811;// level 9
assign po2739 = ~w2704;// level 9
assign po2740 = ~w3622;// level 9
assign po2741 = ~w12468;// level 9
assign po2742 = ~w6053;// level 9
assign po2743 = ~w8223;// level 9
assign po2744 = ~w10626;// level 9
assign po2745 = ~w17930;// level 9
assign po2746 = ~w9271;// level 9
assign po2747 = ~w1511;// level 9
assign po2748 = ~w5155;// level 9
assign po2749 = ~w16255;// level 9
assign po2750 = ~w11401;// level 9
assign po2751 = ~w12172;// level 9
assign po2752 = ~w3073;// level 9
assign po2753 = ~w11995;// level 9
assign po2754 = ~w3030;// level 9
assign po2755 = ~w12974;// level 9
assign po2756 = ~w13512;// level 9
assign po2757 = ~w14320;// level 9
assign po2758 = ~w15124;// level 9
assign po2759 = ~w12249;// level 9
assign po2760 = ~w4586;// level 9
assign po2761 = ~w16788;// level 9
assign po2762 = ~w10706;// level 9
assign po2763 = ~w7771;// level 9
assign po2764 = ~w16587;// level 9
assign po2765 = ~w16740;// level 9
assign po2766 = ~w12184;// level 9
assign po2767 = w18086;// level 9
assign po2768 = w15453;// level 11
assign po2769 = w4640;// level 10
assign po2770 = w9602;// level 10
assign po2771 = w11736;// level 10
assign po2772 = w14890;// level 10
assign po2773 = w1851;// level 10
assign po2774 = w6942;// level 10
assign po2775 = w2850;// level 10
assign po2776 = w6566;// level 10
assign po2777 = w7587;// level 10
assign po2778 = w12339;// level 10
assign po2779 = w16570;// level 10
assign po2780 = w11379;// level 8
assign po2781 = w15969;// level 8
assign po2782 = w1091;// level 8
assign po2783 = w2524;// level 8
assign po2784 = w7139;// level 8
assign po2785 = w14053;// level 8
assign po2786 = w3189;// level 8
assign po2787 = w11680;// level 8
assign po2788 = w11548;// level 8
assign po2789 = w1514;// level 8
assign po2790 = w9777;// level 8
assign po2791 = w5584;// level 8
assign po2792 = w2854;// level 8
assign po2793 = w14734;// level 8
assign po2794 = w12751;// level 10
assign po2795 = w9290;// level 10
assign po2796 = w2686;// level 10
assign po2797 = w9880;// level 10
assign po2798 = w4808;// level 10
assign po2799 = w10083;// level 10
assign po2800 = w13559;// level 10
assign po2801 = w15787;// level 10
assign po2802 = w12530;// level 10
assign po2803 = w6572;// level 10
assign po2804 = w11353;// level 8
assign po2805 = w15258;// level 10
assign po2806 = w944;// level 10
assign po2807 = w638;// level 10
assign po2808 = w2507;// level 10
assign po2809 = w7563;// level 10
assign po2810 = w11012;// level 10
assign po2811 = w8778;// level 10
assign po2812 = w6658;// level 10
assign po2813 = w10637;// level 10
assign po2814 = w16933;// level 10
assign po2815 = w5149;// level 10
assign po2816 = w3793;// level 8
assign po2817 = w8570;// level 10
assign po2818 = w4171;// level 8
assign po2819 = w1188;// level 10
assign po2820 = w17046;// level 10
assign po2821 = w8282;// level 10
assign po2822 = w17557;// level 10
assign po2823 = w11253;// level 10
assign po2824 = w9386;// level 10
assign po2825 = w2156;// level 10
assign po2826 = w11566;// level 10
assign po2827 = w1074;// level 10
assign po2828 = w2175;// level 9
assign po2829 = w4606;// level 9
assign po2830 = w16731;// level 9
assign po2831 = w8209;// level 9
assign po2832 = w11895;// level 9
assign po2833 = w14822;// level 9
assign po2834 = w5637;// level 9
assign po2835 = w14130;// level 9
assign po2836 = w6420;// level 9
assign po2837 = w13259;// level 9
assign po2838 = w9283;// level 9
assign po2839 = w2349;// level 10
assign po2840 = w881;// level 10
assign po2841 = w4742;// level 10
assign po2842 = w11330;// level 10
assign po2843 = w6989;// level 10
assign po2844 = w1751;// level 10
assign po2845 = w2190;// level 10
assign po2846 = w2391;// level 10
assign po2847 = w12134;// level 10
assign po2848 = w9276;// level 10
assign po2849 = w4570;// level 10
assign po2850 = w17112;// level 10
assign po2851 = w1211;// level 10
assign po2852 = w16125;// level 10
assign po2853 = w16818;// level 10
assign po2854 = w15416;// level 10
assign po2855 = w14077;// level 10
assign po2856 = w8397;// level 10
assign po2857 = w14034;// level 10
assign po2858 = w2343;// level 10
assign po2859 = w14774;// level 9
assign po2860 = w14740;// level 9
assign po2861 = w1398;// level 10
assign po2862 = w9610;// level 10
assign po2863 = w14002;// level 10
assign po2864 = w15397;// level 8
assign po2865 = w8872;// level 9
assign po2866 = w12498;// level 10
assign po2867 = w1257;// level 10
assign po2868 = w18307;// level 10
assign po2869 = w5906;// level 10
assign po2870 = w18560;// level 10
assign po2871 = w8833;// level 10
assign po2872 = w11145;// level 10
assign po2873 = w3665;// level 10
assign po2874 = w392;// level 10
assign po2875 = w5919;// level 10
assign po2876 = w6031;// level 10
assign po2877 = w11052;// level 10
assign po2878 = w18293;// level 10
assign po2879 = ~w14365;// level 9
assign po2880 = w886;// level 8
assign po2881 = w4889;// level 10
assign po2882 = w5342;// level 10
assign po2883 = w850;// level 10
assign po2884 = w6178;// level 10
assign po2885 = w8776;// level 10
assign po2886 = w538;// level 8
assign po2887 = w966;// level 10
assign po2888 = w6201;// level 10
assign po2889 = w9455;// level 10
assign po2890 = w15385;// level 9
assign po2891 = w9769;// level 10
assign po2892 = w9008;// level 8
assign po2893 = w7160;// level 10
assign po2894 = w278;// level 10
assign po2895 = w5910;// level 10
assign po2896 = w2768;// level 10
assign po2897 = w6063;// level 10
assign po2898 = w11771;// level 10
assign po2899 = w17648;// level 10
assign po2900 = w17006;// level 8
assign po2901 = w6416;// level 8
assign po2902 = w10650;// level 8
assign po2903 = w10711;// level 8
assign po2904 = w3716;// level 10
assign po2905 = w11562;// level 8
assign po2906 = w11535;// level 8
assign po2907 = ~w13482;// level 9
assign po2908 = w3867;// level 8
assign po2909 = w3077;// level 8
assign po2910 = ~w10414;// level 9
assign po2911 = ~w3092;// level 9
assign po2912 = ~w13817;// level 9
assign po2913 = w12859;// level 9
assign po2914 = w14108;// level 10
assign po2915 = w15046;// level 9
assign po2916 = w9454;// level 10
assign po2917 = w4073;// level 10
assign po2918 = w17780;// level 10
assign po2919 = w5461;// level 10
assign po2920 = w14359;// level 10
assign po2921 = w13976;// level 10
assign po2922 = w13698;// level 8
assign po2923 = ~w2113;// level 9
assign po2924 = w6335;// level 10
assign po2925 = w4159;// level 10
assign po2926 = ~w2452;// level 8
assign po2927 = w1848;// level 10
assign po2928 = w109;// level 10
assign po2929 = w66;// level 9
assign po2930 = w16532;// level 10
assign po2931 = ~w7313;// level 7
assign po2932 = ~w18443;// level 9
assign po2933 = w7105;// level 10
assign po2934 = ~w13409;// level 8
assign po2935 = ~w5529;// level 8
assign po2936 = ~w11026;// level 8
assign po2937 = w2339;// level 10
assign po2938 = w5929;// level 10
assign po2939 = ~w15759;// level 8
assign po2940 = ~w10836;// level 8
assign po2941 = ~w8779;// level 8
assign po2942 = w9881;// level 10
assign po2943 = w1788;// level 10
assign po2944 = w13510;// level 10
assign po2945 = w13067;// level 10
assign po2946 = w10420;// level 10
assign po2947 = w18401;// level 10
assign po2948 = w8404;// level 10
assign po2949 = w18246;// level 10
assign po2950 = w13338;// level 9
assign po2951 = w2255;// level 9
assign po2952 = w11555;// level 10
assign po2953 = ~w2837;// level 8
assign po2954 = w13119;// level 10
assign po2955 = w3191;// level 10
assign po2956 = w11309;// level 10
assign po2957 = w17199;// level 10
assign po2958 = w16976;// level 8
assign po2959 = w10956;// level 10
assign po2960 = w4079;// level 10
assign po2961 = ~w419;// level 9
assign po2962 = w15098;// level 10
assign po2963 = w13076;// level 10
assign po2964 = w9542;// level 10
assign po2965 = w9889;// level 10
assign po2966 = w7833;// level 10
assign po2967 = w11794;// level 10
assign po2968 = w11715;// level 10
assign po2969 = ~w556;// level 8
assign po2970 = w12399;// level 9
assign po2971 = w17605;// level 9
assign po2972 = w4678;// level 10
assign po2973 = w1446;// level 10
assign po2974 = w11162;// level 10
assign po2975 = w13939;// level 10
assign po2976 = w10076;// level 10
assign po2977 = w939;// level 10
assign po2978 = w11968;// level 10
assign po2979 = w13293;// level 10
assign po2980 = w13634;// level 10
assign po2981 = w10879;// level 10
assign po2982 = w8972;// level 10
assign po2983 = w11631;// level 10
assign po2984 = w67;// level 10
assign po2985 = w6273;// level 10
assign po2986 = w11823;// level 9
assign po2987 = w873;// level 10
assign po2988 = w1178;// level 10
assign po2989 = w14506;// level 10
assign po2990 = w15294;// level 10
assign po2991 = w14358;// level 9
assign po2992 = ~w11503;// level 8
assign po2993 = ~w1119;// level 8
assign po2994 = w624;// level 9
assign po2995 = w11049;// level 10
assign po2996 = w13941;// level 10
assign po2997 = w6025;// level 9
assign po2998 = w18269;// level 10
assign po2999 = w7424;// level 10
assign po3000 = w12479;// level 10
assign po3001 = w1656;// level 10
assign po3002 = w10156;// level 10
assign po3003 = w11402;// level 10
assign po3004 = w10851;// level 10
assign po3005 = w13972;// level 8
assign po3006 = w3001;// level 10
assign po3007 = w7235;// level 10
assign po3008 = ~w4023;// level 8
assign po3009 = w5423;// level 10
assign po3010 = w7231;// level 10
assign po3011 = w9089;// level 10
assign po3012 = ~w10378;// level 8
assign po3013 = w16436;// level 10
assign po3014 = ~w13445;// level 8
assign po3015 = ~w5066;// level 8
assign po3016 = ~w11238;// level 8
assign po3017 = ~w503;// level 8
assign po3018 = w14646;// level 10
assign po3019 = ~w6174;// level 8
assign po3020 = w145;// level 8
assign po3021 = ~w16809;// level 8
assign po3022 = w13448;// level 8
assign po3023 = ~w1203;// level 8
assign po3024 = ~w10118;// level 8
assign po3025 = w7126;// level 8
assign po3026 = w52;// level 8
assign po3027 = ~w11492;// level 8
assign po3028 = ~w16701;// level 8
assign po3029 = w15105;// level 10
assign po3030 = ~w17841;// level 9
assign po3031 = w4390;// level 10
assign po3032 = ~w4830;// level 8
assign po3033 = ~w17772;// level 8
assign po3034 = w16889;// level 10
assign po3035 = ~w12367;// level 8
assign po3036 = ~w2480;// level 8
assign po3037 = ~w15678;// level 8
assign po3038 = ~w5449;// level 8
assign po3039 = ~w38;// level 8
assign po3040 = ~w10285;// level 8
assign po3041 = ~w9064;// level 8
assign po3042 = ~w5611;// level 8
assign po3043 = ~w10946;// level 8
assign po3044 = ~w4221;// level 8
assign po3045 = ~w11632;// level 8
assign po3046 = ~w6980;// level 8
assign po3047 = w15374;// level 8
assign po3048 = w11532;// level 9
assign po3049 = w17152;// level 10
assign po3050 = w18445;// level 10
assign po3051 = w9826;// level 10
assign po3052 = w719;// level 10
assign po3053 = w1839;// level 10
assign po3054 = w13437;// level 10
assign po3055 = w13848;// level 10
assign po3056 = w10619;// level 10
assign po3057 = w7555;// level 10
assign po3058 = ~w4260;// level 9
assign po3059 = ~w16227;// level 9
assign po3060 = w5427;// level 10
assign po3061 = w17285;// level 10
assign po3062 = ~w3290;// level 9
assign po3063 = ~w18004;// level 9
assign po3064 = w18513;// level 10
assign po3065 = w9845;// level 9
assign po3066 = w16066;// level 10
assign po3067 = w17002;// level 10
assign po3068 = ~w3737;// level 9
assign po3069 = ~w16256;// level 9
assign po3070 = w16985;// level 10
assign po3071 = w17542;// level 10
assign po3072 = w1592;// level 10
assign po3073 = w786;// level 9
assign po3074 = w11938;// level 10
assign po3075 = ~w9297;// level 9
assign po3076 = w5833;// level 10
assign po3077 = w9919;// level 10
assign po3078 = ~w7731;// level 9
assign po3079 = w5884;// level 10
assign po3080 = w17699;// level 8
assign po3081 = ~w8189;// level 8
assign po3082 = w8301;// level 8
assign po3083 = ~w5308;// level 6
assign po3084 = ~w4610;// level 8
assign po3085 = ~w17375;// level 9
assign po3086 = w16633;// level 5
assign po3087 = ~w9347;// level 6
assign po3088 = ~w11352;// level 9
assign po3089 = ~w6905;// level 10
assign po3090 = ~w7586;// level 10
assign po3091 = w3420;// level 7
assign po3092 = w13985;// level 6
assign po3093 = w16946;// level 6
assign po3094 = ~w15167;// level 4
assign po3095 = ~w13110;// level 9
assign po3096 = w10327;// level 7
assign po3097 = ~w16841;// level 8
assign po3098 = w4000;// level 7
assign po3099 = w643;// level 6
assign po3100 = w842;// level 10
assign po3101 = w3500;// level 10
assign po3102 = w5851;// level 10
assign po3103 = w2067;// level 10
assign po3104 = w6128;// level 9
assign po3105 = w7847;// level 10
assign po3106 = w16512;// level 10
assign po3107 = w12107;// level 8
assign po3108 = ~w13723;// level 7
assign po3109 = ~w10024;// level 7
assign po3110 = ~w585;// level 7
assign po3111 = ~w11661;// level 8
assign po3112 = ~w7852;// level 6
assign po3113 = ~w8280;// level 16
assign po3114 = w5632;// level 7
assign po3115 = ~w264;// level 6
assign po3116 = ~w17488;// level 7
assign po3117 = w1061;// level 5
assign po3118 = w8557;// level 5
assign po3119 = ~w3165;// level 7
assign po3120 = w7393;// level 7
assign po3121 = w13251;// level 16
assign po3122 = w960;// level 1
assign po3123 = ~w11929;// level 9
assign po3124 = w9172;// level 3
assign po3125 = ~w589;// level 7
assign po3126 = ~w15387;// level 6
assign po3127 = w4845;// level 9
assign po3128 = ~w8218;// level 7
assign po3129 = ~w1963;// level 6
assign po3130 = ~w5476;// level 7
assign po3131 = w18582;// level 14
assign po3132 = ~w18373;// level 6
assign po3133 = ~w11514;// level 6
assign po3134 = ~w12221;// level 6
assign po3135 = w18346;// level 4
assign po3136 = w13492;// level 13
assign po3137 = ~w6502;// level 6
assign po3138 = w7905;// level 2
assign po3139 = ~w14088;// level 4
assign po3140 = ~w2630;// level 4
assign po3141 = ~w1888;// level 4
assign po3142 = w2081;// level 4
assign po3143 = ~w5976;// level 4
assign po3144 = w18352;// level 12
assign po3145 = w370;// level 4
assign po3146 = w9432;// level 4
assign po3147 = w516;// level 10
assign po3148 = w6789;// level 15
assign po3149 = w14354;// level 5
assign po3150 = w7145;// level 2
assign po3151 = w11333;// level 9
assign po3152 = w782;// level 11
assign po3153 = w14127;// level 6
assign po3154 = ~w5297;// level 4
assign po3155 = ~w10441;// level 4
assign po3156 = ~w2021;// level 4
assign po3157 = w5924;// level 8
assign po3158 = ~w15304;// level 5
assign po3159 = pi3122;// level 0
assign po3160 = w14602;// level 5
assign po3161 = ~w7402;// level 4
assign po3162 = ~w4307;// level 4
assign po3163 = ~w5742;// level 3
assign po3164 = ~w17449;// level 4
assign po3165 = w7599;// level 4
assign po3166 = ~w15879;// level 4
assign po3167 = ~w15872;// level 4
assign po3168 = w16334;// level 3
assign po3169 = ~w9589;// level 4
assign po3170 = ~w14600;// level 4
assign po3171 = ~w928;// level 4
assign po3172 = w10070;// level 7
assign po3173 = w17927;// level 4
assign po3174 = ~w7309;// level 4
assign po3175 = ~w18223;// level 4
assign po3176 = w11468;// level 4
assign po3177 = ~w9910;// level 4
assign po3178 = ~w16848;// level 4
assign po3179 = ~w12735;// level 4
assign po3180 = ~w4622;// level 4
assign po3181 = ~w16757;// level 4
assign po3182 = ~w8827;// level 4
assign po3183 = ~w13599;// level 4
assign po3184 = ~w12777;// level 4
assign po3185 = ~w3205;// level 4
assign po3186 = ~w18038;// level 4
assign po3187 = ~w6008;// level 4
assign po3188 = ~w17041;// level 4
assign po3189 = ~w12861;// level 4
assign po3190 = w13998;// level 4
assign po3191 = ~w3095;// level 4
assign po3192 = w12968;// level 4
assign po3193 = ~w11384;// level 4
assign po3194 = w5380;// level 4
assign po3195 = ~w2713;// level 4
assign po3196 = ~w7379;// level 4
assign po3197 = ~w17025;// level 4
assign po3198 = ~w10979;// level 4
assign po3199 = ~w13291;// level 4
assign po3200 = ~w2234;// level 4
assign po3201 = w3832;// level 5
assign po3202 = ~w17318;// level 4
assign po3203 = ~w5886;// level 4
assign po3204 = ~w18402;// level 4
assign po3205 = ~w17066;// level 4
assign po3206 = ~w8477;// level 4
assign po3207 = ~w7964;// level 4
assign po3208 = w9121;// level 5
assign po3209 = ~w9576;// level 4
assign po3210 = ~w739;// level 4
assign po3211 = ~w12966;// level 4
assign po3212 = ~w4595;// level 4
assign po3213 = ~w3510;// level 4
assign po3214 = ~w1969;// level 4
assign po3215 = ~w15599;// level 4
assign po3216 = ~w4055;// level 4
assign po3217 = ~w10221;// level 4
assign po3218 = ~w2842;// level 4
assign po3219 = w12038;// level 2
assign po3220 = ~w11745;// level 4
assign po3221 = w4248;// level 2
assign po3222 = w7100;// level 2
assign po3223 = w15586;// level 2
assign po3224 = w9081;// level 2
assign po3225 = ~w909;// level 4
assign po3226 = ~w2664;// level 2
assign po3227 = ~w18060;// level 2
assign po3228 = ~w2766;// level 2
assign po3229 = w11073;// level 2
assign po3230 = w5963;// level 2
assign po3231 = w16375;// level 4
assign po3232 = w7540;// level 2
assign po3233 = w2670;// level 2
assign po3234 = w10098;// level 2
assign po3235 = w13952;// level 2
assign po3236 = w6084;// level 2
assign po3237 = ~w3443;// level 4
assign po3238 = w13899;// level 4
assign po3239 = ~w18500;// level 4
assign po3240 = ~w2085;// level 4
assign po3241 = ~w18070;// level 4
assign po3242 = ~w17437;// level 4
assign po3243 = ~w1410;// level 4
assign po3244 = w4123;// level 4
assign po3245 = w3408;// level 5
assign po3246 = ~w7784;// level 4
assign po3247 = ~w2968;// level 4
assign po3248 = ~w16202;// level 4
assign po3249 = ~w426;// level 4
assign po3250 = ~w13911;// level 4
assign po3251 = ~w16121;// level 4
assign po3252 = ~w13842;// level 4
assign po3253 = ~w1950;// level 4
assign po3254 = ~w11741;// level 4
assign po3255 = ~w3511;// level 4
assign po3256 = w2469;// level 3
assign po3257 = w13116;// level 2
assign po3258 = w424;// level 2
assign po3259 = w14479;// level 2
assign po3260 = w16852;// level 2
assign po3261 = w1068;// level 2
assign po3262 = w13936;// level 2
assign po3263 = w2296;// level 2
assign po3264 = ~w1004;// level 2
assign po3265 = w17345;// level 2
assign po3266 = ~w17872;// level 2
assign po3267 = ~w6601;// level 2
assign po3268 = ~w12170;// level 2
assign po3269 = ~w1356;// level 2
assign po3270 = w10337;// level 2
assign po3271 = w8130;// level 2
assign po3272 = w10107;// level 2
assign po3273 = w3551;// level 2
assign po3274 = w474;// level 2
assign po3275 = w6333;// level 2
assign po3276 = ~w620;// level 4
assign po3277 = w5207;// level 1
assign po3278 = ~w13330;// level 4
assign po3279 = ~w1309;// level 4
assign po3280 = ~w4028;// level 4
assign po3281 = ~w1549;// level 4
assign po3282 = ~w11584;// level 4
assign po3283 = ~w1785;// level 4
assign po3284 = ~w9709;// level 4
assign po3285 = ~w2213;// level 4
assign po3286 = ~w1558;// level 4
assign po3287 = ~w16491;// level 4
assign po3288 = ~w12453;// level 4
assign po3289 = ~w8424;// level 4
assign po3290 = ~w11008;// level 4
assign po3291 = w3449;// level 4
assign po3292 = ~w17949;// level 4
assign po3293 = w527;// level 5
assign po3294 = w7876;// level 4
assign po3295 = w9830;// level 1
assign po3296 = w2259;// level 3
assign po3297 = w2453;// level 4
assign po3298 = pi3140;// level 0
assign po3299 = pi3137;// level 0
assign po3300 = ~w7725;// level 3
assign po3301 = ~pi3207;// level 0
assign po3302 = w1913;// level 2
assign po3303 = pi3117;// level 0
assign po3304 = w39;// level 2
assign po3305 = w2374;// level 2
assign po3306 = w6129;// level 2
assign po3307 = w12863;// level 2
assign po3308 = w14850;// level 2
assign po3309 = w11693;// level 2
assign po3310 = ~w7167;// level 3
assign po3311 = w10023;// level 2
assign po3312 = w9521;// level 2
assign po3313 = w10050;// level 4
assign po3314 = w5811;// level 2
assign po3315 = w10688;// level 2
assign po3316 = w14671;// level 2
assign po3317 = pi3173;// level 0
assign po3318 = w5690;// level 2
assign po3319 = w2532;// level 2
assign po3320 = w13360;// level 2
assign po3321 = ~pi3191;// level 0
assign po3322 = pi3181;// level 0
assign po3323 = w16854;// level 2
assign po3324 = w3891;// level 2
assign po3325 = w6152;// level 2
assign po3326 = w3996;// level 2
assign po3327 = w16631;// level 2
assign po3328 = pi3249;// level 0
assign po3329 = w3468;// level 2
assign po3330 = w9049;// level 2
assign po3331 = w13102;// level 2
assign po3332 = ~w10940;// level 1
assign po3333 = w15409;// level 2
assign po3334 = w15077;// level 2
assign po3335 = w249;// level 2
assign po3336 = w8846;// level 2
assign po3337 = w2926;// level 2
assign po3338 = w9657;// level 2
assign po3339 = w15106;// level 1
assign po3340 = w3032;// level 2
assign po3341 = w11443;// level 2
assign po3342 = w16349;// level 2
assign po3343 = w2717;// level 2
assign po3344 = w17842;// level 2
assign po3345 = pi3211;// level 0
assign po3346 = pi3202;// level 0
assign po3347 = pi3196;// level 0
assign po3348 = pi3215;// level 0
assign po3349 = pi3221;// level 0
assign po3350 = pi3212;// level 0
assign po3351 = ~w325;// level 1
assign po3352 = pi3197;// level 0
assign po3353 = pi3160;// level 0
assign po3354 = pi3236;// level 0
assign po3355 = ~pi3160;// level 0
assign po3356 = pi3234;// level 0
assign po3357 = pi3250;// level 0
assign po3358 = pi3248;// level 0
assign po3359 = pi3230;// level 0
assign po3360 = pi3251;// level 0
assign po3361 = pi3231;// level 0
assign po3362 = pi3123;// level 0
assign po3363 = pi3238;// level 0
assign po3364 = pi3267;// level 0
assign po3365 = pi3265;// level 0
assign po3366 = pi3270;// level 0
assign po3367 = ~pi1973;// level 0
assign po3368 = w12525;// level 1
assign po3369 = ~pi1877;// level 0
assign po3370 = pi3257;// level 0
assign po3371 = pi3252;// level 0
assign po3372 = pi1353;// level 0
assign po3373 = pi3027;// level 0
assign po3374 = ~pi0078;// level 0
assign po3375 = ~pi1965;// level 0
assign po3376 = pi3256;// level 0
assign po3377 = pi3264;// level 0
assign po3378 = ~pi1318;// level 0
assign po3379 = ~pi0120;// level 0
assign po3380 = pi3258;// level 0
assign po3381 = pi3261;// level 0
assign po3382 = pi3269;// level 0
assign po3383 = w17801;// level 1
assign po3384 = w368;// level 1
assign po3385 = pi3253;// level 0
assign po3386 = pi3255;// level 0
assign po3387 = w15733;// level 1
assign po3388 = pi3260;// level 0
assign po3389 = pi3266;// level 0
assign po3390 = pi3263;// level 0
assign po3391 = pi3268;// level 0
assign po3392 = pi3259;// level 0
assign po3393 = w5144;// level 1
assign po3394 = pi3262;// level 0
assign po3395 = pi3271;// level 0
assign po3396 = pi3284;// level 0
assign po3397 = pi3331;// level 0
assign po3398 = pi3339;// level 0
assign po3399 = pi1973;// level 0
assign po3400 = pi3302;// level 0
assign po3401 = pi3323;// level 0
assign po3402 = ~pi1374;// level 0
assign po3403 = pi1685;// level 0
assign po3404 = pi3342;// level 0
assign po3405 = pi3324;// level 0
assign po3406 = pi2908;// level 0
assign po3407 = pi3285;// level 0
assign po3408 = ~pi1405;// level 0
assign po3409 = pi3309;// level 0
assign po3410 = pi2918;// level 0
assign po3411 = pi3184;// level 0
assign po3412 = pi3289;// level 0
assign po3413 = pi3317;// level 0
assign po3414 = pi3296;// level 0
assign po3415 = pi3322;// level 0
assign po3416 = pi3319;// level 0
assign po3417 = pi3352;// level 0
assign po3418 = pi3338;// level 0
assign po3419 = pi3308;// level 0
assign po3420 = pi3297;// level 0
assign po3421 = pi3325;// level 0
assign po3422 = pi3345;// level 0
assign po3423 = pi1400;// level 0
assign po3424 = ~pi0319;// level 0
assign po3425 = ~pi1208;// level 0
assign po3426 = pi0076;// level 0
assign po3427 = ~pi1196;// level 0
assign po3428 = ~pi1409;// level 0
assign po3429 = ~pi1248;// level 0
assign po3430 = ~pi0320;// level 0
assign po3431 = ~pi1383;// level 0
assign po3432 = ~pi1986;// level 0
assign po3433 = ~pi1253;// level 0
assign po3434 = ~pi2384;// level 0
assign po3435 = ~pi2907;// level 0
assign po3436 = ~pi0318;// level 0
assign po3437 = ~pi1408;// level 0
assign po3438 = ~pi2594;// level 0
assign po3439 = ~pi1249;// level 0
assign po3440 = ~pi2358;// level 0
assign po3441 = ~pi1406;// level 0
assign po3442 = ~pi1247;// level 0
assign po3443 = ~pi1194;// level 0
assign po3444 = pi3272;// level 0
assign po3445 = pi3273;// level 0
assign po3446 = pi3274;// level 0
assign po3447 = pi3275;// level 0
assign po3448 = pi3276;// level 0
assign po3449 = pi3277;// level 0
assign po3450 = pi3278;// level 0
assign po3451 = pi3279;// level 0
assign po3452 = pi3280;// level 0
assign po3453 = pi3281;// level 0
assign po3454 = pi3282;// level 0
assign po3455 = pi3283;// level 0
assign po3456 = pi1214;// level 0
assign po3457 = pi2936;// level 0
assign po3458 = pi3455;// level 0
assign po3459 = pi3453;// level 0
assign po3460 = pi3452;// level 0
assign po3461 = pi1222;// level 0
assign po3462 = pi3457;// level 0
assign po3463 = pi3291;// level 0
assign po3464 = pi3292;// level 0
assign po3465 = pi3448;// level 0
assign po3466 = pi3294;// level 0
assign po3467 = pi3467;// level 0
assign po3468 = pi1709;// level 0
assign po3469 = pi3182;// level 0
assign po3470 = pi3461;// level 0
assign po3471 = pi3472;// level 0
assign po3472 = pi3300;// level 0
assign po3473 = pi3301;// level 0
assign po3474 = pi1175;// level 0
assign po3475 = pi3303;// level 0
assign po3476 = pi3304;// level 0
assign po3477 = pi3305;// level 0
assign po3478 = pi3306;// level 0
assign po3479 = pi3307;// level 0
assign po3480 = pi1712;// level 0
assign po3481 = pi1172;// level 0
assign po3482 = pi3310;// level 0
assign po3483 = pi3446;// level 0
assign po3484 = pi3312;// level 0
assign po3485 = pi3450;// level 0
assign po3486 = pi3458;// level 0
assign po3487 = pi3459;// level 0
assign po3488 = pi3443;// level 0
assign po3489 = pi3468;// level 0
assign po3490 = pi1589;// level 0
assign po3491 = pi3464;// level 0
assign po3492 = pi1404;// level 0
assign po3493 = pi2945;// level 0
assign po3494 = pi1215;// level 0
assign po3495 = pi2948;// level 0
assign po3496 = pi3465;// level 0
assign po3497 = pi3327;// level 0
assign po3498 = pi3454;// level 0
assign po3499 = pi3329;// level 0
assign po3500 = pi3463;// level 0
assign po3501 = pi2935;// level 0
assign po3502 = pi3332;// level 0
assign po3503 = pi3462;// level 0
assign po3504 = pi3334;// level 0
assign po3505 = pi3451;// level 0
assign po3506 = pi3466;// level 0
assign po3507 = pi3449;// level 0
assign po3508 = pi1362;// level 0
assign po3509 = pi1153;// level 0
assign po3510 = pi3456;// level 0
assign po3511 = pi3473;// level 0
assign po3512 = pi1166;// level 0
assign po3513 = pi3442;// level 0
assign po3514 = pi3344;// level 0
assign po3515 = pi3210;// level 0
assign po3516 = pi3445;// level 0
assign po3517 = pi3460;// level 0
assign po3518 = pi3174;// level 0
assign po3519 = pi3469;// level 0
assign po3520 = pi3470;// level 0
assign po3521 = pi1403;// level 0
assign po3522 = pi3447;// level 0
assign po3523 = pi3471;// level 0
assign po3524 = pi3444;// level 0
assign po3525 = pi3356;// level 0
assign po3526 = pi3357;// level 0
assign po3527 = pi3358;// level 0
endmodule
