module DSP ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204, pi1205,
    pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213, pi1214,
    pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222, pi1223,
    pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231, pi1232,
    pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240, pi1241,
    pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249, pi1250,
    pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258, pi1259,
    pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267, pi1268,
    pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276, pi1277,
    pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285, pi1286,
    pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294, pi1295,
    pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303, pi1304,
    pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312, pi1313,
    pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321, pi1322,
    pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330, pi1331,
    pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339, pi1340,
    pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348, pi1349,
    pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357, pi1358,
    pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366, pi1367,
    pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375, pi1376,
    pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384, pi1385,
    pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393, pi1394,
    pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402, pi1403,
    pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411, pi1412,
    pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420, pi1421,
    pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429, pi1430,
    pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438, pi1439,
    pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447, pi1448,
    pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456, pi1457,
    pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465, pi1466,
    pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474, pi1475,
    pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483, pi1484,
    pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492, pi1493,
    pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501, pi1502,
    pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510, pi1511,
    pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519, pi1520,
    pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528, pi1529,
    pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537, pi1538,
    pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546, pi1547,
    pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555, pi1556,
    pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564, pi1565,
    pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573, pi1574,
    pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582, pi1583,
    pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591, pi1592,
    pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600, pi1601,
    pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609, pi1610,
    pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618, pi1619,
    pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627, pi1628,
    pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636, pi1637,
    pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645, pi1646,
    pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654, pi1655,
    pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663, pi1664,
    pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672, pi1673,
    pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681, pi1682,
    pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690, pi1691,
    pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699, pi1700,
    pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708, pi1709,
    pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717, pi1718,
    pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726, pi1727,
    pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735, pi1736,
    pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744, pi1745,
    pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753, pi1754,
    pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762, pi1763,
    pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771, pi1772,
    pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780, pi1781,
    pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789, pi1790,
    pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798, pi1799,
    pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807, pi1808,
    pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816, pi1817,
    pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825, pi1826,
    pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834, pi1835,
    pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843, pi1844,
    pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852, pi1853,
    pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861, pi1862,
    pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870, pi1871,
    pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879, pi1880,
    pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888, pi1889,
    pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897, pi1898,
    pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906, pi1907,
    pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915, pi1916,
    pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924, pi1925,
    pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933, pi1934,
    pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942, pi1943,
    pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951, pi1952,
    pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960, pi1961,
    pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969, pi1970,
    pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978, pi1979,
    pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987, pi1988,
    pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996, pi1997,
    pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005, pi2006,
    pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014, pi2015,
    pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023, pi2024,
    pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032, pi2033,
    pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041, pi2042,
    pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050, pi2051,
    pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059, pi2060,
    pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068, pi2069,
    pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077, pi2078,
    pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086, pi2087,
    pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095, pi2096,
    pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104, pi2105,
    pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113, pi2114,
    pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122, pi2123,
    pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131, pi2132,
    pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140, pi2141,
    pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149, pi2150,
    pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158, pi2159,
    pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167, pi2168,
    pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176, pi2177,
    pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185, pi2186,
    pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194, pi2195,
    pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203, pi2204,
    pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212, pi2213,
    pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221, pi2222,
    pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230, pi2231,
    pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239, pi2240,
    pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248, pi2249,
    pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257, pi2258,
    pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266, pi2267,
    pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275, pi2276,
    pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284, pi2285,
    pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293, pi2294,
    pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302, pi2303,
    pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311, pi2312,
    pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320, pi2321,
    pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329, pi2330,
    pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338, pi2339,
    pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347, pi2348,
    pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356, pi2357,
    pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365, pi2366,
    pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374, pi2375,
    pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383, pi2384,
    pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392, pi2393,
    pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401, pi2402,
    pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410, pi2411,
    pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419, pi2420,
    pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428, pi2429,
    pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437, pi2438,
    pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446, pi2447,
    pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455, pi2456,
    pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464, pi2465,
    pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473, pi2474,
    pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482, pi2483,
    pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491, pi2492,
    pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500, pi2501,
    pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509, pi2510,
    pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518, pi2519,
    pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527, pi2528,
    pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536, pi2537,
    pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545, pi2546,
    pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554, pi2555,
    pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563, pi2564,
    pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572, pi2573,
    pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581, pi2582,
    pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590, pi2591,
    pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599, pi2600,
    pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608, pi2609,
    pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617, pi2618,
    pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626, pi2627,
    pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635, pi2636,
    pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644, pi2645,
    pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653, pi2654,
    pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662, pi2663,
    pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671, pi2672,
    pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680, pi2681,
    pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689, pi2690,
    pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698, pi2699,
    pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707, pi2708,
    pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716, pi2717,
    pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725, pi2726,
    pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734, pi2735,
    pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743, pi2744,
    pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752, pi2753,
    pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761, pi2762,
    pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770, pi2771,
    pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779, pi2780,
    pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788, pi2789,
    pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797, pi2798,
    pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806, pi2807,
    pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815, pi2816,
    pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824, pi2825,
    pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833, pi2834,
    pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842, pi2843,
    pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851, pi2852,
    pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860, pi2861,
    pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869, pi2870,
    pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878, pi2879,
    pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887, pi2888,
    pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896, pi2897,
    pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905, pi2906,
    pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914, pi2915,
    pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923, pi2924,
    pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932, pi2933,
    pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941, pi2942,
    pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950, pi2951,
    pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959, pi2960,
    pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968, pi2969,
    pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977, pi2978,
    pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986, pi2987,
    pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995, pi2996,
    pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004, pi3005,
    pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013, pi3014,
    pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022, pi3023,
    pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031, pi3032,
    pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040, pi3041,
    pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049, pi3050,
    pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058, pi3059,
    pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067, pi3068,
    pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076, pi3077,
    pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085, pi3086,
    pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094, pi3095,
    pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103, pi3104,
    pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112, pi3113,
    pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121, pi3122,
    pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130, pi3131,
    pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139, pi3140,
    pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148, pi3149,
    pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157, pi3158,
    pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166, pi3167,
    pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175, pi3176,
    pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184, pi3185,
    pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193, pi3194,
    pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202, pi3203,
    pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211, pi3212,
    pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220, pi3221,
    pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229, pi3230,
    pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238, pi3239,
    pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247, pi3248,
    pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256, pi3257,
    pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265, pi3266,
    pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274, pi3275,
    pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283, pi3284,
    pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292, pi3293,
    pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301, pi3302,
    pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310, pi3311,
    pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319, pi3320,
    pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328, pi3329,
    pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337, pi3338,
    pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346, pi3347,
    pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355, pi3356,
    pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364, pi3365,
    pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373, pi3374,
    pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382, pi3383,
    pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391, pi3392,
    pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400, pi3401,
    pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409, pi3410,
    pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418, pi3419,
    pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427, pi3428,
    pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436, pi3437,
    pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445, pi3446,
    pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454, pi3455,
    pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463, pi3464,
    pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472, pi3473,
    pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481, pi3482,
    pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490, pi3491,
    pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499, pi3500,
    pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508, pi3509,
    pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517, pi3518,
    pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526, pi3527,
    pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535, pi3536,
    pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544, pi3545,
    pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553, pi3554,
    pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562, pi3563,
    pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571, pi3572,
    pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580, pi3581,
    pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589, pi3590,
    pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598, pi3599,
    pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607, pi3608,
    pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616, pi3617,
    pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625, pi3626,
    pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634, pi3635,
    pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643, pi3644,
    pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652, pi3653,
    pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661, pi3662,
    pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670, pi3671,
    pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679, pi3680,
    pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688, pi3689,
    pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697, pi3698,
    pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706, pi3707,
    pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715, pi3716,
    pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724, pi3725,
    pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733, pi3734,
    pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742, pi3743,
    pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751, pi3752,
    pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760, pi3761,
    pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769, pi3770,
    pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778, pi3779,
    pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787, pi3788,
    pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796, pi3797,
    pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805, pi3806,
    pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814, pi3815,
    pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823, pi3824,
    pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832, pi3833,
    pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841, pi3842,
    pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850, pi3851,
    pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859, pi3860,
    pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868, pi3869,
    pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877, pi3878,
    pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886, pi3887,
    pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895, pi3896,
    pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904, pi3905,
    pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913, pi3914,
    pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922, pi3923,
    pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931, pi3932,
    pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940, pi3941,
    pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949, pi3950,
    pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958, pi3959,
    pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967, pi3968,
    pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976, pi3977,
    pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985, pi3986,
    pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994, pi3995,
    pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003, pi4004,
    pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012, pi4013,
    pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021, pi4022,
    pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030, pi4031,
    pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039, pi4040,
    pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048, pi4049,
    pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057, pi4058,
    pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066, pi4067,
    pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075, pi4076,
    pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084, pi4085,
    pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093, pi4094,
    pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102, pi4103,
    pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111, pi4112,
    pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120, pi4121,
    pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129, pi4130,
    pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138, pi4139,
    pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147, pi4148,
    pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156, pi4157,
    pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165, pi4166,
    pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174, pi4175,
    pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183, pi4184,
    pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192, pi4193,
    pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201, pi4202,
    pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210, pi4211,
    pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219, pi4220,
    pi4221, pi4222,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231, po1232,
    po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240, po1241,
    po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249, po1250,
    po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258, po1259,
    po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267, po1268,
    po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276, po1277,
    po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285, po1286,
    po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294, po1295,
    po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303, po1304,
    po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312, po1313,
    po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321, po1322,
    po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330, po1331,
    po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339, po1340,
    po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348, po1349,
    po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357, po1358,
    po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366, po1367,
    po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375, po1376,
    po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384, po1385,
    po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393, po1394,
    po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402, po1403,
    po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411, po1412,
    po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420, po1421,
    po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429, po1430,
    po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438, po1439,
    po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447, po1448,
    po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456, po1457,
    po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465, po1466,
    po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474, po1475,
    po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483, po1484,
    po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492, po1493,
    po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501, po1502,
    po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510, po1511,
    po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519, po1520,
    po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528, po1529,
    po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537, po1538,
    po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546, po1547,
    po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555, po1556,
    po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564, po1565,
    po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573, po1574,
    po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582, po1583,
    po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591, po1592,
    po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600, po1601,
    po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609, po1610,
    po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618, po1619,
    po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627, po1628,
    po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636, po1637,
    po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645, po1646,
    po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654, po1655,
    po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663, po1664,
    po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672, po1673,
    po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681, po1682,
    po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690, po1691,
    po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699, po1700,
    po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708, po1709,
    po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717, po1718,
    po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726, po1727,
    po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735, po1736,
    po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744, po1745,
    po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753, po1754,
    po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762, po1763,
    po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771, po1772,
    po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780, po1781,
    po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789, po1790,
    po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798, po1799,
    po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807, po1808,
    po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816, po1817,
    po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825, po1826,
    po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834, po1835,
    po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843, po1844,
    po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852, po1853,
    po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861, po1862,
    po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870, po1871,
    po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879, po1880,
    po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888, po1889,
    po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897, po1898,
    po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906, po1907,
    po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915, po1916,
    po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924, po1925,
    po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933, po1934,
    po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942, po1943,
    po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951, po1952,
    po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960, po1961,
    po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969, po1970,
    po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978, po1979,
    po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987, po1988,
    po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996, po1997,
    po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005, po2006,
    po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014, po2015,
    po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023, po2024,
    po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032, po2033,
    po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041, po2042,
    po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050, po2051,
    po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059, po2060,
    po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068, po2069,
    po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077, po2078,
    po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086, po2087,
    po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095, po2096,
    po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104, po2105,
    po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113, po2114,
    po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122, po2123,
    po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131, po2132,
    po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140, po2141,
    po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149, po2150,
    po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158, po2159,
    po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167, po2168,
    po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176, po2177,
    po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185, po2186,
    po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194, po2195,
    po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203, po2204,
    po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212, po2213,
    po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221, po2222,
    po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230, po2231,
    po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239, po2240,
    po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248, po2249,
    po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257, po2258,
    po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266, po2267,
    po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275, po2276,
    po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284, po2285,
    po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293, po2294,
    po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302, po2303,
    po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311, po2312,
    po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320, po2321,
    po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329, po2330,
    po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338, po2339,
    po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347, po2348,
    po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356, po2357,
    po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365, po2366,
    po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374, po2375,
    po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383, po2384,
    po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392, po2393,
    po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401, po2402,
    po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410, po2411,
    po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419, po2420,
    po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428, po2429,
    po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437, po2438,
    po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446, po2447,
    po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455, po2456,
    po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464, po2465,
    po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473, po2474,
    po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482, po2483,
    po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491, po2492,
    po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500, po2501,
    po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509, po2510,
    po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518, po2519,
    po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527, po2528,
    po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536, po2537,
    po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545, po2546,
    po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554, po2555,
    po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563, po2564,
    po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572, po2573,
    po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581, po2582,
    po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590, po2591,
    po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599, po2600,
    po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608, po2609,
    po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617, po2618,
    po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626, po2627,
    po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635, po2636,
    po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644, po2645,
    po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653, po2654,
    po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662, po2663,
    po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671, po2672,
    po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680, po2681,
    po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689, po2690,
    po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698, po2699,
    po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707, po2708,
    po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716, po2717,
    po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725, po2726,
    po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734, po2735,
    po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743, po2744,
    po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752, po2753,
    po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761, po2762,
    po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770, po2771,
    po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779, po2780,
    po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788, po2789,
    po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797, po2798,
    po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806, po2807,
    po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815, po2816,
    po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824, po2825,
    po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833, po2834,
    po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842, po2843,
    po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851, po2852,
    po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860, po2861,
    po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869, po2870,
    po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878, po2879,
    po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887, po2888,
    po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896, po2897,
    po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905, po2906,
    po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914, po2915,
    po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923, po2924,
    po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932, po2933,
    po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941, po2942,
    po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950, po2951,
    po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959, po2960,
    po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968, po2969,
    po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977, po2978,
    po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986, po2987,
    po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995, po2996,
    po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004, po3005,
    po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013, po3014,
    po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022, po3023,
    po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031, po3032,
    po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040, po3041,
    po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049, po3050,
    po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058, po3059,
    po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067, po3068,
    po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076, po3077,
    po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085, po3086,
    po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094, po3095,
    po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103, po3104,
    po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112, po3113,
    po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121, po3122,
    po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130, po3131,
    po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139, po3140,
    po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148, po3149,
    po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157, po3158,
    po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166, po3167,
    po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175, po3176,
    po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184, po3185,
    po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193, po3194,
    po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202, po3203,
    po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211, po3212,
    po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220, po3221,
    po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229, po3230,
    po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238, po3239,
    po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247, po3248,
    po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256, po3257,
    po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265, po3266,
    po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274, po3275,
    po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283, po3284,
    po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292, po3293,
    po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301, po3302,
    po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310, po3311,
    po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319, po3320,
    po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328, po3329,
    po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337, po3338,
    po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346, po3347,
    po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355, po3356,
    po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364, po3365,
    po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373, po3374,
    po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382, po3383,
    po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391, po3392,
    po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400, po3401,
    po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409, po3410,
    po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418, po3419,
    po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427, po3428,
    po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436, po3437,
    po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445, po3446,
    po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454, po3455,
    po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463, po3464,
    po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472, po3473,
    po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481, po3482,
    po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490, po3491,
    po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499, po3500,
    po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508, po3509,
    po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517, po3518,
    po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526, po3527,
    po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535, po3536,
    po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544, po3545,
    po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553, po3554,
    po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562, po3563,
    po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571, po3572,
    po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580, po3581,
    po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589, po3590,
    po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598, po3599,
    po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607, po3608,
    po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616, po3617,
    po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625, po3626,
    po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634, po3635,
    po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643, po3644,
    po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652, po3653,
    po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661, po3662,
    po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670, po3671,
    po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679, po3680,
    po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688, po3689,
    po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697, po3698,
    po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706, po3707,
    po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715, po3716,
    po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724, po3725,
    po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733, po3734,
    po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742, po3743,
    po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751, po3752,
    po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760, po3761,
    po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769, po3770,
    po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778, po3779,
    po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787, po3788,
    po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796, po3797,
    po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805, po3806,
    po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814, po3815,
    po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823, po3824,
    po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832, po3833,
    po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841, po3842,
    po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850, po3851,
    po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859, po3860,
    po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868, po3869,
    po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877, po3878,
    po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886, po3887,
    po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895, po3896,
    po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904, po3905,
    po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913, po3914,
    po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922, po3923,
    po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931, po3932,
    po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940, po3941,
    po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949, po3950,
    po3951, po3952  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203, pi1204,
    pi1205, pi1206, pi1207, pi1208, pi1209, pi1210, pi1211, pi1212, pi1213,
    pi1214, pi1215, pi1216, pi1217, pi1218, pi1219, pi1220, pi1221, pi1222,
    pi1223, pi1224, pi1225, pi1226, pi1227, pi1228, pi1229, pi1230, pi1231,
    pi1232, pi1233, pi1234, pi1235, pi1236, pi1237, pi1238, pi1239, pi1240,
    pi1241, pi1242, pi1243, pi1244, pi1245, pi1246, pi1247, pi1248, pi1249,
    pi1250, pi1251, pi1252, pi1253, pi1254, pi1255, pi1256, pi1257, pi1258,
    pi1259, pi1260, pi1261, pi1262, pi1263, pi1264, pi1265, pi1266, pi1267,
    pi1268, pi1269, pi1270, pi1271, pi1272, pi1273, pi1274, pi1275, pi1276,
    pi1277, pi1278, pi1279, pi1280, pi1281, pi1282, pi1283, pi1284, pi1285,
    pi1286, pi1287, pi1288, pi1289, pi1290, pi1291, pi1292, pi1293, pi1294,
    pi1295, pi1296, pi1297, pi1298, pi1299, pi1300, pi1301, pi1302, pi1303,
    pi1304, pi1305, pi1306, pi1307, pi1308, pi1309, pi1310, pi1311, pi1312,
    pi1313, pi1314, pi1315, pi1316, pi1317, pi1318, pi1319, pi1320, pi1321,
    pi1322, pi1323, pi1324, pi1325, pi1326, pi1327, pi1328, pi1329, pi1330,
    pi1331, pi1332, pi1333, pi1334, pi1335, pi1336, pi1337, pi1338, pi1339,
    pi1340, pi1341, pi1342, pi1343, pi1344, pi1345, pi1346, pi1347, pi1348,
    pi1349, pi1350, pi1351, pi1352, pi1353, pi1354, pi1355, pi1356, pi1357,
    pi1358, pi1359, pi1360, pi1361, pi1362, pi1363, pi1364, pi1365, pi1366,
    pi1367, pi1368, pi1369, pi1370, pi1371, pi1372, pi1373, pi1374, pi1375,
    pi1376, pi1377, pi1378, pi1379, pi1380, pi1381, pi1382, pi1383, pi1384,
    pi1385, pi1386, pi1387, pi1388, pi1389, pi1390, pi1391, pi1392, pi1393,
    pi1394, pi1395, pi1396, pi1397, pi1398, pi1399, pi1400, pi1401, pi1402,
    pi1403, pi1404, pi1405, pi1406, pi1407, pi1408, pi1409, pi1410, pi1411,
    pi1412, pi1413, pi1414, pi1415, pi1416, pi1417, pi1418, pi1419, pi1420,
    pi1421, pi1422, pi1423, pi1424, pi1425, pi1426, pi1427, pi1428, pi1429,
    pi1430, pi1431, pi1432, pi1433, pi1434, pi1435, pi1436, pi1437, pi1438,
    pi1439, pi1440, pi1441, pi1442, pi1443, pi1444, pi1445, pi1446, pi1447,
    pi1448, pi1449, pi1450, pi1451, pi1452, pi1453, pi1454, pi1455, pi1456,
    pi1457, pi1458, pi1459, pi1460, pi1461, pi1462, pi1463, pi1464, pi1465,
    pi1466, pi1467, pi1468, pi1469, pi1470, pi1471, pi1472, pi1473, pi1474,
    pi1475, pi1476, pi1477, pi1478, pi1479, pi1480, pi1481, pi1482, pi1483,
    pi1484, pi1485, pi1486, pi1487, pi1488, pi1489, pi1490, pi1491, pi1492,
    pi1493, pi1494, pi1495, pi1496, pi1497, pi1498, pi1499, pi1500, pi1501,
    pi1502, pi1503, pi1504, pi1505, pi1506, pi1507, pi1508, pi1509, pi1510,
    pi1511, pi1512, pi1513, pi1514, pi1515, pi1516, pi1517, pi1518, pi1519,
    pi1520, pi1521, pi1522, pi1523, pi1524, pi1525, pi1526, pi1527, pi1528,
    pi1529, pi1530, pi1531, pi1532, pi1533, pi1534, pi1535, pi1536, pi1537,
    pi1538, pi1539, pi1540, pi1541, pi1542, pi1543, pi1544, pi1545, pi1546,
    pi1547, pi1548, pi1549, pi1550, pi1551, pi1552, pi1553, pi1554, pi1555,
    pi1556, pi1557, pi1558, pi1559, pi1560, pi1561, pi1562, pi1563, pi1564,
    pi1565, pi1566, pi1567, pi1568, pi1569, pi1570, pi1571, pi1572, pi1573,
    pi1574, pi1575, pi1576, pi1577, pi1578, pi1579, pi1580, pi1581, pi1582,
    pi1583, pi1584, pi1585, pi1586, pi1587, pi1588, pi1589, pi1590, pi1591,
    pi1592, pi1593, pi1594, pi1595, pi1596, pi1597, pi1598, pi1599, pi1600,
    pi1601, pi1602, pi1603, pi1604, pi1605, pi1606, pi1607, pi1608, pi1609,
    pi1610, pi1611, pi1612, pi1613, pi1614, pi1615, pi1616, pi1617, pi1618,
    pi1619, pi1620, pi1621, pi1622, pi1623, pi1624, pi1625, pi1626, pi1627,
    pi1628, pi1629, pi1630, pi1631, pi1632, pi1633, pi1634, pi1635, pi1636,
    pi1637, pi1638, pi1639, pi1640, pi1641, pi1642, pi1643, pi1644, pi1645,
    pi1646, pi1647, pi1648, pi1649, pi1650, pi1651, pi1652, pi1653, pi1654,
    pi1655, pi1656, pi1657, pi1658, pi1659, pi1660, pi1661, pi1662, pi1663,
    pi1664, pi1665, pi1666, pi1667, pi1668, pi1669, pi1670, pi1671, pi1672,
    pi1673, pi1674, pi1675, pi1676, pi1677, pi1678, pi1679, pi1680, pi1681,
    pi1682, pi1683, pi1684, pi1685, pi1686, pi1687, pi1688, pi1689, pi1690,
    pi1691, pi1692, pi1693, pi1694, pi1695, pi1696, pi1697, pi1698, pi1699,
    pi1700, pi1701, pi1702, pi1703, pi1704, pi1705, pi1706, pi1707, pi1708,
    pi1709, pi1710, pi1711, pi1712, pi1713, pi1714, pi1715, pi1716, pi1717,
    pi1718, pi1719, pi1720, pi1721, pi1722, pi1723, pi1724, pi1725, pi1726,
    pi1727, pi1728, pi1729, pi1730, pi1731, pi1732, pi1733, pi1734, pi1735,
    pi1736, pi1737, pi1738, pi1739, pi1740, pi1741, pi1742, pi1743, pi1744,
    pi1745, pi1746, pi1747, pi1748, pi1749, pi1750, pi1751, pi1752, pi1753,
    pi1754, pi1755, pi1756, pi1757, pi1758, pi1759, pi1760, pi1761, pi1762,
    pi1763, pi1764, pi1765, pi1766, pi1767, pi1768, pi1769, pi1770, pi1771,
    pi1772, pi1773, pi1774, pi1775, pi1776, pi1777, pi1778, pi1779, pi1780,
    pi1781, pi1782, pi1783, pi1784, pi1785, pi1786, pi1787, pi1788, pi1789,
    pi1790, pi1791, pi1792, pi1793, pi1794, pi1795, pi1796, pi1797, pi1798,
    pi1799, pi1800, pi1801, pi1802, pi1803, pi1804, pi1805, pi1806, pi1807,
    pi1808, pi1809, pi1810, pi1811, pi1812, pi1813, pi1814, pi1815, pi1816,
    pi1817, pi1818, pi1819, pi1820, pi1821, pi1822, pi1823, pi1824, pi1825,
    pi1826, pi1827, pi1828, pi1829, pi1830, pi1831, pi1832, pi1833, pi1834,
    pi1835, pi1836, pi1837, pi1838, pi1839, pi1840, pi1841, pi1842, pi1843,
    pi1844, pi1845, pi1846, pi1847, pi1848, pi1849, pi1850, pi1851, pi1852,
    pi1853, pi1854, pi1855, pi1856, pi1857, pi1858, pi1859, pi1860, pi1861,
    pi1862, pi1863, pi1864, pi1865, pi1866, pi1867, pi1868, pi1869, pi1870,
    pi1871, pi1872, pi1873, pi1874, pi1875, pi1876, pi1877, pi1878, pi1879,
    pi1880, pi1881, pi1882, pi1883, pi1884, pi1885, pi1886, pi1887, pi1888,
    pi1889, pi1890, pi1891, pi1892, pi1893, pi1894, pi1895, pi1896, pi1897,
    pi1898, pi1899, pi1900, pi1901, pi1902, pi1903, pi1904, pi1905, pi1906,
    pi1907, pi1908, pi1909, pi1910, pi1911, pi1912, pi1913, pi1914, pi1915,
    pi1916, pi1917, pi1918, pi1919, pi1920, pi1921, pi1922, pi1923, pi1924,
    pi1925, pi1926, pi1927, pi1928, pi1929, pi1930, pi1931, pi1932, pi1933,
    pi1934, pi1935, pi1936, pi1937, pi1938, pi1939, pi1940, pi1941, pi1942,
    pi1943, pi1944, pi1945, pi1946, pi1947, pi1948, pi1949, pi1950, pi1951,
    pi1952, pi1953, pi1954, pi1955, pi1956, pi1957, pi1958, pi1959, pi1960,
    pi1961, pi1962, pi1963, pi1964, pi1965, pi1966, pi1967, pi1968, pi1969,
    pi1970, pi1971, pi1972, pi1973, pi1974, pi1975, pi1976, pi1977, pi1978,
    pi1979, pi1980, pi1981, pi1982, pi1983, pi1984, pi1985, pi1986, pi1987,
    pi1988, pi1989, pi1990, pi1991, pi1992, pi1993, pi1994, pi1995, pi1996,
    pi1997, pi1998, pi1999, pi2000, pi2001, pi2002, pi2003, pi2004, pi2005,
    pi2006, pi2007, pi2008, pi2009, pi2010, pi2011, pi2012, pi2013, pi2014,
    pi2015, pi2016, pi2017, pi2018, pi2019, pi2020, pi2021, pi2022, pi2023,
    pi2024, pi2025, pi2026, pi2027, pi2028, pi2029, pi2030, pi2031, pi2032,
    pi2033, pi2034, pi2035, pi2036, pi2037, pi2038, pi2039, pi2040, pi2041,
    pi2042, pi2043, pi2044, pi2045, pi2046, pi2047, pi2048, pi2049, pi2050,
    pi2051, pi2052, pi2053, pi2054, pi2055, pi2056, pi2057, pi2058, pi2059,
    pi2060, pi2061, pi2062, pi2063, pi2064, pi2065, pi2066, pi2067, pi2068,
    pi2069, pi2070, pi2071, pi2072, pi2073, pi2074, pi2075, pi2076, pi2077,
    pi2078, pi2079, pi2080, pi2081, pi2082, pi2083, pi2084, pi2085, pi2086,
    pi2087, pi2088, pi2089, pi2090, pi2091, pi2092, pi2093, pi2094, pi2095,
    pi2096, pi2097, pi2098, pi2099, pi2100, pi2101, pi2102, pi2103, pi2104,
    pi2105, pi2106, pi2107, pi2108, pi2109, pi2110, pi2111, pi2112, pi2113,
    pi2114, pi2115, pi2116, pi2117, pi2118, pi2119, pi2120, pi2121, pi2122,
    pi2123, pi2124, pi2125, pi2126, pi2127, pi2128, pi2129, pi2130, pi2131,
    pi2132, pi2133, pi2134, pi2135, pi2136, pi2137, pi2138, pi2139, pi2140,
    pi2141, pi2142, pi2143, pi2144, pi2145, pi2146, pi2147, pi2148, pi2149,
    pi2150, pi2151, pi2152, pi2153, pi2154, pi2155, pi2156, pi2157, pi2158,
    pi2159, pi2160, pi2161, pi2162, pi2163, pi2164, pi2165, pi2166, pi2167,
    pi2168, pi2169, pi2170, pi2171, pi2172, pi2173, pi2174, pi2175, pi2176,
    pi2177, pi2178, pi2179, pi2180, pi2181, pi2182, pi2183, pi2184, pi2185,
    pi2186, pi2187, pi2188, pi2189, pi2190, pi2191, pi2192, pi2193, pi2194,
    pi2195, pi2196, pi2197, pi2198, pi2199, pi2200, pi2201, pi2202, pi2203,
    pi2204, pi2205, pi2206, pi2207, pi2208, pi2209, pi2210, pi2211, pi2212,
    pi2213, pi2214, pi2215, pi2216, pi2217, pi2218, pi2219, pi2220, pi2221,
    pi2222, pi2223, pi2224, pi2225, pi2226, pi2227, pi2228, pi2229, pi2230,
    pi2231, pi2232, pi2233, pi2234, pi2235, pi2236, pi2237, pi2238, pi2239,
    pi2240, pi2241, pi2242, pi2243, pi2244, pi2245, pi2246, pi2247, pi2248,
    pi2249, pi2250, pi2251, pi2252, pi2253, pi2254, pi2255, pi2256, pi2257,
    pi2258, pi2259, pi2260, pi2261, pi2262, pi2263, pi2264, pi2265, pi2266,
    pi2267, pi2268, pi2269, pi2270, pi2271, pi2272, pi2273, pi2274, pi2275,
    pi2276, pi2277, pi2278, pi2279, pi2280, pi2281, pi2282, pi2283, pi2284,
    pi2285, pi2286, pi2287, pi2288, pi2289, pi2290, pi2291, pi2292, pi2293,
    pi2294, pi2295, pi2296, pi2297, pi2298, pi2299, pi2300, pi2301, pi2302,
    pi2303, pi2304, pi2305, pi2306, pi2307, pi2308, pi2309, pi2310, pi2311,
    pi2312, pi2313, pi2314, pi2315, pi2316, pi2317, pi2318, pi2319, pi2320,
    pi2321, pi2322, pi2323, pi2324, pi2325, pi2326, pi2327, pi2328, pi2329,
    pi2330, pi2331, pi2332, pi2333, pi2334, pi2335, pi2336, pi2337, pi2338,
    pi2339, pi2340, pi2341, pi2342, pi2343, pi2344, pi2345, pi2346, pi2347,
    pi2348, pi2349, pi2350, pi2351, pi2352, pi2353, pi2354, pi2355, pi2356,
    pi2357, pi2358, pi2359, pi2360, pi2361, pi2362, pi2363, pi2364, pi2365,
    pi2366, pi2367, pi2368, pi2369, pi2370, pi2371, pi2372, pi2373, pi2374,
    pi2375, pi2376, pi2377, pi2378, pi2379, pi2380, pi2381, pi2382, pi2383,
    pi2384, pi2385, pi2386, pi2387, pi2388, pi2389, pi2390, pi2391, pi2392,
    pi2393, pi2394, pi2395, pi2396, pi2397, pi2398, pi2399, pi2400, pi2401,
    pi2402, pi2403, pi2404, pi2405, pi2406, pi2407, pi2408, pi2409, pi2410,
    pi2411, pi2412, pi2413, pi2414, pi2415, pi2416, pi2417, pi2418, pi2419,
    pi2420, pi2421, pi2422, pi2423, pi2424, pi2425, pi2426, pi2427, pi2428,
    pi2429, pi2430, pi2431, pi2432, pi2433, pi2434, pi2435, pi2436, pi2437,
    pi2438, pi2439, pi2440, pi2441, pi2442, pi2443, pi2444, pi2445, pi2446,
    pi2447, pi2448, pi2449, pi2450, pi2451, pi2452, pi2453, pi2454, pi2455,
    pi2456, pi2457, pi2458, pi2459, pi2460, pi2461, pi2462, pi2463, pi2464,
    pi2465, pi2466, pi2467, pi2468, pi2469, pi2470, pi2471, pi2472, pi2473,
    pi2474, pi2475, pi2476, pi2477, pi2478, pi2479, pi2480, pi2481, pi2482,
    pi2483, pi2484, pi2485, pi2486, pi2487, pi2488, pi2489, pi2490, pi2491,
    pi2492, pi2493, pi2494, pi2495, pi2496, pi2497, pi2498, pi2499, pi2500,
    pi2501, pi2502, pi2503, pi2504, pi2505, pi2506, pi2507, pi2508, pi2509,
    pi2510, pi2511, pi2512, pi2513, pi2514, pi2515, pi2516, pi2517, pi2518,
    pi2519, pi2520, pi2521, pi2522, pi2523, pi2524, pi2525, pi2526, pi2527,
    pi2528, pi2529, pi2530, pi2531, pi2532, pi2533, pi2534, pi2535, pi2536,
    pi2537, pi2538, pi2539, pi2540, pi2541, pi2542, pi2543, pi2544, pi2545,
    pi2546, pi2547, pi2548, pi2549, pi2550, pi2551, pi2552, pi2553, pi2554,
    pi2555, pi2556, pi2557, pi2558, pi2559, pi2560, pi2561, pi2562, pi2563,
    pi2564, pi2565, pi2566, pi2567, pi2568, pi2569, pi2570, pi2571, pi2572,
    pi2573, pi2574, pi2575, pi2576, pi2577, pi2578, pi2579, pi2580, pi2581,
    pi2582, pi2583, pi2584, pi2585, pi2586, pi2587, pi2588, pi2589, pi2590,
    pi2591, pi2592, pi2593, pi2594, pi2595, pi2596, pi2597, pi2598, pi2599,
    pi2600, pi2601, pi2602, pi2603, pi2604, pi2605, pi2606, pi2607, pi2608,
    pi2609, pi2610, pi2611, pi2612, pi2613, pi2614, pi2615, pi2616, pi2617,
    pi2618, pi2619, pi2620, pi2621, pi2622, pi2623, pi2624, pi2625, pi2626,
    pi2627, pi2628, pi2629, pi2630, pi2631, pi2632, pi2633, pi2634, pi2635,
    pi2636, pi2637, pi2638, pi2639, pi2640, pi2641, pi2642, pi2643, pi2644,
    pi2645, pi2646, pi2647, pi2648, pi2649, pi2650, pi2651, pi2652, pi2653,
    pi2654, pi2655, pi2656, pi2657, pi2658, pi2659, pi2660, pi2661, pi2662,
    pi2663, pi2664, pi2665, pi2666, pi2667, pi2668, pi2669, pi2670, pi2671,
    pi2672, pi2673, pi2674, pi2675, pi2676, pi2677, pi2678, pi2679, pi2680,
    pi2681, pi2682, pi2683, pi2684, pi2685, pi2686, pi2687, pi2688, pi2689,
    pi2690, pi2691, pi2692, pi2693, pi2694, pi2695, pi2696, pi2697, pi2698,
    pi2699, pi2700, pi2701, pi2702, pi2703, pi2704, pi2705, pi2706, pi2707,
    pi2708, pi2709, pi2710, pi2711, pi2712, pi2713, pi2714, pi2715, pi2716,
    pi2717, pi2718, pi2719, pi2720, pi2721, pi2722, pi2723, pi2724, pi2725,
    pi2726, pi2727, pi2728, pi2729, pi2730, pi2731, pi2732, pi2733, pi2734,
    pi2735, pi2736, pi2737, pi2738, pi2739, pi2740, pi2741, pi2742, pi2743,
    pi2744, pi2745, pi2746, pi2747, pi2748, pi2749, pi2750, pi2751, pi2752,
    pi2753, pi2754, pi2755, pi2756, pi2757, pi2758, pi2759, pi2760, pi2761,
    pi2762, pi2763, pi2764, pi2765, pi2766, pi2767, pi2768, pi2769, pi2770,
    pi2771, pi2772, pi2773, pi2774, pi2775, pi2776, pi2777, pi2778, pi2779,
    pi2780, pi2781, pi2782, pi2783, pi2784, pi2785, pi2786, pi2787, pi2788,
    pi2789, pi2790, pi2791, pi2792, pi2793, pi2794, pi2795, pi2796, pi2797,
    pi2798, pi2799, pi2800, pi2801, pi2802, pi2803, pi2804, pi2805, pi2806,
    pi2807, pi2808, pi2809, pi2810, pi2811, pi2812, pi2813, pi2814, pi2815,
    pi2816, pi2817, pi2818, pi2819, pi2820, pi2821, pi2822, pi2823, pi2824,
    pi2825, pi2826, pi2827, pi2828, pi2829, pi2830, pi2831, pi2832, pi2833,
    pi2834, pi2835, pi2836, pi2837, pi2838, pi2839, pi2840, pi2841, pi2842,
    pi2843, pi2844, pi2845, pi2846, pi2847, pi2848, pi2849, pi2850, pi2851,
    pi2852, pi2853, pi2854, pi2855, pi2856, pi2857, pi2858, pi2859, pi2860,
    pi2861, pi2862, pi2863, pi2864, pi2865, pi2866, pi2867, pi2868, pi2869,
    pi2870, pi2871, pi2872, pi2873, pi2874, pi2875, pi2876, pi2877, pi2878,
    pi2879, pi2880, pi2881, pi2882, pi2883, pi2884, pi2885, pi2886, pi2887,
    pi2888, pi2889, pi2890, pi2891, pi2892, pi2893, pi2894, pi2895, pi2896,
    pi2897, pi2898, pi2899, pi2900, pi2901, pi2902, pi2903, pi2904, pi2905,
    pi2906, pi2907, pi2908, pi2909, pi2910, pi2911, pi2912, pi2913, pi2914,
    pi2915, pi2916, pi2917, pi2918, pi2919, pi2920, pi2921, pi2922, pi2923,
    pi2924, pi2925, pi2926, pi2927, pi2928, pi2929, pi2930, pi2931, pi2932,
    pi2933, pi2934, pi2935, pi2936, pi2937, pi2938, pi2939, pi2940, pi2941,
    pi2942, pi2943, pi2944, pi2945, pi2946, pi2947, pi2948, pi2949, pi2950,
    pi2951, pi2952, pi2953, pi2954, pi2955, pi2956, pi2957, pi2958, pi2959,
    pi2960, pi2961, pi2962, pi2963, pi2964, pi2965, pi2966, pi2967, pi2968,
    pi2969, pi2970, pi2971, pi2972, pi2973, pi2974, pi2975, pi2976, pi2977,
    pi2978, pi2979, pi2980, pi2981, pi2982, pi2983, pi2984, pi2985, pi2986,
    pi2987, pi2988, pi2989, pi2990, pi2991, pi2992, pi2993, pi2994, pi2995,
    pi2996, pi2997, pi2998, pi2999, pi3000, pi3001, pi3002, pi3003, pi3004,
    pi3005, pi3006, pi3007, pi3008, pi3009, pi3010, pi3011, pi3012, pi3013,
    pi3014, pi3015, pi3016, pi3017, pi3018, pi3019, pi3020, pi3021, pi3022,
    pi3023, pi3024, pi3025, pi3026, pi3027, pi3028, pi3029, pi3030, pi3031,
    pi3032, pi3033, pi3034, pi3035, pi3036, pi3037, pi3038, pi3039, pi3040,
    pi3041, pi3042, pi3043, pi3044, pi3045, pi3046, pi3047, pi3048, pi3049,
    pi3050, pi3051, pi3052, pi3053, pi3054, pi3055, pi3056, pi3057, pi3058,
    pi3059, pi3060, pi3061, pi3062, pi3063, pi3064, pi3065, pi3066, pi3067,
    pi3068, pi3069, pi3070, pi3071, pi3072, pi3073, pi3074, pi3075, pi3076,
    pi3077, pi3078, pi3079, pi3080, pi3081, pi3082, pi3083, pi3084, pi3085,
    pi3086, pi3087, pi3088, pi3089, pi3090, pi3091, pi3092, pi3093, pi3094,
    pi3095, pi3096, pi3097, pi3098, pi3099, pi3100, pi3101, pi3102, pi3103,
    pi3104, pi3105, pi3106, pi3107, pi3108, pi3109, pi3110, pi3111, pi3112,
    pi3113, pi3114, pi3115, pi3116, pi3117, pi3118, pi3119, pi3120, pi3121,
    pi3122, pi3123, pi3124, pi3125, pi3126, pi3127, pi3128, pi3129, pi3130,
    pi3131, pi3132, pi3133, pi3134, pi3135, pi3136, pi3137, pi3138, pi3139,
    pi3140, pi3141, pi3142, pi3143, pi3144, pi3145, pi3146, pi3147, pi3148,
    pi3149, pi3150, pi3151, pi3152, pi3153, pi3154, pi3155, pi3156, pi3157,
    pi3158, pi3159, pi3160, pi3161, pi3162, pi3163, pi3164, pi3165, pi3166,
    pi3167, pi3168, pi3169, pi3170, pi3171, pi3172, pi3173, pi3174, pi3175,
    pi3176, pi3177, pi3178, pi3179, pi3180, pi3181, pi3182, pi3183, pi3184,
    pi3185, pi3186, pi3187, pi3188, pi3189, pi3190, pi3191, pi3192, pi3193,
    pi3194, pi3195, pi3196, pi3197, pi3198, pi3199, pi3200, pi3201, pi3202,
    pi3203, pi3204, pi3205, pi3206, pi3207, pi3208, pi3209, pi3210, pi3211,
    pi3212, pi3213, pi3214, pi3215, pi3216, pi3217, pi3218, pi3219, pi3220,
    pi3221, pi3222, pi3223, pi3224, pi3225, pi3226, pi3227, pi3228, pi3229,
    pi3230, pi3231, pi3232, pi3233, pi3234, pi3235, pi3236, pi3237, pi3238,
    pi3239, pi3240, pi3241, pi3242, pi3243, pi3244, pi3245, pi3246, pi3247,
    pi3248, pi3249, pi3250, pi3251, pi3252, pi3253, pi3254, pi3255, pi3256,
    pi3257, pi3258, pi3259, pi3260, pi3261, pi3262, pi3263, pi3264, pi3265,
    pi3266, pi3267, pi3268, pi3269, pi3270, pi3271, pi3272, pi3273, pi3274,
    pi3275, pi3276, pi3277, pi3278, pi3279, pi3280, pi3281, pi3282, pi3283,
    pi3284, pi3285, pi3286, pi3287, pi3288, pi3289, pi3290, pi3291, pi3292,
    pi3293, pi3294, pi3295, pi3296, pi3297, pi3298, pi3299, pi3300, pi3301,
    pi3302, pi3303, pi3304, pi3305, pi3306, pi3307, pi3308, pi3309, pi3310,
    pi3311, pi3312, pi3313, pi3314, pi3315, pi3316, pi3317, pi3318, pi3319,
    pi3320, pi3321, pi3322, pi3323, pi3324, pi3325, pi3326, pi3327, pi3328,
    pi3329, pi3330, pi3331, pi3332, pi3333, pi3334, pi3335, pi3336, pi3337,
    pi3338, pi3339, pi3340, pi3341, pi3342, pi3343, pi3344, pi3345, pi3346,
    pi3347, pi3348, pi3349, pi3350, pi3351, pi3352, pi3353, pi3354, pi3355,
    pi3356, pi3357, pi3358, pi3359, pi3360, pi3361, pi3362, pi3363, pi3364,
    pi3365, pi3366, pi3367, pi3368, pi3369, pi3370, pi3371, pi3372, pi3373,
    pi3374, pi3375, pi3376, pi3377, pi3378, pi3379, pi3380, pi3381, pi3382,
    pi3383, pi3384, pi3385, pi3386, pi3387, pi3388, pi3389, pi3390, pi3391,
    pi3392, pi3393, pi3394, pi3395, pi3396, pi3397, pi3398, pi3399, pi3400,
    pi3401, pi3402, pi3403, pi3404, pi3405, pi3406, pi3407, pi3408, pi3409,
    pi3410, pi3411, pi3412, pi3413, pi3414, pi3415, pi3416, pi3417, pi3418,
    pi3419, pi3420, pi3421, pi3422, pi3423, pi3424, pi3425, pi3426, pi3427,
    pi3428, pi3429, pi3430, pi3431, pi3432, pi3433, pi3434, pi3435, pi3436,
    pi3437, pi3438, pi3439, pi3440, pi3441, pi3442, pi3443, pi3444, pi3445,
    pi3446, pi3447, pi3448, pi3449, pi3450, pi3451, pi3452, pi3453, pi3454,
    pi3455, pi3456, pi3457, pi3458, pi3459, pi3460, pi3461, pi3462, pi3463,
    pi3464, pi3465, pi3466, pi3467, pi3468, pi3469, pi3470, pi3471, pi3472,
    pi3473, pi3474, pi3475, pi3476, pi3477, pi3478, pi3479, pi3480, pi3481,
    pi3482, pi3483, pi3484, pi3485, pi3486, pi3487, pi3488, pi3489, pi3490,
    pi3491, pi3492, pi3493, pi3494, pi3495, pi3496, pi3497, pi3498, pi3499,
    pi3500, pi3501, pi3502, pi3503, pi3504, pi3505, pi3506, pi3507, pi3508,
    pi3509, pi3510, pi3511, pi3512, pi3513, pi3514, pi3515, pi3516, pi3517,
    pi3518, pi3519, pi3520, pi3521, pi3522, pi3523, pi3524, pi3525, pi3526,
    pi3527, pi3528, pi3529, pi3530, pi3531, pi3532, pi3533, pi3534, pi3535,
    pi3536, pi3537, pi3538, pi3539, pi3540, pi3541, pi3542, pi3543, pi3544,
    pi3545, pi3546, pi3547, pi3548, pi3549, pi3550, pi3551, pi3552, pi3553,
    pi3554, pi3555, pi3556, pi3557, pi3558, pi3559, pi3560, pi3561, pi3562,
    pi3563, pi3564, pi3565, pi3566, pi3567, pi3568, pi3569, pi3570, pi3571,
    pi3572, pi3573, pi3574, pi3575, pi3576, pi3577, pi3578, pi3579, pi3580,
    pi3581, pi3582, pi3583, pi3584, pi3585, pi3586, pi3587, pi3588, pi3589,
    pi3590, pi3591, pi3592, pi3593, pi3594, pi3595, pi3596, pi3597, pi3598,
    pi3599, pi3600, pi3601, pi3602, pi3603, pi3604, pi3605, pi3606, pi3607,
    pi3608, pi3609, pi3610, pi3611, pi3612, pi3613, pi3614, pi3615, pi3616,
    pi3617, pi3618, pi3619, pi3620, pi3621, pi3622, pi3623, pi3624, pi3625,
    pi3626, pi3627, pi3628, pi3629, pi3630, pi3631, pi3632, pi3633, pi3634,
    pi3635, pi3636, pi3637, pi3638, pi3639, pi3640, pi3641, pi3642, pi3643,
    pi3644, pi3645, pi3646, pi3647, pi3648, pi3649, pi3650, pi3651, pi3652,
    pi3653, pi3654, pi3655, pi3656, pi3657, pi3658, pi3659, pi3660, pi3661,
    pi3662, pi3663, pi3664, pi3665, pi3666, pi3667, pi3668, pi3669, pi3670,
    pi3671, pi3672, pi3673, pi3674, pi3675, pi3676, pi3677, pi3678, pi3679,
    pi3680, pi3681, pi3682, pi3683, pi3684, pi3685, pi3686, pi3687, pi3688,
    pi3689, pi3690, pi3691, pi3692, pi3693, pi3694, pi3695, pi3696, pi3697,
    pi3698, pi3699, pi3700, pi3701, pi3702, pi3703, pi3704, pi3705, pi3706,
    pi3707, pi3708, pi3709, pi3710, pi3711, pi3712, pi3713, pi3714, pi3715,
    pi3716, pi3717, pi3718, pi3719, pi3720, pi3721, pi3722, pi3723, pi3724,
    pi3725, pi3726, pi3727, pi3728, pi3729, pi3730, pi3731, pi3732, pi3733,
    pi3734, pi3735, pi3736, pi3737, pi3738, pi3739, pi3740, pi3741, pi3742,
    pi3743, pi3744, pi3745, pi3746, pi3747, pi3748, pi3749, pi3750, pi3751,
    pi3752, pi3753, pi3754, pi3755, pi3756, pi3757, pi3758, pi3759, pi3760,
    pi3761, pi3762, pi3763, pi3764, pi3765, pi3766, pi3767, pi3768, pi3769,
    pi3770, pi3771, pi3772, pi3773, pi3774, pi3775, pi3776, pi3777, pi3778,
    pi3779, pi3780, pi3781, pi3782, pi3783, pi3784, pi3785, pi3786, pi3787,
    pi3788, pi3789, pi3790, pi3791, pi3792, pi3793, pi3794, pi3795, pi3796,
    pi3797, pi3798, pi3799, pi3800, pi3801, pi3802, pi3803, pi3804, pi3805,
    pi3806, pi3807, pi3808, pi3809, pi3810, pi3811, pi3812, pi3813, pi3814,
    pi3815, pi3816, pi3817, pi3818, pi3819, pi3820, pi3821, pi3822, pi3823,
    pi3824, pi3825, pi3826, pi3827, pi3828, pi3829, pi3830, pi3831, pi3832,
    pi3833, pi3834, pi3835, pi3836, pi3837, pi3838, pi3839, pi3840, pi3841,
    pi3842, pi3843, pi3844, pi3845, pi3846, pi3847, pi3848, pi3849, pi3850,
    pi3851, pi3852, pi3853, pi3854, pi3855, pi3856, pi3857, pi3858, pi3859,
    pi3860, pi3861, pi3862, pi3863, pi3864, pi3865, pi3866, pi3867, pi3868,
    pi3869, pi3870, pi3871, pi3872, pi3873, pi3874, pi3875, pi3876, pi3877,
    pi3878, pi3879, pi3880, pi3881, pi3882, pi3883, pi3884, pi3885, pi3886,
    pi3887, pi3888, pi3889, pi3890, pi3891, pi3892, pi3893, pi3894, pi3895,
    pi3896, pi3897, pi3898, pi3899, pi3900, pi3901, pi3902, pi3903, pi3904,
    pi3905, pi3906, pi3907, pi3908, pi3909, pi3910, pi3911, pi3912, pi3913,
    pi3914, pi3915, pi3916, pi3917, pi3918, pi3919, pi3920, pi3921, pi3922,
    pi3923, pi3924, pi3925, pi3926, pi3927, pi3928, pi3929, pi3930, pi3931,
    pi3932, pi3933, pi3934, pi3935, pi3936, pi3937, pi3938, pi3939, pi3940,
    pi3941, pi3942, pi3943, pi3944, pi3945, pi3946, pi3947, pi3948, pi3949,
    pi3950, pi3951, pi3952, pi3953, pi3954, pi3955, pi3956, pi3957, pi3958,
    pi3959, pi3960, pi3961, pi3962, pi3963, pi3964, pi3965, pi3966, pi3967,
    pi3968, pi3969, pi3970, pi3971, pi3972, pi3973, pi3974, pi3975, pi3976,
    pi3977, pi3978, pi3979, pi3980, pi3981, pi3982, pi3983, pi3984, pi3985,
    pi3986, pi3987, pi3988, pi3989, pi3990, pi3991, pi3992, pi3993, pi3994,
    pi3995, pi3996, pi3997, pi3998, pi3999, pi4000, pi4001, pi4002, pi4003,
    pi4004, pi4005, pi4006, pi4007, pi4008, pi4009, pi4010, pi4011, pi4012,
    pi4013, pi4014, pi4015, pi4016, pi4017, pi4018, pi4019, pi4020, pi4021,
    pi4022, pi4023, pi4024, pi4025, pi4026, pi4027, pi4028, pi4029, pi4030,
    pi4031, pi4032, pi4033, pi4034, pi4035, pi4036, pi4037, pi4038, pi4039,
    pi4040, pi4041, pi4042, pi4043, pi4044, pi4045, pi4046, pi4047, pi4048,
    pi4049, pi4050, pi4051, pi4052, pi4053, pi4054, pi4055, pi4056, pi4057,
    pi4058, pi4059, pi4060, pi4061, pi4062, pi4063, pi4064, pi4065, pi4066,
    pi4067, pi4068, pi4069, pi4070, pi4071, pi4072, pi4073, pi4074, pi4075,
    pi4076, pi4077, pi4078, pi4079, pi4080, pi4081, pi4082, pi4083, pi4084,
    pi4085, pi4086, pi4087, pi4088, pi4089, pi4090, pi4091, pi4092, pi4093,
    pi4094, pi4095, pi4096, pi4097, pi4098, pi4099, pi4100, pi4101, pi4102,
    pi4103, pi4104, pi4105, pi4106, pi4107, pi4108, pi4109, pi4110, pi4111,
    pi4112, pi4113, pi4114, pi4115, pi4116, pi4117, pi4118, pi4119, pi4120,
    pi4121, pi4122, pi4123, pi4124, pi4125, pi4126, pi4127, pi4128, pi4129,
    pi4130, pi4131, pi4132, pi4133, pi4134, pi4135, pi4136, pi4137, pi4138,
    pi4139, pi4140, pi4141, pi4142, pi4143, pi4144, pi4145, pi4146, pi4147,
    pi4148, pi4149, pi4150, pi4151, pi4152, pi4153, pi4154, pi4155, pi4156,
    pi4157, pi4158, pi4159, pi4160, pi4161, pi4162, pi4163, pi4164, pi4165,
    pi4166, pi4167, pi4168, pi4169, pi4170, pi4171, pi4172, pi4173, pi4174,
    pi4175, pi4176, pi4177, pi4178, pi4179, pi4180, pi4181, pi4182, pi4183,
    pi4184, pi4185, pi4186, pi4187, pi4188, pi4189, pi4190, pi4191, pi4192,
    pi4193, pi4194, pi4195, pi4196, pi4197, pi4198, pi4199, pi4200, pi4201,
    pi4202, pi4203, pi4204, pi4205, pi4206, pi4207, pi4208, pi4209, pi4210,
    pi4211, pi4212, pi4213, pi4214, pi4215, pi4216, pi4217, pi4218, pi4219,
    pi4220, pi4221, pi4222;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230, po1231,
    po1232, po1233, po1234, po1235, po1236, po1237, po1238, po1239, po1240,
    po1241, po1242, po1243, po1244, po1245, po1246, po1247, po1248, po1249,
    po1250, po1251, po1252, po1253, po1254, po1255, po1256, po1257, po1258,
    po1259, po1260, po1261, po1262, po1263, po1264, po1265, po1266, po1267,
    po1268, po1269, po1270, po1271, po1272, po1273, po1274, po1275, po1276,
    po1277, po1278, po1279, po1280, po1281, po1282, po1283, po1284, po1285,
    po1286, po1287, po1288, po1289, po1290, po1291, po1292, po1293, po1294,
    po1295, po1296, po1297, po1298, po1299, po1300, po1301, po1302, po1303,
    po1304, po1305, po1306, po1307, po1308, po1309, po1310, po1311, po1312,
    po1313, po1314, po1315, po1316, po1317, po1318, po1319, po1320, po1321,
    po1322, po1323, po1324, po1325, po1326, po1327, po1328, po1329, po1330,
    po1331, po1332, po1333, po1334, po1335, po1336, po1337, po1338, po1339,
    po1340, po1341, po1342, po1343, po1344, po1345, po1346, po1347, po1348,
    po1349, po1350, po1351, po1352, po1353, po1354, po1355, po1356, po1357,
    po1358, po1359, po1360, po1361, po1362, po1363, po1364, po1365, po1366,
    po1367, po1368, po1369, po1370, po1371, po1372, po1373, po1374, po1375,
    po1376, po1377, po1378, po1379, po1380, po1381, po1382, po1383, po1384,
    po1385, po1386, po1387, po1388, po1389, po1390, po1391, po1392, po1393,
    po1394, po1395, po1396, po1397, po1398, po1399, po1400, po1401, po1402,
    po1403, po1404, po1405, po1406, po1407, po1408, po1409, po1410, po1411,
    po1412, po1413, po1414, po1415, po1416, po1417, po1418, po1419, po1420,
    po1421, po1422, po1423, po1424, po1425, po1426, po1427, po1428, po1429,
    po1430, po1431, po1432, po1433, po1434, po1435, po1436, po1437, po1438,
    po1439, po1440, po1441, po1442, po1443, po1444, po1445, po1446, po1447,
    po1448, po1449, po1450, po1451, po1452, po1453, po1454, po1455, po1456,
    po1457, po1458, po1459, po1460, po1461, po1462, po1463, po1464, po1465,
    po1466, po1467, po1468, po1469, po1470, po1471, po1472, po1473, po1474,
    po1475, po1476, po1477, po1478, po1479, po1480, po1481, po1482, po1483,
    po1484, po1485, po1486, po1487, po1488, po1489, po1490, po1491, po1492,
    po1493, po1494, po1495, po1496, po1497, po1498, po1499, po1500, po1501,
    po1502, po1503, po1504, po1505, po1506, po1507, po1508, po1509, po1510,
    po1511, po1512, po1513, po1514, po1515, po1516, po1517, po1518, po1519,
    po1520, po1521, po1522, po1523, po1524, po1525, po1526, po1527, po1528,
    po1529, po1530, po1531, po1532, po1533, po1534, po1535, po1536, po1537,
    po1538, po1539, po1540, po1541, po1542, po1543, po1544, po1545, po1546,
    po1547, po1548, po1549, po1550, po1551, po1552, po1553, po1554, po1555,
    po1556, po1557, po1558, po1559, po1560, po1561, po1562, po1563, po1564,
    po1565, po1566, po1567, po1568, po1569, po1570, po1571, po1572, po1573,
    po1574, po1575, po1576, po1577, po1578, po1579, po1580, po1581, po1582,
    po1583, po1584, po1585, po1586, po1587, po1588, po1589, po1590, po1591,
    po1592, po1593, po1594, po1595, po1596, po1597, po1598, po1599, po1600,
    po1601, po1602, po1603, po1604, po1605, po1606, po1607, po1608, po1609,
    po1610, po1611, po1612, po1613, po1614, po1615, po1616, po1617, po1618,
    po1619, po1620, po1621, po1622, po1623, po1624, po1625, po1626, po1627,
    po1628, po1629, po1630, po1631, po1632, po1633, po1634, po1635, po1636,
    po1637, po1638, po1639, po1640, po1641, po1642, po1643, po1644, po1645,
    po1646, po1647, po1648, po1649, po1650, po1651, po1652, po1653, po1654,
    po1655, po1656, po1657, po1658, po1659, po1660, po1661, po1662, po1663,
    po1664, po1665, po1666, po1667, po1668, po1669, po1670, po1671, po1672,
    po1673, po1674, po1675, po1676, po1677, po1678, po1679, po1680, po1681,
    po1682, po1683, po1684, po1685, po1686, po1687, po1688, po1689, po1690,
    po1691, po1692, po1693, po1694, po1695, po1696, po1697, po1698, po1699,
    po1700, po1701, po1702, po1703, po1704, po1705, po1706, po1707, po1708,
    po1709, po1710, po1711, po1712, po1713, po1714, po1715, po1716, po1717,
    po1718, po1719, po1720, po1721, po1722, po1723, po1724, po1725, po1726,
    po1727, po1728, po1729, po1730, po1731, po1732, po1733, po1734, po1735,
    po1736, po1737, po1738, po1739, po1740, po1741, po1742, po1743, po1744,
    po1745, po1746, po1747, po1748, po1749, po1750, po1751, po1752, po1753,
    po1754, po1755, po1756, po1757, po1758, po1759, po1760, po1761, po1762,
    po1763, po1764, po1765, po1766, po1767, po1768, po1769, po1770, po1771,
    po1772, po1773, po1774, po1775, po1776, po1777, po1778, po1779, po1780,
    po1781, po1782, po1783, po1784, po1785, po1786, po1787, po1788, po1789,
    po1790, po1791, po1792, po1793, po1794, po1795, po1796, po1797, po1798,
    po1799, po1800, po1801, po1802, po1803, po1804, po1805, po1806, po1807,
    po1808, po1809, po1810, po1811, po1812, po1813, po1814, po1815, po1816,
    po1817, po1818, po1819, po1820, po1821, po1822, po1823, po1824, po1825,
    po1826, po1827, po1828, po1829, po1830, po1831, po1832, po1833, po1834,
    po1835, po1836, po1837, po1838, po1839, po1840, po1841, po1842, po1843,
    po1844, po1845, po1846, po1847, po1848, po1849, po1850, po1851, po1852,
    po1853, po1854, po1855, po1856, po1857, po1858, po1859, po1860, po1861,
    po1862, po1863, po1864, po1865, po1866, po1867, po1868, po1869, po1870,
    po1871, po1872, po1873, po1874, po1875, po1876, po1877, po1878, po1879,
    po1880, po1881, po1882, po1883, po1884, po1885, po1886, po1887, po1888,
    po1889, po1890, po1891, po1892, po1893, po1894, po1895, po1896, po1897,
    po1898, po1899, po1900, po1901, po1902, po1903, po1904, po1905, po1906,
    po1907, po1908, po1909, po1910, po1911, po1912, po1913, po1914, po1915,
    po1916, po1917, po1918, po1919, po1920, po1921, po1922, po1923, po1924,
    po1925, po1926, po1927, po1928, po1929, po1930, po1931, po1932, po1933,
    po1934, po1935, po1936, po1937, po1938, po1939, po1940, po1941, po1942,
    po1943, po1944, po1945, po1946, po1947, po1948, po1949, po1950, po1951,
    po1952, po1953, po1954, po1955, po1956, po1957, po1958, po1959, po1960,
    po1961, po1962, po1963, po1964, po1965, po1966, po1967, po1968, po1969,
    po1970, po1971, po1972, po1973, po1974, po1975, po1976, po1977, po1978,
    po1979, po1980, po1981, po1982, po1983, po1984, po1985, po1986, po1987,
    po1988, po1989, po1990, po1991, po1992, po1993, po1994, po1995, po1996,
    po1997, po1998, po1999, po2000, po2001, po2002, po2003, po2004, po2005,
    po2006, po2007, po2008, po2009, po2010, po2011, po2012, po2013, po2014,
    po2015, po2016, po2017, po2018, po2019, po2020, po2021, po2022, po2023,
    po2024, po2025, po2026, po2027, po2028, po2029, po2030, po2031, po2032,
    po2033, po2034, po2035, po2036, po2037, po2038, po2039, po2040, po2041,
    po2042, po2043, po2044, po2045, po2046, po2047, po2048, po2049, po2050,
    po2051, po2052, po2053, po2054, po2055, po2056, po2057, po2058, po2059,
    po2060, po2061, po2062, po2063, po2064, po2065, po2066, po2067, po2068,
    po2069, po2070, po2071, po2072, po2073, po2074, po2075, po2076, po2077,
    po2078, po2079, po2080, po2081, po2082, po2083, po2084, po2085, po2086,
    po2087, po2088, po2089, po2090, po2091, po2092, po2093, po2094, po2095,
    po2096, po2097, po2098, po2099, po2100, po2101, po2102, po2103, po2104,
    po2105, po2106, po2107, po2108, po2109, po2110, po2111, po2112, po2113,
    po2114, po2115, po2116, po2117, po2118, po2119, po2120, po2121, po2122,
    po2123, po2124, po2125, po2126, po2127, po2128, po2129, po2130, po2131,
    po2132, po2133, po2134, po2135, po2136, po2137, po2138, po2139, po2140,
    po2141, po2142, po2143, po2144, po2145, po2146, po2147, po2148, po2149,
    po2150, po2151, po2152, po2153, po2154, po2155, po2156, po2157, po2158,
    po2159, po2160, po2161, po2162, po2163, po2164, po2165, po2166, po2167,
    po2168, po2169, po2170, po2171, po2172, po2173, po2174, po2175, po2176,
    po2177, po2178, po2179, po2180, po2181, po2182, po2183, po2184, po2185,
    po2186, po2187, po2188, po2189, po2190, po2191, po2192, po2193, po2194,
    po2195, po2196, po2197, po2198, po2199, po2200, po2201, po2202, po2203,
    po2204, po2205, po2206, po2207, po2208, po2209, po2210, po2211, po2212,
    po2213, po2214, po2215, po2216, po2217, po2218, po2219, po2220, po2221,
    po2222, po2223, po2224, po2225, po2226, po2227, po2228, po2229, po2230,
    po2231, po2232, po2233, po2234, po2235, po2236, po2237, po2238, po2239,
    po2240, po2241, po2242, po2243, po2244, po2245, po2246, po2247, po2248,
    po2249, po2250, po2251, po2252, po2253, po2254, po2255, po2256, po2257,
    po2258, po2259, po2260, po2261, po2262, po2263, po2264, po2265, po2266,
    po2267, po2268, po2269, po2270, po2271, po2272, po2273, po2274, po2275,
    po2276, po2277, po2278, po2279, po2280, po2281, po2282, po2283, po2284,
    po2285, po2286, po2287, po2288, po2289, po2290, po2291, po2292, po2293,
    po2294, po2295, po2296, po2297, po2298, po2299, po2300, po2301, po2302,
    po2303, po2304, po2305, po2306, po2307, po2308, po2309, po2310, po2311,
    po2312, po2313, po2314, po2315, po2316, po2317, po2318, po2319, po2320,
    po2321, po2322, po2323, po2324, po2325, po2326, po2327, po2328, po2329,
    po2330, po2331, po2332, po2333, po2334, po2335, po2336, po2337, po2338,
    po2339, po2340, po2341, po2342, po2343, po2344, po2345, po2346, po2347,
    po2348, po2349, po2350, po2351, po2352, po2353, po2354, po2355, po2356,
    po2357, po2358, po2359, po2360, po2361, po2362, po2363, po2364, po2365,
    po2366, po2367, po2368, po2369, po2370, po2371, po2372, po2373, po2374,
    po2375, po2376, po2377, po2378, po2379, po2380, po2381, po2382, po2383,
    po2384, po2385, po2386, po2387, po2388, po2389, po2390, po2391, po2392,
    po2393, po2394, po2395, po2396, po2397, po2398, po2399, po2400, po2401,
    po2402, po2403, po2404, po2405, po2406, po2407, po2408, po2409, po2410,
    po2411, po2412, po2413, po2414, po2415, po2416, po2417, po2418, po2419,
    po2420, po2421, po2422, po2423, po2424, po2425, po2426, po2427, po2428,
    po2429, po2430, po2431, po2432, po2433, po2434, po2435, po2436, po2437,
    po2438, po2439, po2440, po2441, po2442, po2443, po2444, po2445, po2446,
    po2447, po2448, po2449, po2450, po2451, po2452, po2453, po2454, po2455,
    po2456, po2457, po2458, po2459, po2460, po2461, po2462, po2463, po2464,
    po2465, po2466, po2467, po2468, po2469, po2470, po2471, po2472, po2473,
    po2474, po2475, po2476, po2477, po2478, po2479, po2480, po2481, po2482,
    po2483, po2484, po2485, po2486, po2487, po2488, po2489, po2490, po2491,
    po2492, po2493, po2494, po2495, po2496, po2497, po2498, po2499, po2500,
    po2501, po2502, po2503, po2504, po2505, po2506, po2507, po2508, po2509,
    po2510, po2511, po2512, po2513, po2514, po2515, po2516, po2517, po2518,
    po2519, po2520, po2521, po2522, po2523, po2524, po2525, po2526, po2527,
    po2528, po2529, po2530, po2531, po2532, po2533, po2534, po2535, po2536,
    po2537, po2538, po2539, po2540, po2541, po2542, po2543, po2544, po2545,
    po2546, po2547, po2548, po2549, po2550, po2551, po2552, po2553, po2554,
    po2555, po2556, po2557, po2558, po2559, po2560, po2561, po2562, po2563,
    po2564, po2565, po2566, po2567, po2568, po2569, po2570, po2571, po2572,
    po2573, po2574, po2575, po2576, po2577, po2578, po2579, po2580, po2581,
    po2582, po2583, po2584, po2585, po2586, po2587, po2588, po2589, po2590,
    po2591, po2592, po2593, po2594, po2595, po2596, po2597, po2598, po2599,
    po2600, po2601, po2602, po2603, po2604, po2605, po2606, po2607, po2608,
    po2609, po2610, po2611, po2612, po2613, po2614, po2615, po2616, po2617,
    po2618, po2619, po2620, po2621, po2622, po2623, po2624, po2625, po2626,
    po2627, po2628, po2629, po2630, po2631, po2632, po2633, po2634, po2635,
    po2636, po2637, po2638, po2639, po2640, po2641, po2642, po2643, po2644,
    po2645, po2646, po2647, po2648, po2649, po2650, po2651, po2652, po2653,
    po2654, po2655, po2656, po2657, po2658, po2659, po2660, po2661, po2662,
    po2663, po2664, po2665, po2666, po2667, po2668, po2669, po2670, po2671,
    po2672, po2673, po2674, po2675, po2676, po2677, po2678, po2679, po2680,
    po2681, po2682, po2683, po2684, po2685, po2686, po2687, po2688, po2689,
    po2690, po2691, po2692, po2693, po2694, po2695, po2696, po2697, po2698,
    po2699, po2700, po2701, po2702, po2703, po2704, po2705, po2706, po2707,
    po2708, po2709, po2710, po2711, po2712, po2713, po2714, po2715, po2716,
    po2717, po2718, po2719, po2720, po2721, po2722, po2723, po2724, po2725,
    po2726, po2727, po2728, po2729, po2730, po2731, po2732, po2733, po2734,
    po2735, po2736, po2737, po2738, po2739, po2740, po2741, po2742, po2743,
    po2744, po2745, po2746, po2747, po2748, po2749, po2750, po2751, po2752,
    po2753, po2754, po2755, po2756, po2757, po2758, po2759, po2760, po2761,
    po2762, po2763, po2764, po2765, po2766, po2767, po2768, po2769, po2770,
    po2771, po2772, po2773, po2774, po2775, po2776, po2777, po2778, po2779,
    po2780, po2781, po2782, po2783, po2784, po2785, po2786, po2787, po2788,
    po2789, po2790, po2791, po2792, po2793, po2794, po2795, po2796, po2797,
    po2798, po2799, po2800, po2801, po2802, po2803, po2804, po2805, po2806,
    po2807, po2808, po2809, po2810, po2811, po2812, po2813, po2814, po2815,
    po2816, po2817, po2818, po2819, po2820, po2821, po2822, po2823, po2824,
    po2825, po2826, po2827, po2828, po2829, po2830, po2831, po2832, po2833,
    po2834, po2835, po2836, po2837, po2838, po2839, po2840, po2841, po2842,
    po2843, po2844, po2845, po2846, po2847, po2848, po2849, po2850, po2851,
    po2852, po2853, po2854, po2855, po2856, po2857, po2858, po2859, po2860,
    po2861, po2862, po2863, po2864, po2865, po2866, po2867, po2868, po2869,
    po2870, po2871, po2872, po2873, po2874, po2875, po2876, po2877, po2878,
    po2879, po2880, po2881, po2882, po2883, po2884, po2885, po2886, po2887,
    po2888, po2889, po2890, po2891, po2892, po2893, po2894, po2895, po2896,
    po2897, po2898, po2899, po2900, po2901, po2902, po2903, po2904, po2905,
    po2906, po2907, po2908, po2909, po2910, po2911, po2912, po2913, po2914,
    po2915, po2916, po2917, po2918, po2919, po2920, po2921, po2922, po2923,
    po2924, po2925, po2926, po2927, po2928, po2929, po2930, po2931, po2932,
    po2933, po2934, po2935, po2936, po2937, po2938, po2939, po2940, po2941,
    po2942, po2943, po2944, po2945, po2946, po2947, po2948, po2949, po2950,
    po2951, po2952, po2953, po2954, po2955, po2956, po2957, po2958, po2959,
    po2960, po2961, po2962, po2963, po2964, po2965, po2966, po2967, po2968,
    po2969, po2970, po2971, po2972, po2973, po2974, po2975, po2976, po2977,
    po2978, po2979, po2980, po2981, po2982, po2983, po2984, po2985, po2986,
    po2987, po2988, po2989, po2990, po2991, po2992, po2993, po2994, po2995,
    po2996, po2997, po2998, po2999, po3000, po3001, po3002, po3003, po3004,
    po3005, po3006, po3007, po3008, po3009, po3010, po3011, po3012, po3013,
    po3014, po3015, po3016, po3017, po3018, po3019, po3020, po3021, po3022,
    po3023, po3024, po3025, po3026, po3027, po3028, po3029, po3030, po3031,
    po3032, po3033, po3034, po3035, po3036, po3037, po3038, po3039, po3040,
    po3041, po3042, po3043, po3044, po3045, po3046, po3047, po3048, po3049,
    po3050, po3051, po3052, po3053, po3054, po3055, po3056, po3057, po3058,
    po3059, po3060, po3061, po3062, po3063, po3064, po3065, po3066, po3067,
    po3068, po3069, po3070, po3071, po3072, po3073, po3074, po3075, po3076,
    po3077, po3078, po3079, po3080, po3081, po3082, po3083, po3084, po3085,
    po3086, po3087, po3088, po3089, po3090, po3091, po3092, po3093, po3094,
    po3095, po3096, po3097, po3098, po3099, po3100, po3101, po3102, po3103,
    po3104, po3105, po3106, po3107, po3108, po3109, po3110, po3111, po3112,
    po3113, po3114, po3115, po3116, po3117, po3118, po3119, po3120, po3121,
    po3122, po3123, po3124, po3125, po3126, po3127, po3128, po3129, po3130,
    po3131, po3132, po3133, po3134, po3135, po3136, po3137, po3138, po3139,
    po3140, po3141, po3142, po3143, po3144, po3145, po3146, po3147, po3148,
    po3149, po3150, po3151, po3152, po3153, po3154, po3155, po3156, po3157,
    po3158, po3159, po3160, po3161, po3162, po3163, po3164, po3165, po3166,
    po3167, po3168, po3169, po3170, po3171, po3172, po3173, po3174, po3175,
    po3176, po3177, po3178, po3179, po3180, po3181, po3182, po3183, po3184,
    po3185, po3186, po3187, po3188, po3189, po3190, po3191, po3192, po3193,
    po3194, po3195, po3196, po3197, po3198, po3199, po3200, po3201, po3202,
    po3203, po3204, po3205, po3206, po3207, po3208, po3209, po3210, po3211,
    po3212, po3213, po3214, po3215, po3216, po3217, po3218, po3219, po3220,
    po3221, po3222, po3223, po3224, po3225, po3226, po3227, po3228, po3229,
    po3230, po3231, po3232, po3233, po3234, po3235, po3236, po3237, po3238,
    po3239, po3240, po3241, po3242, po3243, po3244, po3245, po3246, po3247,
    po3248, po3249, po3250, po3251, po3252, po3253, po3254, po3255, po3256,
    po3257, po3258, po3259, po3260, po3261, po3262, po3263, po3264, po3265,
    po3266, po3267, po3268, po3269, po3270, po3271, po3272, po3273, po3274,
    po3275, po3276, po3277, po3278, po3279, po3280, po3281, po3282, po3283,
    po3284, po3285, po3286, po3287, po3288, po3289, po3290, po3291, po3292,
    po3293, po3294, po3295, po3296, po3297, po3298, po3299, po3300, po3301,
    po3302, po3303, po3304, po3305, po3306, po3307, po3308, po3309, po3310,
    po3311, po3312, po3313, po3314, po3315, po3316, po3317, po3318, po3319,
    po3320, po3321, po3322, po3323, po3324, po3325, po3326, po3327, po3328,
    po3329, po3330, po3331, po3332, po3333, po3334, po3335, po3336, po3337,
    po3338, po3339, po3340, po3341, po3342, po3343, po3344, po3345, po3346,
    po3347, po3348, po3349, po3350, po3351, po3352, po3353, po3354, po3355,
    po3356, po3357, po3358, po3359, po3360, po3361, po3362, po3363, po3364,
    po3365, po3366, po3367, po3368, po3369, po3370, po3371, po3372, po3373,
    po3374, po3375, po3376, po3377, po3378, po3379, po3380, po3381, po3382,
    po3383, po3384, po3385, po3386, po3387, po3388, po3389, po3390, po3391,
    po3392, po3393, po3394, po3395, po3396, po3397, po3398, po3399, po3400,
    po3401, po3402, po3403, po3404, po3405, po3406, po3407, po3408, po3409,
    po3410, po3411, po3412, po3413, po3414, po3415, po3416, po3417, po3418,
    po3419, po3420, po3421, po3422, po3423, po3424, po3425, po3426, po3427,
    po3428, po3429, po3430, po3431, po3432, po3433, po3434, po3435, po3436,
    po3437, po3438, po3439, po3440, po3441, po3442, po3443, po3444, po3445,
    po3446, po3447, po3448, po3449, po3450, po3451, po3452, po3453, po3454,
    po3455, po3456, po3457, po3458, po3459, po3460, po3461, po3462, po3463,
    po3464, po3465, po3466, po3467, po3468, po3469, po3470, po3471, po3472,
    po3473, po3474, po3475, po3476, po3477, po3478, po3479, po3480, po3481,
    po3482, po3483, po3484, po3485, po3486, po3487, po3488, po3489, po3490,
    po3491, po3492, po3493, po3494, po3495, po3496, po3497, po3498, po3499,
    po3500, po3501, po3502, po3503, po3504, po3505, po3506, po3507, po3508,
    po3509, po3510, po3511, po3512, po3513, po3514, po3515, po3516, po3517,
    po3518, po3519, po3520, po3521, po3522, po3523, po3524, po3525, po3526,
    po3527, po3528, po3529, po3530, po3531, po3532, po3533, po3534, po3535,
    po3536, po3537, po3538, po3539, po3540, po3541, po3542, po3543, po3544,
    po3545, po3546, po3547, po3548, po3549, po3550, po3551, po3552, po3553,
    po3554, po3555, po3556, po3557, po3558, po3559, po3560, po3561, po3562,
    po3563, po3564, po3565, po3566, po3567, po3568, po3569, po3570, po3571,
    po3572, po3573, po3574, po3575, po3576, po3577, po3578, po3579, po3580,
    po3581, po3582, po3583, po3584, po3585, po3586, po3587, po3588, po3589,
    po3590, po3591, po3592, po3593, po3594, po3595, po3596, po3597, po3598,
    po3599, po3600, po3601, po3602, po3603, po3604, po3605, po3606, po3607,
    po3608, po3609, po3610, po3611, po3612, po3613, po3614, po3615, po3616,
    po3617, po3618, po3619, po3620, po3621, po3622, po3623, po3624, po3625,
    po3626, po3627, po3628, po3629, po3630, po3631, po3632, po3633, po3634,
    po3635, po3636, po3637, po3638, po3639, po3640, po3641, po3642, po3643,
    po3644, po3645, po3646, po3647, po3648, po3649, po3650, po3651, po3652,
    po3653, po3654, po3655, po3656, po3657, po3658, po3659, po3660, po3661,
    po3662, po3663, po3664, po3665, po3666, po3667, po3668, po3669, po3670,
    po3671, po3672, po3673, po3674, po3675, po3676, po3677, po3678, po3679,
    po3680, po3681, po3682, po3683, po3684, po3685, po3686, po3687, po3688,
    po3689, po3690, po3691, po3692, po3693, po3694, po3695, po3696, po3697,
    po3698, po3699, po3700, po3701, po3702, po3703, po3704, po3705, po3706,
    po3707, po3708, po3709, po3710, po3711, po3712, po3713, po3714, po3715,
    po3716, po3717, po3718, po3719, po3720, po3721, po3722, po3723, po3724,
    po3725, po3726, po3727, po3728, po3729, po3730, po3731, po3732, po3733,
    po3734, po3735, po3736, po3737, po3738, po3739, po3740, po3741, po3742,
    po3743, po3744, po3745, po3746, po3747, po3748, po3749, po3750, po3751,
    po3752, po3753, po3754, po3755, po3756, po3757, po3758, po3759, po3760,
    po3761, po3762, po3763, po3764, po3765, po3766, po3767, po3768, po3769,
    po3770, po3771, po3772, po3773, po3774, po3775, po3776, po3777, po3778,
    po3779, po3780, po3781, po3782, po3783, po3784, po3785, po3786, po3787,
    po3788, po3789, po3790, po3791, po3792, po3793, po3794, po3795, po3796,
    po3797, po3798, po3799, po3800, po3801, po3802, po3803, po3804, po3805,
    po3806, po3807, po3808, po3809, po3810, po3811, po3812, po3813, po3814,
    po3815, po3816, po3817, po3818, po3819, po3820, po3821, po3822, po3823,
    po3824, po3825, po3826, po3827, po3828, po3829, po3830, po3831, po3832,
    po3833, po3834, po3835, po3836, po3837, po3838, po3839, po3840, po3841,
    po3842, po3843, po3844, po3845, po3846, po3847, po3848, po3849, po3850,
    po3851, po3852, po3853, po3854, po3855, po3856, po3857, po3858, po3859,
    po3860, po3861, po3862, po3863, po3864, po3865, po3866, po3867, po3868,
    po3869, po3870, po3871, po3872, po3873, po3874, po3875, po3876, po3877,
    po3878, po3879, po3880, po3881, po3882, po3883, po3884, po3885, po3886,
    po3887, po3888, po3889, po3890, po3891, po3892, po3893, po3894, po3895,
    po3896, po3897, po3898, po3899, po3900, po3901, po3902, po3903, po3904,
    po3905, po3906, po3907, po3908, po3909, po3910, po3911, po3912, po3913,
    po3914, po3915, po3916, po3917, po3918, po3919, po3920, po3921, po3922,
    po3923, po3924, po3925, po3926, po3927, po3928, po3929, po3930, po3931,
    po3932, po3933, po3934, po3935, po3936, po3937, po3938, po3939, po3940,
    po3941, po3942, po3943, po3944, po3945, po3946, po3947, po3948, po3949,
    po3950, po3951, po3952;
  wire n8179, n8180, n8181, n8182, n8185, n8186, n8188, n8191, n8192, n8193,
    n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
    n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
    n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310, n8312, n8313, n8314, n8315,
    n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
    n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
    n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372, n8374, n8375, n8376, n8377,
    n8379, n8380, n8381, n8382, n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8395, n8396, n8397, n8398, n8400, n8401, n8405,
    n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8456, n8457,
    n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467,
    n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487,
    n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497,
    n8498, n8499, n8500, n8501, n8502, n8503, n8505, n8506, n8508, n8509,
    n8511, n8512, n8513, n8514, n8516, n8517, n8518, n8520, n8521, n8522,
    n8523, n8525, n8526, n8527, n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8557,
    n8558, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
    n8630, n8631, n8632, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
    n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
    n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
    n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
    n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9475, n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501,
    n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531,
    n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561,
    n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581,
    n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591,
    n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
    n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
    n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
    n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711,
    n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721,
    n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731,
    n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741,
    n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751,
    n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761,
    n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771,
    n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781,
    n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791,
    n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801,
    n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811,
    n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831,
    n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841,
    n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851,
    n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861,
    n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878, n9880, n9881, n9882, n9883,
    n9884, n9886, n9887, n9888, n9889, n9890, n9892, n9893, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9903, n9904, n9905, n9906, n9907,
    n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917,
    n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927,
    n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937,
    n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947,
    n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957,
    n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967,
    n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977,
    n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987,
    n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997,
    n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006,
    n10007, n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
    n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
    n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
    n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
    n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
    n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
    n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
    n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077, n10078,
    n10079, n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
    n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
    n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
    n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
    n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
    n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149, n10150,
    n10151, n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
    n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
    n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
    n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221, n10222,
    n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
    n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
    n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
    n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
    n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
    n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
    n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
    n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
    n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
    n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
    n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
    n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10698, n10699, n10701, n10702, n10704,
    n10706, n10707, n10708, n10709, n10711, n10712, n10713, n10715, n10717,
    n10719, n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
    n10728, n10729, n10730, n10732, n10733, n10734, n10735, n10736, n10737,
    n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
    n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
    n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763, n10764,
    n10765, n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
    n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781, n10782,
    n10783, n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
    n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
    n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
    n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
    n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
    n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
    n10837, n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
    n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10854,
    n10855, n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
    n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
    n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
    n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
    n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
    n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
    n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
    n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925, n10926,
    n10927, n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
    n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
    n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
    n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
    n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
    n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
    n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
    n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
    n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
    n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
    n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
    n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
    n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
    n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
    n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
    n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
    n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
    n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213, n11214,
    n11215, n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
    n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
    n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
    n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
    n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
    n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
    n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
    n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285, n11286,
    n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
    n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
    n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
    n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
    n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
    n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
    n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
    n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
    n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
    n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
    n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
    n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
    n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502,
    n11503, n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
    n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
    n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
    n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
    n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
    n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
    n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
    n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
    n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
    n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
    n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
    n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
    n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
    n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
    n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
    n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
    n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
    n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
    n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717, n11718,
    n11719, n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
    n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
    n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
    n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
    n11755, n11756, n11757, n11759, n11760, n11761, n11762, n11763, n11764,
    n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
    n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781, n11782,
    n11783, n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
    n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
    n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
    n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
    n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
    n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
    n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853, n11854,
    n11855, n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
    n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
    n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
    n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925, n11926,
    n11927, n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
    n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
    n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
    n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
    n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997, n11998,
    n11999, n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
    n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
    n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
    n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
    n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
    n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
    n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069, n12070,
    n12071, n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
    n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
    n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
    n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
    n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
    n12125, n12126, n12127, n12128, n12129, n12130, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
    n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
    n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
    n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
    n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
    n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
    n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
    n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
    n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
    n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
    n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
    n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
    n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
    n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
    n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
    n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
    n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
    n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
    n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
    n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
    n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
    n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
    n12757, n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
    n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773, n12774,
    n12775, n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
    n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
    n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
    n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
    n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
    n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827, n12828,
    n12829, n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
    n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845, n12846,
    n12847, n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
    n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
    n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
    n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
    n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
    n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899, n12900,
    n12901, n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
    n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917, n12918,
    n12919, n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
    n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
    n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
    n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
    n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
    n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971, n12972,
    n12973, n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
    n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989, n12990,
    n12991, n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
    n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
    n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
    n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
    n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
    n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043, n13044,
    n13045, n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
    n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061, n13062,
    n13063, n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
    n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
    n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
    n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
    n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
    n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115, n13116,
    n13117, n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
    n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134,
    n13135, n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
    n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
    n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
    n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
    n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
    n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205, n13206,
    n13207, n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
    n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
    n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
    n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
    n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259, n13260,
    n13261, n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
    n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277, n13278,
    n13279, n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
    n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
    n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
    n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
    n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
    n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331, n13332,
    n13333, n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
    n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
    n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
    n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13408, n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
    n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
    n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
    n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467, n13468,
    n13469, n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
    n13478, n13479, n13480, n13482, n13483, n13484, n13485, n13486, n13487,
    n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
    n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
    n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
    n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
    n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
    n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
    n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
    n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
    n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
    n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
    n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
    n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
    n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
    n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
    n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
    n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
    n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
    n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
    n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
    n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
    n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
    n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
    n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
    n14182, n14183, n14184, n14185, n14186, n14187, n14189, n14190, n14191,
    n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
    n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
    n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
    n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, n14236,
    n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
    n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254,
    n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
    n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
    n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
    n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
    n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
    n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, n14308,
    n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
    n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, n14326,
    n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
    n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
    n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
    n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
    n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
    n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, n14380,
    n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
    n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, n14398,
    n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
    n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
    n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
    n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
    n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
    n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, n14452,
    n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, n14470,
    n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
    n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
    n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, n14524,
    n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, n14542,
    n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
    n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
    n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, n14596,
    n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, n14614,
    n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
    n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
    n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, n14668,
    n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, n14686,
    n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
    n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
    n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, n14740,
    n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, n14758,
    n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
    n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
    n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, n14812,
    n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
    n14823, n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
    n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
    n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
    n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
    n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
    n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
    n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
    n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
    n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
    n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
    n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
    n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
    n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
    n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
    n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
    n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
    n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
    n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
    n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
    n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
    n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
    n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
    n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
    n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
    n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
    n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
    n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
    n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
    n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
    n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
    n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
    n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
    n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
    n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
    n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458, n15460, n15461, n15462,
    n15463, n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
    n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
    n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15496, n15497, n15499, n15500, n15501,
    n15502, n15504, n15506, n15507, n15508, n15510, n15511, n15513, n15515,
    n15517, n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
    n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15534, n15535,
    n15536, n15537, n15538, n15539, n15540, n15542, n15543, n15546, n15547,
    n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555, n15556,
    n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
    n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573, n15574,
    n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
    n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
    n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
    n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
    n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
    n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627, n15628,
    n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
    n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
    n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
    n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
    n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717, n15718,
    n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
    n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
    n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
    n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
    n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771, n15772,
    n15773, n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
    n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789, n15790,
    n15791, n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
    n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
    n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
    n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
    n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
    n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
    n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
    n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
    n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
    n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
    n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
    n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987, n15988,
    n15989, n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
    n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006,
    n16007, n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
    n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
    n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
    n16034, n16035, n16036, n16037, n16039, n16040, n16041, n16042, n16043,
    n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
    n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062,
    n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
    n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
    n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
    n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
    n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
    n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116,
    n16117, n16118, n16119, n16120, n16121, n16123, n16124, n16125, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
    n16138, n16139, n16140, n16141, n16142, n16143, n16145, n16146, n16147,
    n16148, n16149, n16150, n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16187, n16189, n16190, n16192, n16194, n16195, n16196, n16197,
    n16199, n16201, n16202, n16204, n16206, n16207, n16208, n16209, n16210,
    n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245, n16247, n16248, n16249,
    n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16259,
    n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278,
    n16279, n16280, n16281, n16283, n16284, n16285, n16286, n16287, n16288,
    n16289, n16290, n16291, n16292, n16293, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16307, n16308,
    n16309, n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
    n16319, n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
    n16328, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
    n16338, n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
    n16348, n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
    n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
    n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
    n16404, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422,
    n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
    n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
    n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
    n16451, n16452, n16453, n16454, n16455, n16456, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
    n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
    n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
    n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538, n16540, n16541, n16542,
    n16543, n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
    n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
    n16570, n16571, n16572, n16573, n16574, n16576, n16577, n16578, n16579,
    n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587, n16588,
    n16589, n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
    n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16608, n16609, n16610, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
    n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
    n16644, n16645, n16646, n16648, n16649, n16650, n16651, n16652, n16653,
    n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661, n16662,
    n16663, n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
    n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
    n16681, n16682, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
    n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707, n16708,
    n16709, n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
    n16718, n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
    n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
    n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
    n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764,
    n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
    n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782,
    n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16792,
    n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
    n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16828, n16829,
    n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862, n16864, n16865, n16866,
    n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
    n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883, n16884,
    n16885, n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
    n16894, n16895, n16896, n16897, n16898, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
    n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
    n16931, n16932, n16933, n16934, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
    n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
    n16968, n16969, n16970, n16972, n16973, n16974, n16975, n16976, n16977,
    n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
    n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
    n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003, n17004,
    n17005, n17006, n17008, n17009, n17010, n17011, n17012, n17013, n17014,
    n17015, n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
    n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
    n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
    n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
    n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
    n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067, n17068,
    n17069, n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
    n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085, n17086,
    n17087, n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
    n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
    n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
    n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
    n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139, n17140,
    n17141, n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
    n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157, n17158,
    n17159, n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
    n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
    n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
    n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
    n17204, n17205, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
    n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
    n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
    n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
    n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
    n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
    n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
    n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
    n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
    n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
    n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
    n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17402, n17403,
    n17404, n17405, n17407, n17408, n17409, n17411, n17412, n17413, n17415,
    n17416, n17417, n17419, n17420, n17421, n17423, n17424, n17425, n17427,
    n17428, n17429, n17431, n17432, n17433, n17435, n17438, n17442, n17445,
    n17447, n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17456,
    n17457, n17458, n17459, n17460, n17461, n17463, n17464, n17465, n17466,
    n17467, n17468, n17470, n17471, n17472, n17473, n17474, n17475, n17477,
    n17478, n17479, n17480, n17481, n17482, n17484, n17485, n17486, n17487,
    n17488, n17489, n17491, n17492, n17493, n17494, n17495, n17496, n17498,
    n17499, n17500, n17501, n17502, n17503, n17505, n17506, n17507, n17508,
    n17509, n17510, n17512, n17513, n17514, n17515, n17516, n17517, n17519,
    n17520, n17521, n17522, n17523, n17524, n17526, n17527, n17528, n17529,
    n17530, n17531, n17533, n17534, n17535, n17536, n17537, n17538, n17540,
    n17541, n17542, n17543, n17544, n17545, n17547, n17548, n17549, n17550,
    n17551, n17552, n17554, n17555, n17556, n17557, n17558, n17559, n17561,
    n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576, n17578, n17579, n17580,
    n17581, n17582, n17583, n17584, n17585, n17586, n17588, n17589, n17590,
    n17591, n17592, n17593, n17594, n17595, n17596, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606, n17608, n17609, n17610,
    n17611, n17612, n17613, n17614, n17615, n17616, n17618, n17619, n17620,
    n17621, n17622, n17623, n17624, n17625, n17626, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636, n17638, n17639, n17640,
    n17641, n17642, n17643, n17644, n17645, n17646, n17648, n17649, n17650,
    n17651, n17652, n17653, n17654, n17655, n17656, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666, n17668, n17669, n17670,
    n17671, n17672, n17673, n17674, n17675, n17676, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696, n17698, n17699, n17700,
    n17701, n17702, n17703, n17704, n17705, n17706, n17708, n17709, n17710,
    n17711, n17712, n17713, n17714, n17715, n17716, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726, n17728, n17729, n17730,
    n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
    n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747, n17748,
    n17749, n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
    n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
    n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
    n17776, n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
    n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
    n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
    n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
    n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
    n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
    n17886, n17887, n17888, n17889, n17890, n17891, n17893, n17894, n17895,
    n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
    n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
    n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
    n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
    n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939, n17940,
    n17941, n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
    n17950, n17951, n17952, n17954, n17955, n17956, n17957, n17958, n17959,
    n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
    n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
    n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
    n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003, n18004,
    n18005, n18006, n18007, n18008, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
    n18024, n18025, n18026, n18027, n18029, n18030, n18031, n18032, n18033,
    n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
    n18043, n18044, n18045, n18046, n18048, n18049, n18050, n18051, n18052,
    n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
    n18062, n18063, n18064, n18065, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18086, n18087, n18088, n18089, n18090,
    n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
    n18100, n18101, n18102, n18103, n18105, n18106, n18107, n18108, n18109,
    n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
    n18138, n18139, n18140, n18141, n18143, n18144, n18145, n18146, n18147,
    n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
    n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173, n18174,
    n18175, n18176, n18177, n18178, n18179, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
    n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
    n18212, n18213, n18214, n18215, n18216, n18217, n18219, n18220, n18221,
    n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
    n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18257, n18258,
    n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
    n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276,
    n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
    n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18295,
    n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
    n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
    n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
    n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
    n18333, n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
    n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
    n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
    n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18390, n18391, n18392, n18393, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405, n18406,
    n18407, n18408, n18409, n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
    n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
    n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18458, n18459, n18460, n18461,
    n18463, n18464, n18465, n18466, n18467, n18468, n18469, n18470, n18471,
    n18472, n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
    n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
    n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
    n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
    n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515, n18516,
    n18517, n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
    n18526, n18527, n18528, n18529, n18530, n18532, n18533, n18534, n18535,
    n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18603, n18605, n18606, n18607, n18608, n18610,
    n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627, n18628,
    n18629, n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645, n18646,
    n18647, n18648, n18649, n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
    n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18676, n18677, n18678, n18679, n18681, n18682, n18683, n18684,
    n18685, n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
    n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702,
    n18703, n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711,
    n18712, n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
    n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
    n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
    n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18748,
    n18749, n18750, n18751, n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
    n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
    n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
    n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, n18812,
    n18813, n18814, n18815, n18816, n18818, n18819, n18820, n18821, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
    n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
    n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867, n18868,
    n18869, n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885, n18886,
    n18888, n18889, n18890, n18891, n18893, n18894, n18895, n18896, n18897,
    n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
    n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
    n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923, n18924,
    n18925, n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
    n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948, n18949, n18950, n18951,
    n18952, n18953, n18954, n18956, n18957, n18958, n18959, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
    n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
    n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004, n19005, n19006, n19007,
    n19008, n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022, n19024, n19025, n19026,
    n19027, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036,
    n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
    n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054,
    n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063,
    n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
    n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
    n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
    n19091, n19092, n19093, n19094, n19095, n19096, n19098, n19099, n19100,
    n19101, n19103, n19104, n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116, n19117, n19118, n19119,
    n19120, n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
    n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
    n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
    n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
    n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163, n19164,
    n19165, n19166, n19167, n19168, n19169, n19171, n19172, n19173, n19174,
    n19176, n19177, n19178, n19179, n19180, n19182, n19183, n19184, n19185,
    n19186, n19188, n19189, n19190, n19191, n19192, n19194, n19195, n19196,
    n19197, n19198, n19200, n19201, n19202, n19203, n19204, n19206, n19207,
    n19208, n19209, n19210, n19212, n19213, n19214, n19215, n19216, n19218,
    n19219, n19220, n19221, n19222, n19224, n19225, n19226, n19227, n19228,
    n19230, n19231, n19232, n19233, n19234, n19236, n19237, n19238, n19239,
    n19240, n19242, n19243, n19244, n19245, n19246, n19248, n19249, n19250,
    n19251, n19252, n19254, n19255, n19256, n19257, n19258, n19260, n19261,
    n19262, n19263, n19264, n19266, n19267, n19268, n19269, n19270, n19272,
    n19273, n19274, n19275, n19276, n19278, n19279, n19280, n19281, n19282,
    n19284, n19285, n19286, n19287, n19288, n19290, n19291, n19292, n19293,
    n19294, n19296, n19297, n19298, n19299, n19300, n19302, n19303, n19304,
    n19305, n19306, n19308, n19309, n19310, n19311, n19312, n19314, n19315,
    n19316, n19317, n19318, n19320, n19321, n19323, n19324, n19326, n19327,
    n19329, n19330, n19332, n19333, n19335, n19336, n19337, n19339, n19340,
    n19341, n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350,
    n19351, n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359,
    n19360, n19361, n19362, n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
    n19380, n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
    n19391, n19392, n19393, n19394, n19395, n19396, n19397, n19398, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19409, n19410,
    n19411, n19412, n19413, n19414, n19415, n19416, n19418, n19419, n19420,
    n19421, n19422, n19423, n19424, n19425, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19436, n19437, n19438, n19439, n19440,
    n19441, n19442, n19443, n19445, n19446, n19448, n19450, n19451, n19452,
    n19453, n19454, n19455, n19456, n19457, n19458, n19459, n19461, n19462,
    n19463, n19464, n19465, n19467, n19468, n19469, n19470, n19471, n19473,
    n19474, n19475, n19476, n19477, n19479, n19480, n19481, n19482, n19483,
    n19485, n19486, n19487, n19488, n19489, n19491, n19492, n19493, n19494,
    n19495, n19497, n19498, n19499, n19500, n19501, n19503, n19504, n19505,
    n19506, n19507, n19509, n19510, n19511, n19512, n19513, n19515, n19516,
    n19517, n19518, n19519, n19521, n19522, n19523, n19524, n19525, n19527,
    n19528, n19529, n19530, n19531, n19533, n19534, n19535, n19536, n19537,
    n19539, n19540, n19542, n19543, n19544, n19545, n19546, n19547, n19548,
    n19549, n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
    n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566,
    n19567, n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
    n19576, n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
    n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
    n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
    n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
    n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620,
    n19621, n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
    n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
    n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647,
    n19648, n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
    n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
    n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
    n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
    n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692,
    n19693, n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
    n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710,
    n19711, n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719,
    n19720, n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
    n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
    n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
    n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
    n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764,
    n19765, n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
    n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782,
    n19783, n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791,
    n19792, n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
    n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
    n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
    n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
    n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836,
    n19837, n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
    n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854,
    n19855, n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
    n19864, n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
    n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
    n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
    n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
    n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908,
    n19909, n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
    n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926,
    n19927, n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935,
    n19936, n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944,
    n19945, n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
    n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
    n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
    n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980,
    n19981, n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
    n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998,
    n19999, n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007,
    n20008, n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016,
    n20017, n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
    n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
    n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
    n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052,
    n20053, n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
    n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
    n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079,
    n20080, n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088,
    n20089, n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
    n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
    n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
    n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124,
    n20125, n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
    n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142,
    n20143, n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151,
    n20152, n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160,
    n20161, n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
    n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
    n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
    n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196,
    n20197, n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
    n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214,
    n20215, n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223,
    n20224, n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232,
    n20233, n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
    n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
    n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
    n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
    n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286,
    n20287, n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295,
    n20296, n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304,
    n20305, n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
    n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
    n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
    n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340,
    n20341, n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
    n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358,
    n20359, n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367,
    n20368, n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376,
    n20377, n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
    n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
    n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
    n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412,
    n20413, n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
    n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430,
    n20431, n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439,
    n20440, n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448,
    n20449, n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
    n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
    n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
    n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484,
    n20485, n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
    n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502,
    n20503, n20504, n20505, n20506, n20507, n20508, n20509, n20512, n20513,
    n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
    n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
    n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, n20567,
    n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
    n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
    n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
    n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, n20639,
    n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
    n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
    n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
    n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, n20711,
    n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
    n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
    n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
    n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, n20783,
    n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
    n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
    n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
    n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, n20855,
    n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
    n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
    n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
    n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, n20927,
    n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
    n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
    n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
    n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, n20999,
    n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
    n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
    n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
    n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, n21071,
    n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
    n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
    n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
    n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, n21143,
    n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
    n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
    n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
    n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, n21215,
    n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
    n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
    n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
    n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, n21287,
    n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
    n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
    n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
    n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, n21359,
    n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
    n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
    n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, n21431,
    n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
    n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
    n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, n21503,
    n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
    n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
    n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
    n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, n21575,
    n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
    n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
    n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, n21620,
    n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
    n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, n21647,
    n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
    n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
    n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, n21692,
    n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
    n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, n21710,
    n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, n21719,
    n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, n21728,
    n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
    n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
    n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
    n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, n21764,
    n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
    n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, n21782,
    n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, n21791,
    n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, n21800,
    n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
    n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
    n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, n21836,
    n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
    n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, n21854,
    n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, n21863,
    n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, n21872,
    n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
    n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
    n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
    n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, n21908,
    n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
    n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, n21935,
    n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
    n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
    n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
    n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
    n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, n22007,
    n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
    n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
    n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
    n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, n22079,
    n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
    n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
    n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133,
    n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, n22151,
    n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, n22160,
    n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
    n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
    n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
    n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, n22214,
    n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, n22223,
    n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, n22232,
    n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
    n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
    n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
    n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277,
    n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, n22295,
    n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
    n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
    n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
    n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, n22358,
    n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, n22367,
    n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
    n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
    n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421,
    n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, n22439,
    n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, n22448,
    n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
    n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
    n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, n22484,
    n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493,
    n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, n22502,
    n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, n22511,
    n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
    n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
    n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
    n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580, n22581, n22582, n22583,
    n22584, n22585, n22586, n22587, n22588, n22589, n22590, n22591, n22592,
    n22593, n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
    n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
    n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
    n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645, n22646,
    n22647, n22648, n22649, n22650, n22651, n22652, n22653, n22654, n22655,
    n22656, n22657, n22658, n22659, n22660, n22661, n22662, n22663, n22664,
    n22665, n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
    n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
    n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
    n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
    n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
    n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
    n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
    n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
    n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
    n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
    n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
    n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
    n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868, n22869, n22870, n22871,
    n22872, n22873, n22874, n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
    n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
    n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
    n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940, n22941, n22942, n22943,
    n22944, n22945, n22946, n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
    n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
    n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
    n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012, n23013, n23014, n23015,
    n23016, n23017, n23018, n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
    n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
    n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
    n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086, n23087,
    n23088, n23089, n23090, n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
    n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
    n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
    n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158, n23159,
    n23160, n23161, n23162, n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
    n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
    n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
    n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230, n23231,
    n23232, n23233, n23234, n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
    n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
    n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
    n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302, n23303,
    n23304, n23305, n23306, n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
    n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
    n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
    n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374, n23375,
    n23376, n23377, n23378, n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
    n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
    n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429,
    n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446, n23447,
    n23448, n23449, n23450, n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
    n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
    n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
    n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518, n23519,
    n23520, n23521, n23522, n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
    n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
    n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563, n23564,
    n23565, n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
    n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582,
    n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590, n23591,
    n23592, n23593, n23594, n23595, n23596, n23597, n23598, n23599, n23600,
    n23601, n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
    n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
    n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
    n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662, n23663,
    n23664, n23665, n23666, n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
    n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
    n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
    n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734, n23735,
    n23736, n23737, n23738, n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
    n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
    n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
    n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806, n23807,
    n23808, n23809, n23810, n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
    n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
    n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
    n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878, n23879,
    n23880, n23881, n23882, n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
    n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
    n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
    n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948, n23949, n23950, n23951,
    n23952, n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
    n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
    n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
    n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020, n24021, n24022, n24023,
    n24024, n24025, n24026, n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
    n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
    n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
    n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092, n24093, n24094, n24095,
    n24096, n24097, n24098, n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
    n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
    n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
    n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164, n24165, n24166, n24167,
    n24168, n24169, n24170, n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
    n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
    n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
    n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238, n24239,
    n24240, n24241, n24242, n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
    n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24275, n24276,
    n24277, n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285,
    n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294,
    n24295, n24296, n24298, n24299, n24300, n24301, n24302, n24303, n24304,
    n24305, n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
    n24323, n24324, n24325, n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338, n24340, n24341, n24342,
    n24344, n24345, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
    n24426, n24427, n24428, n24430, n24431, n24432, n24433, n24434, n24435,
    n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443, n24444,
    n24445, n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
    n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462, n24463,
    n24464, n24465, n24466, n24468, n24469, n24471, n24472, n24473, n24474,
    n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
    n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491, n24492,
    n24493, n24494, n24495, n24497, n24498, n24499, n24500, n24501, n24502,
    n24503, n24504, n24505, n24506, n24507, n24508, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
    n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
    n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547, n24548,
    n24549, n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
    n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
    n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574, n24575,
    n24576, n24577, n24578, n24579, n24580, n24581, n24582, n24583, n24584,
    n24585, n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
    n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
    n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
    n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619, n24620,
    n24621, n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
    n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637, n24638,
    n24639, n24640, n24641, n24642, n24643, n24644, n24645, n24646, n24647,
    n24648, n24649, n24650, n24651, n24652, n24653, n24654, n24655, n24656,
    n24657, n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691, n24692,
    n24693, n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
    n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709, n24710,
    n24711, n24712, n24713, n24714, n24715, n24716, n24717, n24718, n24719,
    n24720, n24721, n24722, n24723, n24724, n24725, n24726, n24727, n24728,
    n24729, n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
    n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
    n24747, n24748, n24749, n24750, n24751, n24753, n24754, n24755, n24756,
    n24757, n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765,
    n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773, n24774,
    n24775, n24776, n24778, n24779, n24780, n24781, n24782, n24783, n24784,
    n24785, n24786, n24787, n24788, n24789, n24791, n24792, n24793, n24794,
    n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24804,
    n24805, n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
    n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821, n24822,
    n24823, n24824, n24825, n24826, n24827, n24828, n24829, n24830, n24831,
    n24832, n24833, n24834, n24835, n24836, n24837, n24838, n24839, n24840,
    n24841, n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
    n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
    n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
    n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875, n24876,
    n24877, n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
    n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893, n24894,
    n24895, n24896, n24897, n24898, n24899, n24900, n24901, n24902, n24903,
    n24904, n24905, n24906, n24907, n24908, n24909, n24910, n24911, n24912,
    n24913, n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
    n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
    n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
    n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947, n24948,
    n24949, n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957,
    n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972, n24973, n24974, n24975,
    n24976, n24977, n24978, n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
    n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
    n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019, n25020,
    n25021, n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029,
    n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037, n25038,
    n25039, n25040, n25041, n25042, n25043, n25044, n25045, n25046, n25047,
    n25048, n25049, n25050, n25051, n25052, n25053, n25054, n25055, n25056,
    n25057, n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
    n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
    n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
    n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091, n25092,
    n25093, n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
    n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109, n25110,
    n25111, n25112, n25113, n25114, n25115, n25116, n25117, n25118, n25119,
    n25120, n25121, n25122, n25123, n25124, n25125, n25126, n25127, n25128,
    n25129, n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
    n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
    n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
    n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163, n25164,
    n25165, n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
    n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181, n25182,
    n25183, n25184, n25185, n25186, n25187, n25188, n25189, n25190, n25191,
    n25192, n25193, n25194, n25195, n25196, n25197, n25198, n25199, n25200,
    n25201, n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
    n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
    n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
    n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235, n25236,
    n25237, n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245,
    n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253, n25254,
    n25255, n25256, n25257, n25258, n25259, n25260, n25261, n25262, n25263,
    n25264, n25265, n25266, n25267, n25268, n25269, n25270, n25271, n25272,
    n25273, n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
    n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
    n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
    n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307, n25308,
    n25309, n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317,
    n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325, n25326,
    n25327, n25328, n25329, n25330, n25331, n25332, n25333, n25334, n25335,
    n25336, n25337, n25338, n25339, n25340, n25341, n25342, n25343, n25344,
    n25345, n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
    n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
    n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
    n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379, n25380,
    n25381, n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389,
    n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397, n25398,
    n25399, n25400, n25401, n25402, n25403, n25404, n25405, n25406, n25407,
    n25408, n25409, n25410, n25411, n25412, n25413, n25414, n25415, n25416,
    n25417, n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
    n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
    n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
    n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451, n25452,
    n25453, n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461,
    n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469, n25470,
    n25471, n25472, n25473, n25474, n25475, n25476, n25477, n25478, n25479,
    n25480, n25481, n25482, n25483, n25484, n25485, n25486, n25487, n25488,
    n25489, n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
    n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
    n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
    n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523, n25524,
    n25525, n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
    n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541, n25542,
    n25543, n25544, n25545, n25546, n25547, n25548, n25549, n25550, n25551,
    n25552, n25553, n25554, n25555, n25556, n25557, n25558, n25559, n25560,
    n25561, n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
    n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
    n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
    n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595, n25596,
    n25597, n25598, n25599, n25600, n25601, n25602, n25603, n25604, n25605,
    n25606, n25607, n25608, n25609, n25610, n25611, n25612, n25613, n25614,
    n25615, n25616, n25617, n25618, n25620, n25621, n25622, n25623, n25624,
    n25625, n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25634,
    n25635, n25637, n25638, n25639, n25640, n25641, n25642, n25643, n25644,
    n25645, n25646, n25647, n25648, n25649, n25650, n25651, n25652, n25653,
    n25654, n25655, n25656, n25657, n25658, n25659, n25660, n25661, n25663,
    n25664, n25665, n25666, n25667, n25668, n25669, n25670, n25671, n25672,
    n25673, n25675, n25676, n25678, n25679, n25681, n25682, n25683, n25684,
    n25685, n25686, n25687, n25688, n25689, n25690, n25691, n25692, n25693,
    n25694, n25695, n25696, n25697, n25698, n25699, n25700, n25701, n25702,
    n25703, n25704, n25705, n25706, n25708, n25709, n25710, n25711, n25712,
    n25713, n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
    n25722, n25723, n25724, n25725, n25727, n25728, n25729, n25730, n25731,
    n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749, n25750,
    n25751, n25753, n25754, n25755, n25756, n25757, n25758, n25759, n25760,
    n25761, n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
    n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
    n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
    n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795, n25796,
    n25797, n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
    n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813, n25814,
    n25815, n25816, n25817, n25818, n25819, n25820, n25821, n25822, n25823,
    n25824, n25825, n25826, n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
    n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
    n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867, n25868,
    n25869, n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
    n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892, n25893, n25894, n25895,
    n25896, n25897, n25898, n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
    n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
    n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
    n25950, n25951, n25952, n25953, n25954, n25955, n25956, n25957, n25958,
    n25959, n25960, n25961, n25962, n25963, n25964, n25965, n25966, n25967,
    n25968, n25969, n25970, n25971, n25972, n25973, n25974, n25975, n25976,
    n25977, n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25986,
    n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25995, n25996,
    n25997, n25998, n25999, n26000, n26001, n26002, n26003, n26004, n26005,
    n26006, n26007, n26008, n26009, n26010, n26011, n26012, n26013, n26014,
    n26015, n26016, n26017, n26018, n26019, n26020, n26021, n26022, n26023,
    n26024, n26025, n26026, n26027, n26028, n26029, n26030, n26031, n26032,
    n26033, n26034, n26035, n26037, n26038, n26039, n26040, n26041, n26042,
    n26043, n26044, n26045, n26046, n26047, n26048, n26050, n26051, n26052,
    n26053, n26055, n26056, n26057, n26058, n26060, n26062, n26063, n26064,
    n26065, n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
    n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
    n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
    n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099, n26100,
    n26101, n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
    n26110, n26111, n26112, n26113, n26114, n26115, n26116, n26117, n26118,
    n26119, n26120, n26121, n26122, n26123, n26124, n26125, n26126, n26127,
    n26128, n26129, n26130, n26131, n26132, n26133, n26134, n26135, n26136,
    n26137, n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
    n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
    n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
    n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171, n26172,
    n26173, n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
    n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189, n26190,
    n26191, n26192, n26193, n26194, n26195, n26196, n26197, n26198, n26199,
    n26200, n26201, n26202, n26203, n26204, n26205, n26206, n26207, n26208,
    n26209, n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
    n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
    n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
    n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243, n26244,
    n26245, n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
    n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261, n26262,
    n26263, n26264, n26265, n26266, n26267, n26268, n26269, n26270, n26271,
    n26272, n26273, n26274, n26275, n26276, n26277, n26278, n26279, n26280,
    n26281, n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
    n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
    n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
    n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315, n26316,
    n26317, n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
    n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333, n26334,
    n26335, n26336, n26337, n26338, n26339, n26340, n26341, n26342, n26343,
    n26344, n26345, n26346, n26347, n26348, n26349, n26350, n26351, n26352,
    n26353, n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
    n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
    n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
    n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26388, n26389,
    n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397, n26398,
    n26399, n26400, n26401, n26402, n26403, n26404, n26405, n26406, n26407,
    n26408, n26409, n26410, n26411, n26412, n26413, n26414, n26415, n26416,
    n26417, n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
    n26426, n26427, n26428, n26429, n26430, n26432, n26433, n26434, n26435,
    n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443, n26444,
    n26445, n26446, n26447, n26448, n26449, n26450, n26451, n26452, n26453,
    n26454, n26455, n26456, n26457, n26458, n26459, n26460, n26461, n26462,
    n26463, n26464, n26465, n26466, n26467, n26468, n26469, n26470, n26471,
    n26472, n26473, n26474, n26475, n26476, n26477, n26478, n26479, n26480,
    n26481, n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
    n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
    n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
    n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515, n26516,
    n26517, n26518, n26519, n26520, n26521, n26522, n26523, n26524, n26525,
    n26526, n26527, n26528, n26529, n26530, n26531, n26532, n26533, n26534,
    n26535, n26536, n26537, n26538, n26539, n26540, n26541, n26542, n26543,
    n26544, n26545, n26546, n26547, n26548, n26549, n26550, n26551, n26552,
    n26553, n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
    n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
    n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
    n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587, n26588,
    n26589, n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
    n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605, n26606,
    n26607, n26608, n26609, n26610, n26611, n26612, n26613, n26614, n26615,
    n26616, n26617, n26618, n26619, n26620, n26621, n26622, n26623, n26624,
    n26625, n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
    n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
    n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
    n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659, n26660,
    n26661, n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669,
    n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677, n26678,
    n26679, n26680, n26681, n26682, n26683, n26684, n26685, n26686, n26687,
    n26688, n26689, n26690, n26691, n26692, n26693, n26694, n26695, n26696,
    n26697, n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
    n26706, n26707, n26708, n26709, n26710, n26712, n26713, n26714, n26715,
    n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723, n26724,
    n26725, n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
    n26734, n26735, n26736, n26737, n26738, n26739, n26740, n26741, n26742,
    n26743, n26744, n26745, n26746, n26747, n26748, n26749, n26750, n26751,
    n26752, n26753, n26754, n26755, n26756, n26757, n26758, n26759, n26760,
    n26761, n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
    n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
    n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
    n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795, n26796,
    n26797, n26798, n26799, n26800, n26801, n26802, n26803, n26804, n26805,
    n26806, n26807, n26808, n26809, n26810, n26811, n26812, n26813, n26814,
    n26815, n26816, n26817, n26818, n26819, n26820, n26821, n26822, n26823,
    n26824, n26825, n26826, n26827, n26828, n26829, n26830, n26831, n26832,
    n26833, n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
    n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
    n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
    n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867, n26868,
    n26869, n26870, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
    n26878, n26879, n26880, n26881, n26882, n26883, n26884, n26885, n26886,
    n26887, n26888, n26889, n26890, n26891, n26892, n26893, n26894, n26895,
    n26896, n26897, n26898, n26899, n26900, n26901, n26902, n26903, n26904,
    n26905, n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
    n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
    n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
    n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939, n26940,
    n26941, n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
    n26950, n26952, n26953, n26954, n26955, n26956, n26957, n26958, n26959,
    n26960, n26961, n26962, n26963, n26964, n26965, n26966, n26967, n26968,
    n26969, n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
    n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
    n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
    n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003, n27004,
    n27005, n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
    n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021, n27022,
    n27023, n27024, n27025, n27026, n27027, n27028, n27029, n27030, n27031,
    n27032, n27033, n27034, n27035, n27036, n27037, n27038, n27039, n27040,
    n27041, n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
    n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
    n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
    n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075, n27076,
    n27077, n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
    n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093, n27094,
    n27095, n27096, n27097, n27098, n27099, n27100, n27101, n27102, n27103,
    n27104, n27105, n27106, n27107, n27108, n27109, n27110, n27111, n27112,
    n27113, n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
    n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
    n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
    n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147, n27148,
    n27149, n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
    n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165, n27166,
    n27167, n27168, n27169, n27170, n27171, n27172, n27173, n27174, n27175,
    n27176, n27177, n27178, n27179, n27180, n27181, n27182, n27183, n27184,
    n27185, n27186, n27187, n27189, n27190, n27191, n27192, n27193, n27194,
    n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
    n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211, n27212,
    n27213, n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
    n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229, n27230,
    n27231, n27232, n27233, n27234, n27235, n27236, n27237, n27238, n27239,
    n27240, n27241, n27242, n27243, n27244, n27245, n27246, n27247, n27248,
    n27249, n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
    n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
    n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
    n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283, n27284,
    n27285, n27286, n27287, n27288, n27289, n27290, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301, n27302,
    n27303, n27304, n27305, n27306, n27307, n27308, n27309, n27310, n27311,
    n27312, n27313, n27314, n27315, n27316, n27317, n27318, n27319, n27320,
    n27321, n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
    n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
    n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
    n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355, n27356,
    n27357, n27358, n27359, n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371, n27372, n27373, n27374,
    n27375, n27376, n27377, n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389, n27390, n27391, n27392,
    n27393, n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
    n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427, n27428,
    n27429, n27430, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443, n27444, n27445, n27446,
    n27447, n27448, n27449, n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461, n27462, n27463, n27464,
    n27465, n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
    n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
    n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
    n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499, n27500,
    n27501, n27502, n27503, n27504, n27505, n27506, n27508, n27509, n27510,
    n27511, n27512, n27513, n27514, n27515, n27517, n27518, n27519, n27520,
    n27521, n27522, n27523, n27524, n27526, n27527, n27528, n27529, n27530,
    n27531, n27532, n27533, n27535, n27536, n27537, n27538, n27539, n27540,
    n27541, n27542, n27544, n27545, n27547, n27548, n27550, n27551, n27553,
    n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
    n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
    n27572, n27573, n27574, n27575, n27576, n27578, n27579, n27580, n27581,
    n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589, n27590,
    n27591, n27592, n27593, n27594, n27595, n27596, n27597, n27598, n27599,
    n27600, n27601, n27602, n27603, n27604, n27605, n27606, n27607, n27608,
    n27609, n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
    n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
    n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
    n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643, n27644,
    n27645, n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
    n27654, n27655, n27656, n27657, n27658, n27659, n27660, n27661, n27662,
    n27663, n27664, n27665, n27666, n27667, n27668, n27669, n27670, n27671,
    n27672, n27673, n27674, n27675, n27676, n27677, n27678, n27679, n27680,
    n27681, n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
    n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
    n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
    n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715, n27716,
    n27717, n27718, n27719, n27720, n27721, n27722, n27723, n27724, n27725,
    n27726, n27727, n27728, n27729, n27730, n27731, n27732, n27733, n27734,
    n27735, n27736, n27737, n27738, n27739, n27740, n27741, n27742, n27743,
    n27744, n27745, n27746, n27747, n27748, n27749, n27750, n27751, n27752,
    n27753, n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27762,
    n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27772,
    n27773, n27774, n27775, n27776, n27777, n27778, n27779, n27780, n27782,
    n27783, n27785, n27786, n27788, n27789, n27791, n27792, n27794, n27795,
    n27797, n27798, n27800, n27801, n27802, n27803, n27804, n27805, n27806,
    n27807, n27808, n27809, n27810, n27811, n27812, n27813, n27814, n27815,
    n27816, n27817, n27818, n27819, n27820, n27821, n27822, n27823, n27824,
    n27825, n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
    n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
    n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
    n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859, n27860,
    n27861, n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
    n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27881, n27882, n27883, n27884, n27885, n27886, n27887,
    n27888, n27889, n27890, n27891, n27892, n27893, n27894, n27895, n27896,
    n27897, n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
    n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
    n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
    n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931, n27932,
    n27933, n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
    n27942, n27943, n27944, n27945, n27946, n27947, n27948, n27949, n27950,
    n27951, n27952, n27953, n27954, n27955, n27956, n27957, n27958, n27959,
    n27960, n27961, n27962, n27963, n27964, n27965, n27966, n27967, n27968,
    n27969, n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
    n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
    n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
    n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003, n28004,
    n28005, n28006, n28007, n28008, n28009, n28010, n28011, n28012, n28013,
    n28014, n28015, n28016, n28017, n28018, n28019, n28020, n28021, n28022,
    n28023, n28024, n28025, n28026, n28027, n28028, n28029, n28030, n28031,
    n28032, n28033, n28034, n28035, n28036, n28037, n28038, n28039, n28040,
    n28041, n28042, n28043, n28044, n28045, n28046, n28047, n28049, n28050,
    n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
    n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067, n28068,
    n28069, n28070, n28071, n28072, n28073, n28074, n28075, n28076, n28077,
    n28078, n28079, n28080, n28081, n28082, n28083, n28084, n28085, n28086,
    n28087, n28088, n28089, n28090, n28091, n28092, n28093, n28094, n28095,
    n28096, n28097, n28098, n28099, n28100, n28101, n28102, n28103, n28104,
    n28105, n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
    n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
    n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
    n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139, n28140,
    n28141, n28142, n28143, n28144, n28145, n28146, n28147, n28148, n28149,
    n28150, n28151, n28152, n28153, n28154, n28155, n28156, n28157, n28158,
    n28159, n28160, n28161, n28162, n28163, n28164, n28165, n28166, n28167,
    n28168, n28169, n28170, n28171, n28172, n28173, n28174, n28175, n28176,
    n28177, n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
    n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
    n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
    n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211, n28212,
    n28213, n28214, n28215, n28216, n28217, n28218, n28219, n28220, n28221,
    n28222, n28223, n28224, n28225, n28226, n28227, n28228, n28229, n28230,
    n28231, n28232, n28233, n28234, n28235, n28236, n28237, n28238, n28239,
    n28240, n28241, n28242, n28243, n28244, n28245, n28246, n28247, n28248,
    n28249, n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
    n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
    n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
    n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283, n28284,
    n28285, n28286, n28287, n28288, n28289, n28290, n28291, n28292, n28294,
    n28295, n28296, n28297, n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309, n28310, n28311, n28312,
    n28313, n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
    n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347, n28348,
    n28349, n28350, n28351, n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28361, n28362, n28363, n28364, n28365, n28366,
    n28367, n28368, n28369, n28370, n28371, n28372, n28373, n28374, n28375,
    n28376, n28377, n28378, n28379, n28380, n28381, n28382, n28383, n28384,
    n28385, n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
    n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
    n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
    n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419, n28420,
    n28421, n28422, n28423, n28424, n28425, n28426, n28427, n28428, n28429,
    n28430, n28431, n28432, n28433, n28434, n28435, n28436, n28437, n28438,
    n28439, n28440, n28441, n28442, n28443, n28444, n28445, n28446, n28447,
    n28448, n28449, n28450, n28451, n28452, n28453, n28454, n28455, n28456,
    n28457, n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
    n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
    n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
    n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491, n28492,
    n28493, n28494, n28495, n28496, n28497, n28498, n28499, n28500, n28501,
    n28502, n28503, n28504, n28505, n28506, n28507, n28508, n28509, n28510,
    n28511, n28512, n28513, n28514, n28515, n28516, n28517, n28518, n28519,
    n28520, n28521, n28522, n28523, n28524, n28525, n28526, n28527, n28528,
    n28529, n28530, n28531, n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
    n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562, n28563, n28564, n28565,
    n28566, n28567, n28568, n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580, n28581, n28582, n28583,
    n28584, n28585, n28586, n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
    n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
    n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634, n28635, n28636, n28637,
    n28638, n28639, n28640, n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652, n28653, n28654, n28655,
    n28656, n28657, n28658, n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
    n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
    n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706, n28707, n28708, n28709,
    n28710, n28711, n28712, n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724, n28725, n28726, n28727,
    n28728, n28729, n28730, n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
    n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
    n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778, n28779, n28780, n28781,
    n28782, n28783, n28785, n28786, n28787, n28788, n28789, n28790, n28791,
    n28792, n28793, n28794, n28795, n28796, n28797, n28798, n28799, n28800,
    n28801, n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
    n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
    n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
    n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835, n28836,
    n28837, n28838, n28839, n28840, n28841, n28842, n28843, n28844, n28845,
    n28846, n28847, n28848, n28849, n28850, n28851, n28852, n28853, n28854,
    n28855, n28856, n28857, n28858, n28859, n28860, n28861, n28862, n28863,
    n28864, n28865, n28866, n28867, n28868, n28869, n28870, n28871, n28872,
    n28873, n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
    n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
    n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
    n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907, n28908,
    n28909, n28910, n28911, n28912, n28913, n28914, n28915, n28916, n28917,
    n28918, n28919, n28920, n28921, n28922, n28923, n28924, n28925, n28926,
    n28927, n28928, n28929, n28930, n28931, n28932, n28933, n28934, n28935,
    n28936, n28937, n28938, n28939, n28940, n28941, n28942, n28943, n28944,
    n28945, n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
    n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
    n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
    n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979, n28980,
    n28981, n28982, n28983, n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995, n28996, n28997, n28998,
    n28999, n29000, n29001, n29002, n29003, n29004, n29005, n29006, n29007,
    n29008, n29009, n29010, n29011, n29012, n29013, n29014, n29015, n29016,
    n29017, n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
    n29026, n29027, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
    n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043, n29044,
    n29045, n29046, n29047, n29048, n29049, n29050, n29051, n29052, n29053,
    n29054, n29055, n29056, n29057, n29058, n29059, n29060, n29061, n29062,
    n29063, n29064, n29065, n29066, n29067, n29068, n29069, n29070, n29071,
    n29072, n29073, n29074, n29075, n29076, n29077, n29078, n29079, n29080,
    n29081, n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
    n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
    n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
    n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115, n29116,
    n29117, n29118, n29119, n29120, n29121, n29122, n29123, n29124, n29125,
    n29126, n29127, n29128, n29129, n29130, n29131, n29132, n29133, n29134,
    n29135, n29136, n29137, n29138, n29139, n29140, n29141, n29142, n29143,
    n29144, n29145, n29146, n29147, n29148, n29149, n29150, n29151, n29152,
    n29153, n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
    n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
    n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
    n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187, n29188,
    n29189, n29190, n29191, n29192, n29193, n29194, n29195, n29196, n29197,
    n29198, n29199, n29200, n29201, n29202, n29203, n29204, n29205, n29206,
    n29207, n29208, n29209, n29210, n29211, n29212, n29213, n29214, n29215,
    n29216, n29217, n29218, n29219, n29220, n29221, n29222, n29223, n29224,
    n29225, n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
    n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
    n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
    n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259, n29260,
    n29261, n29262, n29263, n29264, n29265, n29266, n29267, n29268, n29269,
    n29270, n29271, n29272, n29273, n29274, n29276, n29277, n29278, n29279,
    n29280, n29281, n29282, n29283, n29284, n29285, n29286, n29287, n29288,
    n29289, n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
    n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
    n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
    n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323, n29324,
    n29325, n29326, n29327, n29328, n29329, n29330, n29331, n29332, n29333,
    n29334, n29335, n29336, n29337, n29338, n29339, n29340, n29341, n29342,
    n29343, n29344, n29345, n29346, n29347, n29348, n29349, n29350, n29351,
    n29352, n29353, n29354, n29355, n29356, n29357, n29358, n29359, n29360,
    n29361, n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
    n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
    n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
    n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395, n29396,
    n29397, n29398, n29399, n29400, n29401, n29402, n29403, n29404, n29405,
    n29406, n29407, n29408, n29409, n29410, n29411, n29412, n29413, n29414,
    n29415, n29416, n29417, n29418, n29419, n29420, n29421, n29422, n29423,
    n29424, n29425, n29426, n29427, n29428, n29429, n29430, n29431, n29432,
    n29433, n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
    n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
    n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
    n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467, n29468,
    n29469, n29470, n29471, n29472, n29473, n29474, n29475, n29476, n29477,
    n29478, n29479, n29480, n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492, n29493, n29494, n29495,
    n29496, n29497, n29498, n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
    n29514, n29515, n29516, n29518, n29519, n29520, n29521, n29522, n29523,
    n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531, n29532,
    n29533, n29534, n29535, n29536, n29537, n29538, n29539, n29540, n29541,
    n29542, n29543, n29544, n29545, n29546, n29547, n29548, n29549, n29550,
    n29551, n29552, n29553, n29554, n29555, n29556, n29557, n29558, n29559,
    n29560, n29561, n29562, n29563, n29564, n29565, n29566, n29567, n29568,
    n29569, n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
    n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
    n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
    n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603, n29604,
    n29605, n29606, n29607, n29608, n29609, n29610, n29611, n29612, n29613,
    n29614, n29615, n29616, n29617, n29618, n29619, n29620, n29621, n29622,
    n29623, n29624, n29625, n29626, n29627, n29628, n29629, n29630, n29631,
    n29632, n29633, n29634, n29635, n29636, n29637, n29638, n29639, n29640,
    n29641, n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
    n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
    n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
    n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675, n29676,
    n29677, n29678, n29679, n29680, n29681, n29682, n29683, n29684, n29685,
    n29686, n29687, n29688, n29689, n29690, n29691, n29692, n29693, n29694,
    n29695, n29696, n29697, n29698, n29699, n29700, n29701, n29702, n29703,
    n29704, n29705, n29706, n29707, n29708, n29709, n29710, n29711, n29712,
    n29713, n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
    n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
    n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
    n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747, n29748,
    n29749, n29750, n29751, n29752, n29753, n29754, n29755, n29756, n29757,
    n29758, n29759, n29760, n29761, n29762, n29763, n29764, n29765, n29766,
    n29768, n29769, n29770, n29771, n29772, n29773, n29774, n29775, n29776,
    n29777, n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
    n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
    n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
    n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811, n29812,
    n29813, n29814, n29815, n29816, n29817, n29818, n29819, n29820, n29821,
    n29822, n29823, n29824, n29825, n29826, n29827, n29828, n29829, n29830,
    n29831, n29832, n29833, n29834, n29835, n29836, n29837, n29838, n29839,
    n29840, n29841, n29842, n29843, n29844, n29845, n29846, n29847, n29848,
    n29849, n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
    n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
    n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
    n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883, n29884,
    n29885, n29886, n29887, n29888, n29889, n29890, n29891, n29892, n29893,
    n29894, n29895, n29896, n29897, n29898, n29899, n29900, n29901, n29902,
    n29903, n29904, n29905, n29906, n29907, n29908, n29909, n29910, n29911,
    n29912, n29913, n29914, n29915, n29916, n29917, n29918, n29919, n29920,
    n29921, n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
    n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
    n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
    n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955, n29956,
    n29957, n29958, n29959, n29960, n29961, n29962, n29963, n29964, n29965,
    n29966, n29967, n29968, n29969, n29970, n29971, n29972, n29973, n29974,
    n29975, n29976, n29977, n29978, n29979, n29980, n29981, n29982, n29983,
    n29984, n29985, n29986, n29987, n29988, n29989, n29990, n29991, n29992,
    n29993, n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
    n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
    n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30019, n30020,
    n30021, n30022, n30023, n30024, n30025, n30026, n30027, n30028, n30029,
    n30030, n30031, n30032, n30033, n30034, n30035, n30036, n30037, n30038,
    n30039, n30040, n30041, n30042, n30043, n30044, n30045, n30046, n30047,
    n30048, n30049, n30050, n30051, n30052, n30053, n30054, n30055, n30056,
    n30057, n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
    n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
    n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
    n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091, n30092,
    n30093, n30094, n30095, n30096, n30097, n30098, n30099, n30100, n30101,
    n30102, n30103, n30104, n30105, n30106, n30107, n30108, n30109, n30110,
    n30111, n30112, n30113, n30114, n30115, n30116, n30117, n30118, n30119,
    n30120, n30121, n30122, n30123, n30124, n30125, n30126, n30127, n30128,
    n30129, n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
    n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
    n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
    n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163, n30164,
    n30165, n30166, n30167, n30168, n30169, n30170, n30171, n30172, n30173,
    n30174, n30175, n30176, n30177, n30178, n30179, n30180, n30181, n30182,
    n30183, n30184, n30185, n30186, n30187, n30188, n30189, n30190, n30191,
    n30192, n30193, n30194, n30195, n30196, n30197, n30198, n30199, n30200,
    n30201, n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
    n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
    n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
    n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235, n30236,
    n30237, n30238, n30239, n30240, n30241, n30242, n30243, n30244, n30245,
    n30246, n30247, n30248, n30249, n30250, n30251, n30252, n30253, n30254,
    n30255, n30256, n30257, n30258, n30259, n30260, n30262, n30263, n30264,
    n30265, n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30274,
    n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30283, n30284,
    n30285, n30286, n30287, n30288, n30289, n30290, n30291, n30292, n30293,
    n30295, n30296, n30297, n30298, n30299, n30300, n30301, n30302, n30304,
    n30305, n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
    n30314, n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
    n30324, n30325, n30326, n30328, n30329, n30330, n30331, n30332, n30333,
    n30334, n30335, n30336, n30337, n30338, n30340, n30341, n30342, n30343,
    n30344, n30345, n30346, n30347, n30349, n30350, n30351, n30352, n30353,
    n30354, n30355, n30356, n30358, n30359, n30360, n30361, n30362, n30363,
    n30364, n30365, n30367, n30368, n30369, n30370, n30371, n30372, n30373,
    n30374, n30375, n30376, n30377, n30378, n30379, n30380, n30381, n30382,
    n30384, n30385, n30386, n30387, n30388, n30389, n30390, n30391, n30392,
    n30393, n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
    n30402, n30403, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
    n30412, n30413, n30414, n30415, n30416, n30418, n30419, n30420, n30421,
    n30422, n30423, n30424, n30425, n30426, n30428, n30429, n30430, n30431,
    n30432, n30433, n30434, n30435, n30436, n30438, n30439, n30440, n30441,
    n30442, n30443, n30444, n30445, n30446, n30448, n30449, n30451, n30452,
    n30454, n30455, n30457, n30458, n30460, n30461, n30463, n30464, n30466,
    n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
    n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483, n30484,
    n30485, n30486, n30487, n30488, n30489, n30490, n30491, n30492, n30493,
    n30494, n30495, n30496, n30497, n30499, n30500, n30501, n30502, n30503,
    n30504, n30505, n30506, n30507, n30508, n30509, n30510, n30511, n30512,
    n30513, n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
    n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
    n30531, n30532, n30534, n30535, n30536, n30537, n30538, n30539, n30540,
    n30541, n30542, n30543, n30544, n30545, n30546, n30547, n30548, n30549,
    n30550, n30551, n30552, n30553, n30554, n30555, n30556, n30557, n30559,
    n30560, n30561, n30562, n30563, n30564, n30565, n30566, n30567, n30568,
    n30569, n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
    n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
    n30587, n30588, n30590, n30591, n30592, n30593, n30594, n30595, n30596,
    n30597, n30598, n30600, n30601, n30603, n30604, n30606, n30607, n30608,
    n30609, n30613, n30614, n30615, n30616, n30617, n30618, n30619, n30620,
    n30621, n30622, n30623, n30624, n30625, n30626, n30627, n30628, n30629,
    n30630, n30632, n30633, n30634, n30635, n30636, n30637, n30638, n30639,
    n30640, n30641, n30642, n30643, n30644, n30645, n30646, n30647, n30649,
    n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30659,
    n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667, n30669,
    n30670, n30672, n30673, n30675, n30676, n30678, n30679, n30681, n30682,
    n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699, n30700,
    n30701, n30702, n30703, n30704, n30705, n30707, n30708, n30709, n30710,
    n30711, n30713, n30714, n30715, n30716, n30717, n30718, n30719, n30720,
    n30721, n30722, n30723, n30724, n30726, n30727, n30728, n30729, n30730,
    n30731, n30732, n30733, n30734, n30736, n30737, n30739, n30740, n30742,
    n30743, n30744, n30745, n30746, n30747, n30748, n30749, n30750, n30751,
    n30752, n30753, n30754, n30755, n30756, n30757, n30758, n30759, n30760,
    n30761, n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
    n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
    n30779, n30781, n30782, n30783, n30784, n30785, n30786, n30787, n30788,
    n30789, n30791, n30792, n30793, n30794, n30796, n30797, n30798, n30800,
    n30801, n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30810,
    n30811, n30812, n30813, n30814, n30815, n30817, n30818, n30819, n30820,
    n30821, n30822, n30824, n30825, n30826, n30827, n30828, n30829, n30831,
    n30832, n30833, n30834, n30835, n30836, n30838, n30839, n30840, n30841,
    n30842, n30843, n30845, n30846, n30847, n30848, n30849, n30850, n30852,
    n30853, n30854, n30855, n30856, n30857, n30859, n30860, n30861, n30862,
    n30863, n30864, n30866, n30867, n30868, n30869, n30870, n30871, n30873,
    n30874, n30875, n30876, n30877, n30878, n30880, n30881, n30882, n30883,
    n30884, n30885, n30887, n30888, n30889, n30890, n30891, n30892, n30894,
    n30895, n30896, n30897, n30898, n30899, n30901, n30902, n30904, n30905,
    n30907, n30908, n30910, n30911, n30913, n30914, n30916, n30917, n30919,
    n30920, n30922, n30923, n30924, n30925, n30926, n30927, n30929, n30930,
    n30932, n30933, n30935, n30936, n30938, n30939, n30941, n30942, n30944,
    n30945, n30947, n30948, n30950, n30951, n30953, n30954, n30955, n30956,
    n30957, n30958, n30959, n30960, n30962, n30963, n30964, n30965, n30966,
    n30967, n30968, n30970, n30971, n30972, n30973, n30974, n30975, n30976,
    n30977, n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
    n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994,
    n30995, n30997, n30998, n30999, n31000, n31001, n31002, n31003, n31004,
    n31005, n31007, n31008, n31010, n31011, n31013, n31014, n31016, n31017,
    n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
    n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
    n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043, n31044,
    n31045, n31046, n31047, n31048, n31049, n31050, n31051, n31052, n31053,
    n31054, n31055, n31056, n31057, n31058, n31059, n31060, n31061, n31062,
    n31063, n31064, n31065, n31066, n31067, n31068, n31069, n31070, n31071,
    n31072, n31073, n31074, n31075, n31076, n31077, n31078, n31079, n31080,
    n31081, n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
    n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
    n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
    n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115, n31116,
    n31117, n31118, n31119, n31120, n31121, n31122, n31123, n31124, n31125,
    n31126, n31127, n31128, n31129, n31130, n31131, n31132, n31133, n31134,
    n31135, n31136, n31137, n31138, n31139, n31140, n31141, n31142, n31143,
    n31144, n31145, n31146, n31147, n31148, n31149, n31150, n31151, n31152,
    n31153, n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
    n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170,
    n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
    n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187, n31188,
    n31189, n31190, n31191, n31192, n31193, n31194, n31195, n31196, n31197,
    n31198, n31199, n31200, n31201, n31202, n31203, n31204, n31205, n31206,
    n31207, n31208, n31209, n31210, n31211, n31212, n31213, n31214, n31215,
    n31216, n31217, n31218, n31219, n31220, n31221, n31222, n31223, n31224,
    n31225, n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
    n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242,
    n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
    n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259, n31260,
    n31261, n31262, n31263, n31264, n31265, n31266, n31267, n31268, n31269,
    n31270, n31271, n31272, n31273, n31274, n31275, n31276, n31277, n31278,
    n31279, n31280, n31281, n31282, n31283, n31284, n31285, n31286, n31287,
    n31288, n31289, n31290, n31291, n31292, n31293, n31294, n31295, n31296,
    n31297, n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
    n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
    n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
    n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331, n31332,
    n31333, n31334, n31335, n31336, n31337, n31338, n31339, n31340, n31341,
    n31342, n31343, n31344, n31345, n31346, n31347, n31348, n31349, n31350,
    n31351, n31352, n31353, n31355, n31356, n31357, n31358, n31359, n31360,
    n31361, n31362, n31363, n31364, n31365, n31366, n31368, n31369, n31370,
    n31371, n31372, n31373, n31374, n31375, n31376, n31378, n31379, n31380,
    n31381, n31382, n31383, n31384, n31385, n31386, n31387, n31388, n31389,
    n31390, n31391, n31392, n31393, n31394, n31396, n31397, n31398, n31399,
    n31400, n31401, n31402, n31403, n31404, n31405, n31406, n31407, n31408,
    n31409, n31410, n31411, n31412, n31414, n31415, n31417, n31418, n31420,
    n31421, n31422, n31424, n31425, n31426, n31427, n31428, n31430, n31431,
    n31433, n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
    n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450,
    n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
    n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467, n31468,
    n31469, n31470, n31471, n31472, n31473, n31474, n31475, n31476, n31477,
    n31478, n31479, n31480, n31481, n31482, n31483, n31484, n31485, n31486,
    n31487, n31488, n31489, n31490, n31491, n31492, n31493, n31494, n31495,
    n31496, n31497, n31498, n31499, n31500, n31501, n31502, n31503, n31504,
    n31505, n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
    n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
    n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
    n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539, n31540,
    n31541, n31542, n31543, n31544, n31545, n31546, n31547, n31548, n31549,
    n31550, n31551, n31552, n31553, n31554, n31555, n31556, n31557, n31558,
    n31559, n31560, n31561, n31562, n31563, n31564, n31565, n31566, n31567,
    n31568, n31569, n31570, n31571, n31572, n31573, n31574, n31575, n31576,
    n31577, n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
    n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594,
    n31595, n31597, n31598, n31599, n31600, n31601, n31603, n31604, n31605,
    n31606, n31607, n31609, n31610, n31611, n31612, n31613, n31615, n31616,
    n31617, n31619, n31620, n31622, n31623, n31624, n31625, n31626, n31628,
    n31629, n31631, n31632, n31634, n31635, n31637, n31638, n31639, n31640,
    n31641, n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
    n31650, n31651, n31652, n31653, n31654, n31656, n31657, n31658, n31659,
    n31660, n31661, n31662, n31663, n31664, n31666, n31667, n31668, n31669,
    n31670, n31671, n31672, n31673, n31674, n31676, n31677, n31678, n31679,
    n31680, n31681, n31682, n31683, n31684, n31686, n31687, n31689, n31690,
    n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699, n31700,
    n31701, n31702, n31703, n31704, n31705, n31706, n31707, n31708, n31709,
    n31710, n31711, n31713, n31714, n31715, n31716, n31717, n31718, n31719,
    n31720, n31721, n31722, n31723, n31724, n31726, n31727, n31728, n31729,
    n31730, n31731, n31732, n31733, n31734, n31736, n31737, n31738, n31739,
    n31740, n31741, n31742, n31743, n31744, n31746, n31747, n31749, n31750,
    n31752, n31753, n31755, n31756, n31758, n31759, n31761, n31762, n31763,
    n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771, n31772,
    n31773, n31774, n31775, n31776, n31777, n31778, n31779, n31780, n31781,
    n31782, n31783, n31784, n31785, n31786, n31787, n31788, n31789, n31790,
    n31791, n31792, n31793, n31794, n31795, n31796, n31797, n31798, n31799,
    n31800, n31801, n31802, n31803, n31804, n31805, n31806, n31807, n31808,
    n31809, n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
    n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
    n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
    n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843, n31844,
    n31845, n31846, n31847, n31848, n31849, n31850, n31851, n31852, n31853,
    n31854, n31855, n31856, n31857, n31858, n31859, n31860, n31861, n31862,
    n31863, n31864, n31865, n31866, n31867, n31868, n31869, n31870, n31872,
    n31873, n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
    n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890,
    n31891, n31892, n31893, n31894, n31896, n31897, n31898, n31899, n31900,
    n31901, n31902, n31903, n31904, n31905, n31906, n31907, n31908, n31909,
    n31910, n31911, n31912, n31913, n31914, n31915, n31917, n31918, n31919,
    n31920, n31921, n31923, n31924, n31926, n31927, n31928, n31929, n31930,
    n31931, n31932, n31933, n31934, n31936, n31937, n31938, n31939, n31940,
    n31941, n31942, n31943, n31944, n31946, n31947, n31948, n31949, n31950,
    n31951, n31952, n31953, n31955, n31956, n31957, n31959, n31960, n31961,
    n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
    n31971, n31972, n31973, n31974, n31976, n31977, n31978, n31979, n31980,
    n31982, n31983, n31985, n31986, n31987, n31988, n31989, n31990, n31991,
    n31993, n31994, n31995, n31996, n31997, n31999, n32000, n32001, n32002,
    n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
    n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019, n32020,
    n32022, n32023, n32024, n32025, n32026, n32028, n32029, n32031, n32032,
    n32033, n32034, n32035, n32036, n32037, n32038, n32039, n32041, n32042,
    n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32051, n32052,
    n32053, n32054, n32055, n32057, n32058, n32059, n32060, n32061, n32063,
    n32064, n32066, n32067, n32069, n32070, n32071, n32072, n32073, n32074,
    n32075, n32076, n32077, n32078, n32079, n32080, n32082, n32083, n32084,
    n32085, n32086, n32087, n32088, n32089, n32090, n32091, n32092, n32093,
    n32094, n32095, n32096, n32097, n32099, n32100, n32101, n32102, n32103,
    n32104, n32105, n32106, n32107, n32108, n32109, n32110, n32111, n32112,
    n32113, n32114, n32116, n32117, n32118, n32119, n32120, n32122, n32123,
    n32124, n32125, n32126, n32128, n32129, n32130, n32131, n32132, n32134,
    n32135, n32137, n32138, n32140, n32141, n32143, n32144, n32145, n32146,
    n32147, n32148, n32149, n32150, n32151, n32153, n32154, n32155, n32156,
    n32157, n32158, n32159, n32160, n32161, n32163, n32164, n32165, n32166,
    n32167, n32168, n32169, n32170, n32171, n32173, n32174, n32175, n32176,
    n32177, n32178, n32179, n32180, n32181, n32183, n32184, n32185, n32186,
    n32187, n32189, n32190, n32191, n32192, n32193, n32195, n32196, n32197,
    n32198, n32199, n32201, n32202, n32203, n32204, n32205, n32207, n32208,
    n32210, n32211, n32213, n32214, n32216, n32217, n32219, n32220, n32221,
    n32222, n32223, n32224, n32225, n32226, n32227, n32229, n32230, n32231,
    n32232, n32233, n32234, n32235, n32236, n32237, n32239, n32240, n32241,
    n32242, n32243, n32245, n32246, n32248, n32249, n32250, n32251, n32252,
    n32254, n32255, n32257, n32258, n32259, n32260, n32261, n32263, n32264,
    n32265, n32266, n32267, n32269, n32270, n32272, n32273, n32275, n32276,
    n32277, n32278, n32279, n32280, n32281, n32282, n32283, n32284, n32285,
    n32287, n32288, n32289, n32290, n32291, n32292, n32293, n32294, n32295,
    n32296, n32297, n32298, n32299, n32300, n32301, n32302, n32303, n32305,
    n32306, n32307, n32308, n32309, n32311, n32312, n32314, n32315, n32316,
    n32317, n32318, n32320, n32321, n32322, n32323, n32324, n32326, n32327,
    n32329, n32330, n32332, n32333, n32334, n32335, n32336, n32338, n32339,
    n32341, n32342, n32343, n32344, n32345, n32347, n32348, n32349, n32350,
    n32351, n32353, n32354, n32355, n32356, n32357, n32359, n32360, n32362,
    n32363, n32365, n32366, n32368, n32369, n32370, n32371, n32372, n32373,
    n32374, n32375, n32376, n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32388, n32389, n32390, n32391, n32392, n32394,
    n32395, n32397, n32398, n32399, n32400, n32401, n32403, n32404, n32406,
    n32407, n32408, n32409, n32410, n32412, n32413, n32415, n32416, n32417,
    n32418, n32419, n32421, n32422, n32424, n32425, n32426, n32427, n32428,
    n32429, n32430, n32431, n32432, n32433, n32434, n32436, n32437, n32438,
    n32439, n32440, n32442, n32443, n32444, n32445, n32446, n32448, n32449,
    n32451, n32452, n32454, n32455, n32456, n32457, n32458, n32460, n32461,
    n32462, n32463, n32464, n32466, n32467, n32469, n32470, n32472, n32473,
    n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32482, n32483,
    n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32492, n32493,
    n32494, n32495, n32496, n32497, n32498, n32499, n32501, n32502, n32503,
    n32504, n32505, n32507, n32508, n32510, n32511, n32512, n32513, n32514,
    n32516, n32517, n32518, n32519, n32520, n32522, n32523, n32525, n32526,
    n32528, n32529, n32530, n32531, n32532, n32534, n32535, n32537, n32538,
    n32539, n32540, n32541, n32543, n32544, n32546, n32547, n32548, n32549,
    n32550, n32552, n32553, n32555, n32556, n32557, n32558, n32559, n32560,
    n32561, n32562, n32563, n32565, n32566, n32567, n32568, n32569, n32570,
    n32571, n32572, n32573, n32575, n32576, n32577, n32578, n32579, n32580,
    n32581, n32582, n32583, n32584, n32585, n32586, n32587, n32588, n32589,
    n32590, n32591, n32593, n32594, n32595, n32596, n32597, n32599, n32600,
    n32601, n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
    n32610, n32611, n32612, n32613, n32614, n32616, n32617, n32618, n32619,
    n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627, n32628,
    n32629, n32630, n32631, n32632, n32633, n32635, n32636, n32637, n32639,
    n32640, n32641, n32642, n32643, n32644, n32645, n32646, n32647, n32649,
    n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32659,
    n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667, n32668,
    n32669, n32670, n32671, n32673, n32674, n32675, n32676, n32677, n32679,
    n32680, n32681, n32682, n32683, n32685, n32686, n32688, n32689, n32691,
    n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699, n32700,
    n32701, n32702, n32703, n32704, n32705, n32706, n32707, n32708, n32709,
    n32710, n32711, n32713, n32714, n32715, n32716, n32718, n32719, n32720,
    n32721, n32723, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
    n32732, n32733, n32735, n32736, n32737, n32738, n32739, n32740, n32741,
    n32742, n32743, n32745, n32746, n32747, n32748, n32749, n32751, n32752,
    n32753, n32754, n32755, n32757, n32758, n32760, n32761, n32763, n32764,
    n32765, n32766, n32767, n32768, n32769, n32770, n32771, n32772, n32773,
    n32774, n32775, n32776, n32777, n32778, n32780, n32781, n32782, n32783,
    n32784, n32785, n32786, n32787, n32788, n32789, n32790, n32791, n32792,
    n32793, n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
    n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
    n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
    n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827, n32828,
    n32829, n32830, n32831, n32832, n32833, n32834, n32835, n32836, n32837,
    n32838, n32839, n32840, n32841, n32842, n32843, n32844, n32845, n32846,
    n32847, n32848, n32849, n32850, n32851, n32852, n32853, n32854, n32855,
    n32856, n32857, n32858, n32859, n32860, n32861, n32862, n32864, n32865,
    n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
    n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883,
    n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891, n32893,
    n32894, n32895, n32896, n32897, n32898, n32899, n32900, n32901, n32902,
    n32903, n32904, n32905, n32906, n32907, n32908, n32909, n32910, n32911,
    n32912, n32913, n32914, n32915, n32916, n32917, n32918, n32919, n32920,
    n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
    n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
    n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947, n32948,
    n32949, n32951, n32952, n32953, n32954, n32955, n32956, n32957, n32958,
    n32959, n32960, n32961, n32962, n32963, n32964, n32965, n32966, n32967,
    n32968, n32969, n32970, n32971, n32972, n32973, n32974, n32975, n32976,
    n32977, n32978, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
    n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
    n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003, n33004,
    n33005, n33006, n33007, n33009, n33010, n33011, n33012, n33013, n33014,
    n33015, n33016, n33017, n33018, n33019, n33020, n33021, n33022, n33023,
    n33024, n33025, n33026, n33027, n33028, n33029, n33030, n33031, n33032,
    n33033, n33034, n33035, n33036, n33038, n33039, n33040, n33041, n33042,
    n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
    n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059, n33060,
    n33061, n33062, n33063, n33064, n33065, n33067, n33068, n33069, n33070,
    n33071, n33072, n33073, n33074, n33075, n33076, n33077, n33078, n33079,
    n33080, n33081, n33082, n33083, n33084, n33085, n33086, n33087, n33088,
    n33089, n33090, n33091, n33092, n33093, n33094, n33096, n33097, n33098,
    n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
    n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115, n33116,
    n33117, n33118, n33119, n33120, n33121, n33122, n33123, n33125, n33126,
    n33127, n33128, n33129, n33130, n33131, n33132, n33133, n33134, n33135,
    n33136, n33137, n33138, n33139, n33140, n33141, n33142, n33143, n33144,
    n33145, n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33154,
    n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
    n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171, n33172,
    n33173, n33174, n33175, n33176, n33177, n33178, n33179, n33180, n33181,
    n33183, n33184, n33185, n33186, n33187, n33188, n33189, n33190, n33191,
    n33192, n33193, n33194, n33195, n33196, n33197, n33198, n33199, n33200,
    n33201, n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
    n33210, n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
    n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227, n33228,
    n33229, n33230, n33231, n33232, n33233, n33234, n33235, n33236, n33237,
    n33238, n33239, n33241, n33242, n33243, n33244, n33245, n33246, n33247,
    n33248, n33249, n33250, n33251, n33252, n33253, n33254, n33255, n33256,
    n33257, n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
    n33266, n33267, n33268, n33270, n33271, n33272, n33273, n33274, n33275,
    n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283, n33284,
    n33285, n33286, n33287, n33288, n33289, n33290, n33291, n33292, n33293,
    n33294, n33295, n33296, n33297, n33299, n33300, n33301, n33302, n33303,
    n33304, n33305, n33306, n33307, n33308, n33309, n33311, n33312, n33313,
    n33314, n33315, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
    n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331, n33332,
    n33333, n33334, n33335, n33336, n33337, n33338, n33339, n33341, n33342,
    n33343, n33344, n33345, n33346, n33347, n33348, n33349, n33350, n33351,
    n33352, n33353, n33354, n33355, n33356, n33358, n33359, n33360, n33361,
    n33362, n33363, n33364, n33365, n33367, n33368, n33369, n33370, n33371,
    n33372, n33373, n33374, n33376, n33377, n33378, n33379, n33380, n33381,
    n33382, n33383, n33385, n33386, n33387, n33388, n33389, n33390, n33391,
    n33392, n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
    n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
    n33412, n33413, n33415, n33416, n33417, n33418, n33419, n33420, n33421,
    n33422, n33423, n33424, n33425, n33427, n33428, n33429, n33430, n33431,
    n33432, n33433, n33434, n33435, n33436, n33437, n33439, n33440, n33441,
    n33442, n33443, n33444, n33445, n33446, n33448, n33449, n33450, n33451,
    n33452, n33453, n33454, n33455, n33457, n33458, n33459, n33460, n33461,
    n33462, n33463, n33464, n33465, n33466, n33467, n33469, n33470, n33471,
    n33472, n33473, n33474, n33475, n33476, n33477, n33478, n33479, n33481,
    n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
    n33491, n33493, n33494, n33495, n33496, n33497, n33498, n33499, n33500,
    n33501, n33502, n33503, n33504, n33505, n33506, n33507, n33508, n33509,
    n33510, n33511, n33512, n33513, n33514, n33515, n33516, n33517, n33518,
    n33519, n33520, n33522, n33523, n33524, n33525, n33526, n33527, n33528,
    n33529, n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
    n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546,
    n33547, n33548, n33549, n33551, n33552, n33553, n33554, n33555, n33556,
    n33557, n33558, n33559, n33560, n33561, n33562, n33563, n33564, n33565,
    n33566, n33567, n33568, n33569, n33570, n33571, n33572, n33573, n33574,
    n33575, n33576, n33577, n33578, n33580, n33581, n33582, n33583, n33584,
    n33585, n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
    n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
    n33603, n33604, n33605, n33606, n33607, n33609, n33610, n33611, n33612,
    n33613, n33614, n33615, n33616, n33617, n33618, n33619, n33620, n33621,
    n33622, n33623, n33624, n33625, n33626, n33627, n33628, n33629, n33630,
    n33631, n33632, n33633, n33634, n33635, n33636, n33638, n33639, n33640,
    n33641, n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
    n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658,
    n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33667, n33668,
    n33669, n33670, n33671, n33672, n33673, n33674, n33675, n33676, n33677,
    n33678, n33679, n33680, n33681, n33682, n33683, n33684, n33685, n33686,
    n33687, n33688, n33689, n33690, n33691, n33692, n33693, n33694, n33696,
    n33697, n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
    n33706, n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
    n33716, n33717, n33718, n33720, n33721, n33722, n33723, n33724, n33725,
    n33726, n33727, n33728, n33729, n33730, n33731, n33732, n33733, n33734,
    n33735, n33736, n33737, n33738, n33739, n33740, n33741, n33742, n33743,
    n33744, n33745, n33746, n33747, n33749, n33750, n33751, n33752, n33753,
    n33755, n33756, n33758, n33759, n33760, n33761, n33762, n33763, n33764,
    n33765, n33766, n33768, n33769, n33770, n33771, n33772, n33773, n33774,
    n33775, n33776, n33778, n33779, n33780, n33781, n33782, n33783, n33784,
    n33785, n33786, n33787, n33788, n33790, n33791, n33792, n33793, n33794,
    n33796, n33797, n33799, n33800, n33801, n33802, n33803, n33805, n33806,
    n33808, n33809, n33810, n33811, n33813, n33814, n33815, n33816, n33817,
    n33818, n33819, n33820, n33822, n33823, n33824, n33825, n33826, n33827,
    n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835, n33836,
    n33837, n33838, n33839, n33840, n33841, n33842, n33843, n33844, n33845,
    n33846, n33847, n33848, n33849, n33850, n33851, n33852, n33853, n33854,
    n33855, n33856, n33857, n33858, n33859, n33860, n33861, n33862, n33863,
    n33864, n33865, n33866, n33867, n33868, n33869, n33870, n33871, n33872,
    n33873, n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
    n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890,
    n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
    n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907, n33908,
    n33909, n33910, n33911, n33912, n33913, n33914, n33915, n33916, n33917,
    n33918, n33919, n33920, n33921, n33922, n33923, n33924, n33925, n33926,
    n33927, n33928, n33929, n33930, n33931, n33932, n33933, n33934, n33935,
    n33936, n33937, n33938, n33939, n33940, n33941, n33942, n33943, n33944,
    n33945, n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
    n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962,
    n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
    n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979, n33980,
    n33981, n33982, n33983, n33984, n33985, n33986, n33987, n33988, n33989,
    n33990, n33991, n33992, n33993, n33994, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004, n34005, n34006, n34007,
    n34008, n34009, n34010, n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
    n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
    n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051, n34052,
    n34053, n34054, n34055, n34056, n34057, n34058, n34059, n34060, n34061,
    n34062, n34063, n34064, n34065, n34066, n34067, n34068, n34069, n34070,
    n34071, n34072, n34073, n34074, n34075, n34076, n34077, n34078, n34079,
    n34080, n34081, n34082, n34083, n34084, n34085, n34086, n34087, n34088,
    n34089, n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
    n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
    n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
    n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123, n34124,
    n34125, n34126, n34127, n34128, n34129, n34130, n34131, n34132, n34133,
    n34134, n34135, n34136, n34137, n34138, n34139, n34140, n34141, n34142,
    n34143, n34144, n34145, n34146, n34147, n34148, n34149, n34150, n34151,
    n34152, n34153, n34154, n34155, n34156, n34157, n34158, n34159, n34160,
    n34161, n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
    n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
    n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
    n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195, n34196,
    n34197, n34198, n34199, n34200, n34201, n34202, n34203, n34204, n34205,
    n34206, n34207, n34208, n34209, n34210, n34211, n34212, n34213, n34214,
    n34215, n34216, n34217, n34218, n34219, n34220, n34221, n34222, n34223,
    n34224, n34225, n34226, n34227, n34228, n34229, n34230, n34231, n34232,
    n34233, n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
    n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
    n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
    n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267, n34268,
    n34269, n34270, n34271, n34272, n34273, n34274, n34275, n34276, n34277,
    n34278, n34279, n34280, n34281, n34282, n34283, n34284, n34285, n34286,
    n34287, n34288, n34289, n34290, n34291, n34292, n34293, n34294, n34295,
    n34296, n34297, n34298, n34299, n34300, n34301, n34302, n34303, n34304,
    n34305, n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
    n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
    n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
    n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339, n34340,
    n34341, n34342, n34343, n34344, n34345, n34346, n34347, n34348, n34349,
    n34350, n34351, n34352, n34353, n34354, n34355, n34356, n34357, n34358,
    n34359, n34360, n34361, n34362, n34363, n34364, n34365, n34366, n34367,
    n34368, n34369, n34370, n34371, n34372, n34373, n34374, n34375, n34376,
    n34377, n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
    n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
    n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
    n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411, n34412,
    n34413, n34414, n34415, n34416, n34417, n34418, n34419, n34420, n34421,
    n34422, n34423, n34424, n34425, n34426, n34427, n34428, n34429, n34430,
    n34431, n34432, n34433, n34434, n34435, n34436, n34437, n34438, n34439,
    n34440, n34441, n34442, n34443, n34444, n34445, n34446, n34447, n34448,
    n34449, n34450, n34451, n34453, n34454, n34455, n34456, n34457, n34459,
    n34460, n34461, n34462, n34463, n34465, n34466, n34467, n34468, n34469,
    n34471, n34472, n34473, n34474, n34475, n34477, n34478, n34479, n34480,
    n34481, n34483, n34484, n34485, n34486, n34487, n34489, n34490, n34491,
    n34492, n34493, n34495, n34496, n34497, n34498, n34499, n34501, n34502,
    n34503, n34504, n34505, n34507, n34508, n34509, n34510, n34511, n34513,
    n34514, n34515, n34516, n34517, n34519, n34520, n34521, n34522, n34523,
    n34525, n34526, n34527, n34528, n34529, n34531, n34532, n34533, n34534,
    n34535, n34537, n34538, n34539, n34540, n34541, n34543, n34544, n34545,
    n34546, n34547, n34549, n34550, n34551, n34552, n34553, n34555, n34556,
    n34557, n34558, n34559, n34561, n34562, n34563, n34564, n34565, n34567,
    n34568, n34569, n34570, n34571, n34573, n34574, n34575, n34576, n34577,
    n34579, n34580, n34581, n34582, n34583, n34585, n34586, n34587, n34588,
    n34589, n34591, n34592, n34593, n34594, n34595, n34596, n34597, n34598,
    n34599, n34600, n34601, n34602, n34604, n34605, n34606, n34607, n34609,
    n34610, n34611, n34612, n34614, n34615, n34616, n34617, n34619, n34620,
    n34621, n34622, n34624, n34625, n34626, n34627, n34629, n34630, n34631,
    n34632, n34634, n34635, n34636, n34637, n34639, n34640, n34641, n34642,
    n34643, n34645, n34646, n34648, n34649, n34650, n34651, n34652, n34653,
    n34654, n34655, n34656, n34657, n34659, n34660, n34661, n34662, n34663,
    n34664, n34665, n34666, n34668, n34669, n34670, n34671, n34672, n34674,
    n34675, n34676, n34677, n34678, n34680, n34681, n34682, n34683, n34684,
    n34686, n34687, n34688, n34689, n34690, n34692, n34693, n34694, n34695,
    n34696, n34698, n34699, n34700, n34701, n34702, n34704, n34705, n34706,
    n34707, n34708, n34710, n34711, n34712, n34713, n34714, n34716, n34717,
    n34718, n34719, n34720, n34722, n34723, n34724, n34725, n34726, n34728,
    n34729, n34730, n34731, n34732, n34734, n34735, n34736, n34737, n34738,
    n34740, n34741, n34742, n34743, n34744, n34746, n34747, n34748, n34749,
    n34750, n34751, n34752, n34753, n34755, n34756, n34757, n34758, n34759,
    n34760, n34761, n34762, n34764, n34765, n34766, n34767, n34768, n34769,
    n34770, n34771, n34773, n34774, n34775, n34776, n34777, n34778, n34779,
    n34780, n34782, n34783, n34784, n34785, n34786, n34787, n34788, n34789,
    n34791, n34792, n34793, n34794, n34795, n34796, n34797, n34798, n34799,
    n34800, n34801, n34803, n34804, n34805, n34806, n34807, n34809, n34810,
    n34811, n34812, n34813, n34815, n34816, n34817, n34818, n34819, n34820,
    n34821, n34822, n34824, n34825, n34826, n34827, n34828, n34830, n34831,
    n34832, n34833, n34834, n34836, n34837, n34839, n34840, n34841, n34842,
    n34843, n34845, n34846, n34847, n34848, n34849, n34850, n34851, n34852,
    n34853, n34854, n34855, n34858, n34859, n34860, n34861, n34862, n34863,
    n34864, n34865, n34866, n34867, n34868, n34869, n34870, n34871, n34872,
    n34873, n34874, n34875, n34876, n34877, n34878, n34880, n34881, n34882,
    n34883, n34885, n34886, n34887, n34888, n34890, n34891, n34892, n34893,
    n34895, n34896, n34897, n34898, n34900, n34901, n34902, n34903, n34905,
    n34906, n34907, n34908, n34910, n34911, n34912, n34913, n34915, n34916,
    n34917, n34918, n34920, n34921, n34922, n34923, n34925, n34926, n34927,
    n34928, n34930, n34931, n34932, n34933, n34935, n34936, n34937, n34938,
    n34940, n34941, n34942, n34944, n34945, n34946, n34947, n34948, n34949,
    n34950, n34951, n34952, n34953, n34954, n34956, n34957, n34958, n34959,
    n34960, n34962, n34963, n34965, n34966, n34967, n34968, n34969, n34970,
    n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
    n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987, n34988,
    n34989, n34990, n34991, n34992, n34993, n34994, n34995, n34996, n34997,
    n34998, n34999, n35000, n35001, n35002, n35003, n35004, n35005, n35006,
    n35007, n35008, n35009, n35010, n35011, n35012, n35013, n35014, n35015,
    n35016, n35017, n35018, n35019, n35020, n35021, n35022, n35023, n35024,
    n35025, n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
    n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042,
    n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
    n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059, n35060,
    n35061, n35062, n35063, n35064, n35065, n35066, n35067, n35068, n35069,
    n35070, n35071, n35072, n35073, n35074, n35075, n35076, n35077, n35078,
    n35079, n35080, n35081, n35082, n35083, n35084, n35085, n35086, n35087,
    n35088, n35089, n35090, n35091, n35092, n35093, n35094, n35095, n35096,
    n35097, n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
    n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114,
    n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
    n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131, n35132,
    n35133, n35134, n35135, n35136, n35137, n35138, n35139, n35140, n35141,
    n35142, n35143, n35144, n35145, n35146, n35147, n35148, n35149, n35150,
    n35151, n35152, n35153, n35154, n35155, n35156, n35157, n35158, n35159,
    n35160, n35161, n35162, n35163, n35164, n35165, n35166, n35167, n35168,
    n35169, n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
    n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186,
    n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
    n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203, n35204,
    n35205, n35206, n35207, n35208, n35209, n35210, n35211, n35212, n35213,
    n35214, n35215, n35216, n35217, n35218, n35219, n35220, n35221, n35222,
    n35223, n35224, n35225, n35226, n35227, n35228, n35229, n35230, n35231,
    n35232, n35233, n35234, n35235, n35236, n35237, n35238, n35239, n35240,
    n35241, n35242, n35243, n35244, n35245, n35247, n35248, n35249, n35250,
    n35251, n35252, n35253, n35254, n35256, n35257, n35258, n35259, n35261,
    n35262, n35263, n35264, n35266, n35267, n35269, n35270, n35272, n35273,
    n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
    n35285, n35286, n35287, n35288, n35289, n35290, n35291, n35292, n35293,
    n35295, n35296, n35297, n35298, n35299, n35300, n35302, n35303, n35304,
    n35305, n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
    n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322,
    n35323, n35324, n35327, n35328, n35329, n35330, n35331, n35332, n35333,
    n35334, n35336, n35337, n35338, n35339, n35340, n35342, n35343, n35344,
    n35345, n35346, n35348, n35349, n35351, n35352, n35353, n35354, n35355,
    n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363, n35365,
    n35366, n35367, n35368, n35369, n35371, n35372, n35373, n35375, n35376,
    n35377, n35378, n35379, n35381, n35382, n35383, n35384, n35385, n35386,
    n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35396, n35397,
    n35398, n35399, n35400, n35401, n35402, n35403, n35404, n35405, n35406,
    n35407, n35408, n35409, n35410, n35411, n35412, n35413, n35414, n35415,
    n35416, n35417, n35418, n35419, n35420, n35421, n35422, n35423, n35424,
    n35425, n35426, n35427, n35430, n35431, n35432, n35433, n35435, n35436,
    n35437, n35438, n35439, n35441, n35442, n35443, n35444, n35445, n35447,
    n35448, n35449, n35450, n35451, n35453, n35454, n35455, n35457, n35458,
    n35459, n35460, n35461, n35463, n35464, n35465, n35466, n35467, n35468,
    n35469, n35470, n35471, n35472, n35473, n35474, n35475, n35476, n35477,
    n35478, n35479, n35480, n35481, n35482, n35483, n35484, n35485, n35486,
    n35487, n35488, n35489, n35490, n35491, n35492, n35493, n35494, n35495,
    n35496, n35497, n35498, n35499, n35500, n35501, n35502, n35503, n35504,
    n35505, n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
    n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
    n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
    n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539, n35540,
    n35541, n35543, n35544, n35545, n35546, n35547, n35548, n35549, n35550,
    n35551, n35552, n35553, n35554, n35555, n35557, n35558, n35559, n35560,
    n35561, n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
    n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579,
    n35580, n35581, n35582, n35583, n35585, n35586, n35587, n35588, n35589,
    n35590, n35591, n35592, n35593, n35594, n35595, n35596, n35597, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605, n35606, n35607, n35608,
    n35609, n35610, n35611, n35613, n35614, n35615, n35616, n35617, n35618,
    n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
    n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635, n35636,
    n35637, n35638, n35639, n35640, n35641, n35642, n35643, n35644, n35645,
    n35646, n35647, n35648, n35649, n35650, n35651, n35652, n35653, n35654,
    n35655, n35656, n35657, n35658, n35659, n35660, n35661, n35662, n35664,
    n35665, n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
    n35674, n35675, n35676, n35678, n35679, n35680, n35681, n35682, n35683,
    n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35692, n35693,
    n35694, n35695, n35696, n35697, n35698, n35699, n35700, n35701, n35702,
    n35703, n35704, n35706, n35707, n35708, n35709, n35710, n35711, n35712,
    n35713, n35714, n35715, n35716, n35717, n35718, n35720, n35721, n35722,
    n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
    n35732, n35734, n35735, n35736, n35737, n35738, n35739, n35740, n35741,
    n35742, n35743, n35744, n35745, n35746, n35748, n35749, n35750, n35751,
    n35752, n35753, n35754, n35755, n35756, n35757, n35758, n35759, n35760,
    n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770,
    n35771, n35772, n35773, n35774, n35776, n35777, n35778, n35779, n35780,
    n35781, n35782, n35783, n35784, n35785, n35786, n35787, n35788, n35790,
    n35791, n35792, n35793, n35794, n35795, n35796, n35797, n35798, n35799,
    n35800, n35801, n35802, n35804, n35805, n35806, n35807, n35808, n35809,
    n35810, n35811, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
    n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827, n35828,
    n35829, n35830, n35831, n35832, n35833, n35834, n35835, n35836, n35837,
    n35838, n35839, n35840, n35841, n35842, n35843, n35844, n35845, n35846,
    n35847, n35848, n35849, n35850, n35851, n35852, n35853, n35854, n35855,
    n35856, n35857, n35858, n35859, n35860, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
    n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
    n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35891, n35892,
    n35893, n35895, n35896, n35897, n35898, n35899, n35901, n35902, n35904,
    n35905, n35906, n35908, n35909, n35910, n35911, n35912, n35913, n35914,
    n35915, n35918, n35919, n35920, n35921, n35924, n35925, n35927, n35928,
    n35929, n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
    n35938, n35939, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
    n35948, n35949, n35950, n35951, n35952, n35953, n35955, n35956, n35957,
    n35958, n35959, n35960, n35961, n35962, n35963, n35964, n35965, n35966,
    n35967, n35969, n35970, n35971, n35972, n35973, n35974, n35975, n35976,
    n35977, n35978, n35979, n35980, n35981, n35983, n35984, n35985, n35986,
    n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
    n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003, n36004,
    n36005, n36007, n36008, n36010, n36011, n36012, n36013, n36014, n36015,
    n36016, n36017, n36018, n36019, n36020, n36021, n36022, n36023, n36024,
    n36025, n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
    n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042,
    n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
    n36052, n36053, n36054, n36055, n36056, n36057, n36059, n36060, n36061,
    n36062, n36063, n36064, n36065, n36066, n36067, n36068, n36069, n36070,
    n36071, n36072, n36073, n36074, n36075, n36076, n36077, n36078, n36079,
    n36080, n36081, n36082, n36083, n36084, n36085, n36086, n36087, n36088,
    n36089, n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
    n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106,
    n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
    n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123, n36124,
    n36125, n36126, n36127, n36128, n36129, n36131, n36132, n36133, n36134,
    n36135, n36136, n36137, n36138, n36139, n36140, n36141, n36142, n36144,
    n36145, n36146, n36147, n36148, n36150, n36151, n36152, n36154, n36155,
    n36157, n36158, n36159, n36160, n36161, n36162, n36163, n36164, n36166,
    n36167, n36168, n36169, n36170, n36171, n36172, n36173, n36174, n36175,
    n36176, n36177, n36178, n36179, n36180, n36181, n36182, n36183, n36184,
    n36185, n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
    n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
    n36203, n36205, n36206, n36207, n36208, n36209, n36210, n36211, n36212,
    n36213, n36214, n36216, n36217, n36218, n36219, n36220, n36221, n36222,
    n36223, n36224, n36225, n36226, n36227, n36228, n36230, n36231, n36232,
    n36233, n36234, n36235, n36236, n36237, n36238, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36252,
    n36253, n36254, n36255, n36256, n36257, n36258, n36259, n36260, n36262,
    n36263, n36264, n36265, n36266, n36267, n36268, n36270, n36271, n36272,
    n36273, n36274, n36275, n36276, n36278, n36279, n36280, n36281, n36282,
    n36284, n36285, n36286, n36287, n36288, n36290, n36291, n36292, n36293,
    n36294, n36295, n36296, n36297, n36298, n36299, n36300, n36301, n36303,
    n36304, n36305, n36306, n36307, n36308, n36309, n36310, n36311, n36313,
    n36314, n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322,
    n36323, n36325, n36326, n36327, n36328, n36329, n36330, n36331, n36332,
    n36334, n36335, n36336, n36337, n36338, n36339, n36340, n36342, n36343,
    n36344, n36345, n36346, n36347, n36348, n36350, n36351, n36352, n36353,
    n36354, n36356, n36357, n36358, n36360, n36361, n36363, n36364, n36365,
    n36366, n36367, n36368, n36369, n36371, n36372, n36373, n36374, n36375,
    n36376, n36377, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
    n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395, n36396,
    n36397, n36398, n36399, n36400, n36401, n36402, n36403, n36404, n36405,
    n36406, n36407, n36408, n36409, n36410, n36411, n36412, n36413, n36414,
    n36415, n36416, n36417, n36418, n36419, n36420, n36421, n36422, n36423,
    n36424, n36425, n36426, n36427, n36428, n36429, n36430, n36431, n36432,
    n36433, n36434, n36435, n36436, n36437, n36438, n36439, n36440, n36441,
    n36442, n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
    n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
    n36460, n36461, n36463, n36464, n36465, n36466, n36467, n36468, n36469,
    n36470, n36471, n36472, n36473, n36474, n36476, n36477, n36478, n36479,
    n36480, n36481, n36482, n36483, n36484, n36485, n36486, n36488, n36489,
    n36490, n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498,
    n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507, n36508,
    n36509, n36510, n36512, n36513, n36514, n36515, n36516, n36517, n36518,
    n36519, n36520, n36521, n36522, n36524, n36525, n36526, n36527, n36528,
    n36530, n36531, n36533, n36534, n36536, n36537, n36538, n36539, n36540,
    n36541, n36542, n36543, n36544, n36545, n36546, n36547, n36548, n36549,
    n36550, n36551, n36552, n36553, n36554, n36555, n36556, n36558, n36559,
    n36560, n36561, n36562, n36563, n36564, n36565, n36566, n36567, n36568,
    n36569, n36570, n36571, n36572, n36573, n36574, n36575, n36576, n36577,
    n36578, n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
    n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
    n36596, n36597, n36598, n36599, n36600, n36601, n36603, n36604, n36606,
    n36607, n36608, n36609, n36610, n36611, n36612, n36613, n36614, n36615,
    n36616, n36618, n36619, n36621, n36622, n36623, n36624, n36625, n36626,
    n36627, n36628, n36629, n36630, n36631, n36632, n36634, n36635, n36636,
    n36637, n36638, n36639, n36640, n36641, n36642, n36643, n36644, n36646,
    n36647, n36648, n36649, n36650, n36651, n36652, n36653, n36654, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662, n36663, n36664, n36666,
    n36667, n36669, n36670, n36671, n36672, n36673, n36674, n36675, n36676,
    n36677, n36678, n36679, n36680, n36681, n36682, n36683, n36684, n36685,
    n36686, n36687, n36688, n36689, n36690, n36691, n36692, n36693, n36694,
    n36695, n36696, n36697, n36699, n36700, n36701, n36702, n36703, n36704,
    n36705, n36706, n36707, n36708, n36709, n36710, n36712, n36713, n36714,
    n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36724,
    n36725, n36726, n36727, n36728, n36729, n36730, n36731, n36732, n36733,
    n36734, n36736, n36737, n36739, n36740, n36742, n36743, n36745, n36746,
    n36748, n36749, n36751, n36752, n36754, n36755, n36756, n36757, n36758,
    n36759, n36760, n36761, n36763, n36764, n36765, n36766, n36767, n36768,
    n36769, n36770, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
    n36779, n36781, n36782, n36783, n36784, n36785, n36786, n36787, n36789,
    n36790, n36791, n36792, n36793, n36794, n36795, n36796, n36797, n36798,
    n36799, n36800, n36801, n36802, n36803, n36804, n36805, n36806, n36807,
    n36808, n36809, n36810, n36811, n36812, n36813, n36814, n36815, n36816,
    n36817, n36818, n36819, n36820, n36821, n36822, n36823, n36824, n36825,
    n36826, n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834,
    n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
    n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851, n36852,
    n36853, n36854, n36855, n36856, n36857, n36858, n36859, n36860, n36861,
    n36862, n36863, n36864, n36865, n36866, n36867, n36868, n36869, n36870,
    n36871, n36872, n36873, n36874, n36875, n36876, n36877, n36878, n36879,
    n36881, n36882, n36883, n36884, n36885, n36886, n36887, n36888, n36889,
    n36890, n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
    n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
    n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915, n36916,
    n36917, n36918, n36919, n36920, n36921, n36922, n36923, n36924, n36925,
    n36926, n36927, n36928, n36929, n36930, n36931, n36932, n36933, n36934,
    n36935, n36936, n36937, n36938, n36939, n36940, n36941, n36942, n36943,
    n36944, n36945, n36946, n36947, n36948, n36949, n36950, n36951, n36952,
    n36953, n36954, n36955, n36956, n36957, n36958, n36959, n36960, n36961,
    n36962, n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
    n36971, n36973, n36974, n36976, n36977, n36980, n36982, n36983, n36984,
    n36985, n36986, n36987, n36988, n36989, n36990, n36991, n36992, n36993,
    n36994, n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002,
    n37003, n37005, n37006, n37007, n37008, n37009, n37010, n37011, n37012,
    n37013, n37014, n37016, n37017, n37018, n37019, n37020, n37021, n37022,
    n37023, n37024, n37025, n37027, n37028, n37029, n37030, n37031, n37032,
    n37033, n37034, n37035, n37036, n37038, n37039, n37040, n37041, n37042,
    n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
    n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059, n37060,
    n37061, n37062, n37063, n37064, n37065, n37066, n37067, n37068, n37069,
    n37070, n37071, n37072, n37073, n37074, n37075, n37076, n37077, n37078,
    n37079, n37080, n37081, n37082, n37083, n37084, n37085, n37086, n37087,
    n37088, n37089, n37090, n37091, n37092, n37093, n37094, n37095, n37096,
    n37097, n37098, n37099, n37100, n37101, n37102, n37103, n37104, n37105,
    n37106, n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
    n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
    n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131, n37132,
    n37133, n37134, n37135, n37136, n37137, n37138, n37139, n37140, n37141,
    n37142, n37143, n37144, n37145, n37146, n37147, n37148, n37149, n37150,
    n37151, n37152, n37153, n37154, n37155, n37156, n37157, n37158, n37159,
    n37160, n37161, n37162, n37163, n37164, n37165, n37166, n37167, n37168,
    n37169, n37170, n37171, n37172, n37173, n37174, n37175, n37176, n37177,
    n37178, n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
    n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
    n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203, n37204,
    n37205, n37206, n37207, n37208, n37209, n37210, n37211, n37212, n37213,
    n37214, n37215, n37216, n37217, n37218, n37219, n37220, n37221, n37222,
    n37223, n37224, n37225, n37226, n37227, n37228, n37229, n37230, n37231,
    n37232, n37233, n37234, n37235, n37236, n37237, n37238, n37239, n37240,
    n37242, n37243, n37244, n37245, n37247, n37248, n37249, n37250, n37252,
    n37253, n37254, n37255, n37256, n37257, n37258, n37259, n37260, n37261,
    n37262, n37263, n37264, n37265, n37266, n37267, n37268, n37269, n37270,
    n37271, n37272, n37273, n37274, n37275, n37276, n37277, n37278, n37279,
    n37280, n37281, n37282, n37283, n37284, n37285, n37286, n37287, n37288,
    n37289, n37290, n37291, n37292, n37293, n37294, n37296, n37297, n37298,
    n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307,
    n37308, n37310, n37311, n37312, n37313, n37314, n37315, n37316, n37317,
    n37318, n37319, n37320, n37321, n37322, n37324, n37325, n37326, n37327,
    n37328, n37329, n37330, n37331, n37332, n37333, n37334, n37335, n37336,
    n37337, n37338, n37339, n37340, n37341, n37342, n37343, n37344, n37345,
    n37346, n37347, n37349, n37350, n37352, n37353, n37354, n37355, n37356,
    n37357, n37358, n37359, n37360, n37361, n37362, n37363, n37364, n37365,
    n37366, n37367, n37368, n37370, n37371, n37372, n37373, n37374, n37375,
    n37376, n37377, n37378, n37379, n37380, n37381, n37382, n37383, n37384,
    n37385, n37386, n37387, n37389, n37390, n37391, n37392, n37393, n37394,
    n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
    n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411, n37412,
    n37413, n37415, n37416, n37417, n37418, n37419, n37420, n37421, n37422,
    n37423, n37424, n37425, n37427, n37428, n37429, n37431, n37432, n37433,
    n37434, n37436, n37437, n37438, n37439, n37441, n37442, n37443, n37444,
    n37446, n37447, n37448, n37449, n37451, n37452, n37453, n37454, n37456,
    n37457, n37458, n37459, n37461, n37462, n37463, n37464, n37466, n37467,
    n37468, n37469, n37471, n37472, n37473, n37474, n37476, n37477, n37478,
    n37479, n37481, n37482, n37485, n37486, n37487, n37488, n37489, n37490,
    n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37500, n37501,
    n37502, n37503, n37504, n37505, n37506, n37507, n37508, n37509, n37510,
    n37511, n37512, n37514, n37515, n37516, n37517, n37518, n37519, n37520,
    n37521, n37522, n37523, n37524, n37525, n37526, n37528, n37529, n37530,
    n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539,
    n37540, n37542, n37543, n37544, n37545, n37546, n37547, n37548, n37549,
    n37550, n37551, n37552, n37553, n37554, n37556, n37557, n37558, n37559,
    n37560, n37561, n37562, n37563, n37564, n37565, n37566, n37567, n37568,
    n37570, n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578,
    n37579, n37580, n37581, n37582, n37584, n37585, n37586, n37587, n37588,
    n37589, n37590, n37591, n37592, n37593, n37594, n37595, n37596, n37597,
    n37598, n37599, n37600, n37601, n37602, n37603, n37604, n37605, n37606,
    n37607, n37608, n37609, n37611, n37612, n37613, n37614, n37615, n37616,
    n37617, n37618, n37619, n37620, n37621, n37622, n37623, n37624, n37625,
    n37626, n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635,
    n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643, n37644,
    n37645, n37646, n37647, n37648, n37649, n37650, n37651, n37652, n37653,
    n37654, n37655, n37656, n37657, n37658, n37659, n37660, n37661, n37662,
    n37663, n37664, n37665, n37666, n37667, n37668, n37670, n37671, n37672,
    n37673, n37674, n37675, n37676, n37677, n37678, n37679, n37680, n37681,
    n37682, n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
    n37692, n37693, n37694, n37695, n37696, n37698, n37699, n37700, n37701,
    n37702, n37703, n37704, n37706, n37707, n37708, n37709, n37710, n37711,
    n37713, n37714, n37715, n37716, n37717, n37718, n37719, n37720, n37721,
    n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731,
    n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739, n37740,
    n37741, n37742, n37743, n37744, n37745, n37746, n37747, n37748, n37749,
    n37750, n37751, n37752, n37753, n37755, n37756, n37757, n37758, n37759,
    n37760, n37761, n37762, n37764, n37765, n37766, n37767, n37768, n37769,
    n37770, n37771, n37773, n37774, n37775, n37776, n37777, n37778, n37779,
    n37780, n37781, n37782, n37783, n37785, n37786, n37787, n37788, n37789,
    n37790, n37791, n37792, n37793, n37794, n37795, n37796, n37797, n37799,
    n37800, n37801, n37802, n37803, n37804, n37805, n37806, n37807, n37808,
    n37809, n37810, n37811, n37813, n37814, n37815, n37816, n37817, n37818,
    n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37827, n37828,
    n37829, n37831, n37832, n37833, n37834, n37835, n37836, n37837, n37838,
    n37839, n37840, n37841, n37842, n37843, n37844, n37845, n37846, n37848,
    n37849, n37850, n37851, n37852, n37853, n37854, n37855, n37856, n37857,
    n37858, n37859, n37860, n37861, n37862, n37863, n37865, n37866, n37867,
    n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875, n37876,
    n37877, n37878, n37879, n37880, n37882, n37883, n37884, n37885, n37886,
    n37887, n37888, n37889, n37890, n37891, n37892, n37893, n37894, n37895,
    n37896, n37897, n37899, n37900, n37901, n37902, n37903, n37904, n37905,
    n37906, n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914,
    n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923, n37924,
    n37925, n37926, n37927, n37928, n37929, n37930, n37931, n37933, n37934,
    n37935, n37936, n37937, n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37950, n37951, n37952, n37953,
    n37954, n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962,
    n37963, n37964, n37965, n37967, n37968, n37969, n37970, n37971, n37972,
    n37973, n37974, n37975, n37976, n37977, n37978, n37979, n37981, n37982,
    n37983, n37984, n37985, n37986, n37987, n37988, n37989, n37990, n37991,
    n37992, n37993, n37995, n37996, n37997, n37998, n37999, n38000, n38001,
    n38002, n38003, n38004, n38005, n38006, n38007, n38009, n38010, n38011,
    n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019, n38020,
    n38021, n38023, n38024, n38025, n38026, n38027, n38028, n38029, n38030,
    n38031, n38032, n38033, n38034, n38035, n38037, n38038, n38039, n38040,
    n38041, n38042, n38043, n38044, n38045, n38046, n38047, n38048, n38049,
    n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059,
    n38060, n38061, n38062, n38063, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075, n38076, n38077, n38079,
    n38080, n38081, n38082, n38083, n38084, n38085, n38086, n38087, n38088,
    n38089, n38090, n38091, n38093, n38094, n38095, n38096, n38097, n38098,
    n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
    n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115, n38116,
    n38117, n38118, n38120, n38121, n38122, n38123, n38124, n38125, n38126,
    n38127, n38128, n38129, n38130, n38131, n38132, n38133, n38134, n38135,
    n38137, n38138, n38139, n38140, n38141, n38142, n38143, n38144, n38145,
    n38146, n38147, n38148, n38149, n38150, n38151, n38152, n38154, n38155,
    n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163, n38164,
    n38165, n38166, n38167, n38168, n38169, n38171, n38172, n38173, n38174,
    n38175, n38176, n38177, n38178, n38179, n38180, n38181, n38182, n38183,
    n38184, n38185, n38186, n38188, n38189, n38190, n38191, n38192, n38193,
    n38194, n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202,
    n38203, n38205, n38206, n38207, n38208, n38209, n38210, n38211, n38212,
    n38213, n38214, n38215, n38216, n38217, n38218, n38219, n38220, n38222,
    n38223, n38224, n38225, n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237, n38238, n38239, n38240,
    n38241, n38242, n38243, n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
    n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38267, n38268,
    n38269, n38270, n38272, n38273, n38274, n38276, n38277, n38278, n38279,
    n38280, n38281, n38282, n38283, n38284, n38285, n38286, n38287, n38288,
    n38289, n38290, n38291, n38292, n38293, n38294, n38295, n38296, n38297,
    n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307,
    n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315, n38316,
    n38317, n38318, n38319, n38320, n38321, n38322, n38324, n38325, n38326,
    n38327, n38328, n38329, n38330, n38331, n38333, n38334, n38335, n38336,
    n38337, n38338, n38339, n38340, n38342, n38343, n38344, n38345, n38346,
    n38347, n38348, n38349, n38351, n38352, n38354, n38355, n38356, n38357,
    n38358, n38360, n38361, n38363, n38364, n38365, n38366, n38367, n38368,
    n38370, n38371, n38372, n38373, n38374, n38376, n38377, n38379, n38380,
    n38381, n38382, n38383, n38384, n38385, n38386, n38387, n38388, n38389,
    n38391, n38392, n38393, n38394, n38395, n38396, n38397, n38398, n38399,
    n38400, n38401, n38403, n38404, n38405, n38406, n38407, n38408, n38409,
    n38410, n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38419,
    n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427, n38428,
    n38429, n38430, n38431, n38432, n38434, n38435, n38436, n38437, n38438,
    n38439, n38440, n38441, n38442, n38443, n38444, n38445, n38446, n38447,
    n38449, n38450, n38451, n38452, n38453, n38454, n38455, n38456, n38457,
    n38458, n38459, n38460, n38461, n38462, n38464, n38465, n38466, n38467,
    n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475, n38476,
    n38477, n38479, n38480, n38481, n38482, n38483, n38484, n38485, n38486,
    n38487, n38488, n38489, n38490, n38491, n38492, n38494, n38495, n38496,
    n38497, n38498, n38499, n38500, n38501, n38502, n38503, n38504, n38505,
    n38506, n38507, n38509, n38510, n38511, n38512, n38513, n38514, n38515,
    n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523, n38524,
    n38525, n38526, n38527, n38528, n38529, n38530, n38531, n38532, n38533,
    n38534, n38535, n38536, n38537, n38538, n38539, n38541, n38542, n38543,
    n38544, n38545, n38546, n38548, n38549, n38550, n38551, n38553, n38554,
    n38555, n38556, n38557, n38559, n38560, n38561, n38563, n38564, n38565,
    n38566, n38568, n38569, n38570, n38572, n38573, n38574, n38576, n38577,
    n38579, n38580, n38582, n38583, n38585, n38586, n38588, n38589, n38591,
    n38592, n38594, n38595, n38596, n38597, n38598, n38599, n38600, n38601,
    n38602, n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
    n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619,
    n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627, n38628,
    n38629, n38631, n38632, n38633, n38634, n38635, n38636, n38637, n38638,
    n38640, n38641, n38642, n38643, n38644, n38645, n38646, n38647, n38648,
    n38649, n38650, n38651, n38652, n38653, n38655, n38656, n38657, n38658,
    n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667,
    n38669, n38670, n38671, n38672, n38673, n38674, n38675, n38676, n38677,
    n38678, n38680, n38681, n38682, n38683, n38684, n38685, n38686, n38687,
    n38688, n38689, n38690, n38692, n38693, n38694, n38695, n38696, n38697,
    n38698, n38699, n38700, n38701, n38702, n38703, n38705, n38706, n38707,
    n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715, n38716,
    n38717, n38718, n38719, n38720, n38721, n38722, n38723, n38724, n38725,
    n38726, n38727, n38728, n38729, n38730, n38731, n38732, n38733, n38734,
    n38735, n38736, n38737, n38738, n38739, n38740, n38741, n38742, n38743,
    n38744, n38745, n38746, n38747, n38748, n38749, n38750, n38751, n38752,
    n38753, n38754, n38755, n38756, n38757, n38758, n38759, n38760, n38761,
    n38762, n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
    n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779,
    n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787, n38788,
    n38789, n38790, n38791, n38792, n38793, n38794, n38795, n38796, n38797,
    n38798, n38799, n38800, n38801, n38802, n38803, n38804, n38805, n38806,
    n38808, n38809, n38810, n38811, n38812, n38813, n38814, n38815, n38816,
    n38817, n38818, n38819, n38820, n38821, n38822, n38823, n38824, n38825,
    n38826, n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
    n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
    n38845, n38846, n38847, n38848, n38849, n38850, n38851, n38852, n38854,
    n38855, n38856, n38857, n38858, n38859, n38860, n38861, n38863, n38864,
    n38865, n38866, n38867, n38868, n38870, n38871, n38872, n38873, n38874,
    n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38883, n38884,
    n38885, n38886, n38887, n38888, n38889, n38890, n38891, n38892, n38893,
    n38895, n38896, n38897, n38898, n38899, n38900, n38901, n38902, n38903,
    n38904, n38905, n38906, n38907, n38908, n38909, n38910, n38911, n38912,
    n38913, n38915, n38916, n38917, n38918, n38919, n38920, n38922, n38923,
    n38924, n38926, n38927, n38928, n38930, n38931, n38932, n38934, n38935,
    n38936, n38938, n38939, n38940, n38942, n38943, n38944, n38946, n38947,
    n38948, n38950, n38951, n38952, n38954, n38955, n38956, n38958, n38959,
    n38960, n38962, n38963, n38964, n38965, n38966, n38967, n38969, n38970,
    n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38979, n38980,
    n38981, n38982, n38983, n38984, n38985, n38986, n38987, n38989, n38990,
    n38991, n38992, n38993, n38994, n38995, n38996, n38997, n38998, n38999,
    n39000, n39001, n39002, n39003, n39004, n39005, n39006, n39007, n39008,
    n39010, n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018,
    n39019, n39020, n39022, n39023, n39024, n39025, n39026, n39027, n39028,
    n39029, n39030, n39031, n39032, n39033, n39034, n39035, n39036, n39038,
    n39039, n39040, n39041, n39042, n39043, n39044, n39045, n39046, n39047,
    n39048, n39049, n39050, n39051, n39053, n39054, n39055, n39056, n39057,
    n39058, n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066,
    n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075, n39076,
    n39077, n39078, n39079, n39080, n39081, n39083, n39084, n39085, n39086,
    n39087, n39088, n39090, n39091, n39093, n39094, n39095, n39096, n39097,
    n39098, n39099, n39100, n39102, n39103, n39105, n39106, n39107, n39108,
    n39109, n39110, n39111, n39112, n39113, n39114, n39116, n39117, n39119,
    n39120, n39122, n39123, n39125, n39126, n39128, n39129, n39131, n39132,
    n39134, n39135, n39136, n39137, n39138, n39139, n39140, n39141, n39143,
    n39144, n39145, n39146, n39147, n39148, n39149, n39150, n39152, n39154,
    n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39164, n39165,
    n39166, n39167, n39168, n39169, n39170, n39172, n39173, n39174, n39175,
    n39176, n39177, n39178, n39179, n39180, n39181, n39182, n39183, n39184,
    n39186, n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39195,
    n39196, n39197, n39198, n39199, n39200, n39201, n39203, n39204, n39205,
    n39206, n39207, n39208, n39209, n39211, n39212, n39213, n39214, n39215,
    n39216, n39217, n39219, n39220, n39221, n39222, n39223, n39224, n39225,
    n39226, n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235,
    n39236, n39237, n39238, n39239, n39240, n39241, n39243, n39244, n39245,
    n39246, n39247, n39248, n39249, n39250, n39251, n39252, n39253, n39254,
    n39256, n39257, n39258, n39259, n39260, n39261, n39262, n39263, n39264,
    n39265, n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39275,
    n39276, n39279, n39280, n39281, n39282, n39283, n39284, n39285, n39286,
    n39287, n39288, n39289, n39290, n39291, n39292, n39293, n39294, n39295,
    n39296, n39297, n39298, n39299, n39300, n39301, n39302, n39303, n39304,
    n39305, n39306, n39307, n39308, n39309, n39310, n39311, n39312, n39313,
    n39314, n39315, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
    n39324, n39326, n39327, n39328, n39329, n39330, n39332, n39333, n39334,
    n39335, n39336, n39337, n39338, n39340, n39341, n39342, n39344, n39345,
    n39346, n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355,
    n39356, n39357, n39358, n39359, n39361, n39362, n39363, n39365, n39366,
    n39367, n39369, n39370, n39371, n39373, n39374, n39375, n39376, n39377,
    n39378, n39380, n39381, n39382, n39384, n39385, n39386, n39388, n39389,
    n39390, n39392, n39393, n39394, n39395, n39396, n39397, n39399, n39400,
    n39401, n39403, n39404, n39405, n39407, n39408, n39409, n39411, n39412,
    n39413, n39415, n39416, n39417, n39419, n39420, n39421, n39422, n39423,
    n39425, n39426, n39427, n39428, n39429, n39431, n39432, n39433, n39434,
    n39435, n39437, n39438, n39439, n39440, n39441, n39443, n39444, n39445,
    n39446, n39447, n39449, n39450, n39451, n39452, n39453, n39455, n39456,
    n39457, n39458, n39459, n39461, n39462, n39463, n39464, n39465, n39467,
    n39468, n39469, n39470, n39471, n39473, n39474, n39475, n39476, n39477,
    n39479, n39480, n39481, n39482, n39483, n39485, n39486, n39487, n39488,
    n39489, n39491, n39492, n39493, n39494, n39495, n39497, n39498, n39499,
    n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507, n39508,
    n39509, n39510, n39511, n39512, n39513, n39514, n39515, n39516, n39517,
    n39518, n39519, n39520, n39521, n39522, n39523, n39524, n39525, n39526,
    n39527, n39528, n39529, n39530, n39531, n39532, n39533, n39534, n39535,
    n39536, n39537, n39539, n39540, n39541, n39542, n39543, n39544, n39545,
    n39546, n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
    n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563, n39564,
    n39565, n39566, n39567, n39568, n39569, n39570, n39571, n39572, n39573,
    n39574, n39575, n39576, n39577, n39578, n39579, n39580, n39581, n39582,
    n39583, n39584, n39585, n39586, n39588, n39589, n39590, n39591, n39592,
    n39593, n39594, n39595, n39596, n39597, n39598, n39599, n39600, n39602,
    n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611,
    n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619, n39620,
    n39621, n39622, n39623, n39624, n39625, n39626, n39627, n39628, n39629,
    n39630, n39631, n39632, n39633, n39634, n39635, n39636, n39638, n39639,
    n39640, n39641, n39642, n39643, n39644, n39645, n39646, n39647, n39648,
    n39649, n39650, n39651, n39652, n39653, n39654, n39655, n39656, n39657,
    n39658, n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
    n39667, n39668, n39669, n39670, n39671, n39673, n39674, n39675, n39676,
    n39677, n39678, n39679, n39680, n39681, n39682, n39683, n39684, n39685,
    n39686, n39687, n39688, n39689, n39690, n39691, n39692, n39693, n39694,
    n39695, n39696, n39697, n39698, n39699, n39700, n39701, n39702, n39703,
    n39704, n39705, n39706, n39707, n39708, n39709, n39710, n39712, n39713,
    n39714, n39715, n39716, n39718, n39719, n39720, n39721, n39722, n39723,
    n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731, n39732,
    n39733, n39734, n39735, n39736, n39737, n39738, n39739, n39740, n39741,
    n39743, n39744, n39745, n39746, n39747, n39748, n39749, n39750, n39751,
    n39752, n39753, n39754, n39755, n39756, n39757, n39758, n39759, n39760,
    n39761, n39762, n39763, n39764, n39765, n39766, n39768, n39769, n39770,
    n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
    n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787, n39788,
    n39789, n39790, n39791, n39793, n39794, n39795, n39796, n39797, n39798,
    n39799, n39800, n39801, n39802, n39803, n39804, n39805, n39806, n39807,
    n39808, n39809, n39810, n39811, n39812, n39813, n39814, n39815, n39817,
    n39818, n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
    n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
    n39836, n39837, n39838, n39839, n39840, n39842, n39843, n39844, n39845,
    n39846, n39847, n39849, n39850, n39851, n39852, n39853, n39854, n39856,
    n39857, n39858, n39859, n39861, n39862, n39863, n39864, n39866, n39867,
    n39868, n39870, n39871, n39873, n39874, n39876, n39877, n39879, n39880,
    n39881, n39882, n39883, n39884, n39885, n39886, n39887, n39888, n39889,
    n39890, n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
    n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
    n39908, n39909, n39910, n39912, n39913, n39914, n39915, n39916, n39918,
    n39919, n39920, n39921, n39922, n39924, n39925, n39926, n39927, n39928,
    n39930, n39931, n39932, n39933, n39934, n39936, n39937, n39938, n39939,
    n39940, n39941, n39943, n39944, n39945, n39946, n39947, n39948, n39949,
    n39950, n39951, n39952, n39954, n39955, n39956, n39958, n39959, n39960,
    n39961, n39962, n39963, n39964, n39965, n39967, n39968, n39969, n39970,
    n39971, n39972, n39973, n39974, n39976, n39977, n39978, n39979, n39980,
    n39981, n39982, n39983, n39984, n39985, n39986, n39988, n39989, n39990,
    n39992, n39993, n39994, n39995, n39996, n39997, n39998, n39999, n40000,
    n40001, n40002, n40003, n40004, n40005, n40006, n40007, n40008, n40009,
    n40010, n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
    n40019, n40020, n40021, n40022, n40024, n40025, n40026, n40027, n40028,
    n40029, n40030, n40031, n40032, n40033, n40034, n40035, n40036, n40037,
    n40038, n40039, n40040, n40041, n40042, n40043, n40044, n40045, n40046,
    n40047, n40048, n40049, n40050, n40051, n40052, n40053, n40054, n40056,
    n40057, n40058, n40059, n40060, n40061, n40062, n40063, n40064, n40065,
    n40066, n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
    n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083,
    n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091, n40092,
    n40093, n40095, n40096, n40097, n40098, n40099, n40100, n40101, n40102,
    n40103, n40104, n40105, n40106, n40107, n40108, n40109, n40110, n40111,
    n40112, n40113, n40114, n40115, n40116, n40117, n40118, n40119, n40120,
    n40121, n40122, n40123, n40124, n40125, n40126, n40127, n40128, n40129,
    n40130, n40131, n40132, n40134, n40135, n40136, n40137, n40138, n40139,
    n40140, n40141, n40142, n40143, n40145, n40146, n40147, n40148, n40149,
    n40150, n40151, n40152, n40153, n40154, n40155, n40156, n40157, n40158,
    n40159, n40160, n40161, n40162, n40163, n40164, n40165, n40166, n40167,
    n40168, n40169, n40170, n40171, n40172, n40174, n40175, n40176, n40177,
    n40178, n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
    n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
    n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203, n40204,
    n40205, n40206, n40207, n40208, n40209, n40210, n40211, n40213, n40214,
    n40215, n40216, n40217, n40218, n40219, n40220, n40221, n40222, n40223,
    n40224, n40225, n40226, n40227, n40228, n40229, n40230, n40231, n40232,
    n40233, n40234, n40235, n40236, n40237, n40238, n40239, n40240, n40241,
    n40242, n40243, n40244, n40245, n40246, n40248, n40249, n40250, n40251,
    n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259, n40260,
    n40261, n40262, n40263, n40264, n40265, n40266, n40267, n40268, n40269,
    n40270, n40271, n40272, n40273, n40274, n40275, n40276, n40277, n40278,
    n40279, n40280, n40281, n40283, n40284, n40285, n40286, n40287, n40288,
    n40289, n40290, n40291, n40292, n40293, n40294, n40295, n40296, n40297,
    n40298, n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306,
    n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315,
    n40316, n40318, n40319, n40320, n40321, n40322, n40323, n40324, n40325,
    n40326, n40327, n40328, n40329, n40330, n40331, n40332, n40333, n40334,
    n40335, n40336, n40337, n40338, n40339, n40340, n40341, n40342, n40343,
    n40344, n40345, n40346, n40347, n40348, n40350, n40351, n40352, n40353,
    n40354, n40355, n40356, n40357, n40359, n40360, n40361, n40362, n40363,
    n40364, n40365, n40366, n40368, n40369, n40370, n40371, n40372, n40373,
    n40374, n40375, n40376, n40377, n40378, n40380, n40381, n40382, n40383,
    n40384, n40386, n40387, n40388, n40389, n40390, n40392, n40393, n40395,
    n40396, n40397, n40398, n40400, n40401, n40402, n40403, n40404, n40405,
    n40406, n40407, n40408, n40409, n40410, n40411, n40412, n40413, n40414,
    n40415, n40416, n40417, n40418, n40419, n40420, n40421, n40422, n40424,
    n40425, n40426, n40428, n40429, n40430, n40432, n40433, n40435, n40436,
    n40437, n40439, n40440, n40441, n40442, n40443, n40444, n40445, n40446,
    n40448, n40449, n40450, n40451, n40452, n40453, n40454, n40455, n40456,
    n40457, n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466,
    n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475,
    n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483, n40484,
    n40485, n40487, n40488, n40489, n40490, n40491, n40492, n40493, n40494,
    n40495, n40496, n40497, n40502, n40503, n40504, n40506, n40507, n40508,
    n40510, n40511, n40512, n40514, n40515, n40516, n40518, n40519, n40520,
    n40522, n40523, n40525, n40526, n40527, n40529, n40530, n40531, n40533,
    n40534, n40536, n40537, n40538, n40540, n40541, n40542, n40543, n40544,
    n40545, n40547, n40548, n40549, n40551, n40552, n40553, n40555, n40556,
    n40557, n40559, n40560, n40562, n40563, n40565, n40566, n40568, n40569,
    n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
    n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587, n40588,
    n40589, n40590, n40591, n40592, n40593, n40594, n40595, n40596, n40597,
    n40598, n40599, n40600, n40601, n40602, n40603, n40604, n40605, n40606,
    n40607, n40608, n40609, n40610, n40611, n40612, n40613, n40614, n40615,
    n40616, n40617, n40618, n40619, n40620, n40621, n40622, n40623, n40624,
    n40625, n40626, n40627, n40628, n40629, n40630, n40631, n40632, n40633,
    n40634, n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
    n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
    n40653, n40654, n40655, n40657, n40658, n40659, n40661, n40662, n40663,
    n40664, n40665, n40666, n40667, n40668, n40669, n40670, n40671, n40672,
    n40673, n40674, n40675, n40676, n40677, n40678, n40679, n40680, n40681,
    n40682, n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
    n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
    n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707, n40708,
    n40709, n40710, n40711, n40712, n40713, n40714, n40715, n40716, n40717,
    n40718, n40719, n40720, n40721, n40722, n40723, n40724, n40725, n40726,
    n40727, n40728, n40729, n40730, n40731, n40732, n40733, n40734, n40735,
    n40736, n40737, n40738, n40739, n40740, n40741, n40743, n40744, n40745,
    n40746, n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
    n40755, n40756, n40757, n40758, n40759, n40760, n40762, n40763, n40764,
    n40765, n40766, n40767, n40768, n40769, n40770, n40771, n40772, n40774,
    n40775, n40776, n40777, n40778, n40779, n40780, n40781, n40782, n40783,
    n40784, n40786, n40787, n40788, n40789, n40790, n40791, n40792, n40793,
    n40794, n40795, n40796, n40797, n40799, n40800, n40801, n40802, n40803,
    n40804, n40805, n40806, n40807, n40808, n40810, n40811, n40812, n40813,
    n40814, n40815, n40816, n40817, n40818, n40819, n40821, n40822, n40823,
    n40824, n40825, n40826, n40827, n40828, n40829, n40830, n40831, n40833,
    n40834, n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842,
    n40843, n40844, n40845, n40846, n40847, n40848, n40850, n40851, n40852,
    n40853, n40854, n40855, n40856, n40857, n40858, n40859, n40860, n40861,
    n40862, n40864, n40865, n40866, n40867, n40868, n40869, n40870, n40871,
    n40872, n40873, n40874, n40875, n40876, n40877, n40879, n40880, n40881,
    n40882, n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
    n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
    n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907, n40908,
    n40909, n40910, n40911, n40912, n40914, n40915, n40916, n40917, n40918,
    n40919, n40920, n40921, n40922, n40923, n40924, n40925, n40926, n40927,
    n40928, n40929, n40930, n40931, n40932, n40933, n40934, n40935, n40936,
    n40937, n40938, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
    n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
    n40956, n40957, n40958, n40959, n40960, n40961, n40963, n40964, n40965,
    n40966, n40967, n40968, n40969, n40970, n40971, n40972, n40973, n40974,
    n40975, n40976, n40977, n40978, n40979, n40980, n40981, n40982, n40983,
    n40984, n40985, n40987, n40988, n40989, n40990, n40991, n40992, n40993,
    n40994, n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
    n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41012,
    n41013, n41014, n41015, n41016, n41017, n41018, n41019, n41020, n41021,
    n41022, n41023, n41024, n41025, n41026, n41027, n41028, n41029, n41030,
    n41031, n41032, n41033, n41035, n41036, n41037, n41038, n41039, n41040,
    n41041, n41042, n41043, n41044, n41045, n41046, n41047, n41048, n41049,
    n41050, n41051, n41052, n41053, n41054, n41055, n41056, n41058, n41059,
    n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067, n41068,
    n41069, n41070, n41071, n41072, n41073, n41074, n41075, n41076, n41077,
    n41078, n41079, n41081, n41082, n41083, n41084, n41085, n41086, n41088,
    n41089, n41090, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
    n41099, n41100, n41101, n41102, n41104, n41105, n41106, n41107, n41108,
    n41109, n41110, n41111, n41113, n41114, n41115, n41116, n41117, n41118,
    n41119, n41120, n41122, n41123, n41124, n41125, n41126, n41127, n41128,
    n41129, n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
    n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147, n41149,
    n41150, n41151, n41152, n41153, n41154, n41155, n41156, n41158, n41159,
    n41160, n41161, n41162, n41163, n41164, n41165, n41166, n41167, n41168,
    n41169, n41170, n41171, n41172, n41173, n41174, n41175, n41176, n41177,
    n41178, n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
    n41188, n41189, n41190, n41191, n41192, n41194, n41195, n41196, n41197,
    n41198, n41200, n41201, n41202, n41203, n41204, n41205, n41206, n41207,
    n41209, n41210, n41211, n41212, n41213, n41215, n41216, n41217, n41218,
    n41219, n41220, n41221, n41222, n41224, n41225, n41226, n41227, n41228,
    n41229, n41230, n41231, n41234, n41235, n41236, n41237, n41238, n41239,
    n41240, n41241, n41242, n41243, n41244, n41245, n41246, n41247, n41248,
    n41249, n41250, n41251, n41252, n41253, n41254, n41255, n41256, n41257,
    n41258, n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
    n41267, n41268, n41269, n41270, n41272, n41273, n41274, n41275, n41276,
    n41277, n41278, n41279, n41280, n41281, n41282, n41283, n41284, n41285,
    n41286, n41287, n41288, n41289, n41290, n41292, n41293, n41294, n41295,
    n41296, n41297, n41298, n41299, n41300, n41301, n41302, n41303, n41304,
    n41305, n41306, n41307, n41308, n41309, n41310, n41311, n41312, n41313,
    n41314, n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322,
    n41323, n41324, n41325, n41326, n41327, n41329, n41331, n41332, n41333,
    n41334, n41335, n41336, n41337, n41338, n41340, n41341, n41342, n41343,
    n41344, n41345, n41346, n41347, n41349, n41350, n41351, n41353, n41354,
    n41355, n41356, n41357, n41358, n41359, n41360, n41362, n41363, n41364,
    n41365, n41366, n41367, n41368, n41369, n41371, n41372, n41373, n41375,
    n41376, n41377, n41378, n41379, n41380, n41382, n41383, n41384, n41385,
    n41386, n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394,
    n41396, n41397, n41399, n41400, n41402, n41403, n41405, n41406, n41408,
    n41409, n41411, n41412, n41413, n41415, n41416, n41417, n41419, n41420,
    n41421, n41423, n41424, n41425, n41427, n41428, n41429, n41431, n41432,
    n41433, n41435, n41436, n41437, n41439, n41440, n41441, n41443, n41444,
    n41445, n41447, n41448, n41449, n41451, n41452, n41454, n41455, n41457,
    n41458, n41460, n41461, n41463, n41464, n41465, n41467, n41468, n41469,
    n41471, n41472, n41473, n41475, n41476, n41478, n41479, n41481, n41482,
    n41483, n41485, n41486, n41488, n41489, n41490, n41491, n41492, n41493,
    n41494, n41495, n41496, n41497, n41498, n41499, n41500, n41502, n41503,
    n41504, n41505, n41506, n41507, n41508, n41509, n41510, n41511, n41512,
    n41513, n41514, n41515, n41517, n41518, n41519, n41520, n41521, n41522,
    n41523, n41524, n41525, n41527, n41528, n41529, n41530, n41531, n41532,
    n41533, n41534, n41535, n41536, n41537, n41538, n41539, n41540, n41541,
    n41542, n41543, n41544, n41545, n41546, n41547, n41548, n41549, n41550,
    n41551, n41552, n41553, n41554, n41556, n41557, n41559, n41560, n41562,
    n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
    n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579, n41580,
    n41581, n41582, n41584, n41585, n41586, n41587, n41588, n41589, n41590,
    n41591, n41592, n41593, n41594, n41595, n41596, n41597, n41598, n41599,
    n41600, n41601, n41602, n41604, n41605, n41607, n41608, n41609, n41610,
    n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41620, n41621,
    n41622, n41624, n41625, n41626, n41627, n41629, n41630, n41631, n41632,
    n41633, n41635, n41636, n41637, n41638, n41640, n41641, n41642, n41643,
    n41645, n41646, n41647, n41648, n41650, n41651, n41652, n41653, n41655,
    n41656, n41657, n41659, n41660, n41661, n41663, n41664, n41665, n41667,
    n41668, n41669, n41671, n41672, n41673, n41674, n41675, n41677, n41678,
    n41679, n41680, n41682, n41683, n41684, n41686, n41687, n41688, n41690,
    n41691, n41692, n41694, n41695, n41696, n41698, n41699, n41700, n41701,
    n41702, n41703, n41704, n41705, n41706, n41707, n41708, n41709, n41710,
    n41711, n41712, n41713, n41714, n41715, n41716, n41717, n41718, n41719,
    n41720, n41721, n41722, n41723, n41724, n41726, n41727, n41728, n41729,
    n41730, n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
    n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747,
    n41748, n41749, n41750, n41751, n41752, n41756, n41757, n41758, n41759,
    n41760, n41761, n41762, n41763, n41764, n41765, n41766, n41767, n41768,
    n41769, n41770, n41771, n41772, n41773, n41774, n41775, n41776, n41777,
    n41778, n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
    n41787, n41788, n41790, n41791, n41792, n41793, n41794, n41795, n41796,
    n41797, n41798, n41799, n41800, n41801, n41802, n41803, n41804, n41805,
    n41806, n41807, n41808, n41809, n41810, n41811, n41813, n41814, n41815,
    n41816, n41817, n41818, n41819, n41820, n41821, n41822, n41823, n41825,
    n41826, n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
    n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843,
    n41844, n41845, n41847, n41848, n41850, n41851, n41852, n41853, n41855,
    n41856, n41858, n41859, n41860, n41862, n41863, n41864, n41865, n41867,
    n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875, n41876,
    n41877, n41878, n41879, n41880, n41881, n41882, n41883, n41884, n41885,
    n41886, n41887, n41888, n41889, n41890, n41891, n41892, n41893, n41894,
    n41895, n41896, n41898, n41899, n41901, n41902, n41903, n41904, n41905,
    n41906, n41907, n41908, n41910, n41911, n41912, n41913, n41914, n41915,
    n41916, n41917, n41918, n41919, n41920, n41922, n41923, n41924, n41926,
    n41927, n41929, n41930, n41931, n41933, n41934, n41935, n41936, n41937,
    n41938, n41939, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
    n41948, n41949, n41950, n41952, n41953, n41954, n41955, n41956, n41957,
    n41958, n41959, n41960, n41961, n41963, n41964, n41965, n41966, n41967,
    n41968, n41969, n41970, n41971, n41972, n41974, n41975, n41976, n41977,
    n41978, n41979, n41980, n41981, n41982, n41983, n41985, n41986, n41987,
    n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41996, n41997,
    n41998, n41999, n42000, n42001, n42002, n42003, n42004, n42005, n42006,
    n42007, n42008, n42009, n42010, n42011, n42012, n42013, n42015, n42016,
    n42017, n42018, n42019, n42020, n42021, n42022, n42023, n42024, n42025,
    n42026, n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42036,
    n42037, n42039, n42040, n42042, n42043, n42045, n42046, n42048, n42049,
    n42050, n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
    n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
    n42068, n42069, n42070, n42071, n42072, n42073, n42075, n42076, n42077,
    n42078, n42079, n42080, n42081, n42082, n42083, n42084, n42085, n42086,
    n42087, n42088, n42089, n42090, n42091, n42092, n42093, n42094, n42095,
    n42096, n42097, n42098, n42099, n42100, n42102, n42103, n42104, n42105,
    n42106, n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
    n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123,
    n42124, n42125, n42126, n42127, n42129, n42130, n42132, n42133, n42135,
    n42136, n42138, n42139, n42141, n42142, n42143, n42144, n42145, n42146,
    n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
    n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163, n42164,
    n42165, n42166, n42168, n42169, n42170, n42171, n42172, n42173, n42174,
    n42175, n42177, n42178, n42179, n42180, n42181, n42182, n42183, n42184,
    n42185, n42186, n42187, n42188, n42189, n42190, n42191, n42192, n42193,
    n42194, n42195, n42197, n42198, n42200, n42201, n42202, n42203, n42204,
    n42205, n42206, n42208, n42209, n42210, n42211, n42212, n42213, n42214,
    n42216, n42217, n42218, n42219, n42220, n42221, n42222, n42223, n42224,
    n42225, n42226, n42227, n42228, n42229, n42230, n42232, n42233, n42235,
    n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243, n42244,
    n42246, n42247, n42248, n42249, n42250, n42251, n42252, n42253, n42255,
    n42256, n42257, n42258, n42259, n42260, n42261, n42262, n42263, n42264,
    n42266, n42267, n42268, n42270, n42271, n42272, n42273, n42275, n42276,
    n42277, n42278, n42279, n42280, n42281, n42282, n42283, n42284, n42285,
    n42286, n42287, n42288, n42289, n42291, n42292, n42294, n42295, n42297,
    n42298, n42300, n42301, n42303, n42304, n42306, n42307, n42309, n42310,
    n42312, n42313, n42314, n42315, n42316, n42317, n42319, n42320, n42321,
    n42322, n42323, n42324, n42326, n42327, n42328, n42329, n42330, n42331,
    n42333, n42334, n42335, n42336, n42337, n42338, n42340, n42341, n42342,
    n42343, n42344, n42345, n42347, n42348, n42349, n42350, n42351, n42352,
    n42354, n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
    n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371, n42373,
    n42374, n42375, n42376, n42377, n42378, n42379, n42381, n42382, n42383,
    n42384, n42385, n42386, n42387, n42388, n42390, n42391, n42392, n42393,
    n42394, n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
    n42403, n42405, n42406, n42407, n42408, n42409, n42410, n42411, n42412,
    n42414, n42415, n42416, n42417, n42418, n42419, n42420, n42421, n42423,
    n42424, n42425, n42426, n42427, n42428, n42429, n42430, n42431, n42433,
    n42434, n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
    n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451,
    n42452, n42453, n42454, n42455, n42456, n42458, n42459, n42461, n42462,
    n42463, n42464, n42465, n42466, n42467, n42468, n42469, n42470, n42471,
    n42472, n42473, n42474, n42476, n42477, n42478, n42479, n42480, n42481,
    n42482, n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
    n42491, n42492, n42493, n42494, n42495, n42497, n42498, n42499, n42500,
    n42501, n42502, n42503, n42504, n42505, n42506, n42507, n42509, n42510,
    n42511, n42512, n42513, n42514, n42515, n42516, n42518, n42519, n42520,
    n42521, n42522, n42523, n42524, n42525, n42526, n42527, n42528, n42529,
    n42530, n42531, n42532, n42535, n42536, n42537, n42538, n42539, n42540,
    n42541, n42542, n42543, n42544, n42545, n42546, n42547, n42548, n42550,
    n42551, n42552, n42553, n42554, n42555, n42556, n42557, n42558, n42559,
    n42560, n42561, n42562, n42563, n42564, n42566, n42567, n42568, n42569,
    n42570, n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42579,
    n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587, n42588,
    n42589, n42591, n42592, n42593, n42594, n42595, n42596, n42597, n42598,
    n42599, n42600, n42601, n42603, n42604, n42605, n42606, n42607, n42608,
    n42609, n42610, n42611, n42612, n42613, n42614, n42615, n42616, n42617,
    n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627,
    n42628, n42629, n42631, n42632, n42633, n42634, n42635, n42636, n42637,
    n42638, n42640, n42641, n42642, n42643, n42644, n42645, n42647, n42648,
    n42649, n42650, n42651, n42652, n42653, n42654, n42655, n42656, n42657,
    n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42668,
    n42669, n42670, n42671, n42672, n42673, n42675, n42676, n42677, n42678,
    n42679, n42680, n42681, n42683, n42684, n42685, n42687, n42688, n42689,
    n42691, n42692, n42693, n42694, n42695, n42696, n42698, n42699, n42700,
    n42701, n42702, n42703, n42705, n42706, n42707, n42708, n42709, n42710,
    n42711, n42713, n42714, n42715, n42716, n42717, n42718, n42719, n42721,
    n42722, n42723, n42724, n42725, n42726, n42727, n42729, n42730, n42731,
    n42732, n42733, n42734, n42735, n42737, n42738, n42739, n42740, n42741,
    n42742, n42743, n42745, n42746, n42747, n42748, n42749, n42750, n42751,
    n42752, n42753, n42754, n42755, n42756, n42757, n42758, n42759, n42760,
    n42762, n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771,
    n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779, n42780,
    n42781, n42782, n42783, n42784, n42785, n42786, n42787, n42790, n42791,
    n42792, n42793, n42795, n42796, n42797, n42798, n42799, n42801, n42802,
    n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811,
    n42812, n42813, n42814, n42816, n42817, n42818, n42819, n42820, n42821,
    n42822, n42823, n42824, n42825, n42826, n42828, n42829, n42830, n42831,
    n42832, n42833, n42834, n42835, n42836, n42837, n42838, n42840, n42841,
    n42842, n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
    n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859, n42860,
    n42861, n42862, n42864, n42865, n42866, n42867, n42868, n42869, n42870,
    n42871, n42872, n42873, n42874, n42876, n42877, n42878, n42879, n42880,
    n42881, n42882, n42883, n42884, n42885, n42886, n42888, n42889, n42890,
    n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42900,
    n42901, n42902, n42903, n42904, n42905, n42906, n42907, n42908, n42909,
    n42910, n42912, n42913, n42914, n42915, n42916, n42917, n42918, n42919,
    n42920, n42921, n42922, n42924, n42925, n42926, n42927, n42928, n42929,
    n42930, n42931, n42932, n42933, n42934, n42936, n42937, n42938, n42939,
    n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42948, n42949,
    n42950, n42951, n42952, n42953, n42954, n42955, n42956, n42957, n42958,
    n42960, n42961, n42962, n42963, n42964, n42965, n42966, n42967, n42968,
    n42969, n42970, n42972, n42973, n42974, n42975, n42976, n42977, n42978,
    n42980, n42981, n42982, n42983, n42984, n42986, n42987, n42988, n42989,
    n42990, n42992, n42993, n42994, n42995, n42996, n42998, n42999, n43000,
    n43001, n43002, n43004, n43005, n43006, n43007, n43008, n43010, n43011,
    n43012, n43013, n43014, n43016, n43017, n43018, n43019, n43020, n43022,
    n43023, n43024, n43025, n43026, n43028, n43029, n43030, n43031, n43032,
    n43034, n43035, n43036, n43037, n43038, n43040, n43041, n43042, n43043,
    n43044, n43046, n43047, n43048, n43049, n43050, n43052, n43053, n43054,
    n43055, n43056, n43058, n43059, n43060, n43061, n43062, n43063, n43064,
    n43065, n43067, n43068, n43069, n43070, n43071, n43073, n43074, n43075,
    n43076, n43077, n43079, n43080, n43081, n43082, n43083, n43085, n43086,
    n43087, n43088, n43089, n43091, n43092, n43093, n43094, n43095, n43097,
    n43098, n43099, n43100, n43101, n43103, n43104, n43105, n43106, n43107,
    n43109, n43110, n43111, n43112, n43113, n43115, n43116, n43117, n43118,
    n43119, n43121, n43122, n43123, n43124, n43125, n43127, n43128, n43129,
    n43130, n43131, n43133, n43134, n43135, n43136, n43137, n43139, n43140,
    n43141, n43142, n43143, n43145, n43146, n43147, n43148, n43149, n43150,
    n43151, n43153, n43154, n43155, n43156, n43157, n43159, n43160, n43161,
    n43162, n43163, n43165, n43166, n43167, n43168, n43169, n43171, n43172,
    n43173, n43174, n43175, n43177, n43178, n43179, n43180, n43181, n43183,
    n43184, n43185, n43186, n43187, n43189, n43190, n43191, n43192, n43193,
    n43195, n43196, n43197, n43198, n43199, n43201, n43202, n43203, n43204,
    n43205, n43207, n43208, n43209, n43210, n43211, n43213, n43214, n43215,
    n43216, n43217, n43219, n43220, n43221, n43222, n43223, n43225, n43226,
    n43227, n43228, n43229, n43231, n43232, n43233, n43234, n43235, n43236,
    n43237, n43239, n43240, n43241, n43242, n43243, n43245, n43246, n43247,
    n43248, n43249, n43251, n43252, n43253, n43254, n43255, n43257, n43258,
    n43259, n43260, n43261, n43263, n43264, n43265, n43266, n43267, n43269,
    n43270, n43271, n43272, n43273, n43275, n43276, n43277, n43278, n43279,
    n43281, n43282, n43283, n43284, n43285, n43287, n43288, n43289, n43290,
    n43291, n43293, n43294, n43295, n43296, n43297, n43299, n43300, n43301,
    n43302, n43303, n43305, n43306, n43307, n43308, n43309, n43311, n43312,
    n43313, n43314, n43315, n43317, n43318, n43319, n43320, n43321, n43322,
    n43324, n43325, n43326, n43327, n43328, n43330, n43331, n43332, n43333,
    n43334, n43336, n43337, n43338, n43339, n43340, n43342, n43343, n43344,
    n43345, n43346, n43348, n43349, n43350, n43351, n43352, n43354, n43355,
    n43356, n43357, n43358, n43360, n43361, n43362, n43363, n43364, n43366,
    n43367, n43368, n43369, n43370, n43372, n43373, n43374, n43375, n43376,
    n43378, n43379, n43380, n43381, n43382, n43384, n43385, n43386, n43387,
    n43388, n43390, n43391, n43392, n43393, n43394, n43396, n43397, n43398,
    n43399, n43400, n43402, n43403, n43404, n43405, n43406, n43407, n43408,
    n43410, n43411, n43412, n43413, n43414, n43416, n43417, n43418, n43419,
    n43420, n43422, n43423, n43424, n43425, n43426, n43428, n43429, n43430,
    n43431, n43432, n43434, n43435, n43436, n43437, n43438, n43440, n43441,
    n43442, n43443, n43444, n43446, n43447, n43448, n43449, n43450, n43452,
    n43453, n43454, n43455, n43456, n43458, n43459, n43460, n43461, n43462,
    n43464, n43465, n43466, n43467, n43468, n43470, n43471, n43472, n43473,
    n43474, n43476, n43477, n43478, n43479, n43480, n43482, n43483, n43484,
    n43485, n43486, n43488, n43489, n43490, n43491, n43492, n43493, n43495,
    n43496, n43497, n43498, n43499, n43501, n43502, n43503, n43504, n43505,
    n43507, n43508, n43509, n43510, n43511, n43513, n43514, n43515, n43516,
    n43517, n43519, n43520, n43521, n43522, n43523, n43525, n43526, n43527,
    n43528, n43529, n43531, n43532, n43533, n43534, n43535, n43537, n43538,
    n43539, n43540, n43541, n43543, n43544, n43545, n43546, n43547, n43549,
    n43550, n43551, n43552, n43553, n43555, n43556, n43557, n43558, n43559,
    n43561, n43562, n43563, n43564, n43565, n43567, n43568, n43569, n43570,
    n43571, n43573, n43574, n43575, n43576, n43577, n43578, n43580, n43581,
    n43582, n43583, n43584, n43586, n43587, n43588, n43589, n43590, n43592,
    n43593, n43594, n43595, n43596, n43598, n43599, n43600, n43601, n43602,
    n43604, n43605, n43606, n43607, n43608, n43610, n43611, n43612, n43613,
    n43614, n43616, n43617, n43618, n43619, n43620, n43622, n43623, n43624,
    n43625, n43626, n43628, n43629, n43630, n43631, n43632, n43634, n43635,
    n43636, n43637, n43638, n43640, n43641, n43642, n43643, n43644, n43646,
    n43647, n43648, n43649, n43650, n43652, n43653, n43654, n43655, n43656,
    n43658, n43659, n43660, n43661, n43662, n43663, n43665, n43666, n43667,
    n43668, n43669, n43671, n43672, n43673, n43674, n43675, n43677, n43678,
    n43679, n43680, n43681, n43683, n43684, n43685, n43686, n43687, n43689,
    n43690, n43691, n43692, n43693, n43695, n43696, n43697, n43698, n43699,
    n43701, n43702, n43703, n43704, n43705, n43707, n43708, n43709, n43710,
    n43711, n43713, n43714, n43715, n43716, n43717, n43719, n43720, n43721,
    n43722, n43723, n43725, n43726, n43727, n43728, n43729, n43731, n43732,
    n43733, n43734, n43735, n43737, n43738, n43739, n43740, n43741, n43743,
    n43744, n43745, n43746, n43747, n43748, n43750, n43751, n43752, n43753,
    n43754, n43756, n43757, n43758, n43759, n43760, n43762, n43763, n43764,
    n43765, n43766, n43768, n43769, n43770, n43771, n43772, n43774, n43775,
    n43776, n43777, n43778, n43780, n43781, n43782, n43783, n43784, n43786,
    n43787, n43788, n43789, n43790, n43792, n43793, n43794, n43795, n43796,
    n43798, n43799, n43800, n43801, n43802, n43804, n43805, n43806, n43807,
    n43808, n43810, n43811, n43812, n43813, n43814, n43816, n43817, n43818,
    n43819, n43820, n43822, n43823, n43824, n43825, n43826, n43828, n43829,
    n43830, n43831, n43832, n43833, n43835, n43836, n43837, n43838, n43839,
    n43841, n43842, n43843, n43844, n43845, n43847, n43848, n43849, n43850,
    n43851, n43853, n43854, n43855, n43856, n43857, n43859, n43860, n43861,
    n43862, n43863, n43865, n43866, n43867, n43868, n43869, n43871, n43872,
    n43873, n43874, n43875, n43877, n43878, n43879, n43880, n43881, n43883,
    n43884, n43885, n43886, n43887, n43889, n43890, n43891, n43892, n43893,
    n43895, n43896, n43897, n43898, n43899, n43901, n43902, n43903, n43904,
    n43905, n43907, n43908, n43909, n43910, n43911, n43913, n43914, n43915,
    n43916, n43917, n43918, n43920, n43921, n43922, n43923, n43924, n43926,
    n43927, n43928, n43929, n43930, n43932, n43933, n43934, n43935, n43936,
    n43938, n43939, n43940, n43941, n43942, n43944, n43945, n43946, n43947,
    n43948, n43950, n43951, n43952, n43953, n43954, n43956, n43957, n43958,
    n43959, n43960, n43962, n43963, n43964, n43965, n43966, n43968, n43969,
    n43970, n43971, n43972, n43974, n43975, n43976, n43977, n43978, n43980,
    n43981, n43982, n43983, n43984, n43986, n43987, n43988, n43989, n43990,
    n43992, n43993, n43994, n43995, n43996, n43998, n43999, n44000, n44001,
    n44002, n44003, n44005, n44006, n44007, n44008, n44009, n44011, n44012,
    n44013, n44014, n44015, n44017, n44018, n44019, n44020, n44021, n44023,
    n44024, n44025, n44026, n44027, n44029, n44030, n44031, n44032, n44033,
    n44035, n44036, n44037, n44038, n44039, n44041, n44042, n44043, n44044,
    n44045, n44047, n44048, n44049, n44050, n44051, n44053, n44054, n44055,
    n44056, n44057, n44059, n44060, n44061, n44062, n44063, n44065, n44066,
    n44067, n44068, n44069, n44071, n44072, n44073, n44074, n44075, n44077,
    n44078, n44079, n44080, n44081, n44083, n44084, n44085, n44086, n44087,
    n44088, n44090, n44091, n44092, n44093, n44094, n44096, n44097, n44098,
    n44099, n44100, n44102, n44103, n44104, n44105, n44106, n44108, n44109,
    n44110, n44111, n44112, n44114, n44115, n44116, n44117, n44118, n44120,
    n44121, n44122, n44123, n44124, n44126, n44127, n44128, n44129, n44130,
    n44132, n44133, n44134, n44135, n44136, n44138, n44139, n44140, n44141,
    n44142, n44144, n44145, n44146, n44147, n44148, n44150, n44151, n44152,
    n44153, n44154, n44156, n44157, n44158, n44159, n44160, n44162, n44163,
    n44164, n44165, n44166, n44168, n44169, n44170, n44171, n44172, n44173,
    n44175, n44176, n44177, n44178, n44179, n44181, n44182, n44183, n44184,
    n44185, n44187, n44188, n44189, n44190, n44191, n44193, n44194, n44195,
    n44196, n44197, n44199, n44200, n44201, n44202, n44203, n44205, n44206,
    n44207, n44208, n44209, n44211, n44212, n44213, n44214, n44215, n44217,
    n44218, n44219, n44220, n44221, n44223, n44224, n44225, n44226, n44227,
    n44229, n44230, n44231, n44232, n44233, n44235, n44236, n44237, n44238,
    n44239, n44241, n44242, n44243, n44244, n44245, n44247, n44248, n44249,
    n44250, n44251, n44253, n44254, n44255, n44256, n44257, n44258, n44259,
    n44260, n44261, n44263, n44264, n44266, n44267, n44269, n44270, n44272,
    n44273, n44275, n44276, n44278, n44279, n44281, n44282, n44284, n44285,
    n44287, n44288, n44290, n44291, n44293, n44294, n44296, n44297, n44299,
    n44300, n44302, n44303, n44305, n44306, n44308, n44309, n44311, n44312,
    n44314, n44315, n44317, n44318, n44320, n44321, n44323, n44324, n44326,
    n44327, n44329, n44330, n44332, n44333, n44335, n44336, n44338, n44339,
    n44341, n44342, n44344, n44345, n44347, n44348, n44350, n44351, n44353,
    n44354, n44355, n44356, n44357, n44359, n44360, n44361, n44362, n44363,
    n44364, n44366, n44367, n44368, n44369, n44370, n44371, n44373, n44374,
    n44375, n44376, n44377, n44378, n44380, n44381, n44382, n44383, n44384,
    n44385, n44386, n44388, n44389, n44390, n44391, n44392, n44393, n44395,
    n44396, n44397, n44398, n44399, n44401, n44402, n44403, n44404, n44405,
    n44407, n44408, n44409, n44410, n44411, n44413, n44414, n44415, n44416,
    n44417, n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426,
    n44427, n44429, n44430, n44431, n44432, n44433, n44435, n44436, n44437,
    n44439, n44440, n44441, n44442, n44443, n44444, n44445, n44446, n44447,
    n44448, n44449, n44450, n44451, n44452, n44453, n44454, n44455, n44456,
    n44457, n44459, n44461, n44462, n44463, n44464, n44465, n44466, n44467,
    n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475, n44476,
    n44477, n44478, n44479, n44480, n44481, n44482, n44483, n44484, n44487,
    n44488, n44489, n44490, n44492, n44493, n44494, n44495, n44496, n44498,
    n44499, n44500, n44501, n44502, n44504, n44505, n44506, n44508, n44509,
    n44510, n44511, n44512, n44513, n44514, n44515, n44516, n44517, n44518,
    n44519, n44520, n44521, n44522, n44523, n44524, n44525, n44526, n44527,
    n44528, n44529, n44530, n44531, n44532, n44533, n44534, n44535, n44536,
    n44537, n44538, n44539, n44540, n44541, n44542, n44543, n44544, n44545,
    n44546, n44547, n44548, n44549, n44550, n44552, n44553, n44554, n44555,
    n44556, n44557, n44558, n44559, n44560, n44561, n44563, n44564, n44565,
    n44566, n44567, n44568, n44569, n44571, n44572, n44573, n44574, n44575,
    n44577, n44578, n44579, n44580, n44581, n44583, n44584, n44585, n44586,
    n44587, n44589, n44590, n44591, n44592, n44593, n44595, n44596, n44597,
    n44598, n44599, n44600, n44602, n44603, n44604, n44605, n44606, n44608,
    n44609, n44610, n44611, n44612, n44613, n44614, n44616, n44617, n44618,
    n44619, n44620, n44622, n44623, n44624, n44625, n44626, n44627, n44629,
    n44630, n44631, n44632, n44633, n44634, n44635, n44637, n44638, n44639,
    n44640, n44641, n44642, n44644, n44645, n44646, n44647, n44648, n44649,
    n44650, n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44660,
    n44661, n44662, n44663, n44664, n44666, n44667, n44668, n44669, n44670,
    n44671, n44673, n44674, n44675, n44676, n44677, n44679, n44680, n44681,
    n44682, n44683, n44685, n44686, n44687, n44688, n44689, n44691, n44692,
    n44693, n44694, n44695, n44697, n44698, n44699, n44700, n44701, n44703,
    n44704, n44705, n44706, n44707, n44709, n44710, n44711, n44712, n44713,
    n44715, n44716, n44717, n44718, n44719, n44721, n44722, n44723, n44724,
    n44725, n44727, n44728, n44729, n44730, n44731, n44733, n44734, n44735,
    n44736, n44737, n44739, n44740, n44741, n44742, n44743, n44744, n44745,
    n44747, n44748, n44749, n44750, n44751, n44753, n44754, n44755, n44756,
    n44757, n44759, n44760, n44761, n44762, n44763, n44765, n44766, n44767,
    n44768, n44769, n44771, n44772, n44773, n44774, n44775, n44777, n44778,
    n44779, n44780, n44781, n44783, n44784, n44785, n44786, n44787, n44789,
    n44790, n44791, n44792, n44793, n44795, n44796, n44797, n44798, n44799,
    n44801, n44802, n44803, n44804, n44805, n44807, n44808, n44809, n44810,
    n44811, n44812, n44813, n44815, n44816, n44817, n44818, n44819, n44821,
    n44822, n44823, n44824, n44825, n44827, n44828, n44829, n44830, n44831,
    n44833, n44834, n44835, n44836, n44837, n44839, n44840, n44841, n44842,
    n44843, n44845, n44847, n44849, n44850, n44851, n44853, n44854, n44855,
    n44857, n44858, n44860, n44861, n44863, n44864, n44866, n44867, n44869,
    n44870, n44872, n44873, n44875, n44876, n44878, n44879, n44881, n44882,
    n44883, n44885, n44886, n44887, n44888, n44890, n44891, n44893, n44894,
    n44896, n44897, n44899, n44900, n44902, n44903, n44905, n44906, n44908,
    n44909, n44911, n44912, n44914, n44915, n44917, n44918, n44920, n44921,
    n44923, n44924, n44925, n44927, n44930, n44931, n44932, n44933, n44934,
    n44935, n44936, n44937, n44938, n44939, n44940, n44941, n44942, n44943,
    n44944, n44946, n44947, n44948, n44950, n44951, n44953, n44954, n44956,
    n44957, n44959, n44960, n44962, n44963, n44965, n44966, n44968, n44969,
    n44971, n44972, n44974, n44975, n44977, n44978, n44980, n44981, n44983,
    n44984, n44985, n44986, n44987, n44988, n44989, n44990, n44991, n44992,
    n44993, n44994, n44995, n44996, n44997, n44998, n44999, n45000, n45001,
    n45002, n45003, n45004, n45005, n45006, n45008, n45009, n45010, n45011,
    n45012, n45014, n45015, n45016, n45017, n45018, n45020, n45021, n45022,
    n45023, n45024, n45025, n45027, n45028, n45029, n45030, n45031, n45033,
    n45034, n45035, n45036, n45037, n45038, n45039, n45040, n45042, n45044,
    n45046, n45048, n45050, n45051, n45052, n45053, n45054, n45055, n45057,
    n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45068,
    n45069, n45070, n45071, n45072, n45074, n45075, n45076, n45077, n45078,
    n45080, n45081, n45082, n45083, n45084, n45086, n45087, n45088, n45089,
    n45090, n45092, n45093, n45094, n45095, n45096, n45098, n45099, n45100,
    n45101, n45102, n45104, n45105, n45106, n45107, n45108, n45110, n45111,
    n45112, n45113, n45114, n45116, n45117, n45118, n45119, n45120, n45122,
    n45123, n45124, n45125, n45126, n45128, n45129, n45130, n45131, n45132,
    n45134, n45135, n45136, n45137, n45138, n45140, n45141, n45142, n45143,
    n45144, n45146, n45147, n45148, n45149, n45150, n45152, n45153, n45154,
    n45155, n45156, n45158, n45159, n45160, n45161, n45162, n45164, n45165,
    n45166, n45167, n45168, n45170, n45171, n45172, n45173, n45174, n45176,
    n45177, n45178, n45179, n45180, n45182, n45183, n45184, n45185, n45186,
    n45188, n45189, n45190, n45191, n45192, n45194, n45195, n45196, n45197,
    n45198, n45200, n45201, n45202, n45203, n45204, n45206, n45207, n45208,
    n45209, n45210, n45212, n45213, n45214, n45215, n45216, n45218, n45219,
    n45220, n45221, n45222, n45224, n45225, n45226, n45227, n45228, n45230,
    n45231, n45232, n45233, n45234, n45236, n45237, n45238, n45239, n45240,
    n45242, n45243, n45244, n45245, n45246, n45248, n45249, n45250, n45251,
    n45252, n45254, n45255, n45256, n45257, n45258, n45260, n45261, n45262,
    n45263, n45264, n45266, n45267, n45268, n45269, n45270, n45272, n45273,
    n45274, n45275, n45276, n45278, n45279, n45280, n45281, n45282, n45284,
    n45285, n45286, n45287, n45288, n45290, n45291, n45292, n45293, n45294,
    n45296, n45297, n45298, n45299, n45300, n45302, n45303, n45304, n45305,
    n45306, n45308, n45309, n45310, n45311, n45312, n45314, n45315, n45316,
    n45317, n45318, n45320, n45321, n45322, n45323, n45324, n45326, n45327,
    n45328, n45329, n45330, n45332, n45333, n45334, n45335, n45336, n45338,
    n45339, n45340, n45341, n45342, n45344, n45345, n45346, n45347, n45348,
    n45350, n45351, n45352, n45353, n45354, n45356, n45357, n45358, n45359,
    n45360, n45362, n45363, n45364, n45365, n45366, n45368, n45369, n45370,
    n45371, n45372, n45374, n45375, n45376, n45377, n45378, n45380, n45381,
    n45382, n45383, n45384, n45386, n45387, n45388, n45389, n45390, n45392,
    n45393, n45394, n45395, n45396, n45398, n45399, n45400, n45401, n45402,
    n45404, n45405, n45406, n45407, n45408, n45410, n45411, n45412, n45413,
    n45414, n45416, n45417, n45418, n45419, n45420, n45422, n45423, n45424,
    n45425, n45426, n45428, n45429, n45430, n45431, n45432, n45434, n45435,
    n45436, n45437, n45438, n45440, n45441, n45442, n45443, n45444, n45446,
    n45447, n45448, n45449, n45450, n45452, n45453, n45454, n45455, n45456,
    n45458, n45459, n45460, n45461, n45462, n45464, n45465, n45466, n45467,
    n45468, n45470, n45471, n45472, n45473, n45474, n45476, n45477, n45478,
    n45479, n45480, n45482, n45483, n45484, n45485, n45486, n45488, n45489,
    n45490, n45491, n45492, n45494, n45495, n45496, n45497, n45498, n45500,
    n45501, n45502, n45503, n45504, n45506, n45507, n45508, n45509, n45510,
    n45512, n45513, n45514, n45515, n45516, n45518, n45519, n45520, n45521,
    n45522, n45524, n45525, n45526, n45527, n45528, n45530, n45531, n45532,
    n45533, n45534, n45536, n45537, n45538, n45539, n45540, n45542, n45543,
    n45544, n45545, n45546, n45548, n45549, n45550, n45551, n45552, n45554,
    n45555, n45556, n45557, n45558, n45560, n45561, n45562, n45563, n45564,
    n45566, n45567, n45568, n45569, n45570, n45572, n45573, n45574, n45575,
    n45576, n45578, n45579, n45580, n45581, n45582, n45584, n45585, n45586,
    n45587, n45588, n45590, n45591, n45592, n45593, n45594, n45596, n45597,
    n45598, n45599, n45600, n45602, n45603, n45604, n45605, n45606, n45608,
    n45609, n45610, n45611, n45612, n45614, n45615, n45616, n45617, n45618,
    n45620, n45621, n45622, n45623, n45624, n45626, n45627, n45628, n45629,
    n45630, n45632, n45633, n45634, n45635, n45636, n45638, n45639, n45640,
    n45641, n45642, n45644, n45645, n45646, n45647, n45648, n45650, n45651,
    n45652, n45653, n45654, n45656, n45657, n45658, n45659, n45660, n45662,
    n45663, n45664, n45665, n45666, n45668, n45669, n45670, n45671, n45672,
    n45674, n45675, n45676, n45677, n45678, n45680, n45681, n45682, n45683,
    n45684, n45686, n45687, n45688, n45689, n45690, n45692, n45693, n45694,
    n45695, n45696, n45698, n45699, n45700, n45701, n45702, n45704, n45705,
    n45706, n45707, n45708, n45710, n45711, n45712, n45713, n45714, n45716,
    n45717, n45718, n45719, n45720, n45722, n45723, n45724, n45725, n45726,
    n45728, n45729, n45730, n45731, n45732, n45734, n45735, n45736, n45737,
    n45738, n45740, n45741, n45742, n45743, n45744, n45746, n45747, n45748,
    n45749, n45750, n45752, n45753, n45754, n45755, n45756, n45758, n45759,
    n45760, n45761, n45762, n45764, n45765, n45766, n45767, n45768, n45770,
    n45771, n45772, n45773, n45774, n45776, n45777, n45778, n45779, n45780,
    n45782, n45783, n45784, n45785, n45786, n45788, n45789, n45790, n45791,
    n45792, n45794, n45795, n45796, n45798, n45799, n45800, n45802, n45803,
    n45804, n45805, n45806, n45807, n45809, n45810, n45812, n45813, n45815,
    n45816, n45817, n45818, n45819, n45820, n45821, n45822, n45823, n45824,
    n45825, n45826, n45827, n45828, n45829, n45830, n45831, n45832, n45833,
    n45834, n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
    n45843, n45844, n45845, n45846, n45848, n45849, n45850, n45851, n45852,
    n45853, n45854, n45855, n45857, n45858, n45859, n45860, n45861, n45862,
    n45863, n45864, n45866, n45867, n45868, n45869, n45870, n45871, n45873,
    n45874, n45875, n45876, n45877, n45879, n45880, n45881, n45882, n45883,
    n45884, n45885, n45886, n45888, n45889, n45890, n45891, n45892, n45893,
    n45894, n45895, n45896, n45897, n45898, n45899, n45901, n45902, n45903,
    n45904, n45905, n45906, n45907, n45908, n45909, n45910, n45911, n45912,
    n45914, n45915, n45917, n45918, n45919, n45920, n45921, n45922, n45923,
    n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931, n45932,
    n45934, n45935, n45936, n45937, n45938, n45940, n45941, n45942, n45943,
    n45944, n45946, n45947, n45948, n45949, n45950, n45952, n45953, n45954,
    n45955, n45956, n45958, n45959, n45960, n45961, n45962, n45964, n45965,
    n45966, n45967, n45968, n45970, n45971, n45972, n45973, n45974, n45976,
    n45977, n45978, n45979, n45980, n45982, n45983, n45984, n45985, n45986,
    n45988, n45989, n45990, n45991, n45992, n45994, n45995, n45996, n45997,
    n45998, n46000, n46001, n46002, n46003, n46004, n46006, n46007, n46008,
    n46009, n46010, n46012, n46013, n46014, n46015, n46016, n46018, n46019,
    n46020, n46021, n46022, n46024, n46025, n46026, n46027, n46028, n46030,
    n46031, n46032, n46033, n46034, n46036, n46037, n46038, n46039, n46040,
    n46042, n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46051,
    n46052, n46053, n46054, n46055, n46056, n46058, n46059, n46060, n46061,
    n46062, n46064, n46065, n46066, n46067, n46068, n46070, n46071, n46072,
    n46073, n46074, n46076, n46077, n46078, n46079, n46080, n46081, n46083,
    n46084, n46085, n46086, n46087, n46089, n46090, n46091, n46092, n46093,
    n46095, n46096, n46097, n46098, n46099, n46101, n46102, n46103, n46104,
    n46105, n46107, n46108, n46109, n46110, n46111, n46113, n46114, n46115,
    n46118, n46119, n46120, n46121, n46123, n46124, n46126, n46127, n46128,
    n46129, n46130, n46131, n46132, n46133, n46134, n46135, n46137, n46138,
    n46139, n46140, n46141, n46144, n46145, n46146, n46148, n46149, n46150,
    n46151, n46152, n46153, n46154, n46155, n46156, n46157, n46159, n46160,
    n46161, n46162, n46163, n46164, n46165, n46167, n46168, n46169, n46170,
    n46171, n46173, n46174, n46175, n46176, n46177, n46179, n46180, n46181,
    n46182, n46183, n46185, n46186, n46187, n46188, n46189, n46191, n46192,
    n46193, n46194, n46195, n46197, n46198, n46199, n46200, n46201, n46203,
    n46204, n46205, n46206, n46207, n46209, n46210, n46211, n46212, n46213,
    n46215, n46216, n46217, n46218, n46219, n46221, n46222, n46223, n46224,
    n46225, n46227, n46228, n46229, n46230, n46231, n46233, n46234, n46235,
    n46236, n46237, n46239, n46240, n46241, n46242, n46243, n46245, n46246,
    n46247, n46248, n46249, n46251, n46252, n46253, n46254, n46255, n46257,
    n46258, n46259, n46260, n46261, n46263, n46264, n46265, n46266, n46268,
    n46269, n46270, n46271, n46273, n46274, n46275, n46276, n46277, n46279,
    n46280, n46281, n46282, n46283, n46284, n46286, n46287, n46289, n46290,
    n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299,
    n46300, n46301, n46302, n46304, n46305, n46306, n46307, n46308, n46309,
    n46310, n46311, n46313, n46314, n46315, n46316, n46317, n46318, n46319,
    n46320, n46321, n46323, n46324, n46325, n46326, n46327, n46328, n46329,
    n46330, n46332, n46333, n46334, n46335, n46336, n46338, n46339, n46340,
    n46341, n46342, n46344, n46345, n46346, n46347, n46348, n46350, n46351,
    n46352, n46353, n46354, n46356, n46357, n46358, n46359, n46360, n46362,
    n46363, n46364, n46365, n46366, n46368, n46369, n46370, n46371, n46372,
    n46373, n46374, n46375, n46377, n46378, n46379, n46380, n46381, n46382,
    n46383, n46384, n46385, n46386, n46387, n46388, n46389, n46391, n46392,
    n46393, n46394, n46395, n46396, n46397, n46398, n46399, n46400, n46402,
    n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46412, n46413,
    n46414, n46415, n46416, n46417, n46418, n46419, n46420, n46421, n46422,
    n46423, n46425, n46426, n46427, n46428, n46429, n46430, n46431, n46432,
    n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443,
    n46445, n46446, n46447, n46448, n46449, n46450, n46452, n46453, n46454,
    n46455, n46457, n46458, n46459, n46461, n46462, n46464, n46465, n46467,
    n46468, n46469, n46470, n46471, n46473, n46474, n46475, n46476, n46477,
    n46479, n46480, n46481, n46482, n46483, n46485, n46486, n46487, n46488,
    n46489, n46490, n46492, n46493, n46494, n46495, n46496, n46498, n46499,
    n46500, n46501, n46502, n46503, n46504, n46505, n46507, n46508, n46509,
    n46510, n46511, n46512, n46513, n46514, n46515, n46517, n46518, n46519,
    n46520, n46521, n46522, n46523, n46524, n46526, n46527, n46528, n46529,
    n46530, n46532, n46533, n46534, n46535, n46536, n46538, n46539, n46540,
    n46541, n46542, n46543, n46545, n46546, n46547, n46548, n46549, n46551,
    n46552, n46553, n46554, n46555, n46557, n46558, n46559, n46560, n46561,
    n46562, n46564, n46565, n46566, n46567, n46568, n46570, n46571, n46572,
    n46573, n46574, n46576, n46577, n46578, n46579, n46580, n46581, n46582,
    n46583, n46584, n46585, n46586, n46587, n46588, n46589, n46590, n46591,
    n46592, n46593, n46595, n46596, n46597, n46598, n46599, n46600, n46602,
    n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611,
    n46612, n46613, n46614, n46616, n46617, n46619, n46620, n46622, n46623,
    n46625, n46626, n46628, n46629, n46631, n46632, n46634, n46635, n46637,
    n46638, n46640, n46641, n46643, n46644, n46646, n46647, n46649, n46650,
    n46651, n46652, n46653, n46654, n46655, n46657, n46658, n46660, n46661,
    n46663, n46664, n46666, n46667, n46669, n46670, n46672, n46673, n46675,
    n46676, n46678, n46679, n46681, n46682, n46684, n46685, n46687, n46688,
    n46690, n46691, n46693, n46694, n46695, n46697, n46698, n46699, n46700,
    n46702, n46703, n46704, n46705, n46707, n46708, n46709, n46710, n46712,
    n46713, n46714, n46715, n46717, n46718, n46719, n46720, n46722, n46723,
    n46725, n46726, n46727, n46728, n46729, n46730, n46731, n46732, n46733,
    n46734, n46735, n46736, n46737, n46739, n46740, n46741, n46743, n46744,
    n46745, n46747, n46748, n46750, n46751, n46753, n46754, n46756, n46757,
    n46759, n46760, n46762, n46763, n46765, n46766, n46768, n46769, n46771,
    n46772, n46774, n46775, n46777, n46778, n46780, n46781, n46782, n46784,
    n46785, n46787, n46788, n46790, n46791, n46793, n46794, n46796, n46797,
    n46799, n46800, n46802, n46803, n46805, n46806, n46808, n46809, n46810,
    n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
    n46821, n46822, n46823, n46825, n46826, n46827, n46828, n46829, n46831,
    n46832, n46834, n46835, n46837, n46838, n46840, n46841, n46843, n46844,
    n46846, n46847, n46849, n46850, n46852, n46853, n46855, n46856, n46858,
    n46859, n46861, n46862, n46864, n46865, n46867, n46868, n46870, n46871,
    n46873, n46874, n46875, n46876, n46877, n46878, n46880, n46881, n46882,
    n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891,
    n46893, n46895, n46896, n46897, n46898, n46899, n46900, n46901, n46902,
    n46904, n46905, n46906, n46907, n46908, n46909, n46910, n46911, n46913,
    n46914, n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923,
    n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931, n46932,
    n46934, n46935, n46936, n46937, n46938, n46939, n46940, n46942, n46943,
    n46944, n46945, n46946, n46947, n46948, n46949, n46950, n46952, n46953,
    n46954, n46955, n46956, n46958, n46959, n46960, n46961, n46962, n46963,
    n46964, n46965, n46966, n46967, n46969, n46970, n46972, n46973, n46974,
    n46975, n46976, n46977, n46979, n46980, n46981, n46982, n46983, n46984,
    n46986, n46987, n46988, n46989, n46990, n46992, n46993, n46994, n46995,
    n46996, n46998, n46999, n47000, n47001, n47002, n47004, n47005, n47006,
    n47007, n47008, n47010, n47011, n47012, n47013, n47014, n47016, n47017,
    n47018, n47019, n47020, n47022, n47023, n47024, n47025, n47026, n47028,
    n47029, n47030, n47031, n47032, n47034, n47035, n47036, n47037, n47038,
    n47040, n47041, n47042, n47043, n47044, n47046, n47047, n47048, n47049,
    n47050, n47052, n47053, n47054, n47055, n47056, n47058, n47059, n47060,
    n47061, n47062, n47064, n47065, n47066, n47067, n47068, n47070, n47071,
    n47072, n47073, n47074, n47076, n47077, n47078, n47079, n47080, n47082,
    n47083, n47084, n47085, n47086, n47088, n47089, n47090, n47091, n47092,
    n47094, n47095, n47096, n47097, n47098, n47100, n47101, n47102, n47103,
    n47104, n47106, n47107, n47108, n47109, n47110, n47112, n47113, n47114,
    n47115, n47116, n47118, n47119, n47120, n47122, n47123, n47124, n47125,
    n47126, n47127, n47128, n47129, n47130, n47131, n47132, n47133, n47134,
    n47135, n47136, n47137, n47139, n47140, n47141, n47142, n47144, n47145,
    n47146, n47148, n47149, n47150, n47152, n47153, n47155, n47156, n47158,
    n47159, n47161, n47162, n47164, n47165, n47167, n47168, n47170, n47171,
    n47173, n47174, n47176, n47177, n47179, n47180, n47182, n47183, n47185,
    n47186, n47188, n47189, n47190, n47191, n47192, n47193, n47195, n47196,
    n47197, n47198, n47199, n47200, n47201, n47202, n47204, n47205, n47206,
    n47207, n47208, n47209, n47210, n47211, n47212, n47213, n47215, n47216,
    n47217, n47218, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
    n47227, n47228, n47229, n47231, n47232, n47233, n47234, n47236, n47237,
    n47238, n47239, n47240, n47241, n47242, n47244, n47245, n47246, n47247,
    n47248, n47250, n47251, n47252, n47253, n47254, n47256, n47257, n47258,
    n47259, n47260, n47261, n47262, n47264, n47265, n47266, n47268, n47269,
    n47270, n47271, n47272, n47274, n47275, n47277, n47278, n47280, n47281,
    n47283, n47284, n47285, n47286, n47287, n47289, n47290, n47291, n47292,
    n47293, n47295, n47296, n47298, n47299, n47301, n47302, n47303, n47304,
    n47305, n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315,
    n47316, n47317, n47318, n47319, n47321, n47322, n47323, n47325, n47326,
    n47327, n47329, n47330, n47332, n47333, n47334, n47335, n47336, n47338,
    n47339, n47340, n47341, n47342, n47344, n47345, n47346, n47348, n47349,
    n47350, n47352, n47353, n47355, n47356, n47358, n47359, n47360, n47362,
    n47363, n47365, n47366, n47367, n47369, n47370, n47372, n47373, n47375,
    n47376, n47379, n47380, n47382, n47383, n47385, n47386, n47388, n47389,
    n47391, n47392, n47393, n47395, n47396, n47397, n47401, n47402, n47404,
    n47405, n47407, n47408, n47410, n47411, n47413, n47414, n47416, n47417,
    n47419, n47420, n47422, n47423, n47425, n47426, n47428, n47429, n47431,
    n47432, n47433, n47435, n47436, n47438, n47439, n47442, n47443, n47444,
    n47446, n47447, n47448, n47450, n47451, n47453, n47454, n47456, n47457,
    n47459, n47460, n47462, n47463, n47465, n47466, n47468, n47469, n47471,
    n47472, n47474, n47475, n47477, n47478, n47480, n47481, n47483, n47484,
    n47485, n47487, n47488, n47490, n47491, n47493, n47494, n47496, n47497,
    n47499, n47500, n47501, n47503, n47504, n47505, n47507, n47508, n47510,
    n47511, n47512, n47514, n47515, n47517, n47518, n47520, n47521, n47523,
    n47524, n47526, n47527, n47529, n47530, n47532, n47533, n47535, n47536,
    n47538, n47539, n47541, n47542, n47544, n47545, n47547, n47548, n47550,
    n47551, n47553, n47554, n47556, n47557, n47559, n47560, n47561, n47562,
    n47563, n47564, n47566, n47567, n47568, n47569, n47570, n47571, n47572,
    n47573, n47574, n47576, n47577, n47578, n47579, n47580, n47582, n47583,
    n47584, n47585, n47586, n47587, n47588, n47589, n47591, n47592, n47593,
    n47594, n47596, n47597, n47599, n47600, n47602, n47603, n47605, n47606,
    n47608, n47609, n47611, n47612, n47614, n47615, n47617, n47618, n47619,
    n47620, n47621, n47622, n47624, n47625, n47627, n47628, n47630, n47631,
    n47633, n47634, n47636, n47637, n47639, n47640, n47642, n47643, n47644,
    n47645, n47647, n47648, n47650, n47651, n47652, n47653, n47654, n47655,
    n47656, n47657, n47659, n47660, n47661, n47662, n47663, n47664, n47665,
    n47666, n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675,
    n47677, n47678, n47679, n47680, n47681, n47682, n47683, n47684, n47686,
    n47687, n47688, n47689, n47690, n47691, n47692, n47693, n47695, n47696,
    n47697, n47698, n47699, n47700, n47701, n47702, n47704, n47705, n47706,
    n47707, n47708, n47709, n47710, n47711, n47713, n47714, n47715, n47716,
    n47717, n47718, n47719, n47720, n47722, n47723, n47724, n47725, n47726,
    n47727, n47728, n47729, n47731, n47732, n47733, n47734, n47735, n47736,
    n47737, n47738, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
    n47747, n47749, n47750, n47751, n47752, n47753, n47754, n47755, n47756,
    n47758, n47759, n47760, n47761, n47762, n47763, n47764, n47765, n47767,
    n47768, n47770, n47771, n47773, n47774, n47776, n47777, n47778, n47779,
    n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787, n47788,
    n47789, n47791, n47792, n47794, n47795, n47797, n47798, n47800, n47801,
    n47803, n47804, n47805, n47806, n47807, n47808, n47810, n47811, n47813,
    n47814, n47816, n47817, n47819, n47820, n47822, n47823, n47825, n47826,
    n47828, n47829, n47831, n47832, n47834, n47835, n47837, n47838, n47839,
    n47840, n47841, n47843, n47844, n47845, n47846, n47847, n47849, n47850,
    n47851, n47852, n47853, n47855, n47856, n47857, n47858, n47859, n47861,
    n47862, n47863, n47864, n47865, n47867, n47868, n47869, n47870, n47871,
    n47873, n47874, n47875, n47876, n47877, n47879, n47880, n47881, n47882,
    n47883, n47885, n47886, n47887, n47888, n47889, n47891, n47892, n47893,
    n47894, n47895, n47897, n47898, n47899, n47900, n47901, n47902, n47904,
    n47905, n47906, n47907, n47908, n47910, n47911, n47912, n47913, n47914,
    n47916, n47917, n47918, n47919, n47920, n47922, n47923, n47924, n47925,
    n47926, n47928, n47929, n47930, n47931, n47932, n47934, n47935, n47936,
    n47937, n47938, n47940, n47941, n47942, n47943, n47944, n47946, n47947,
    n47948, n47949, n47950, n47952, n47953, n47954, n47955, n47956, n47958,
    n47959, n47960, n47961, n47962, n47964, n47965, n47966, n47967, n47968,
    n47970, n47971, n47972, n47973, n47974, n47975, n47977, n47978, n47979,
    n47980, n47981, n47983, n47984, n47985, n47986, n47987, n47988, n47989,
    n47990, n47991, n47992, n47993, n47994, n47995, n47997, n47998, n47999,
    n48000, n48001, n48002, n48003, n48004, n48005, n48006, n48007, n48008,
    n48009, n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
    n48019, n48020, n48021, n48022, n48023, n48025, n48026, n48027, n48028,
    n48029, n48030, n48031, n48032, n48033, n48034, n48035, n48036, n48037,
    n48039, n48040, n48041, n48042, n48043, n48044, n48045, n48046, n48047,
    n48048, n48049, n48050, n48051, n48053, n48054, n48055, n48056, n48057,
    n48058, n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48067,
    n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075, n48076,
    n48077, n48078, n48079, n48081, n48082, n48083, n48085, n48086, n48087,
    n48088, n48090, n48091, n48092, n48093, n48094, n48096, n48097, n48098,
    n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107, n48108,
    n48110, n48111, n48113, n48114, n48116, n48117, n48119, n48120, n48122,
    n48123, n48125, n48126, n48128, n48129, n48131, n48132, n48134, n48135,
    n48137, n48138, n48140, n48141, n48143, n48144, n48146, n48147, n48149,
    n48150, n48152, n48153, n48155, n48156, n48158, n48159, n48161, n48162,
    n48164, n48165, n48167, n48168, n48170, n48171, n48173, n48174, n48176,
    n48177, n48179, n48180, n48182, n48183, n48185, n48186, n48188, n48189,
    n48190, n48192, n48193, n48194, n48195, n48196, n48197, n48198, n48199,
    n48200, n48201, n48203, n48204, n48206, n48207, n48209, n48210, n48212,
    n48213, n48215, n48216, n48218, n48219, n48221, n48222, n48223, n48224,
    n48225, n48226, n48227, n48229, n48230, n48232, n48233, n48234, n48235,
    n48236, n48237, n48238, n48240, n48241, n48242, n48243, n48244, n48245,
    n48246, n48248, n48249, n48251, n48252, n48253, n48254, n48255, n48256,
    n48257, n48258, n48259, n48261, n48262, n48264, n48265, n48267, n48268,
    n48270, n48271, n48273, n48274, n48276, n48277, n48278, n48279, n48281,
    n48282, n48283, n48284, n48286, n48287, n48288, n48289, n48290, n48292,
    n48293, n48294, n48295, n48296, n48298, n48299, n48300, n48301, n48302,
    n48304, n48305, n48306, n48307, n48308, n48310, n48311, n48312, n48313,
    n48314, n48316, n48317, n48318, n48319, n48320, n48322, n48323, n48324,
    n48325, n48326, n48328, n48329, n48330, n48331, n48332, n48334, n48335,
    n48336, n48337, n48338, n48340, n48341, n48343, n48344, n48345, n48346,
    n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355,
    n48356, n48358, n48359, n48360, n48361, n48362, n48363, n48364, n48365,
    n48366, n48367, n48368, n48369, n48371, n48372, n48373, n48374, n48375,
    n48376, n48377, n48378, n48380, n48381, n48382, n48383, n48384, n48385,
    n48386, n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
    n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403,
    n48404, n48405, n48406, n48407, n48408, n48409, n48411, n48412, n48413,
    n48414, n48415, n48416, n48417, n48418, n48419, n48420, n48422, n48423,
    n48424, n48425, n48427, n48428, n48429, n48430, n48432, n48433, n48434,
    n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48443, n48444,
    n48446, n48447, n48449, n48450, n48452, n48453, n48455, n48456, n48458,
    n48459, n48461, n48462, n48464, n48465, n48467, n48468, n48470, n48471,
    n48473, n48474, n48476, n48477, n48482, n48483, n48484, n48485, n48486,
    n48487, n48488, n48489, n48490, n48492, n48493, n48494, n48495, n48496,
    n48497, n48498, n48499, n48501, n48502, n48503, n48504, n48505, n48506,
    n48507, n48508, n48510, n48511, n48512, n48513, n48514, n48515, n48516,
    n48517, n48519, n48520, n48521, n48522, n48523, n48524, n48525, n48526,
    n48528, n48529, n48530, n48531, n48532, n48533, n48534, n48535, n48537,
    n48538, n48539, n48540, n48541, n48542, n48543, n48544, n48546, n48547,
    n48548, n48549, n48550, n48551, n48552, n48553, n48555, n48556, n48557,
    n48558, n48559, n48560, n48561, n48562, n48564, n48565, n48566, n48567,
    n48568, n48569, n48570, n48571, n48573, n48574, n48576, n48578, n48579,
    n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587, n48588,
    n48590, n48591, n48592, n48593, n48594, n48595, n48596, n48597, n48598,
    n48599, n48600, n48601, n48602, n48603, n48605, n48606, n48608, n48609,
    n48611, n48612, n48614, n48615, n48617, n48618, n48620, n48621, n48623,
    n48624, n48626, n48627, n48629, n48630, n48631, n48632, n48633, n48634,
    n48635, n48636, n48638, n48639, n48640, n48641, n48643, n48644, n48646,
    n48647, n48649, n48650, n48652, n48653, n48655, n48656, n48658, n48659,
    n48661, n48662, n48664, n48665, n48667, n48668, n48670, n48671, n48673,
    n48674, n48676, n48677, n48679, n48680, n48682, n48683, n48685, n48686,
    n48688, n48689, n48690, n48692, n48693, n48694, n48695, n48696, n48697,
    n48698, n48699, n48701, n48702, n48704, n48706, n48708, n48709, n48711,
    n48712, n48714, n48715, n48717, n48718, n48720, n48721, n48723, n48724,
    n48726, n48727, n48729, n48730, n48732, n48733, n48735, n48736, n48738,
    n48739, n48741, n48742, n48744, n48745, n48747, n48748, n48750, n48751,
    n48753, n48754, n48756, n48757, n48759, n48760, n48761, n48762, n48764,
    n48765, n48767, n48768, n48770, n48771, n48773, n48774, n48776, n48777,
    n48779, n48780, n48782, n48783, n48785, n48786, n48788, n48789, n48791,
    n48792, n48794, n48795, n48797, n48798, n48800, n48801, n48803, n48804,
    n48806, n48807, n48809, n48810, n48811, n48812, n48814, n48815, n48817,
    n48818, n48820, n48821, n48823, n48824, n48826, n48827, n48829, n48830,
    n48832, n48833, n48835, n48836, n48838, n48839, n48841, n48842, n48844,
    n48845, n48847, n48848, n48850, n48851, n48853, n48854, n48856, n48857,
    n48859, n48860, n48861, n48862, n48863, n48865, n48866, n48867, n48868,
    n48869, n48871, n48872, n48873, n48874, n48875, n48876, n48877, n48878,
    n48879, n48880, n48882, n48883, n48884, n48885, n48886, n48888, n48889,
    n48890, n48891, n48892, n48894, n48895, n48896, n48897, n48898, n48899,
    n48900, n48901, n48902, n48904, n48905, n48906, n48907, n48908, n48910,
    n48911, n48912, n48913, n48914, n48915, n48917, n48918, n48919, n48920,
    n48922, n48923, n48925, n48926, n48928, n48929, n48931, n48932, n48934,
    n48935, n48937, n48938, n48940, n48941, n48943, n48944, n48946, n48947,
    n48949, n48950, n48952, n48953, n48955, n48956, n48958, n48959, n48961,
    n48962, n48963, n48964, n48966, n48967, n48969, n48970, n48972, n48973,
    n48975, n48976, n48978, n48979, n48981, n48982, n48984, n48985, n48987,
    n48988, n48990, n48991, n48993, n48994, n48996, n48997, n48999, n49000,
    n49002, n49003, n49005, n49006, n49007, n49008, n49010, n49011, n49013,
    n49014, n49016, n49017, n49019, n49020, n49022, n49023, n49025, n49026,
    n49028, n49029, n49031, n49032, n49034, n49035, n49037, n49038, n49040,
    n49041, n49043, n49044, n49046, n49047, n49049, n49050, n49051, n49052,
    n49054, n49055, n49057, n49058, n49060, n49061, n49063, n49064, n49066,
    n49067, n49069, n49070, n49072, n49073, n49075, n49076, n49078, n49079,
    n49081, n49082, n49084, n49085, n49087, n49088, n49090, n49091, n49093,
    n49094, n49095, n49096, n49097, n49098, n49100, n49101, n49103, n49104,
    n49106, n49107, n49109, n49110, n49111, n49112, n49113, n49114, n49116,
    n49117, n49119, n49120, n49122, n49123, n49125, n49126, n49128, n49129,
    n49131, n49132, n49134, n49135, n49137, n49138, n49140, n49141, n49143,
    n49144, n49145, n49146, n49147, n49148, n49150, n49151, n49153, n49154,
    n49156, n49157, n49159, n49160, n49162, n49163, n49165, n49166, n49168,
    n49169, n49171, n49172, n49174, n49175, n49177, n49178, n49180, n49181,
    n49183, n49184, n49186, n49187, n49189, n49190, n49192, n49193, n49195,
    n49196, n49198, n49199, n49201, n49202, n49204, n49205, n49207, n49208,
    n49210, n49211, n49213, n49214, n49216, n49217, n49219, n49220, n49222,
    n49223, n49225, n49226, n49228, n49229, n49231, n49232, n49234, n49235,
    n49237, n49238, n49240, n49241, n49243, n49244, n49246, n49247, n49249,
    n49250, n49252, n49253, n49255, n49256, n49258, n49259, n49261, n49262,
    n49264, n49265, n49267, n49268, n49270, n49271, n49273, n49274, n49276,
    n49277, n49278, n49279, n49281, n49282, n49284, n49285, n49287, n49288,
    n49290, n49291, n49293, n49294, n49296, n49297, n49299, n49300, n49302,
    n49303, n49305, n49306, n49308, n49309, n49311, n49312, n49314, n49315,
    n49317, n49318, n49320, n49321, n49322, n49323, n49324, n49326, n49327,
    n49328, n49329, n49330, n49332, n49333, n49334, n49335, n49336, n49338,
    n49339, n49340, n49341, n49342, n49344, n49345, n49346, n49347, n49348,
    n49350, n49351, n49352, n49353, n49354, n49356, n49357, n49358, n49359,
    n49360, n49362, n49363, n49364, n49365, n49366, n49368, n49369, n49370,
    n49371, n49372, n49374, n49375, n49376, n49377, n49378, n49380, n49381,
    n49382, n49383, n49384, n49386, n49387, n49388, n49389, n49390, n49392,
    n49393, n49394, n49395, n49396, n49398, n49399, n49400, n49401, n49402,
    n49404, n49405, n49406, n49407, n49408, n49410, n49411, n49412, n49413,
    n49414, n49416, n49417, n49418, n49419, n49420, n49422, n49423, n49424,
    n49425, n49426, n49428, n49429, n49430, n49431, n49432, n49434, n49435,
    n49436, n49437, n49438, n49440, n49441, n49442, n49443, n49444, n49446,
    n49447, n49448, n49449, n49450, n49452, n49453, n49454, n49455, n49456,
    n49458, n49459, n49460, n49461, n49462, n49464, n49465, n49466, n49467,
    n49468, n49470, n49471, n49472, n49473, n49474, n49476, n49477, n49478,
    n49479, n49480, n49482, n49483, n49484, n49485, n49486, n49488, n49489,
    n49490, n49491, n49492, n49494, n49495, n49496, n49497, n49498, n49500,
    n49501, n49502, n49503, n49504, n49506, n49507, n49508, n49509, n49510,
    n49512, n49513, n49514, n49515, n49516, n49518, n49519, n49520, n49521,
    n49522, n49524, n49525, n49526, n49527, n49528, n49530, n49531, n49532,
    n49533, n49534, n49536, n49537, n49538, n49539, n49540, n49542, n49543,
    n49544, n49545, n49546, n49548, n49549, n49550, n49551, n49552, n49554,
    n49555, n49556, n49557, n49558, n49560, n49561, n49562, n49563, n49564,
    n49566, n49567, n49568, n49569, n49570, n49572, n49573, n49574, n49575,
    n49576, n49578, n49579, n49580, n49581, n49582, n49584, n49585, n49586,
    n49587, n49588, n49590, n49591, n49592, n49593, n49594, n49595, n49596,
    n49597, n49598, n49599, n49600, n49601, n49602, n49604, n49605, n49606,
    n49607, n49608, n49609, n49610, n49611, n49612, n49613, n49614, n49615,
    n49616, n49618, n49619, n49620, n49621, n49622, n49624, n49625, n49626,
    n49627, n49628, n49630, n49631, n49632, n49633, n49634, n49635, n49636,
    n49637, n49638, n49639, n49640, n49641, n49642, n49644, n49645, n49646,
    n49647, n49648, n49649, n49650, n49651, n49652, n49653, n49654, n49655,
    n49656, n49658, n49659, n49660, n49662, n49663, n49664, n49665, n49666,
    n49667, n49668, n49669, n49670, n49672, n49673, n49674, n49675, n49676,
    n49677, n49678, n49679, n49680, n49681, n49682, n49683, n49685, n49686,
    n49687, n49688, n49689, n49690, n49691, n49693, n49694, n49695, n49696,
    n49697, n49699, n49700, n49702, n49703, n49704, n49705, n49706, n49708,
    n49709, n49710, n49713, n49714, n49715, n49716, n49717, n49718, n49719,
    n49720, n49721, n49722, n49723, n49724, n49725, n49726, n49727, n49728,
    n49729, n49730, n49731, n49732, n49733, n49734, n49735, n49736, n49737,
    n49738, n49739, n49740, n49741, n49743, n49744, n49745, n49746, n49747,
    n49749, n49750, n49751, n49752, n49753, n49755, n49756, n49757, n49758,
    n49759, n49761, n49762, n49763, n49764, n49765, n49767, n49768, n49769,
    n49770, n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
    n49779, n49781, n49782, n49784, n49785, n49787, n49788, n49790, n49791,
    n49793, n49794, n49796, n49797, n49799, n49800, n49801, n49802, n49803,
    n49804, n49805, n49807, n49808, n49809, n49810, n49811, n49812, n49813,
    n49814, n49815, n49816, n49817, n49818, n49820, n49821, n49822, n49823,
    n49825, n49826, n49827, n49828, n49829, n49830, n49831, n49832, n49833,
    n49834, n49835, n49836, n49838, n49839, n49840, n49841, n49842, n49843,
    n49845, n49846, n49848, n49849, n49850, n49851, n49852, n49854, n49855,
    n49856, n49857, n49858, n49860, n49861, n49863, n49864, n49866, n49867,
    n49868, n49869, n49870, n49871, n49873, n49874, n49876, n49877, n49879,
    n49880, n49882, n49883, n49885, n49886, n49887, n49888, n49889, n49890,
    n49891, n49892, n49893, n49895, n49896, n49897, n49898, n49899, n49900,
    n49902, n49903, n49905, n49906, n49908, n49909, n49911, n49912, n49914,
    n49915, n49917, n49918, n49920, n49921, n49923, n49924, n49926, n49927,
    n49929, n49930, n49932, n49933, n49935, n49936, n49938, n49939, n49941,
    n49942, n49944, n49945, n49947, n49948, n49950, n49951, n49953, n49954,
    n49956, n49957, n49959, n49960, n49962, n49963, n49965, n49966, n49968,
    n49969, n49971, n49972, n49974, n49975, n49977, n49978, n49980, n49981,
    n49983, n49984, n49986, n49987, n49989, n49990, n49992, n49993, n49995,
    n49996, n49997, n49998, n49999, n50001, n50002, n50003, n50004, n50005,
    n50007, n50008, n50009, n50010, n50011, n50013, n50014, n50015, n50016,
    n50017, n50019, n50020, n50021, n50022, n50023, n50024, n50026, n50027,
    n50029, n50030, n50032, n50033, n50035, n50036, n50038, n50039, n50041,
    n50042, n50044, n50045, n50047, n50048, n50050, n50051, n50053, n50054,
    n50056, n50057, n50059, n50060, n50062, n50063, n50065, n50066, n50068,
    n50069, n50071, n50072, n50074, n50075, n50077, n50078, n50080, n50081,
    n50082, n50083, n50084, n50086, n50087, n50089, n50090, n50092, n50093,
    n50095, n50096, n50098, n50099, n50101, n50102, n50104, n50105, n50107,
    n50108, n50110, n50111, n50113, n50114, n50116, n50117, n50119, n50120,
    n50122, n50123, n50125, n50126, n50128, n50129, n50130, n50132, n50133,
    n50135, n50136, n50137, n50139, n50140, n50141, n50142, n50143, n50144,
    n50145, n50147, n50148, n50149, n50150, n50151, n50152, n50154, n50155,
    n50156, n50157, n50158, n50159, n50161, n50162, n50163, n50166, n50167,
    n50168, n50170, n50171, n50172, n50174, n50175, n50177, n50178, n50180,
    n50181, n50183, n50184, n50186, n50187, n50189, n50190, n50192, n50193,
    n50195, n50196, n50198, n50199, n50201, n50202, n50203, n50204, n50205,
    n50206, n50207, n50208, n50210, n50211, n50212, n50214, n50215, n50216,
    n50218, n50219, n50220, n50221, n50223, n50224, n50225, n50226, n50227,
    n50228, n50230, n50231, n50232, n50233, n50234, n50236, n50237, n50239,
    n50240, n50242, n50243, n50245, n50246, n50248, n50250, n50251, n50253,
    n50254, n50256, n50257, n50259, n50260, n50261, n50262, n50263, n50265,
    n50266, n50268, n50269, n50270, n50273, n50274, n50276, n50277, n50279,
    n50280, n50282, n50283, n50285, n50286, n50287, n50288, n50290, n50291,
    n50292, n50293, n50295, n50296, n50297, n50298, n50299, n50300, n50302,
    n50303, n50305, n50306, n50307, n50308, n50310, n50311, n50312, n50313,
    n50314, n50315, n50317, n50318, n50320, n50321, n50323, n50324, n50326,
    n50327, n50328, n50330, n50331, n50333, n50334, n50336, n50337, n50339,
    n50340, n50342, n50343, n50344, n50345, n50347, n50348, n50350, n50351,
    n50353, n50354, n50356, n50357, n50359, n50360, n50362, n50363, n50365,
    n50366, n50368, n50369, n50370, n50371, n50373, n50374, n50376, n50377,
    n50378, n50379, n50381, n50382, n50384, n50385, n50386, n50387, n50388,
    n50391, n50392, n50393, n50394, n50395, n50397, n50398, n50399, n50400,
    n50401, n50403, n50404, n50405, n50406, n50407, n50409, n50410, n50411,
    n50412, n50413, n50415, n50416, n50418, n50419, n50421, n50422, n50423,
    n50424, n50426, n50427, n50429, n50430, n50432, n50433, n50435, n50436,
    n50437, n50438, n50440, n50441, n50443, n50444, n50446, n50447, n50449,
    n50450, n50452, n50453, n50455, n50456, n50458, n50459, n50461, n50462,
    n50464, n50465, n50467, n50468, n50470, n50471, n50473, n50474, n50476,
    n50477, n50479, n50480, n50482, n50483, n50484, n50485, n50486, n50487,
    n50488, n50489, n50491, n50492, n50493, n50494, n50495, n50497, n50498,
    n50499, n50500, n50501, n50503, n50504, n50505, n50506, n50507, n50509,
    n50510, n50511, n50512, n50513, n50515, n50516, n50517, n50518, n50519,
    n50521, n50522, n50523, n50524, n50525, n50527, n50528, n50529, n50530,
    n50531, n50533, n50534, n50535, n50536, n50537, n50539, n50540, n50541,
    n50542, n50543, n50545, n50546, n50547, n50548, n50549, n50551, n50552,
    n50553, n50554, n50555, n50557, n50558, n50559, n50560, n50561, n50563,
    n50564, n50565, n50566, n50567, n50569, n50570, n50571, n50572, n50573,
    n50576, n50577, n50579, n50580, n50581, n50582, n50583, n50584, n50585,
    n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50596, n50597,
    n50599, n50600, n50601, n50602, n50605, n50606, n50608, n50609, n50610,
    n50612, n50613, n50615, n50616, n50618, n50619, n50621, n50622, n50624,
    n50625, n50627, n50628, n50629, n50631, n50632, n50634, n50635, n50637,
    n50638, n50640, n50641, n50643, n50644, n50646, n50647, n50649, n50650,
    n50651, n50653, n50654, n50656, n50657, n50659, n50660, n50662, n50663,
    n50665, n50666, n50668, n50669, n50670, n50672, n50673, n50675, n50676,
    n50678, n50679, n50681, n50682, n50684, n50685, n50687, n50688, n50690,
    n50691, n50693, n50694, n50696, n50697, n50699, n50700, n50702, n50703,
    n50705, n50706, n50708, n50709, n50711, n50712, n50714, n50715, n50717,
    n50718, n50720, n50721, n50723, n50724, n50726, n50727, n50728, n50730,
    n50731, n50733, n50734, n50736, n50737, n50739, n50740, n50742, n50743,
    n50745, n50746, n50748, n50749, n50751, n50752, n50754, n50755, n50757,
    n50758, n50760, n50761, n50763, n50764, n50766, n50767, n50769, n50770,
    n50772, n50773, n50775, n50776, n50778, n50779, n50781, n50782, n50783,
    n50784, n50786, n50787, n50789, n50790, n50792, n50793, n50795, n50796,
    n50798, n50799, n50801, n50802, n50804, n50805, n50807, n50808, n50810,
    n50811, n50813, n50814, n50816, n50817, n50819, n50820, n50822, n50823,
    n50825, n50826, n50828, n50829, n50831, n50832, n50834, n50835, n50837,
    n50838, n50840, n50841, n50843, n50844, n50846, n50847, n50849, n50850,
    n50852, n50853, n50855, n50856, n50858, n50859, n50861, n50862, n50864,
    n50865, n50867, n50868, n50870, n50871, n50873, n50874, n50876, n50877,
    n50879, n50880, n50882, n50883, n50885, n50886, n50888, n50889, n50891,
    n50892, n50894, n50895, n50897, n50898, n50900, n50901, n50903, n50904,
    n50906, n50907, n50909, n50910, n50912, n50913, n50914, n50915, n50916,
    n50918, n50919, n50920, n50921, n50922, n50924, n50925, n50926, n50927,
    n50928, n50930, n50931, n50932, n50933, n50934, n50936, n50937, n50939,
    n50940, n50942, n50943, n50945, n50946, n50948, n50949, n50951, n50952,
    n50954, n50955, n50957, n50958, n50960, n50961, n50963, n50964, n50966,
    n50967, n50969, n50970, n50972, n50973, n50975, n50976, n50978, n50979,
    n50981, n50982, n50984, n50985, n50987, n50988, n50990, n50991, n50993,
    n50994, n50996, n50997, n50999, n51000, n51002, n51003, n51005, n51006,
    n51008, n51009, n51011, n51012, n51014, n51015, n51017, n51018, n51020,
    n51021, n51023, n51024, n51026, n51027, n51029, n51030, n51032, n51033,
    n51035, n51036, n51038, n51039, n51041, n51042, n51044, n51045, n51047,
    n51048, n51050, n51051, n51053, n51054, n51056, n51057, n51059, n51060,
    n51062, n51063, n51065, n51066, n51068, n51069, n51071, n51072, n51074,
    n51075, n51077, n51078, n51080, n51081, n51083, n51084, n51085, n51086,
    n51087, n51089, n51090, n51092, n51093, n51094, n51095, n51096, n51097,
    n51098, n51100, n51101, n51102, n51104, n51105, n51107, n51108, n51110,
    n51111, n51113, n51114, n51115, n51116, n51117, n51119, n51121, n51122,
    n51123, n51124, n51126, n51127, n51129, n51131, n51132, n51133, n51134,
    n51135, n51136, n51138, n51139, n51140, n51142, n51143, n51144, n51145,
    n51147, n51148, n51150, n51151, n51153, n51154, n51155, n51157, n51158,
    n51160, n51161, n51162, n51164, n51165, n51166, n51167, n51169, n51170,
    n51171, n51172, n51174, n51175, n51177, n51178, n51180, n51181, n51183,
    n51184, n51185, n51186, n51188, n51189, n51191, n51192, n51193, n51194,
    n51196, n51197, n51198, n51200, n51201, n51203, n51204, n51206, n51207,
    n51209, n51210, n51211, n51213, n51214, n51215, n51217, n51218, n51219,
    n51221, n51222, n51223, n51224, n51226, n51227, n51229, n51230, n51232,
    n51233, n51235, n51236, n51238, n51239, n51240, n51242, n51243, n51244,
    n51245, n51246, n51248, n51250, n51251, n51253, n51254, n51256, n51257,
    n51259, n51260, n51262, n51263, n51265, n51266, n51268, n51269, n51271,
    n51272, n51274, n51275, n51277, n51278, n51280, n51281, n51283, n51284,
    n51285, n51287, n51288, n51289, n51290, n51291, n51292, n51293, n51294,
    n51295, n51296, n51298, n51299, n51301, n51302, n51303, n51304, n51305,
    n51306, n51307, n51309, n51310, n51312, n51313, n51315, n51316, n51318,
    n51319, n51321, n51322, n51323, n51325, n51326, n51328, n51329, n51331,
    n51332, n51333, n51334, n51335, n51337, n51338, n51339, n51340, n51341,
    n51342, n51344, n51345, n51347, n51348, n51350, n51351, n51353, n51354,
    n51356, n51357, n51359, n51360, n51362, n51363, n51365, n51366, n51368,
    n51369, n51371, n51372, n51374, n51375, n51377, n51378, n51380, n51381,
    n51383, n51384, n51386, n51387, n51388, n51390, n51391, n51392, n51393,
    n51395, n51396, n51398, n51399, n51401, n51402, n51404, n51405, n51407,
    n51408, n51410, n51411, n51413, n51414, n51416, n51417, n51419, n51420,
    n51422, n51423, n51425, n51426, n51428, n51429, n51431, n51432, n51434,
    n51435, n51437, n51438, n51440, n51441, n51443, n51444, n51446, n51447,
    n51448, n51450, n51451, n51452, n51453, n51454, n51456, n51457, n51459,
    n51460, n51462, n51463, n51465, n51466, n51468, n51469, n51471, n51472,
    n51474, n51475, n51477, n51478, n51480, n51481, n51483, n51484, n51486,
    n51487, n51489, n51490, n51492, n51493, n51495, n51496, n51498, n51499,
    n51501, n51502, n51504, n51505, n51507, n51508, n51510, n51511, n51513,
    n51514, n51516, n51517, n51519, n51520, n51522, n51523, n51525, n51526,
    n51528, n51529, n51531, n51532, n51534, n51535, n51536, n51538, n51539,
    n51541, n51542, n51544, n51545, n51547, n51548, n51550, n51551, n51553,
    n51554, n51556, n51557, n51559, n51560, n51562, n51563, n51565, n51566,
    n51568, n51569, n51571, n51572, n51574, n51575, n51577, n51578, n51580,
    n51581, n51583, n51584, n51586, n51587, n51589, n51590, n51592, n51593,
    n51595, n51596, n51598, n51599, n51601, n51602, n51604, n51605, n51607,
    n51608, n51609, n51611, n51612, n51613, n51615, n51616, n51617, n51619,
    n51620, n51622, n51623, n51625, n51626, n51628, n51629, n51631, n51632,
    n51634, n51635, n51637, n51638, n51640, n51641, n51643, n51644, n51646,
    n51647, n51649, n51650, n51652, n51653, n51655, n51656, n51658, n51659,
    n51661, n51662, n51664, n51665, n51667, n51668, n51670, n51671, n51673,
    n51674, n51676, n51677, n51679, n51680, n51682, n51683, n51685, n51686,
    n51688, n51689, n51691, n51692, n51694, n51695, n51697, n51698, n51700,
    n51701, n51703, n51704, n51706, n51707, n51709, n51710, n51712, n51713,
    n51715, n51716, n51718, n51719, n51721, n51722, n51724, n51725, n51727,
    n51728, n51730, n51731, n51732, n51733, n51735, n51736, n51737, n51739,
    n51740, n51742, n51743, n51745, n51746, n51748, n51749, n51751, n51752,
    n51754, n51755, n51757, n51758, n51760, n51761, n51763, n51764, n51766,
    n51767, n51769, n51770, n51772, n51773, n51775, n51776, n51778, n51779,
    n51781, n51782, n51784, n51785, n51787, n51788, n51790, n51791, n51793,
    n51794, n51796, n51797, n51799, n51800, n51802, n51803, n51804, n51805,
    n51807, n51808, n51809, n51811, n51812, n51813, n51815, n51816, n51818,
    n51819, n51820, n51822, n51823, n51825, n51826, n51828, n51829, n51831,
    n51832, n51833, n51835, n51836, n51837, n51838, n51839, n51841, n51842,
    n51844, n51845, n51847, n51848, n51850, n51851, n51853, n51854, n51856,
    n51857, n51859, n51860, n51862, n51863, n51865, n51866, n51868, n51869,
    n51871, n51872, n51874, n51875, n51877, n51878, n51880, n51881, n51883,
    n51884, n51886, n51887, n51889, n51890, n51892, n51893, n51895, n51896,
    n51898, n51899, n51901, n51902, n51904, n51905, n51907, n51908, n51910,
    n51911, n51913, n51914, n51916, n51917, n51919, n51920, n51922, n51923,
    n51925, n51926, n51928, n51929, n51931, n51932, n51934, n51935, n51937,
    n51938, n51940, n51941, n51943, n51944, n51946, n51947, n51949, n51950,
    n51952, n51953, n51955, n51956, n51958, n51959, n51961, n51962, n51964,
    n51965, n51967, n51968, n51970, n51971, n51973, n51974, n51976, n51977,
    n51979, n51980, n51982, n51983, n51985, n51986, n51988, n51989, n51991,
    n51992, n51994, n51995, n51997, n51998, n52000, n52001, n52003, n52004,
    n52006, n52007, n52009, n52010, n52012, n52013, n52015, n52016, n52018,
    n52019, n52021, n52022, n52024, n52025, n52027, n52028, n52030, n52031,
    n52033, n52034, n52036, n52037, n52039, n52040, n52042, n52043, n52045,
    n52046, n52048, n52049, n52051, n52052, n52054, n52055, n52057, n52058,
    n52060, n52061, n52063, n52064, n52066, n52067, n52069, n52070, n52072,
    n52073, n52075, n52076, n52078, n52079, n52081, n52082, n52084, n52085,
    n52087, n52088, n52089, n52091, n52092, n52094, n52095, n52097, n52098,
    n52100, n52101, n52103, n52104, n52106, n52107, n52109, n52110, n52112,
    n52113, n52114, n52116, n52117, n52119, n52120, n52122, n52123, n52125,
    n52126, n52128, n52129, n52131, n52132, n52134, n52135, n52137, n52138,
    n52140, n52141, n52143, n52144, n52146, n52147, n52149, n52150, n52152,
    n52153, n52155, n52156, n52158, n52159, n52161, n52162, n52164, n52165,
    n52167, n52168, n52170, n52171, n52173, n52174, n52176, n52177, n52179,
    n52180, n52182, n52183, n52185, n52186, n52188, n52189, n52191, n52192,
    n52194, n52195, n52197, n52198, n52200, n52201, n52203, n52204, n52206,
    n52207, n52209, n52210, n52212, n52213, n52215, n52216, n52218, n52219,
    n52221, n52222, n52224, n52225, n52227, n52228, n52229, n52230, n52231,
    n52233, n52234, n52235, n52237, n52238, n52239, n52241, n52242, n52243,
    n52245, n52246, n52247, n52248, n52249, n52251, n52252, n52253, n52255,
    n52256, n52258, n52259, n52261, n52262, n52264, n52265, n52267, n52268,
    n52269, n52271, n52272, n52274, n52275, n52277, n52278, n52279, n52281,
    n52282, n52284, n52285, n52287, n52288, n52290, n52291, n52293, n52294,
    n52296, n52297, n52299, n52300, n52301, n52303, n52304, n52305, n52306,
    n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314, n52315,
    n52316, n52317, n52318, n52319, n52320, n52321, n52322, n52323, n52324,
    n52326, n52328, n52329, n52330, n52332, n52333, n52335, n52336, n52338,
    n52339, n52341, n52343, n52345, n52346, n52347, n52348, n52349, n52351,
    n52352, n52354, n52355, n52357, n52358, n52360, n52361, n52363, n52364,
    n52366, n52367, n52369, n52370, n52372, n52373, n52375, n52376, n52378,
    n52379, n52381, n52382, n52384, n52385, n52387, n52388, n52390, n52391,
    n52393, n52394, n52396, n52397, n52399, n52400, n52402, n52403, n52405,
    n52406, n52408, n52409, n52411, n52412, n52414, n52415, n52417, n52418,
    n52420, n52421, n52423, n52424, n52426, n52427, n52429, n52430, n52432,
    n52433, n52435, n52436, n52438, n52439, n52441, n52442, n52444, n52445,
    n52447, n52448, n52450, n52451, n52453, n52454, n52456, n52457, n52459,
    n52460, n52462, n52463, n52464, n52466, n52467, n52468, n52470, n52472,
    n52473, n52474, n52476, n52477, n52478, n52479, n52480, n52482, n52483,
    n52485, n52486, n52487, n52489, n52490, n52491, n52493, n52494, n52495,
    n52497, n52498, n52499, n52501, n52502, n52503, n52505, n52506, n52507,
    n52509, n52510, n52511, n52513, n52514, n52515, n52516, n52517, n52519,
    n52521, n52522, n52524, n52525, n52527, n52528, n52529, n52530, n52532,
    n52533, n52534, n52536, n52538, n52539, n52540, n52541, n52542, n52544,
    n52545, n52546, n52547, n52548, n52550, n52551, n52552, n52553, n52554,
    n52556, n52557, n52558, n52559, n52560, n52562, n52563, n52564, n52566,
    n52567, n52569, n52570, n52571, n52573, n52574, n52575, n52577, n52578,
    n52579, n52581, n52582, n52583, n52584, n52585, n52586, n52587, n52589,
    n52590, n52592, n52593, n52594, n52596, n52597, n52598, n52599, n52600,
    n52601, n52603, n52604, n52605, n52606, n52607, n52608, n52610, n52611,
    n52612, n52613, n52614, n52615, n52617, n52618, n52619, n52620, n52621,
    n52622, n52624, n52625, n52626, n52627, n52628, n52629, n52631, n52632,
    n52633, n52634, n52635, n52636, n52638, n52639, n52640, n52641, n52642,
    n52643, n52645, n52646, n52647, n52648, n52649, n52650, n52652, n52653,
    n52654, n52656, n52657, n52658, n52660, n52661, n52662, n52663, n52664,
    n52666, n52667, n52668, n52669, n52670, n52672, n52673, n52674, n52675,
    n52676, n52678, n52679, n52680, n52681, n52682, n52684, n52685, n52686,
    n52688, n52689, n52691, n52692, n52693, n52694, n52695, n52697, n52698,
    n52699, n52700, n52701, n52703, n52704, n52705, n52706, n52707, n52709,
    n52710, n52711, n52713, n52714, n52715, n52717, n52718, n52719, n52721,
    n52722, n52723, n52724, n52725, n52726, n52728, n52729, n52730, n52731,
    n52732, n52733, n52735, n52736, n52737, n52738, n52739, n52740, n52742,
    n52743, n52744, n52745, n52746, n52747, n52749, n52750, n52752, n52753,
    n52755, n52756, n52757, n52758, n52760, n52761, n52762, n52763, n52764,
    n52766, n52767, n52768, n52770, n52771, n52772, n52773, n52774, n52776,
    n52777, n52778, n52779, n52781, n52782, n52784, n52786, n52788, n52789,
    n52791, n52792, n52794, n52795, n52797, n52798, n52800, n52801, n52803,
    n52804, n52806, n52807, n52809, n52810, n52812, n52813, n52815, n52816,
    n52817, n52819, n52820, n52821, n52823, n52824, n52827, n52828, n52829,
    n52831, n52833, n52835, n52836, n52838, n52839, n52841, n52842, n52844,
    n52845, n52847, n52848, n52850, n52851, n52853, n52854, n52857, n52858,
    n52859, n52861, n52863, n52865, n52866, n52868, n52869, n52871, n52872,
    n52873, n52874, n52875, n52876, n52878, n52879, n52881, n52882, n52884,
    n52885, n52887, n52888, n52889, n52891, n52892, n52894, n52895, n52897,
    n52898, n52900, n52901, n52903, n52904, n52906, n52907, n52908, n52909,
    n52911, n52912, n52914, n52915, n52916, n52918, n52919, n52920, n52921,
    n52922, n52923, n52925, n52926, n52927, n52928, n52929, n52931, n52932,
    n52933, n52934, n52935, n52937, n52938, n52939, n52940, n52941, n52943,
    n52944, n52945, n52947, n52948, n52951, n52952, n52954, n52955, n52956,
    n52958, n52959, n52960, n52961, n52962, n52964, n52965, n52966, n52967,
    n52968, n52970, n52971, n52972, n52973, n52974, n52976, n52977, n52978,
    n52979, n52980, n52982, n52983, n52984, n52985, n52986, n52988, n52989,
    n52990, n52991, n52992, n52994, n52995, n52996, n52997, n52998, n53000,
    n53001, n53002, n53003, n53004, n53006, n53007, n53008, n53009, n53010,
    n53012, n53013, n53014, n53015, n53016, n53018, n53019, n53020, n53021,
    n53022, n53024, n53026, n53028, n53029, n53031, n53033, n53034, n53036,
    n53037, n53039, n53040, n53041, n53043, n53044, n53046, n53047, n53049,
    n53050, n53052, n53054, n53055, n53056, n53058, n53059, n53061, n53062,
    n53064, n53065, n53067, n53068, n53070, n53071, n53073, n53074, n53075,
    n53076, n53077, n53079, n53080, n53082, n53083, n53085, n53086, n53088,
    n53089, n53091, n53092, n53094, n53095, n53096, n53098, n53099, n53101,
    n53102, n53104, n53106, n53107, n53109, n53111, n53112, n53114, n53115,
    n53118, n53120, n53121, n53123, n53124, n53126, n53127, n53129, n53130,
    n53132, n53133, n53135, n53137, n53138, n53139, n53140, n53141, n53143,
    n53144, n53146, n53147, n53149, n53150, n53155, n53156, n53158, n53159,
    n53163, n53164, n53165, n53167, n53168, n53169, n53175, n53176, n53178,
    n53179, n53181, n53182, n53188, n53196, n53197, n53199, n53200, n53202,
    n53203, n53205, n53207, n53208, n53210, n53212, n53213, n53215, n53216,
    n53218, n53219, n53221, n53224, n53225, n53227, n53228, n53230, n53231,
    n53233, n53234, n53236, n53237, n53239, n53240, n53242, n53243, n53246,
    n53247, n53249, n53251, n53252, n53254, n53255, n53256, n53258, n53259,
    n53261, n53262, n53264, n53265, n53267, n53268, n53269, n53270, n53272,
    n53274, n53275, n53277, n53278, n53280, n53281, n53283, n53284, n53285,
    n53287, n53288, n53289, n53292, n53293, n53295, n53296, n53297, n53299,
    n53300, n53302, n53303, n53304, n53306, n53307, n53309, n53310, n53312,
    n53313, n53315, n53316, n53318, n53319, n53321, n53323, n53324, n53326,
    n53327, n53329, n53330, n53332, n53333, n53335, n53336, n53338, n53339,
    n53341, n53342, n53344, n53346, n53347, n53349, n53350, n53352, n53353,
    n53355, n53356, n53358, n53359, n53361, n53362, n53364, n53365, n53367,
    n53368, n53370, n53371, n53373, n53374, n53376, n53377, n53379, n53380,
    n53382, n53383, n53385, n53386, n53388, n53389, n53391, n53392, n53394,
    n53395, n53397, n53398, n53400, n53401, n53403, n53404, n53406, n53407,
    n53410, n53412, n53413, n53415, n53416, n53418, n53419, n53421, n53422,
    n53424, n53425, n53427, n53428, n53430, n53431, n53433, n53434, n53436,
    n53437, n53439, n53440, n53442, n53443, n53446, n53447, n53451, n53452,
    n53453, n53454, n53455, n53457, n53458, n53460, n53461, n53463, n53464,
    n53466, n53467, n53469, n53470, n53472, n53473, n53475, n53476, n53478,
    n53479, n53481, n53482, n53484, n53485, n53487, n53488, n53490, n53491,
    n53493, n53494, n53496, n53497, n53499, n53500, n53502, n53503, n53505,
    n53506, n53508, n53509, n53511, n53512, n53514, n53515, n53517, n53518,
    n53520, n53521, n53523, n53524, n53526, n53527, n53529, n53530, n53532,
    n53533, n53536, n53537, n53539, n53540, n53541, n53542, n53543, n53544,
    n53546, n53547, n53548, n53549, n53551, n53553, n53554, n53555, n53556,
    n53557, n53558, n53559, n53560, n53561, n53563, n53564, n53567, n53568,
    n53570, n53571, n53572, n53573, n53577, n53578, n53579, n53580, n53581,
    n53582, n53583, n53584, n53585, n53586, n53587, n53588, n53589, n53590,
    n53591, n53592, n53593, n53594, n53595;
  assign po0767 = pi3649 & pi3650;
  assign n8179 = pi0939 & po0767;
  assign n8180 = pi3654 & ~pi3655;
  assign n8181 = pi3653 & pi3655;
  assign n8182 = ~n8180 & ~n8181;
  assign po0011 = ~pi2604 | ~po0767;
  assign po1235 = ~n8182 & po0011;
  assign n8185 = ~n8179 & po1235;
  assign n8186 = pi1609 & n8179;
  assign po3741 = n8185 | n8186;
  assign n8188 = pi3415 & po0767;
  assign po3853 = ~po3741 & ~n8188;
  assign po0009 = ~pi1835 & pi2386;
  assign n8191 = ~pi3294 & ~pi3322;
  assign n8192 = pi3323 & pi3324;
  assign n8193 = n8191 & n8192;
  assign n8194 = pi3323 & ~pi3324;
  assign n8195 = pi3294 & ~pi3322;
  assign n8196 = n8194 & n8195;
  assign n8197 = ~pi3323 & ~pi3324;
  assign n8198 = pi3294 & pi3322;
  assign n8199 = n8197 & n8198;
  assign n8200 = ~pi3294 & pi3322;
  assign n8201 = n8194 & n8200;
  assign n8202 = ~pi3419 & n8200;
  assign n8203 = n8192 & n8202;
  assign n8204 = n8194 & n8198;
  assign n8205 = pi1860 & n8204;
  assign n8206 = ~n8203 & ~n8205;
  assign n8207 = ~n8201 & n8206;
  assign n8208 = ~n8199 & n8207;
  assign n8209 = n8197 & n8200;
  assign n8210 = ~pi3323 & pi3324;
  assign n8211 = n8200 & n8210;
  assign n8212 = ~n8209 & ~n8211;
  assign n8213 = n8191 & n8210;
  assign n8214 = ~n8193 & ~n8213;
  assign n8215 = pi3682 & ~n8214;
  assign n8216 = ~pi1462 & ~pi2785;
  assign n8217 = ~pi2813 & n8216;
  assign n8218 = pi3631 & pi3682;
  assign n8219 = ~pi2114 & n8218;
  assign n8220 = n8217 & n8219;
  assign n8221 = ~pi3631 & n8216;
  assign n8222 = ~pi3682 & n8221;
  assign n8223 = pi0783 & n8222;
  assign n8224 = ~pi2114 & ~pi2813;
  assign n8225 = n8223 & n8224;
  assign n8226 = ~n8220 & ~n8225;
  assign n8227 = n8191 & n8197;
  assign n8228 = ~n8226 & n8227;
  assign n8229 = ~n8215 & ~n8228;
  assign n8230 = n8212 & n8229;
  assign po3645 = ~n8208 | ~n8230;
  assign n8232 = n8195 & n8197;
  assign n8233 = ~n8199 & ~n8232;
  assign n8234 = ~n8196 & n8233;
  assign n8235 = pi1928 & ~pi2785;
  assign n8236 = pi1780 & pi2785;
  assign n8237 = ~n8235 & ~n8236;
  assign n8238 = ~pi1462 & ~n8237;
  assign n8239 = pi1462 & pi1772;
  assign n8240 = ~n8238 & ~n8239;
  assign n8241 = ~pi2114 & ~n8240;
  assign n8242 = pi1776 & pi2114;
  assign n8243 = ~n8241 & ~n8242;
  assign n8244 = pi2825 & ~n8243;
  assign n8245 = ~pi2825 & n8243;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = pi1944 & ~pi2785;
  assign n8248 = pi1778 & pi2785;
  assign n8249 = ~n8247 & ~n8248;
  assign n8250 = ~pi1462 & ~n8249;
  assign n8251 = pi1462 & pi1784;
  assign n8252 = ~n8250 & ~n8251;
  assign n8253 = ~pi2114 & ~n8252;
  assign n8254 = pi1774 & pi2114;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = pi2600 & ~n8255;
  assign n8257 = ~pi2600 & n8255;
  assign n8258 = ~n8256 & ~n8257;
  assign n8259 = ~pi1462 & pi2785;
  assign n8260 = pi1942 & n8259;
  assign n8261 = pi1462 & pi1938;
  assign n8262 = ~n8260 & ~n8261;
  assign n8263 = ~pi2114 & ~n8262;
  assign n8264 = pi1940 & pi2114;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = pi2113 & ~n8265;
  assign n8267 = ~pi2113 & n8265;
  assign n8268 = ~n8266 & ~n8267;
  assign n8269 = pi1929 & ~pi2785;
  assign n8270 = pi1786 & pi2785;
  assign n8271 = ~n8269 & ~n8270;
  assign n8272 = ~pi1462 & ~n8271;
  assign n8273 = pi1462 & pi1773;
  assign n8274 = ~n8272 & ~n8273;
  assign n8275 = ~pi2114 & ~n8274;
  assign n8276 = pi1777 & pi2114;
  assign n8277 = ~n8275 & ~n8276;
  assign n8278 = pi2798 & ~n8277;
  assign n8279 = ~pi2798 & n8277;
  assign n8280 = ~n8278 & ~n8279;
  assign n8281 = pi1945 & ~pi2785;
  assign n8282 = pi1779 & pi2785;
  assign n8283 = ~n8281 & ~n8282;
  assign n8284 = ~pi1462 & ~n8283;
  assign n8285 = pi1462 & pi1785;
  assign n8286 = ~n8284 & ~n8285;
  assign n8287 = ~pi2114 & ~n8286;
  assign n8288 = pi1775 & pi2114;
  assign n8289 = ~n8287 & ~n8288;
  assign n8290 = pi2799 & ~n8289;
  assign n8291 = ~pi2799 & n8289;
  assign n8292 = ~n8290 & ~n8291;
  assign n8293 = ~n8280 & ~n8292;
  assign n8294 = ~n8268 & n8293;
  assign n8295 = ~n8258 & n8294;
  assign n8296 = ~n8246 & n8295;
  assign n8297 = pi1943 & n8259;
  assign n8298 = pi1462 & pi1939;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = ~pi2114 & ~n8299;
  assign n8301 = pi1941 & pi2114;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = ~pi2082 & n8302;
  assign n8304 = n8296 & n8303;
  assign n8305 = pi2082 & ~n8302;
  assign n8306 = n8296 & n8305;
  assign n8307 = ~n8304 & ~n8306;
  assign n8308 = ~n8234 & ~n8307;
  assign n8309 = ~n8203 & ~n8308;
  assign n8310 = ~n8205 & n8309;
  assign po3647 = n8211 | ~n8310;
  assign n8312 = ~po3645 & ~po3647;
  assign n8313 = n8195 & n8210;
  assign n8314 = pi3631 & n8227;
  assign n8315 = ~n8216 & n8314;
  assign n8316 = n8224 & n8315;
  assign n8317 = n8224 & n8227;
  assign n8318 = n8223 & n8317;
  assign n8319 = ~n8316 & ~n8318;
  assign n8320 = ~n8313 & n8319;
  assign n8321 = n8191 & n8194;
  assign n8322 = ~n8201 & ~n8205;
  assign n8323 = ~n8196 & n8322;
  assign n8324 = ~n8203 & n8323;
  assign n8325 = ~n8321 & n8324;
  assign po3646 = ~n8320 | ~n8325;
  assign n8327 = pi2522 & pi3099;
  assign n8328 = pi2504 & ~pi3099;
  assign n8329 = ~n8327 & ~n8328;
  assign n8330 = pi3199 & ~n8329;
  assign n8331 = ~pi3199 & n8329;
  assign n8332 = ~n8330 & ~n8331;
  assign n8333 = pi2503 & ~pi3099;
  assign n8334 = pi2504 & pi3099;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = pi2759 & ~n8335;
  assign n8337 = ~pi2759 & n8335;
  assign n8338 = ~n8336 & ~n8337;
  assign n8339 = ~pi2505 & ~pi3099;
  assign n8340 = ~pi3343 & n8339;
  assign n8341 = pi3343 & ~n8339;
  assign n8342 = ~n8340 & ~n8341;
  assign n8343 = n8201 & ~n8342;
  assign n8344 = ~pi2503 & pi3099;
  assign n8345 = ~pi2049 & ~n8344;
  assign n8346 = pi2049 & n8344;
  assign n8347 = ~n8345 & ~n8346;
  assign n8348 = n8343 & n8347;
  assign n8349 = pi2522 & ~pi3099;
  assign n8350 = pi2505 & pi3099;
  assign n8351 = ~n8349 & ~n8350;
  assign n8352 = pi3281 & ~n8351;
  assign n8353 = ~pi3281 & n8351;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = n8348 & ~n8354;
  assign n8356 = ~n8338 & n8355;
  assign n8357 = ~n8332 & n8356;
  assign n8358 = ~pi1035 & pi2978;
  assign n8359 = pi3344 & n8358;
  assign n8360 = ~n8307 & ~n8359;
  assign n8361 = n8232 & ~n8360;
  assign n8362 = ~pi2114 & n8216;
  assign n8363 = n8227 & ~n8362;
  assign n8364 = ~pi2813 & pi3631;
  assign n8365 = n8363 & n8364;
  assign n8366 = ~n8321 & ~n8365;
  assign n8367 = ~n8196 & ~n8199;
  assign n8368 = n8307 & ~n8367;
  assign n8369 = ~n8212 & ~n8307;
  assign n8370 = ~n8368 & ~n8369;
  assign n8371 = n8366 & n8370;
  assign n8372 = ~n8361 & n8371;
  assign po3616 = n8357 | ~n8372;
  assign n8374 = po3646 & po3616;
  assign n8375 = n8312 & n8374;
  assign n8376 = ~n8196 & ~n8375;
  assign n8377 = ~n8193 & n8376;
  assign po0017 = ~pi2785 | n8377;
  assign n8379 = pi3626 & po0017;
  assign n8380 = n8312 & ~po3646;
  assign n8381 = po3616 & n8380;
  assign n8382 = ~n8213 & ~n8381;
  assign po0014 = ~n8232 & n8382;
  assign po0015 = ~pi1462 | n8377;
  assign n8385 = po0014 & po0015;
  assign n8386 = ~n8209 & n8385;
  assign n8387 = ~n8199 & n8386;
  assign n8388 = n8198 & n8210;
  assign n8389 = ~n8211 & ~n8388;
  assign n8390 = ~pi3305 & pi3390;
  assign n8391 = ~n8389 & n8390;
  assign n8392 = n8387 & ~n8391;
  assign n8393 = n8379 & n8392;
  assign po0013 = ~pi3452 & ~n8393;
  assign n8395 = pi1781 & ~po0017;
  assign n8396 = pi1782 & ~po0015;
  assign n8397 = ~n8395 & ~n8396;
  assign n8398 = pi1783 & ~po0014;
  assign po0018 = n8397 & ~n8398;
  assign n8400 = pi3622 & pi3626;
  assign n8401 = pi1601 & ~pi3626;
  assign po0020 = n8400 | n8401;
  assign po0021 = ~pi3452 & pi3620;
  assign po0022 = ~pi3626 | po0021;
  assign n8405 = pi3099 & ~pi3626;
  assign po0023 = po0021 | n8405;
  assign n8407 = ~pi0795 & pi3609;
  assign n8408 = pi0795 & pi3607;
  assign n8409 = ~n8407 & ~n8408;
  assign n8410 = ~pi0793 & pi1009;
  assign n8411 = ~n8409 & n8410;
  assign n8412 = ~pi0795 & pi3605;
  assign n8413 = pi0795 & pi3603;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = pi0793 & pi1009;
  assign n8416 = ~n8414 & n8415;
  assign n8417 = ~n8411 & ~n8416;
  assign n8418 = ~pi0795 & pi3618;
  assign n8419 = pi0795 & pi3615;
  assign n8420 = ~n8418 & ~n8419;
  assign n8421 = ~pi0793 & ~pi1009;
  assign n8422 = ~n8420 & n8421;
  assign n8423 = ~pi0795 & pi3613;
  assign n8424 = pi0795 & pi3611;
  assign n8425 = ~n8423 & ~n8424;
  assign n8426 = pi0793 & ~pi1009;
  assign n8427 = ~n8425 & n8426;
  assign n8428 = ~n8422 & ~n8427;
  assign n8429 = n8417 & n8428;
  assign n8430 = ~pi0957 & ~n8429;
  assign n8431 = ~pi0795 & pi3595;
  assign n8432 = pi0795 & pi3594;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = n8410 & ~n8433;
  assign n8435 = ~pi0795 & ~pi3593;
  assign n8436 = pi0795 & ~pi3592;
  assign n8437 = ~n8435 & ~n8436;
  assign n8438 = n8415 & ~n8437;
  assign n8439 = ~n8434 & ~n8438;
  assign n8440 = ~pi0795 & pi3598;
  assign n8441 = pi0795 & pi3596;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = n8426 & ~n8442;
  assign n8444 = ~pi0795 & pi3601;
  assign n8445 = pi0795 & pi3599;
  assign n8446 = ~n8444 & ~n8445;
  assign n8447 = n8421 & ~n8446;
  assign n8448 = ~n8443 & ~n8447;
  assign n8449 = n8439 & n8448;
  assign n8450 = pi0957 & ~n8449;
  assign n8451 = ~n8430 & ~n8450;
  assign n8452 = ~pi0799 & ~n8451;
  assign n8453 = pi0799 & ~pi3592;
  assign n8454 = ~n8452 & ~n8453;
  assign po0026 = ~pi0958 & ~n8454;
  assign n8456 = pi0893 & pi3461;
  assign n8457 = pi0739 & ~pi0885;
  assign n8458 = ~pi0741 & pi3617;
  assign n8459 = pi0741 & pi3616;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = n8457 & ~n8460;
  assign n8462 = ~pi0739 & ~pi0885;
  assign n8463 = ~pi0741 & pi3623;
  assign n8464 = pi0741 & pi3619;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = n8462 & ~n8465;
  assign n8467 = ~n8461 & ~n8466;
  assign n8468 = ~pi0739 & pi0885;
  assign n8469 = ~pi0741 & pi3614;
  assign n8470 = pi0741 & pi3612;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = n8468 & ~n8471;
  assign n8473 = pi0739 & pi0885;
  assign n8474 = ~pi0741 & pi3610;
  assign n8475 = pi0741 & pi3608;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = n8473 & ~n8476;
  assign n8478 = ~n8472 & ~n8477;
  assign n8479 = n8467 & n8478;
  assign n8480 = ~pi0884 & ~n8479;
  assign n8481 = ~pi0741 & pi3473;
  assign n8482 = pi0741 & pi3461;
  assign n8483 = ~n8481 & ~n8482;
  assign n8484 = n8473 & ~n8483;
  assign n8485 = ~pi0741 & ~pi3597;
  assign n8486 = pi0741 & pi3471;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = n8468 & ~n8487;
  assign n8489 = ~n8484 & ~n8488;
  assign n8490 = ~pi0741 & pi3602;
  assign n8491 = pi0741 & pi3600;
  assign n8492 = ~n8490 & ~n8491;
  assign n8493 = n8457 & ~n8492;
  assign n8494 = n8489 & ~n8493;
  assign n8495 = ~pi0741 & pi3606;
  assign n8496 = pi0741 & pi3604;
  assign n8497 = ~n8495 & ~n8496;
  assign n8498 = n8462 & ~n8497;
  assign n8499 = n8494 & ~n8498;
  assign n8500 = pi0884 & ~n8499;
  assign n8501 = ~n8480 & ~n8500;
  assign n8502 = ~pi0893 & ~n8501;
  assign n8503 = ~n8456 & ~n8502;
  assign po0027 = ~pi0886 & ~n8503;
  assign n8505 = ~pi0960 & pi1746;
  assign n8506 = pi0960 & ~pi1746;
  assign po0028 = n8505 | n8506;
  assign n8508 = ~pi0888 & pi1739;
  assign n8509 = pi0888 & ~pi1739;
  assign po0030 = n8508 | n8509;
  assign n8511 = pi0954 & ~pi1002;
  assign n8512 = ~pi0954 & pi1002;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = pi0796 & pi0962;
  assign po0032 = ~n8513 | n8514;
  assign n8516 = ~pi0956 & pi1002;
  assign n8517 = pi0956 & ~pi1002;
  assign n8518 = ~n8516 & ~n8517;
  assign po0034 = n8514 | ~n8518;
  assign n8520 = pi0881 & ~pi1001;
  assign n8521 = ~pi0881 & pi1001;
  assign n8522 = ~n8520 & ~n8521;
  assign n8523 = pi0890 & pi0947;
  assign po0036 = ~n8522 | n8523;
  assign n8525 = ~pi0880 & pi1001;
  assign n8526 = pi0880 & ~pi1001;
  assign n8527 = ~n8525 & ~n8526;
  assign po0038 = n8523 | ~n8527;
  assign po0041 = pi2515 | pi3645;
  assign po0043 = ~pi3632 & ~pi3677;
  assign n8531 = ~pi0541 & ~pi0565;
  assign n8532 = ~pi0404 & ~pi3190;
  assign n8533 = ~pi0684 & ~pi3515;
  assign n8534 = n8532 & n8533;
  assign n8535 = ~pi3148 & n8534;
  assign n8536 = pi3528 & n8535;
  assign n8537 = n8531 & n8536;
  assign n8538 = pi2813 & pi3526;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = ~pi0541 & pi3548;
  assign n8541 = ~pi0565 & n8540;
  assign n8542 = ~pi3452 & n8541;
  assign n8543 = ~pi3522 & ~pi3523;
  assign n8544 = ~pi0565 & ~n8543;
  assign n8545 = ~pi3215 & n8531;
  assign n8546 = pi3505 & n8535;
  assign n8547 = n8545 & n8546;
  assign n8548 = ~pi1046 & ~pi2800;
  assign n8549 = pi3416 & ~n8548;
  assign n8550 = ~pi3416 & pi3583;
  assign n8551 = ~n8549 & ~n8550;
  assign n8552 = pi3524 & ~n8551;
  assign n8553 = ~n8547 & ~n8552;
  assign n8554 = ~n8544 & n8553;
  assign n8555 = ~n8542 & n8554;
  assign po3946 = ~n8539 | ~n8555;
  assign n8557 = pi2813 & pi3643;
  assign n8558 = ~pi0565 & pi3547;
  assign po3873 = n8557 | n8558;
  assign po3831 = po3946 | po3873;
  assign n8561 = ~pi3551 & ~po3831;
  assign n8562 = ~pi3515 & n8561;
  assign n8563 = ~pi0784 & ~pi1449;
  assign n8564 = ~pi3416 & n8563;
  assign n8565 = n8562 & n8564;
  assign n8566 = pi3585 & pi3631;
  assign n8567 = n8565 & ~n8566;
  assign n8568 = pi3376 & pi3641;
  assign n8569 = pi1642 & pi3641;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = pi1860 & pi3641;
  assign n8572 = n8570 & n8571;
  assign n8573 = pi3304 & pi3641;
  assign n8574 = pi2598 & pi3641;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = ~pi2601 & n8575;
  assign n8577 = n8572 & n8576;
  assign n8578 = ~pi1840 & ~pi1861;
  assign n8579 = pi3099 & n8578;
  assign n8580 = ~pi2986 & ~pi2990;
  assign n8581 = pi0783 & pi3585;
  assign n8582 = n8580 & n8581;
  assign n8583 = pi0752 & n8582;
  assign n8584 = ~pi0779 & ~pi3680;
  assign n8585 = n8583 & ~n8584;
  assign n8586 = n8579 & n8585;
  assign n8587 = n8577 & n8586;
  assign n8588 = n8570 & n8575;
  assign n8589 = pi2601 & n8588;
  assign n8590 = ~pi0819 & ~pi3680;
  assign n8591 = pi0909 & ~n8590;
  assign n8592 = ~pi1422 & pi2515;
  assign n8593 = n8591 & n8592;
  assign n8594 = n8589 & n8593;
  assign n8595 = ~n8587 & ~n8594;
  assign n8596 = ~pi1840 & pi1861;
  assign n8597 = n8583 & n8596;
  assign n8598 = ~n8584 & n8597;
  assign n8599 = ~pi3099 & n8598;
  assign n8600 = n8577 & n8599;
  assign n8601 = ~pi1422 & pi2769;
  assign n8602 = n8589 & n8601;
  assign n8603 = n8591 & n8602;
  assign n8604 = ~n8600 & ~n8603;
  assign n8605 = n8595 & n8604;
  assign n8606 = ~n8567 & ~n8605;
  assign n8607 = ~pi0419 & ~pi0420;
  assign n8608 = ~pi0416 & ~pi0417;
  assign n8609 = ~pi0403 & n8608;
  assign n8610 = pi0418 & n8609;
  assign n8611 = pi0421 & n8610;
  assign n8612 = n8607 & n8611;
  assign n8613 = ~pi0422 & n8612;
  assign n8614 = pi0403 & ~pi0417;
  assign n8615 = pi0416 & n8614;
  assign n8616 = ~n8613 & ~n8615;
  assign n8617 = pi0417 & ~pi0418;
  assign n8618 = ~pi0416 & n8617;
  assign n8619 = ~pi0403 & n8618;
  assign n8620 = ~pi0419 & n8619;
  assign n8621 = n8616 & ~n8620;
  assign n8622 = ~pi0692 & pi3216;
  assign n8623 = ~pi3426 & n8622;
  assign n8624 = ~n8561 & ~n8623;
  assign n8625 = ~pi3416 & ~po3831;
  assign n8626 = ~pi3515 & ~n8566;
  assign n8627 = n8625 & n8626;
  assign n8628 = n8563 & n8627;
  assign n8629 = ~pi2601 & ~n8574;
  assign n8630 = n8570 & ~n8571;
  assign n8631 = ~n8573 & n8630;
  assign n8632 = n8629 & n8631;
  assign po3841 = ~n8628 & ~n8632;
  assign n8634 = ~pi3299 & ~pi3326;
  assign n8635 = ~pi0149 & n8634;
  assign n8636 = pi3248 & n8635;
  assign n8637 = ~pi3267 & n8636;
  assign n8638 = ~pi0134 & ~pi0152;
  assign n8639 = pi0134 & pi0152;
  assign n8640 = ~n8638 & ~n8639;
  assign n8641 = ~pi0149 & ~n8640;
  assign n8642 = n8634 & n8641;
  assign n8643 = ~pi3248 & n8642;
  assign n8644 = pi3267 & n8643;
  assign n8645 = pi0149 & n8634;
  assign n8646 = ~pi3248 & n8645;
  assign n8647 = ~pi3267 & n8646;
  assign n8648 = ~n8644 & ~n8647;
  assign n8649 = ~pi0038 & n8648;
  assign n8650 = ~n8637 & n8649;
  assign n8651 = n8634 & ~n8641;
  assign n8652 = pi3248 & n8651;
  assign n8653 = pi3267 & n8652;
  assign n8654 = ~pi3248 & pi3326;
  assign n8655 = ~pi0482 & n8654;
  assign n8656 = pi3299 & n8655;
  assign n8657 = pi3267 & n8656;
  assign n8658 = ~pi3267 & pi3299;
  assign n8659 = n8654 & n8658;
  assign n8660 = ~n8657 & ~n8659;
  assign n8661 = ~n8653 & n8660;
  assign n8662 = n8650 & n8661;
  assign n8663 = ~pi3633 & ~n8662;
  assign n8664 = pi3326 & n8658;
  assign n8665 = pi3248 & n8664;
  assign n8666 = n8650 & ~n8657;
  assign n8667 = ~n8653 & n8666;
  assign n8668 = ~n8665 & n8667;
  assign n8669 = pi3633 & ~n8668;
  assign n8670 = ~n8663 & ~n8669;
  assign n8671 = pi2812 & pi2911;
  assign n8672 = ~pi2913 & n8671;
  assign n8673 = ~pi2912 & n8672;
  assign n8674 = ~pi2812 & ~pi2911;
  assign n8675 = pi2912 & n8674;
  assign n8676 = pi2913 & n8675;
  assign n8677 = n8641 & n8676;
  assign n8678 = ~pi2913 & ~n8641;
  assign n8679 = n8675 & n8678;
  assign n8680 = ~pi2912 & n8674;
  assign n8681 = pi0149 & pi2913;
  assign n8682 = n8680 & n8681;
  assign n8683 = ~n8679 & ~n8682;
  assign n8684 = ~pi0149 & ~pi2913;
  assign n8685 = n8680 & n8684;
  assign n8686 = n8683 & ~n8685;
  assign n8687 = ~pi0045 & n8686;
  assign n8688 = pi0482 & n8672;
  assign n8689 = pi2912 & n8688;
  assign n8690 = n8687 & ~n8689;
  assign n8691 = ~n8677 & n8690;
  assign n8692 = ~n8673 & n8691;
  assign n8693 = pi3633 & ~n8692;
  assign n8694 = pi2913 & n8671;
  assign n8695 = ~pi2912 & n8694;
  assign n8696 = n8691 & ~n8695;
  assign n8697 = ~pi3633 & ~n8696;
  assign n8698 = ~n8693 & ~n8697;
  assign n8699 = pi3268 & ~pi3426;
  assign n8700 = ~pi2490 & ~n8699;
  assign n8701 = pi2490 & n8699;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = ~pi1014 & ~pi1043;
  assign n8704 = pi0976 & ~pi1044;
  assign n8705 = n8703 & n8704;
  assign n8706 = pi1227 & n8705;
  assign n8707 = ~pi0976 & ~pi1044;
  assign n8708 = pi1014 & ~pi1043;
  assign n8709 = n8707 & n8708;
  assign n8710 = pi1213 & n8709;
  assign n8711 = ~n8706 & ~n8710;
  assign n8712 = pi0976 & pi1014;
  assign n8713 = pi1044 & n8712;
  assign n8714 = ~pi1043 & n8713;
  assign n8715 = pi1297 & n8714;
  assign n8716 = ~pi1043 & ~pi1044;
  assign n8717 = n8712 & n8716;
  assign n8718 = pi1199 & n8717;
  assign n8719 = ~n8715 & ~n8718;
  assign n8720 = ~pi0976 & pi1044;
  assign n8721 = n8708 & n8720;
  assign n8722 = pi1311 & n8721;
  assign n8723 = pi0976 & pi1044;
  assign n8724 = n8703 & n8723;
  assign n8725 = pi1115 & n8724;
  assign n8726 = ~n8722 & ~n8725;
  assign n8727 = pi1014 & pi1043;
  assign n8728 = n8707 & n8727;
  assign n8729 = pi1157 & n8728;
  assign n8730 = ~pi1014 & pi1043;
  assign n8731 = n8723 & n8730;
  assign n8732 = pi1269 & n8731;
  assign n8733 = ~n8729 & ~n8732;
  assign n8734 = ~pi0976 & ~pi1014;
  assign n8735 = ~pi1044 & n8734;
  assign n8736 = pi1043 & n8735;
  assign n8737 = pi1185 & n8736;
  assign n8738 = pi1043 & n8712;
  assign n8739 = ~pi1044 & n8738;
  assign n8740 = pi1143 & n8739;
  assign n8741 = ~n8737 & ~n8740;
  assign n8742 = ~pi1043 & n8734;
  assign n8743 = ~pi1044 & n8742;
  assign n8744 = pi1325 & n8743;
  assign n8745 = pi1044 & n8738;
  assign n8746 = pi1241 & n8745;
  assign n8747 = ~n8744 & ~n8746;
  assign n8748 = n8741 & n8747;
  assign n8749 = n8733 & n8748;
  assign n8750 = n8726 & n8749;
  assign n8751 = pi1043 & pi1044;
  assign n8752 = n8734 & n8751;
  assign n8753 = pi1283 & n8752;
  assign n8754 = pi1044 & n8742;
  assign n8755 = pi1129 & n8754;
  assign n8756 = ~n8753 & ~n8755;
  assign n8757 = n8750 & n8756;
  assign n8758 = n8704 & n8730;
  assign n8759 = pi1171 & n8758;
  assign n8760 = n8720 & n8727;
  assign n8761 = pi1255 & n8760;
  assign n8762 = ~n8759 & ~n8761;
  assign n8763 = n8757 & n8762;
  assign n8764 = n8719 & n8763;
  assign n8765 = n8711 & n8764;
  assign n8766 = ~pi2763 & ~n8765;
  assign n8767 = pi2375 & pi2763;
  assign n8768 = ~n8766 & ~n8767;
  assign n8769 = ~pi2484 & n8768;
  assign n8770 = pi2484 & ~n8768;
  assign n8771 = ~n8769 & ~n8770;
  assign n8772 = pi1310 & n8721;
  assign n8773 = pi1114 & n8724;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = pi1156 & n8728;
  assign n8776 = pi1268 & n8731;
  assign n8777 = ~n8775 & ~n8776;
  assign n8778 = pi1226 & n8705;
  assign n8779 = pi1212 & n8709;
  assign n8780 = ~n8778 & ~n8779;
  assign n8781 = pi1296 & n8714;
  assign n8782 = pi1198 & n8717;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = pi1282 & n8752;
  assign n8785 = pi1128 & n8754;
  assign n8786 = ~n8784 & ~n8785;
  assign n8787 = pi1170 & n8758;
  assign n8788 = pi1254 & n8760;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = n8786 & n8789;
  assign n8791 = n8783 & n8790;
  assign n8792 = n8780 & n8791;
  assign n8793 = pi1184 & n8736;
  assign n8794 = pi1142 & n8739;
  assign n8795 = ~n8793 & ~n8794;
  assign n8796 = n8792 & n8795;
  assign n8797 = pi1324 & n8743;
  assign n8798 = pi1240 & n8745;
  assign n8799 = ~n8797 & ~n8798;
  assign n8800 = n8796 & n8799;
  assign n8801 = n8777 & n8800;
  assign n8802 = n8774 & n8801;
  assign n8803 = ~pi2763 & ~n8802;
  assign n8804 = pi2015 & pi2763;
  assign n8805 = ~n8803 & ~n8804;
  assign n8806 = pi2483 & ~n8805;
  assign n8807 = ~pi2483 & n8805;
  assign n8808 = ~n8806 & ~n8807;
  assign n8809 = pi1224 & n8705;
  assign n8810 = pi1210 & n8709;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = pi1294 & n8714;
  assign n8813 = pi1196 & n8717;
  assign n8814 = ~n8812 & ~n8813;
  assign n8815 = pi1308 & n8721;
  assign n8816 = pi1112 & n8724;
  assign n8817 = ~n8815 & ~n8816;
  assign n8818 = pi1154 & n8728;
  assign n8819 = pi1266 & n8731;
  assign n8820 = ~n8818 & ~n8819;
  assign n8821 = pi1182 & n8736;
  assign n8822 = pi1140 & n8739;
  assign n8823 = ~n8821 & ~n8822;
  assign n8824 = pi1322 & n8743;
  assign n8825 = pi1238 & n8745;
  assign n8826 = ~n8824 & ~n8825;
  assign n8827 = n8823 & n8826;
  assign n8828 = n8820 & n8827;
  assign n8829 = n8817 & n8828;
  assign n8830 = pi1280 & n8752;
  assign n8831 = pi1126 & n8754;
  assign n8832 = ~n8830 & ~n8831;
  assign n8833 = n8829 & n8832;
  assign n8834 = pi1168 & n8758;
  assign n8835 = pi1252 & n8760;
  assign n8836 = ~n8834 & ~n8835;
  assign n8837 = n8833 & n8836;
  assign n8838 = n8814 & n8837;
  assign n8839 = n8811 & n8838;
  assign n8840 = ~pi2763 & ~n8839;
  assign n8841 = pi2013 & pi2763;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = pi2481 & ~n8842;
  assign n8844 = ~pi2481 & n8842;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = pi1222 & n8705;
  assign n8847 = pi1208 & n8709;
  assign n8848 = ~n8846 & ~n8847;
  assign n8849 = pi1292 & n8714;
  assign n8850 = pi1194 & n8717;
  assign n8851 = ~n8849 & ~n8850;
  assign n8852 = pi1306 & n8721;
  assign n8853 = pi1110 & n8724;
  assign n8854 = ~n8852 & ~n8853;
  assign n8855 = pi1152 & n8728;
  assign n8856 = pi1264 & n8731;
  assign n8857 = ~n8855 & ~n8856;
  assign n8858 = pi1180 & n8736;
  assign n8859 = pi1138 & n8739;
  assign n8860 = ~n8858 & ~n8859;
  assign n8861 = pi1320 & n8743;
  assign n8862 = pi1236 & n8745;
  assign n8863 = ~n8861 & ~n8862;
  assign n8864 = n8860 & n8863;
  assign n8865 = n8857 & n8864;
  assign n8866 = n8854 & n8865;
  assign n8867 = pi1278 & n8752;
  assign n8868 = pi1124 & n8754;
  assign n8869 = ~n8867 & ~n8868;
  assign n8870 = n8866 & n8869;
  assign n8871 = pi1166 & n8758;
  assign n8872 = pi1250 & n8760;
  assign n8873 = ~n8871 & ~n8872;
  assign n8874 = n8870 & n8873;
  assign n8875 = n8851 & n8874;
  assign n8876 = n8848 & n8875;
  assign n8877 = ~pi2763 & ~n8876;
  assign n8878 = pi2011 & pi2763;
  assign n8879 = ~n8877 & ~n8878;
  assign n8880 = pi2479 & ~n8879;
  assign n8881 = ~pi2479 & n8879;
  assign n8882 = ~n8880 & ~n8881;
  assign n8883 = pi1304 & n8721;
  assign n8884 = pi1108 & n8724;
  assign n8885 = ~n8883 & ~n8884;
  assign n8886 = pi1150 & n8728;
  assign n8887 = pi1262 & n8731;
  assign n8888 = ~n8886 & ~n8887;
  assign n8889 = pi1164 & n8758;
  assign n8890 = pi1248 & n8760;
  assign n8891 = ~n8889 & ~n8890;
  assign n8892 = pi1220 & n8705;
  assign n8893 = pi1206 & n8709;
  assign n8894 = ~n8892 & ~n8893;
  assign n8895 = pi1276 & n8752;
  assign n8896 = pi1122 & n8754;
  assign n8897 = ~n8895 & ~n8896;
  assign n8898 = pi1290 & n8714;
  assign n8899 = pi1192 & n8717;
  assign n8900 = ~n8898 & ~n8899;
  assign n8901 = n8897 & n8900;
  assign n8902 = n8894 & n8901;
  assign n8903 = n8891 & n8902;
  assign n8904 = pi1178 & n8736;
  assign n8905 = pi1136 & n8739;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = n8903 & n8906;
  assign n8908 = pi1318 & n8743;
  assign n8909 = pi1234 & n8745;
  assign n8910 = ~n8908 & ~n8909;
  assign n8911 = n8907 & n8910;
  assign n8912 = n8888 & n8911;
  assign n8913 = n8885 & n8912;
  assign n8914 = ~pi2763 & ~n8913;
  assign n8915 = pi2010 & pi2763;
  assign n8916 = ~n8914 & ~n8915;
  assign n8917 = pi2477 & ~n8916;
  assign n8918 = ~pi2477 & n8916;
  assign n8919 = ~n8917 & ~n8918;
  assign n8920 = pi1293 & n8714;
  assign n8921 = pi1195 & n8717;
  assign n8922 = ~n8920 & ~n8921;
  assign n8923 = pi1167 & n8758;
  assign n8924 = pi1251 & n8760;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = pi1153 & n8728;
  assign n8927 = pi1265 & n8731;
  assign n8928 = ~n8926 & ~n8927;
  assign n8929 = pi1307 & n8721;
  assign n8930 = pi1111 & n8724;
  assign n8931 = ~n8929 & ~n8930;
  assign n8932 = pi1321 & n8743;
  assign n8933 = pi1237 & n8745;
  assign n8934 = ~n8932 & ~n8933;
  assign n8935 = pi1181 & n8736;
  assign n8936 = pi1139 & n8739;
  assign n8937 = ~n8935 & ~n8936;
  assign n8938 = n8934 & n8937;
  assign n8939 = n8931 & n8938;
  assign n8940 = n8928 & n8939;
  assign n8941 = pi1279 & n8752;
  assign n8942 = pi1125 & n8754;
  assign n8943 = ~n8941 & ~n8942;
  assign n8944 = n8940 & n8943;
  assign n8945 = pi1223 & n8705;
  assign n8946 = pi1209 & n8709;
  assign n8947 = ~n8945 & ~n8946;
  assign n8948 = n8944 & n8947;
  assign n8949 = n8925 & n8948;
  assign n8950 = n8922 & n8949;
  assign n8951 = ~pi2763 & ~n8950;
  assign n8952 = pi2012 & pi2763;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = pi2480 & ~n8953;
  assign n8955 = ~pi2480 & n8953;
  assign n8956 = ~n8954 & ~n8955;
  assign n8957 = pi1221 & n8705;
  assign n8958 = pi1207 & n8709;
  assign n8959 = ~n8957 & ~n8958;
  assign n8960 = pi1291 & n8714;
  assign n8961 = pi1193 & n8717;
  assign n8962 = ~n8960 & ~n8961;
  assign n8963 = pi1305 & n8721;
  assign n8964 = pi1109 & n8724;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = pi1151 & n8728;
  assign n8967 = pi1263 & n8731;
  assign n8968 = ~n8966 & ~n8967;
  assign n8969 = pi1179 & n8736;
  assign n8970 = pi1137 & n8739;
  assign n8971 = ~n8969 & ~n8970;
  assign n8972 = pi1319 & n8743;
  assign n8973 = pi1235 & n8745;
  assign n8974 = ~n8972 & ~n8973;
  assign n8975 = n8971 & n8974;
  assign n8976 = n8968 & n8975;
  assign n8977 = n8965 & n8976;
  assign n8978 = pi1277 & n8752;
  assign n8979 = pi1123 & n8754;
  assign n8980 = ~n8978 & ~n8979;
  assign n8981 = n8977 & n8980;
  assign n8982 = pi1165 & n8758;
  assign n8983 = pi1249 & n8760;
  assign n8984 = ~n8982 & ~n8983;
  assign n8985 = n8981 & n8984;
  assign n8986 = n8962 & n8985;
  assign n8987 = n8959 & n8986;
  assign n8988 = ~pi2763 & ~n8987;
  assign n8989 = pi2374 & pi2763;
  assign n8990 = ~n8988 & ~n8989;
  assign n8991 = pi2478 & ~n8990;
  assign n8992 = ~pi2478 & n8990;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = ~n8956 & ~n8993;
  assign n8995 = ~n8919 & n8994;
  assign n8996 = ~n8882 & n8995;
  assign n8997 = pi2016 & pi2763;
  assign n8998 = pi1315 & n8721;
  assign n8999 = pi1119 & n8724;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = pi1161 & n8728;
  assign n9002 = pi1273 & n8731;
  assign n9003 = ~n9001 & ~n9002;
  assign n9004 = pi1231 & n8705;
  assign n9005 = pi1217 & n8709;
  assign n9006 = ~n9004 & ~n9005;
  assign n9007 = pi1301 & n8714;
  assign n9008 = pi1203 & n8717;
  assign n9009 = ~n9007 & ~n9008;
  assign n9010 = pi1287 & n8752;
  assign n9011 = pi1133 & n8754;
  assign n9012 = ~n9010 & ~n9011;
  assign n9013 = pi1175 & n8758;
  assign n9014 = pi1259 & n8760;
  assign n9015 = ~n9013 & ~n9014;
  assign n9016 = n9012 & n9015;
  assign n9017 = n9009 & n9016;
  assign n9018 = n9006 & n9017;
  assign n9019 = pi1189 & n8736;
  assign n9020 = pi1147 & n8739;
  assign n9021 = ~n9019 & ~n9020;
  assign n9022 = n9018 & n9021;
  assign n9023 = pi1329 & n8743;
  assign n9024 = pi1245 & n8745;
  assign n9025 = ~n9023 & ~n9024;
  assign n9026 = n9022 & n9025;
  assign n9027 = n9003 & n9026;
  assign n9028 = n9000 & n9027;
  assign n9029 = ~pi2763 & ~n9028;
  assign n9030 = ~n8997 & ~n9029;
  assign n9031 = ~pi2516 & ~n9030;
  assign n9032 = pi2516 & n9030;
  assign n9033 = ~n9031 & ~n9032;
  assign n9034 = n8996 & n9033;
  assign n9035 = pi1309 & n8721;
  assign n9036 = pi1113 & n8724;
  assign n9037 = ~n9035 & ~n9036;
  assign n9038 = pi1155 & n8728;
  assign n9039 = pi1267 & n8731;
  assign n9040 = ~n9038 & ~n9039;
  assign n9041 = pi1225 & n8705;
  assign n9042 = pi1211 & n8709;
  assign n9043 = ~n9041 & ~n9042;
  assign n9044 = pi1295 & n8714;
  assign n9045 = pi1197 & n8717;
  assign n9046 = ~n9044 & ~n9045;
  assign n9047 = pi1281 & n8752;
  assign n9048 = pi1127 & n8754;
  assign n9049 = ~n9047 & ~n9048;
  assign n9050 = pi1169 & n8758;
  assign n9051 = pi1253 & n8760;
  assign n9052 = ~n9050 & ~n9051;
  assign n9053 = n9049 & n9052;
  assign n9054 = n9046 & n9053;
  assign n9055 = n9043 & n9054;
  assign n9056 = pi1183 & n8736;
  assign n9057 = pi1141 & n8739;
  assign n9058 = ~n9056 & ~n9057;
  assign n9059 = n9055 & n9058;
  assign n9060 = pi1323 & n8743;
  assign n9061 = pi1239 & n8745;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = n9059 & n9062;
  assign n9064 = n9040 & n9063;
  assign n9065 = n9037 & n9064;
  assign n9066 = ~pi2763 & ~n9065;
  assign n9067 = pi2014 & pi2763;
  assign n9068 = ~n9066 & ~n9067;
  assign n9069 = pi2482 & ~n9068;
  assign n9070 = ~pi2482 & n9068;
  assign n9071 = ~n9069 & ~n9070;
  assign n9072 = n9034 & ~n9071;
  assign n9073 = ~n8845 & n9072;
  assign n9074 = ~n8808 & n9073;
  assign n9075 = pi1302 & n8721;
  assign n9076 = pi1106 & n8724;
  assign n9077 = ~n9075 & ~n9076;
  assign n9078 = pi1148 & n8728;
  assign n9079 = pi1260 & n8731;
  assign n9080 = ~n9078 & ~n9079;
  assign n9081 = pi1218 & n8705;
  assign n9082 = pi1204 & n8709;
  assign n9083 = ~n9081 & ~n9082;
  assign n9084 = pi1288 & n8714;
  assign n9085 = pi1190 & n8717;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = pi1274 & n8752;
  assign n9088 = pi1120 & n8754;
  assign n9089 = ~n9087 & ~n9088;
  assign n9090 = pi1162 & n8758;
  assign n9091 = pi1246 & n8760;
  assign n9092 = ~n9090 & ~n9091;
  assign n9093 = n9089 & n9092;
  assign n9094 = n9086 & n9093;
  assign n9095 = n9083 & n9094;
  assign n9096 = pi1316 & n8743;
  assign n9097 = pi1232 & n8745;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = n9095 & n9098;
  assign n9100 = pi1176 & n8736;
  assign n9101 = pi1134 & n8739;
  assign n9102 = ~n9100 & ~n9101;
  assign n9103 = n9099 & n9102;
  assign n9104 = n9080 & n9103;
  assign n9105 = n9077 & n9104;
  assign n9106 = ~pi2763 & ~n9105;
  assign n9107 = pi2392 & pi2763;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = pi2475 & ~n9108;
  assign n9110 = ~pi2475 & n9108;
  assign n9111 = ~n9109 & ~n9110;
  assign n9112 = pi1303 & n8721;
  assign n9113 = pi1107 & n8724;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = pi1149 & n8728;
  assign n9116 = pi1261 & n8731;
  assign n9117 = ~n9115 & ~n9116;
  assign n9118 = pi1289 & n8714;
  assign n9119 = pi1191 & n8717;
  assign n9120 = ~n9118 & ~n9119;
  assign n9121 = pi1219 & n8705;
  assign n9122 = pi1205 & n8709;
  assign n9123 = ~n9121 & ~n9122;
  assign n9124 = pi1275 & n8752;
  assign n9125 = pi1121 & n8754;
  assign n9126 = ~n9124 & ~n9125;
  assign n9127 = pi1163 & n8758;
  assign n9128 = pi1247 & n8760;
  assign n9129 = ~n9127 & ~n9128;
  assign n9130 = n9126 & n9129;
  assign n9131 = n9123 & n9130;
  assign n9132 = n9120 & n9131;
  assign n9133 = pi1177 & n8736;
  assign n9134 = pi1135 & n8739;
  assign n9135 = ~n9133 & ~n9134;
  assign n9136 = n9132 & n9135;
  assign n9137 = pi1317 & n8743;
  assign n9138 = pi1233 & n8745;
  assign n9139 = ~n9137 & ~n9138;
  assign n9140 = n9136 & n9139;
  assign n9141 = n9117 & n9140;
  assign n9142 = n9114 & n9141;
  assign n9143 = ~pi2763 & ~n9142;
  assign n9144 = pi2373 & pi2763;
  assign n9145 = ~n9143 & ~n9144;
  assign n9146 = pi2476 & ~n9145;
  assign n9147 = ~pi2476 & n9145;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = pi1314 & n8721;
  assign n9150 = pi1118 & n8724;
  assign n9151 = ~n9149 & ~n9150;
  assign n9152 = pi1160 & n8728;
  assign n9153 = pi1272 & n8731;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = pi1230 & n8705;
  assign n9156 = pi1216 & n8709;
  assign n9157 = ~n9155 & ~n9156;
  assign n9158 = pi1300 & n8714;
  assign n9159 = pi1202 & n8717;
  assign n9160 = ~n9158 & ~n9159;
  assign n9161 = pi1286 & n8752;
  assign n9162 = pi1132 & n8754;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = pi1174 & n8758;
  assign n9165 = pi1258 & n8760;
  assign n9166 = ~n9164 & ~n9165;
  assign n9167 = n9163 & n9166;
  assign n9168 = n9160 & n9167;
  assign n9169 = n9157 & n9168;
  assign n9170 = pi1188 & n8736;
  assign n9171 = pi1146 & n8739;
  assign n9172 = ~n9170 & ~n9171;
  assign n9173 = n9169 & n9172;
  assign n9174 = pi1328 & n8743;
  assign n9175 = pi1244 & n8745;
  assign n9176 = ~n9174 & ~n9175;
  assign n9177 = n9173 & n9176;
  assign n9178 = n9154 & n9177;
  assign n9179 = n9151 & n9178;
  assign n9180 = ~pi2763 & ~n9179;
  assign n9181 = pi2378 & pi2763;
  assign n9182 = ~n9180 & ~n9181;
  assign n9183 = pi2517 & ~n9182;
  assign n9184 = ~pi2517 & n9182;
  assign n9185 = ~n9183 & ~n9184;
  assign n9186 = pi1313 & n8721;
  assign n9187 = pi1117 & n8724;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = pi1159 & n8728;
  assign n9190 = pi1271 & n8731;
  assign n9191 = ~n9189 & ~n9190;
  assign n9192 = pi1229 & n8705;
  assign n9193 = pi1215 & n8709;
  assign n9194 = ~n9192 & ~n9193;
  assign n9195 = pi1299 & n8714;
  assign n9196 = pi1201 & n8717;
  assign n9197 = ~n9195 & ~n9196;
  assign n9198 = pi1285 & n8752;
  assign n9199 = pi1131 & n8754;
  assign n9200 = ~n9198 & ~n9199;
  assign n9201 = pi1257 & n8760;
  assign n9202 = pi1173 & n8758;
  assign n9203 = ~n9201 & ~n9202;
  assign n9204 = n9200 & n9203;
  assign n9205 = n9197 & n9204;
  assign n9206 = n9194 & n9205;
  assign n9207 = pi1327 & n8743;
  assign n9208 = pi1243 & n8745;
  assign n9209 = ~n9207 & ~n9208;
  assign n9210 = n9206 & n9209;
  assign n9211 = pi1187 & n8736;
  assign n9212 = pi1145 & n8739;
  assign n9213 = ~n9211 & ~n9212;
  assign n9214 = n9210 & n9213;
  assign n9215 = n9191 & n9214;
  assign n9216 = n9188 & n9215;
  assign n9217 = ~pi2763 & ~n9216;
  assign n9218 = pi2377 & pi2763;
  assign n9219 = ~n9217 & ~n9218;
  assign n9220 = pi2518 & ~n9219;
  assign n9221 = ~pi2518 & n9219;
  assign n9222 = ~n9220 & ~n9221;
  assign n9223 = ~n9185 & ~n9222;
  assign n9224 = ~n9148 & n9223;
  assign n9225 = ~n9111 & n9224;
  assign n9226 = n9074 & n9225;
  assign n9227 = pi1312 & n8721;
  assign n9228 = pi1116 & n8724;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = pi1158 & n8728;
  assign n9231 = pi1270 & n8731;
  assign n9232 = ~n9230 & ~n9231;
  assign n9233 = pi1228 & n8705;
  assign n9234 = pi1214 & n8709;
  assign n9235 = ~n9233 & ~n9234;
  assign n9236 = pi1298 & n8714;
  assign n9237 = pi1200 & n8717;
  assign n9238 = ~n9236 & ~n9237;
  assign n9239 = pi1284 & n8752;
  assign n9240 = pi1130 & n8754;
  assign n9241 = ~n9239 & ~n9240;
  assign n9242 = pi1172 & n8758;
  assign n9243 = pi1256 & n8760;
  assign n9244 = ~n9242 & ~n9243;
  assign n9245 = n9241 & n9244;
  assign n9246 = n9238 & n9245;
  assign n9247 = n9235 & n9246;
  assign n9248 = pi1186 & n8736;
  assign n9249 = pi1144 & n8739;
  assign n9250 = ~n9248 & ~n9249;
  assign n9251 = n9247 & n9250;
  assign n9252 = pi1326 & n8743;
  assign n9253 = pi1242 & n8745;
  assign n9254 = ~n9252 & ~n9253;
  assign n9255 = n9251 & n9254;
  assign n9256 = n9232 & n9255;
  assign n9257 = n9229 & n9256;
  assign n9258 = ~pi2763 & ~n9257;
  assign n9259 = pi2376 & pi2763;
  assign n9260 = ~n9258 & ~n9259;
  assign n9261 = ~pi2485 & n9260;
  assign n9262 = pi2485 & ~n9260;
  assign n9263 = ~n9261 & ~n9262;
  assign n9264 = n9226 & ~n9263;
  assign n9265 = ~n8771 & n9264;
  assign n9266 = ~pi3190 & pi3291;
  assign n9267 = ~pi2489 & n9266;
  assign n9268 = ~n9265 & n9267;
  assign n9269 = ~n8702 & ~n9268;
  assign n9270 = pi2490 & ~n9265;
  assign n9271 = ~pi3210 & ~n9270;
  assign n9272 = n9269 & n9271;
  assign n9273 = n8698 & ~n9272;
  assign n9274 = ~n8702 & ~n9270;
  assign n9275 = ~pi3210 & n9274;
  assign n9276 = ~n9267 & n9275;
  assign n9277 = ~n8698 & ~n9276;
  assign n9278 = ~n9273 & ~n9277;
  assign n9279 = ~n8670 & ~n9278;
  assign n9280 = ~n8699 & ~n9266;
  assign n9281 = ~n8698 & ~n9280;
  assign n9282 = ~pi2485 & n9257;
  assign n9283 = pi2485 & ~n9257;
  assign n9284 = ~n9282 & ~n9283;
  assign n9285 = ~pi2482 & n9065;
  assign n9286 = pi2482 & ~n9065;
  assign n9287 = ~n9285 & ~n9286;
  assign n9288 = ~pi2483 & n8802;
  assign n9289 = pi2483 & ~n8802;
  assign n9290 = ~n9288 & ~n9289;
  assign n9291 = ~pi2480 & n8950;
  assign n9292 = pi2480 & ~n8950;
  assign n9293 = ~n9291 & ~n9292;
  assign n9294 = ~pi2477 & n8913;
  assign n9295 = pi2477 & ~n8913;
  assign n9296 = ~n9294 & ~n9295;
  assign n9297 = ~pi2479 & n8876;
  assign n9298 = pi2479 & ~n8876;
  assign n9299 = ~n9297 & ~n9298;
  assign n9300 = ~pi2478 & n8987;
  assign n9301 = pi2478 & ~n8987;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = ~n9299 & ~n9302;
  assign n9304 = ~n9296 & n9303;
  assign n9305 = ~n9293 & n9304;
  assign n9306 = pi2481 & n8839;
  assign n9307 = ~pi2481 & ~n8839;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = n9305 & n9308;
  assign n9310 = ~pi2516 & n9028;
  assign n9311 = pi2516 & ~n9028;
  assign n9312 = ~n9310 & ~n9311;
  assign n9313 = n9309 & ~n9312;
  assign n9314 = ~n9290 & n9313;
  assign n9315 = ~n9287 & n9314;
  assign n9316 = ~pi2476 & n9142;
  assign n9317 = pi2476 & ~n9142;
  assign n9318 = ~n9316 & ~n9317;
  assign n9319 = ~pi2517 & n9179;
  assign n9320 = pi2517 & ~n9179;
  assign n9321 = ~n9319 & ~n9320;
  assign n9322 = ~pi2518 & n9216;
  assign n9323 = pi2518 & ~n9216;
  assign n9324 = ~n9322 & ~n9323;
  assign n9325 = ~pi2475 & n9105;
  assign n9326 = pi2475 & ~n9105;
  assign n9327 = ~n9325 & ~n9326;
  assign n9328 = ~n9324 & ~n9327;
  assign n9329 = ~n9321 & n9328;
  assign n9330 = ~n9318 & n9329;
  assign n9331 = n9315 & n9330;
  assign n9332 = ~pi2484 & n8765;
  assign n9333 = pi2484 & ~n8765;
  assign n9334 = ~n9332 & ~n9333;
  assign n9335 = n9331 & ~n9334;
  assign n9336 = ~n9284 & n9335;
  assign n9337 = n9266 & ~n9336;
  assign n9338 = ~n8699 & ~n9337;
  assign n9339 = n8698 & ~n9338;
  assign n9340 = ~n9281 & ~n9339;
  assign n9341 = n8670 & ~n9340;
  assign n9342 = ~n9279 & ~n9341;
  assign n9343 = ~pi3408 & n9342;
  assign n9344 = ~pi0540 & n9343;
  assign n9345 = ~pi3371 & n9344;
  assign n9346 = ~po3841 & n9345;
  assign n9347 = n8624 & n9346;
  assign n9348 = ~n8621 & n9347;
  assign n9349 = pi3256 & n8561;
  assign n9350 = ~n9348 & ~n9349;
  assign n9351 = ~n8606 & n9350;
  assign n9352 = ~pi3551 & ~po3946;
  assign n9353 = n8622 & ~n9352;
  assign n9354 = ~po3841 & n9353;
  assign n9355 = pi3370 & n9352;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = n9351 & n9356;
  assign n9358 = ~pi3395 & ~pi3429;
  assign n9359 = ~pi3427 & n9358;
  assign n9360 = ~pi3424 & n9359;
  assign n9361 = ~pi2382 & n9360;
  assign n9362 = pi3436 & pi3451;
  assign n9363 = ~pi3435 & ~n9360;
  assign n9364 = n9362 & n9363;
  assign n9365 = ~pi3426 & ~n9352;
  assign n9366 = pi3367 & ~pi3426;
  assign n9367 = ~pi3391 & n9360;
  assign n9368 = pi2382 & n9367;
  assign n9369 = n9366 & n9368;
  assign n9370 = ~pi0994 & ~n9369;
  assign n9371 = n9365 & ~n9370;
  assign n9372 = ~n9364 & ~n9371;
  assign n9373 = ~pi0418 & n8609;
  assign n9374 = pi0419 & ~pi0421;
  assign n9375 = n9373 & n9374;
  assign n9376 = ~pi0405 & n9375;
  assign n9377 = pi0420 & n9376;
  assign n9378 = ~n8615 & ~n9377;
  assign n9379 = ~pi0415 & n9378;
  assign n9380 = ~pi0412 & ~n9378;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = pi0414 & n9378;
  assign n9383 = pi0411 & ~n9378;
  assign n9384 = ~n9382 & ~n9383;
  assign n9385 = n9381 & n9384;
  assign n9386 = ~n9372 & n9385;
  assign n9387 = pi3435 & ~n9360;
  assign n9388 = n9362 & n9387;
  assign n9389 = pi3391 & n9360;
  assign n9390 = pi2382 & n9389;
  assign n9391 = n9366 & n9390;
  assign n9392 = ~pi0992 & ~n9391;
  assign n9393 = n9365 & ~n9392;
  assign n9394 = ~n9388 & ~n9393;
  assign n9395 = n9381 & ~n9384;
  assign n9396 = ~n9394 & n9395;
  assign n9397 = ~n9386 & ~n9396;
  assign n9398 = ~pi3367 & ~pi3426;
  assign n9399 = n9368 & n9398;
  assign n9400 = ~pi0995 & ~n9399;
  assign n9401 = n9365 & ~n9400;
  assign n9402 = ~pi3436 & pi3451;
  assign n9403 = n9363 & n9402;
  assign n9404 = ~n9401 & ~n9403;
  assign n9405 = ~n9381 & n9384;
  assign n9406 = ~n9404 & n9405;
  assign n9407 = n9387 & n9402;
  assign n9408 = n9390 & n9398;
  assign n9409 = ~pi0993 & ~n9408;
  assign n9410 = n9365 & ~n9409;
  assign n9411 = ~n9407 & ~n9410;
  assign n9412 = ~n9381 & ~n9384;
  assign n9413 = ~n9411 & n9412;
  assign n9414 = ~n9406 & ~n9413;
  assign n9415 = n9397 & n9414;
  assign n9416 = n8624 & ~po3841;
  assign n9417 = ~n9415 & n9416;
  assign n9418 = ~n8573 & n8574;
  assign n9419 = n8570 & n9418;
  assign n9420 = n8570 & n8573;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n8568 & n8569;
  assign n9423 = ~n8568 & ~n9422;
  assign n9424 = n9421 & n9423;
  assign n9425 = ~pi3416 & n8562;
  assign n9426 = ~n9424 & ~n9425;
  assign n9427 = pi1441 & n9422;
  assign n9428 = pi1436 & n8568;
  assign n9429 = ~n9427 & ~n9428;
  assign n9430 = pi1732 & n9419;
  assign n9431 = pi1727 & n9420;
  assign n9432 = ~n9430 & ~n9431;
  assign n9433 = n9429 & n9432;
  assign n9434 = pi1440 & n9422;
  assign n9435 = pi1446 & n8568;
  assign n9436 = ~n9434 & ~n9435;
  assign n9437 = pi1731 & n9419;
  assign n9438 = pi1737 & n9420;
  assign n9439 = ~n9437 & ~n9438;
  assign n9440 = n9436 & n9439;
  assign n9441 = pi1439 & n9422;
  assign n9442 = pi1445 & n8568;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = pi1730 & n9419;
  assign n9445 = pi1736 & n9420;
  assign n9446 = ~n9444 & ~n9445;
  assign n9447 = n9443 & n9446;
  assign n9448 = n9440 & ~n9447;
  assign n9449 = ~n9433 & n9448;
  assign n9450 = ~n9372 & n9449;
  assign n9451 = ~n9440 & ~n9447;
  assign n9452 = ~n9433 & n9451;
  assign n9453 = ~n9394 & n9452;
  assign n9454 = ~n9450 & ~n9453;
  assign n9455 = n9433 & n9448;
  assign n9456 = ~n9404 & n9455;
  assign n9457 = n9433 & n9451;
  assign n9458 = ~n9411 & n9457;
  assign n9459 = ~n9456 & ~n9458;
  assign n9460 = n9454 & n9459;
  assign n9461 = n9426 & ~n9460;
  assign n9462 = ~n9416 & n9461;
  assign n9463 = ~n9417 & ~n9462;
  assign n9464 = n9361 & ~n9463;
  assign n9465 = ~pi3359 & ~pi3363;
  assign n9466 = ~pi3364 & ~pi3385;
  assign n9467 = n9465 & n9466;
  assign n9468 = ~pi3386 & ~pi3387;
  assign n9469 = n9467 & n9468;
  assign n9470 = ~pi3365 & ~pi3388;
  assign n9471 = ~pi3399 & n9470;
  assign n9472 = n9469 & n9471;
  assign n9473 = pi3412 & pi3481;
  assign po3871 = ~pi3515 & n9473;
  assign n9475 = pi0650 & ~po3871;
  assign n9476 = pi1331 & ~n8765;
  assign n9477 = pi3233 & pi3519;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = pi3329 & pi3519;
  assign n9480 = pi0573 & pi1359;
  assign n9481 = pi0378 & pi1057;
  assign n9482 = ~n9480 & ~n9481;
  assign n9483 = ~n9479 & n9482;
  assign n9484 = n9478 & n9483;
  assign n9485 = n9475 & ~n9484;
  assign n9486 = pi0524 & ~po3871;
  assign n9487 = ~pi0979 & pi2613;
  assign n9488 = pi0979 & pi2607;
  assign n9489 = ~n9487 & ~n9488;
  assign n9490 = pi0763 & ~n9489;
  assign n9491 = ~pi0979 & pi2626;
  assign n9492 = pi0979 & pi2620;
  assign n9493 = ~n9491 & ~n9492;
  assign n9494 = pi0764 & ~n9493;
  assign n9495 = ~n9490 & ~n9494;
  assign n9496 = pi0053 & ~pi0979;
  assign n9497 = pi0051 & pi0979;
  assign n9498 = ~n9496 & ~n9497;
  assign n9499 = pi0719 & ~n9498;
  assign n9500 = ~pi0979 & pi2640;
  assign n9501 = pi0979 & pi3173;
  assign n9502 = ~n9500 & ~n9501;
  assign n9503 = pi0765 & ~n9502;
  assign n9504 = ~pi0979 & pi2969;
  assign n9505 = pi0979 & pi3119;
  assign n9506 = ~n9504 & ~n9505;
  assign n9507 = pi0766 & ~n9506;
  assign n9508 = ~n9503 & ~n9507;
  assign n9509 = pi0118 & ~pi0979;
  assign n9510 = pi0116 & pi0979;
  assign n9511 = ~n9509 & ~n9510;
  assign n9512 = pi0720 & ~n9511;
  assign n9513 = pi0229 & ~pi0979;
  assign n9514 = pi0228 & pi0979;
  assign n9515 = ~n9513 & ~n9514;
  assign n9516 = pi0721 & ~n9515;
  assign n9517 = ~n9512 & ~n9516;
  assign n9518 = n9508 & n9517;
  assign n9519 = ~n9499 & n9518;
  assign n9520 = n9495 & n9519;
  assign n9521 = n9486 & ~n9520;
  assign n9522 = ~n9485 & ~n9521;
  assign n9523 = pi0538 & ~po3871;
  assign n9524 = ~pi0979 & pi2852;
  assign n9525 = pi0979 & pi2135;
  assign n9526 = ~n9524 & ~n9525;
  assign n9527 = pi0717 & ~n9526;
  assign n9528 = pi0486 & ~pi0979;
  assign n9529 = pi0483 & pi0979;
  assign n9530 = ~n9528 & ~n9529;
  assign n9531 = pi0718 & ~n9530;
  assign n9532 = pi0203 & ~pi0979;
  assign n9533 = pi0199 & pi0979;
  assign n9534 = ~n9532 & ~n9533;
  assign n9535 = pi1599 & ~n9534;
  assign n9536 = pi0265 & ~pi0979;
  assign n9537 = pi0261 & pi0979;
  assign n9538 = ~n9536 & ~n9537;
  assign n9539 = pi0716 & ~n9538;
  assign n9540 = pi0310 & ~pi0979;
  assign n9541 = pi0308 & pi0979;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = pi0761 & ~n9542;
  assign n9544 = ~n9539 & ~n9543;
  assign n9545 = ~n9535 & n9544;
  assign n9546 = ~n9531 & n9545;
  assign n9547 = ~n9527 & n9546;
  assign n9548 = n9523 & ~n9547;
  assign n9549 = pi0576 & ~po3871;
  assign n9550 = pi0979 & pi2154;
  assign n9551 = ~pi0979 & pi2926;
  assign n9552 = ~n9550 & ~n9551;
  assign n9553 = pi0767 & ~n9552;
  assign n9554 = ~pi0979 & pi2429;
  assign n9555 = pi0979 & pi1964;
  assign n9556 = ~n9554 & ~n9555;
  assign n9557 = pi0768 & ~n9556;
  assign n9558 = ~n9553 & ~n9557;
  assign n9559 = pi0979 & pi2172;
  assign n9560 = ~pi0979 & pi2936;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = pi0836 & ~n9561;
  assign n9563 = ~pi0979 & pi2948;
  assign n9564 = pi0979 & pi2188;
  assign n9565 = ~n9563 & ~n9564;
  assign n9566 = pi0837 & ~n9565;
  assign n9567 = ~n9562 & ~n9566;
  assign n9568 = pi0178 & ~pi0979;
  assign n9569 = pi0163 & pi0979;
  assign n9570 = ~n9568 & ~n9569;
  assign n9571 = pi0838 & ~n9570;
  assign n9572 = n9567 & ~n9571;
  assign n9573 = n9558 & n9572;
  assign n9574 = n9549 & ~n9573;
  assign n9575 = ~n9548 & ~n9574;
  assign n9576 = n9522 & n9575;
  assign n9577 = pi0722 & ~po3871;
  assign n9578 = pi1351 & pi2268;
  assign n9579 = pi1352 & pi2445;
  assign n9580 = ~n9578 & ~n9579;
  assign n9581 = pi1353 & pi1983;
  assign n9582 = n9580 & ~n9581;
  assign n9583 = pi1345 & pi2656;
  assign n9584 = n9582 & ~n9583;
  assign n9585 = pi1348 & pi2694;
  assign n9586 = pi1350 & pi2435;
  assign n9587 = ~n9585 & ~n9586;
  assign n9588 = pi1600 & pi2210;
  assign n9589 = pi1338 & pi2238;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = pi1339 & pi2252;
  assign n9592 = pi1337 & pi2224;
  assign n9593 = ~n9591 & ~n9592;
  assign n9594 = n9590 & n9593;
  assign n9595 = pi1346 & pi2670;
  assign n9596 = pi1347 & pi2684;
  assign n9597 = ~n9595 & ~n9596;
  assign n9598 = n9594 & n9597;
  assign n9599 = n9587 & n9598;
  assign n9600 = n9584 & n9599;
  assign n9601 = n9577 & ~n9600;
  assign n9602 = n9576 & ~n9601;
  assign n9603 = pi1032 & ~pi1033;
  assign n9604 = pi1012 & pi1034;
  assign n9605 = pi1039 & pi2112;
  assign n9606 = n9604 & n9605;
  assign n9607 = n9603 & n9606;
  assign n9608 = ~pi0796 & pi0962;
  assign n9609 = pi0796 & pi1845;
  assign n9610 = ~n9608 & ~n9609;
  assign n9611 = n9607 & ~n9610;
  assign n9612 = ~pi1039 & pi2112;
  assign n9613 = n9604 & n9612;
  assign n9614 = n9603 & n9613;
  assign n9615 = pi0960 & n9614;
  assign n9616 = ~pi1012 & pi1034;
  assign n9617 = n9605 & n9616;
  assign n9618 = n9603 & n9617;
  assign n9619 = pi1905 & n9618;
  assign n9620 = ~n9615 & ~n9619;
  assign n9621 = pi1032 & pi1033;
  assign n9622 = n9606 & n9621;
  assign n9623 = pi1930 & n9622;
  assign n9624 = pi1033 & ~pi1034;
  assign n9625 = ~pi1012 & n9624;
  assign n9626 = ~pi1032 & pi2112;
  assign n9627 = ~pi1039 & n9626;
  assign n9628 = n9625 & n9627;
  assign n9629 = pi2101 & n9628;
  assign n9630 = ~pi1032 & ~pi1033;
  assign n9631 = n9617 & n9630;
  assign n9632 = pi0974 & n9631;
  assign n9633 = ~n9629 & ~n9632;
  assign n9634 = pi1030 & pi1031;
  assign n9635 = ~pi1032 & n9634;
  assign n9636 = pi1013 & n9635;
  assign n9637 = pi1028 & pi1029;
  assign n9638 = pi1037 & n9637;
  assign n9639 = pi1038 & n9638;
  assign n9640 = pi1035 & pi1036;
  assign n9641 = n9639 & n9640;
  assign n9642 = pi1012 & pi1039;
  assign n9643 = ~pi1034 & n9642;
  assign n9644 = ~pi1033 & n9643;
  assign n9645 = n9641 & n9644;
  assign n9646 = n9636 & n9645;
  assign n9647 = pi2112 & n9646;
  assign n9648 = pi2988 & n9647;
  assign n9649 = ~pi1012 & ~pi1039;
  assign n9650 = ~pi1033 & n9649;
  assign n9651 = pi1034 & n9650;
  assign n9652 = n9641 & n9651;
  assign n9653 = n9636 & n9652;
  assign n9654 = pi2112 & n9653;
  assign n9655 = pi0687 & n9654;
  assign n9656 = ~n9648 & ~n9655;
  assign n9657 = n9613 & n9630;
  assign n9658 = pi1761 & n9657;
  assign n9659 = n9606 & n9630;
  assign n9660 = pi1749 & n9659;
  assign n9661 = ~n9658 & ~n9660;
  assign n9662 = n9656 & n9661;
  assign n9663 = n9633 & n9662;
  assign n9664 = ~n9623 & n9663;
  assign n9665 = ~pi1012 & pi1039;
  assign n9666 = ~pi1033 & ~pi1034;
  assign n9667 = n9665 & n9666;
  assign n9668 = n9641 & n9667;
  assign n9669 = n9636 & n9668;
  assign n9670 = pi2112 & n9669;
  assign n9671 = pi0752 & n9670;
  assign n9672 = ~pi1039 & n9666;
  assign n9673 = pi1012 & n9672;
  assign n9674 = n9641 & n9673;
  assign n9675 = n9636 & n9674;
  assign n9676 = pi2112 & n9675;
  assign n9677 = pi0929 & n9676;
  assign n9678 = ~n9671 & ~n9677;
  assign n9679 = n9617 & n9621;
  assign n9680 = pi1879 & n9679;
  assign n9681 = n9612 & n9616;
  assign n9682 = n9621 & n9681;
  assign n9683 = pi0277 & n9682;
  assign n9684 = ~n9680 & ~n9683;
  assign n9685 = n9678 & n9684;
  assign n9686 = n9664 & n9685;
  assign n9687 = n9603 & n9681;
  assign n9688 = pi0981 & n9687;
  assign n9689 = pi1012 & ~pi1034;
  assign n9690 = n9605 & n9689;
  assign n9691 = n9603 & n9690;
  assign n9692 = pi2100 & n9691;
  assign n9693 = ~n9688 & ~n9692;
  assign n9694 = n9686 & n9693;
  assign n9695 = n9620 & n9694;
  assign n9696 = ~n9611 & n9695;
  assign n9697 = n9612 & n9689;
  assign n9698 = n9621 & n9697;
  assign n9699 = pi1836 & n9698;
  assign n9700 = ~pi1012 & ~pi1034;
  assign n9701 = n9612 & n9700;
  assign n9702 = n9621 & n9701;
  assign n9703 = ~pi0890 & pi0947;
  assign n9704 = pi0890 & pi1843;
  assign n9705 = ~n9703 & ~n9704;
  assign n9706 = n9702 & ~n9705;
  assign n9707 = n9603 & n9701;
  assign n9708 = pi0870 & n9707;
  assign n9709 = ~n9706 & ~n9708;
  assign n9710 = n9630 & n9701;
  assign n9711 = pi0909 & n9710;
  assign n9712 = n9613 & n9621;
  assign n9713 = pi1782 & n9712;
  assign n9714 = ~n9711 & ~n9713;
  assign n9715 = n9603 & n9697;
  assign n9716 = pi0888 & n9715;
  assign n9717 = n9605 & n9700;
  assign n9718 = n9603 & n9717;
  assign n9719 = pi1890 & n9718;
  assign n9720 = ~n9716 & ~n9719;
  assign n9721 = n9714 & n9720;
  assign n9722 = n9709 & n9721;
  assign n9723 = ~n9699 & n9722;
  assign n9724 = n9696 & n9723;
  assign n9725 = pi1934 & ~n9724;
  assign n9726 = pi0762 & ~po3871;
  assign n9727 = pi0606 & pi1336;
  assign n9728 = pi1333 & pi1743;
  assign n9729 = ~n9727 & ~n9728;
  assign n9730 = pi1332 & pi2578;
  assign n9731 = pi1335 & pi2593;
  assign n9732 = ~n9730 & ~n9731;
  assign n9733 = n9729 & n9732;
  assign n9734 = n9726 & ~n9733;
  assign n9735 = ~n9725 & ~n9734;
  assign n9736 = pi0539 & ~po3871;
  assign n9737 = pi1355 & pi2458;
  assign n9738 = pi1356 & pi2530;
  assign n9739 = ~n9737 & ~n9738;
  assign n9740 = pi1357 & pi2410;
  assign n9741 = n9739 & ~n9740;
  assign n9742 = pi1054 & pi2716;
  assign n9743 = n9741 & ~n9742;
  assign n9744 = pi1056 & pi2744;
  assign n9745 = pi1354 & pi2748;
  assign n9746 = ~n9744 & ~n9745;
  assign n9747 = pi1340 & pi2287;
  assign n9748 = pi1342 & pi2309;
  assign n9749 = ~n9747 & ~n9748;
  assign n9750 = pi1343 & pi2323;
  assign n9751 = pi1341 & pi2300;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = n9749 & n9752;
  assign n9754 = pi1055 & pi2774;
  assign n9755 = pi1349 & pi2561;
  assign n9756 = ~n9754 & ~n9755;
  assign n9757 = n9753 & n9756;
  assign n9758 = n9746 & n9757;
  assign n9759 = n9743 & n9758;
  assign n9760 = n9736 & ~n9759;
  assign n9761 = n9735 & ~n9760;
  assign n9762 = n9602 & n9761;
  assign n9763 = pi3358 & po3871;
  assign n9764 = n9762 & ~n9763;
  assign n9765 = ~pi1787 & ~n9764;
  assign n9766 = pi1787 & pi2817;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = n9472 & ~n9767;
  assign n9769 = ~pi3387 & n9467;
  assign n9770 = pi3386 & n9471;
  assign n9771 = n9769 & n9770;
  assign n9772 = pi3387 & n9467;
  assign n9773 = ~pi3386 & n9471;
  assign n9774 = n9772 & n9773;
  assign n9775 = ~pi3388 & ~pi3399;
  assign n9776 = n9468 & n9775;
  assign n9777 = ~pi3365 & n9776;
  assign n9778 = ~pi3363 & ~pi3385;
  assign n9779 = n9777 & n9778;
  assign n9780 = pi3359 & ~pi3364;
  assign n9781 = n9779 & n9780;
  assign n9782 = pi3365 & n9776;
  assign n9783 = n9467 & n9782;
  assign n9784 = ~n9781 & ~n9783;
  assign n9785 = ~n9774 & n9784;
  assign n9786 = ~pi3359 & n9777;
  assign n9787 = pi3363 & n9786;
  assign n9788 = n9466 & n9787;
  assign n9789 = ~pi3363 & n9786;
  assign n9790 = ~pi3364 & pi3385;
  assign n9791 = n9789 & n9790;
  assign n9792 = pi3364 & n9778;
  assign n9793 = n9786 & n9792;
  assign n9794 = ~n9791 & ~n9793;
  assign n9795 = ~n9788 & n9794;
  assign n9796 = n9785 & n9795;
  assign n9797 = ~n9771 & n9796;
  assign n9798 = pi3399 & n9470;
  assign n9799 = n9469 & n9798;
  assign n9800 = ~pi3399 & n9469;
  assign n9801 = ~pi3365 & pi3388;
  assign n9802 = n9800 & n9801;
  assign n9803 = ~n9799 & ~n9802;
  assign n9804 = n9797 & n9803;
  assign n9805 = pi3872 & n9804;
  assign n9806 = pi3888 & n9774;
  assign n9807 = ~n9805 & ~n9806;
  assign n9808 = pi3856 & n9802;
  assign n9809 = pi3920 & n9781;
  assign n9810 = pi3904 & n9771;
  assign n9811 = ~n9809 & ~n9810;
  assign n9812 = pi3952 & n9791;
  assign n9813 = pi3936 & n9788;
  assign n9814 = ~n9812 & ~n9813;
  assign n9815 = n9811 & n9814;
  assign n9816 = ~n9808 & n9815;
  assign n9817 = n9807 & n9816;
  assign n9818 = pi3872 & n9799;
  assign n9819 = n9817 & ~n9818;
  assign n9820 = pi3984 & n9783;
  assign n9821 = pi3968 & n9793;
  assign n9822 = ~n9820 & ~n9821;
  assign n9823 = n9819 & n9822;
  assign n9824 = ~n9472 & ~n9823;
  assign n9825 = ~n9768 & ~n9824;
  assign n9826 = n9464 & ~n9825;
  assign n9827 = ~n9416 & ~n9426;
  assign n9828 = n9415 & n9416;
  assign n9829 = ~n9827 & ~n9828;
  assign n9830 = ~n9416 & ~n9461;
  assign n9831 = n9829 & n9830;
  assign n9832 = n9404 & n9455;
  assign n9833 = pi1983 & n9832;
  assign n9834 = n9372 & n9449;
  assign n9835 = pi2445 & n9834;
  assign n9836 = ~n9833 & ~n9835;
  assign n9837 = n9394 & n9452;
  assign n9838 = pi2435 & n9837;
  assign n9839 = n9411 & n9457;
  assign n9840 = pi2268 & n9839;
  assign n9841 = ~n9838 & ~n9840;
  assign n9842 = n9836 & n9841;
  assign n9843 = n9831 & ~n9842;
  assign n9844 = ~n9464 & n9843;
  assign n9845 = ~n9826 & ~n9844;
  assign n9846 = ~n9829 & n9830;
  assign n9847 = ~n9464 & n9846;
  assign n9848 = ~n8586 & ~n8599;
  assign n9849 = n8577 & ~n9848;
  assign n9850 = ~n8567 & n9849;
  assign n9851 = pi2558 & po3871;
  assign n9852 = ~pi1422 & ~n8565;
  assign n9853 = n8589 & n9852;
  assign n9854 = pi0909 & n9853;
  assign n9855 = ~n9851 & ~n9854;
  assign n9856 = pi0565 & n8540;
  assign n9857 = ~pi3452 & n9856;
  assign n9858 = ~pi2813 & pi3362;
  assign n9859 = ~pi0541 & pi0565;
  assign n9860 = n8536 & n9859;
  assign n9861 = pi0565 & pi3546;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = ~pi3215 & n8546;
  assign n9864 = n9859 & n9863;
  assign n9865 = pi0565 & pi3481;
  assign n9866 = ~n9864 & ~n9865;
  assign n9867 = n9862 & n9866;
  assign n9868 = ~n9858 & n9867;
  assign po3852 = n9857 | ~n9868;
  assign n9870 = ~pi3505 & ~pi3545;
  assign n9871 = n8534 & ~n9870;
  assign n9872 = pi3148 & n9871;
  assign n9873 = ~pi3589 & n8563;
  assign n9874 = pi3644 & n9873;
  assign n9875 = ~pi3362 & ~n9874;
  assign n9876 = pi3148 & ~n9875;
  assign n9877 = pi3452 & pi3526;
  assign n9878 = ~n9876 & ~n9877;
  assign po3874 = n9872 | ~n9878;
  assign n9880 = ~po3852 & ~po3874;
  assign n9881 = pi3215 & n8546;
  assign n9882 = n9880 & ~n9881;
  assign n9883 = ~pi3515 & pi3522;
  assign n9884 = ~pi3412 & n9883;
  assign po3855 = pi3548 | n9884;
  assign n9886 = pi0541 & n8535;
  assign n9887 = pi3548 & n9886;
  assign n9888 = ~pi3452 & pi3526;
  assign n9889 = ~n8546 & ~n9888;
  assign n9890 = pi0541 & ~n9889;
  assign po3872 = n9887 | n9890;
  assign n9892 = pi3526 & n9873;
  assign n9893 = pi0565 & n9892;
  assign po3878 = n9858 | n9893;
  assign n9895 = ~po3872 & ~po3878;
  assign n9896 = ~po3855 & n9895;
  assign n9897 = n9882 & n9896;
  assign n9898 = ~n8561 & n8623;
  assign n9899 = ~po3841 & n9898;
  assign n9900 = n9897 & ~n9899;
  assign n9901 = ~pi3236 & pi3523;
  assign po3848 = pi3522 | n9901;
  assign n9903 = n9900 & ~po3848;
  assign n9904 = pi2647 & ~n9903;
  assign n9905 = n9855 & ~n9904;
  assign n9906 = ~n9850 & ~n9905;
  assign n9907 = pi0752 & n9850;
  assign n9908 = ~n9906 & ~n9907;
  assign n9909 = n9847 & ~n9908;
  assign n9910 = n9845 & ~n9909;
  assign n9911 = ~n9464 & ~n9830;
  assign n9912 = ~pi0613 & ~pi0753;
  assign n9913 = pi0614 & ~n9912;
  assign n9914 = pi0613 & pi0753;
  assign n9915 = ~n9913 & ~n9914;
  assign n9916 = ~pi0614 & n9912;
  assign n9917 = ~pi0735 & n9916;
  assign n9918 = ~pi0612 & n9917;
  assign n9919 = ~pi0658 & n9918;
  assign n9920 = ~pi0636 & n9919;
  assign n9921 = ~pi0637 & ~pi0736;
  assign n9922 = n9920 & n9921;
  assign n9923 = ~pi0634 & ~pi0638;
  assign n9924 = n9922 & n9923;
  assign n9925 = ~pi0639 & n9924;
  assign n9926 = pi0640 & ~n9925;
  assign n9927 = ~pi0639 & ~pi0641;
  assign n9928 = ~n9924 & ~n9927;
  assign n9929 = ~pi0639 & ~pi0640;
  assign n9930 = pi0641 & ~n9929;
  assign n9931 = ~n9928 & ~n9930;
  assign n9932 = ~pi0638 & n9922;
  assign n9933 = pi0634 & ~n9932;
  assign n9934 = ~pi0637 & n9920;
  assign n9935 = pi0736 & ~n9934;
  assign n9936 = pi0638 & ~n9922;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = ~n9933 & n9937;
  assign n9939 = n9931 & n9938;
  assign n9940 = ~n9926 & n9939;
  assign n9941 = pi0658 & ~n9918;
  assign n9942 = pi0637 & ~n9920;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = pi0636 & ~n9919;
  assign n9945 = n9943 & ~n9944;
  assign n9946 = n9940 & n9945;
  assign n9947 = pi0612 & ~n9917;
  assign n9948 = pi0735 & ~n9916;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = n9946 & n9949;
  assign n9951 = n9915 & n9950;
  assign n9952 = ~pi0636 & ~pi0637;
  assign n9953 = ~pi0658 & n9952;
  assign n9954 = ~pi0638 & ~pi0736;
  assign n9955 = ~pi0634 & n9954;
  assign n9956 = ~pi0640 & ~pi0641;
  assign n9957 = ~pi0639 & n9956;
  assign n9958 = n9955 & n9957;
  assign n9959 = n9953 & n9958;
  assign n9960 = n9918 & n9959;
  assign n9961 = n9951 & ~n9960;
  assign n9962 = ~pi0753 & ~n9951;
  assign n9963 = ~n9961 & ~n9962;
  assign n9964 = pi0666 & n9963;
  assign n9965 = pi0568 & n9964;
  assign n9966 = ~pi0568 & ~pi0753;
  assign n9967 = pi0568 & pi0753;
  assign n9968 = ~n9966 & ~n9967;
  assign n9969 = ~pi0568 & ~n9964;
  assign n9970 = ~n9968 & ~n9969;
  assign n9971 = ~n9965 & ~n9970;
  assign n9972 = ~pi0614 & ~pi0735;
  assign n9973 = ~pi0612 & n9972;
  assign n9974 = n9955 & n9973;
  assign n9975 = n9957 & n9974;
  assign n9976 = n9953 & n9975;
  assign n9977 = n9951 & ~n9976;
  assign n9978 = n9916 & ~n9951;
  assign n9979 = ~n9977 & ~n9978;
  assign n9980 = pi0756 & n9979;
  assign n9981 = ~pi0535 & ~n9980;
  assign n9982 = pi0535 & n9980;
  assign n9983 = ~n9981 & ~n9982;
  assign n9984 = ~pi0568 & ~pi0614;
  assign n9985 = pi0568 & pi0614;
  assign n9986 = ~n9984 & ~n9985;
  assign n9987 = ~n9983 & ~n9986;
  assign n9988 = n9983 & n9986;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = ~pi0634 & ~pi0639;
  assign n9991 = ~pi0638 & n9990;
  assign n9992 = ~pi0636 & n9921;
  assign n9993 = ~pi0612 & ~pi0658;
  assign n9994 = ~pi0735 & n9993;
  assign n9995 = n9992 & n9994;
  assign n9996 = n9991 & n9995;
  assign n9997 = n9956 & n9996;
  assign n9998 = n9951 & ~n9997;
  assign n9999 = n9917 & ~n9951;
  assign n10000 = ~n9998 & ~n9999;
  assign n10001 = pi0757 & n10000;
  assign n10002 = pi0536 & n10001;
  assign n10003 = ~pi0536 & ~n10001;
  assign n10004 = ~pi0568 & ~pi0735;
  assign n10005 = pi0568 & pi0735;
  assign n10006 = ~n10004 & ~n10005;
  assign n10007 = ~n10003 & ~n10006;
  assign n10008 = ~n10002 & ~n10007;
  assign n10009 = ~n9989 & ~n10008;
  assign n10010 = ~n10002 & ~n10003;
  assign n10011 = ~n10006 & ~n10010;
  assign n10012 = n10006 & n10010;
  assign n10013 = ~n10011 & ~n10012;
  assign n10014 = ~pi0637 & n9954;
  assign n10015 = n9993 & n10014;
  assign n10016 = ~pi0636 & n10015;
  assign n10017 = n9956 & n9990;
  assign n10018 = n10016 & n10017;
  assign n10019 = n9951 & ~n10018;
  assign n10020 = n9918 & ~n9951;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = pi0660 & n10021;
  assign n10023 = pi0533 & n10022;
  assign n10024 = ~pi0533 & ~n10022;
  assign n10025 = ~pi0568 & ~pi0612;
  assign n10026 = pi0568 & pi0612;
  assign n10027 = ~n10025 & ~n10026;
  assign n10028 = ~n10024 & ~n10027;
  assign n10029 = ~n10023 & ~n10028;
  assign n10030 = ~n10013 & ~n10029;
  assign n10031 = n9989 & n10008;
  assign n10032 = n10030 & ~n10031;
  assign n10033 = ~n10009 & ~n10032;
  assign n10034 = ~n10023 & ~n10024;
  assign n10035 = ~n10027 & ~n10034;
  assign n10036 = n10027 & n10034;
  assign n10037 = ~n10035 & ~n10036;
  assign n10038 = n9954 & n10017;
  assign n10039 = n9953 & n10038;
  assign n10040 = n9951 & ~n10039;
  assign n10041 = n9912 & n9972;
  assign n10042 = n9993 & n10041;
  assign n10043 = ~n9951 & n10042;
  assign n10044 = ~n10040 & ~n10043;
  assign n10045 = pi0754 & n10044;
  assign n10046 = pi0566 & n10045;
  assign n10047 = ~pi0566 & ~n10045;
  assign n10048 = ~pi0568 & ~pi0658;
  assign n10049 = pi0568 & pi0658;
  assign n10050 = ~n10048 & ~n10049;
  assign n10051 = ~n10047 & ~n10050;
  assign n10052 = ~n10046 & ~n10051;
  assign n10053 = ~n10037 & ~n10052;
  assign n10054 = n10037 & n10052;
  assign n10055 = ~pi0566 & n10045;
  assign n10056 = pi0566 & ~n10045;
  assign n10057 = ~n10055 & ~n10056;
  assign n10058 = ~n10050 & n10057;
  assign n10059 = n10050 & ~n10057;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = n9952 & n10038;
  assign n10062 = n9951 & ~n10061;
  assign n10063 = n9920 & ~n9951;
  assign n10064 = ~n10062 & ~n10063;
  assign n10065 = pi0755 & n10064;
  assign n10066 = pi0567 & n10065;
  assign n10067 = ~pi0567 & ~n10065;
  assign n10068 = ~pi0568 & ~pi0636;
  assign n10069 = pi0568 & pi0636;
  assign n10070 = ~n10068 & ~n10069;
  assign n10071 = ~n10067 & ~n10070;
  assign n10072 = ~n10066 & ~n10071;
  assign n10073 = ~n10060 & ~n10072;
  assign n10074 = ~n10054 & n10073;
  assign n10075 = ~n10053 & ~n10074;
  assign n10076 = n10013 & n10029;
  assign n10077 = ~n9989 & ~n10076;
  assign n10078 = ~n10008 & ~n10076;
  assign n10079 = ~n10077 & ~n10078;
  assign n10080 = ~n10075 & ~n10079;
  assign n10081 = n10033 & ~n10080;
  assign n10082 = ~n9981 & ~n9986;
  assign n10083 = ~n9982 & ~n10082;
  assign n10084 = n9912 & ~n9951;
  assign n10085 = ~pi0613 & n9975;
  assign n10086 = n9953 & n10085;
  assign n10087 = n9951 & ~n10086;
  assign n10088 = ~n10084 & ~n10087;
  assign n10089 = pi0643 & n10088;
  assign n10090 = ~pi0568 & ~pi0613;
  assign n10091 = pi0568 & pi0613;
  assign n10092 = ~n10090 & ~n10091;
  assign n10093 = ~pi0534 & n10092;
  assign n10094 = n10089 & ~n10093;
  assign n10095 = pi0534 & ~n10092;
  assign n10096 = ~n10094 & ~n10095;
  assign n10097 = ~n9965 & ~n9969;
  assign n10098 = ~n9968 & ~n10097;
  assign n10099 = n9968 & n10097;
  assign n10100 = ~n10098 & ~n10099;
  assign n10101 = n10096 & n10100;
  assign n10102 = ~n10083 & ~n10101;
  assign n10103 = ~pi0534 & n10089;
  assign n10104 = pi0534 & ~n10089;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = ~n10092 & n10105;
  assign n10107 = n10092 & ~n10105;
  assign n10108 = ~n10106 & ~n10107;
  assign n10109 = ~n10101 & ~n10108;
  assign n10110 = ~n10102 & ~n10109;
  assign n10111 = ~n10081 & ~n10110;
  assign n10112 = n10102 & ~n10108;
  assign n10113 = n9916 & n9996;
  assign n10114 = ~pi0640 & n10113;
  assign n10115 = ~n9951 & ~n10114;
  assign n10116 = n9951 & n9956;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = pi0665 & ~n10117;
  assign n10119 = ~pi0568 & ~pi0640;
  assign n10120 = pi0568 & pi0640;
  assign n10121 = ~n10119 & ~n10120;
  assign n10122 = ~pi0510 & n10121;
  assign n10123 = n10118 & ~n10122;
  assign n10124 = pi0510 & ~n10121;
  assign n10125 = ~n10123 & ~n10124;
  assign n10126 = ~pi0568 & ~pi0639;
  assign n10127 = pi0568 & pi0639;
  assign n10128 = ~n10126 & ~n10127;
  assign n10129 = ~pi0641 & n9929;
  assign n10130 = n9951 & ~n10129;
  assign n10131 = n9916 & n9991;
  assign n10132 = n9995 & n10131;
  assign n10133 = ~n9951 & n10132;
  assign n10134 = ~n10130 & ~n10133;
  assign n10135 = pi0664 & n10134;
  assign n10136 = pi0509 & n10135;
  assign n10137 = ~pi0509 & ~n10135;
  assign n10138 = ~n10136 & ~n10137;
  assign n10139 = ~n10128 & n10138;
  assign n10140 = n10128 & ~n10138;
  assign n10141 = ~n10139 & ~n10140;
  assign n10142 = ~n10125 & n10141;
  assign n10143 = ~pi0568 & ~pi0634;
  assign n10144 = pi0568 & pi0634;
  assign n10145 = ~n10143 & ~n10144;
  assign n10146 = n9951 & ~n10017;
  assign n10147 = n9912 & n9953;
  assign n10148 = n9974 & n10147;
  assign n10149 = ~n9951 & n10148;
  assign n10150 = ~n10146 & ~n10149;
  assign n10151 = pi0663 & n10150;
  assign n10152 = ~pi0508 & ~n10151;
  assign n10153 = pi0508 & n10151;
  assign n10154 = ~n10152 & ~n10153;
  assign n10155 = ~n10145 & ~n10154;
  assign n10156 = n10145 & n10154;
  assign n10157 = ~n10155 & ~n10156;
  assign n10158 = ~n10128 & ~n10137;
  assign n10159 = ~n10136 & ~n10158;
  assign n10160 = n10157 & n10159;
  assign n10161 = n10142 & ~n10160;
  assign n10162 = n10014 & n10017;
  assign n10163 = n9994 & n10162;
  assign n10164 = n9916 & n10163;
  assign n10165 = ~pi0636 & n10164;
  assign n10166 = ~n9951 & n10165;
  assign n10167 = pi0641 & n9951;
  assign n10168 = ~n10166 & ~n10167;
  assign n10169 = pi0667 & n10168;
  assign n10170 = ~pi0568 & ~pi0641;
  assign n10171 = pi0568 & pi0641;
  assign n10172 = ~n10170 & ~n10171;
  assign n10173 = ~pi0569 & n10172;
  assign n10174 = n10169 & ~n10173;
  assign n10175 = pi0569 & ~n10172;
  assign n10176 = ~n10174 & ~n10175;
  assign n10177 = ~pi0510 & n10118;
  assign n10178 = pi0510 & ~n10118;
  assign n10179 = ~n10177 & ~n10178;
  assign n10180 = ~n10121 & ~n10179;
  assign n10181 = n10121 & n10179;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = ~n10176 & n10182;
  assign n10184 = n10176 & ~n10182;
  assign n10185 = pi0569 & n10169;
  assign n10186 = ~pi0569 & ~n10169;
  assign n10187 = ~n10185 & ~n10186;
  assign n10188 = ~n10172 & ~n10187;
  assign n10189 = n10172 & n10187;
  assign n10190 = ~n10188 & ~n10189;
  assign n10191 = ~pi0568 & ~n10190;
  assign n10192 = ~n10184 & n10191;
  assign n10193 = ~n10183 & ~n10192;
  assign n10194 = n10141 & ~n10157;
  assign n10195 = ~n10125 & ~n10157;
  assign n10196 = n10125 & ~n10141;
  assign n10197 = ~n10159 & ~n10196;
  assign n10198 = ~n10195 & ~n10197;
  assign n10199 = ~n10194 & n10198;
  assign n10200 = ~n10193 & ~n10199;
  assign n10201 = ~n10157 & ~n10159;
  assign n10202 = ~n10200 & ~n10201;
  assign n10203 = ~n10161 & n10202;
  assign n10204 = ~pi0568 & ~pi0637;
  assign n10205 = pi0568 & pi0637;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = n9921 & n9923;
  assign n10208 = n10129 & n10207;
  assign n10209 = n9951 & ~n10208;
  assign n10210 = n9952 & n10042;
  assign n10211 = ~n9951 & n10210;
  assign n10212 = ~n10209 & ~n10211;
  assign n10213 = pi0642 & n10212;
  assign n10214 = ~pi0505 & n10213;
  assign n10215 = pi0505 & ~n10213;
  assign n10216 = ~n10214 & ~n10215;
  assign n10217 = ~n10206 & n10216;
  assign n10218 = n10206 & ~n10216;
  assign n10219 = ~n10217 & ~n10218;
  assign n10220 = n9951 & ~n10038;
  assign n10221 = n9992 & n10042;
  assign n10222 = ~n9951 & n10221;
  assign n10223 = ~n10220 & ~n10222;
  assign n10224 = pi0661 & n10223;
  assign n10225 = pi0506 & n10224;
  assign n10226 = ~pi0506 & ~n10224;
  assign n10227 = ~pi0568 & ~pi0736;
  assign n10228 = pi0568 & pi0736;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = ~n10226 & ~n10229;
  assign n10231 = ~n10225 & ~n10230;
  assign n10232 = n10219 & n10231;
  assign n10233 = ~n10066 & ~n10067;
  assign n10234 = ~n10070 & ~n10233;
  assign n10235 = n10070 & n10233;
  assign n10236 = ~n10234 & ~n10235;
  assign n10237 = pi0505 & n10213;
  assign n10238 = ~pi0505 & ~n10213;
  assign n10239 = ~n10206 & ~n10238;
  assign n10240 = ~n10237 & ~n10239;
  assign n10241 = n10236 & n10240;
  assign n10242 = ~n10232 & ~n10241;
  assign n10243 = ~pi0568 & ~pi0638;
  assign n10244 = pi0568 & pi0638;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = n9923 & n9957;
  assign n10247 = n9951 & ~n10246;
  assign n10248 = n10016 & n10041;
  assign n10249 = ~n9951 & n10248;
  assign n10250 = ~n10247 & ~n10249;
  assign n10251 = pi0662 & n10250;
  assign n10252 = ~pi0507 & n10251;
  assign n10253 = pi0507 & ~n10251;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = ~n10245 & n10254;
  assign n10256 = n10245 & ~n10254;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = ~n10145 & ~n10152;
  assign n10259 = ~n10153 & ~n10258;
  assign n10260 = n10257 & n10259;
  assign n10261 = pi0507 & n10251;
  assign n10262 = ~pi0507 & ~n10251;
  assign n10263 = ~n10245 & ~n10262;
  assign n10264 = ~n10261 & ~n10263;
  assign n10265 = ~n10225 & ~n10226;
  assign n10266 = ~n10229 & ~n10265;
  assign n10267 = n10229 & n10265;
  assign n10268 = ~n10266 & ~n10267;
  assign n10269 = n10264 & n10268;
  assign n10270 = ~n10260 & ~n10269;
  assign n10271 = n10242 & n10270;
  assign n10272 = ~n10203 & n10271;
  assign n10273 = ~n10257 & ~n10259;
  assign n10274 = n10264 & ~n10273;
  assign n10275 = ~n10268 & ~n10274;
  assign n10276 = ~n10264 & n10273;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = n10242 & ~n10277;
  assign n10279 = ~n10236 & ~n10240;
  assign n10280 = ~n10278 & ~n10279;
  assign n10281 = ~n10219 & ~n10231;
  assign n10282 = ~n10241 & n10281;
  assign n10283 = n10280 & ~n10282;
  assign n10284 = ~n10272 & n10283;
  assign n10285 = n10060 & n10072;
  assign n10286 = ~n10054 & ~n10285;
  assign n10287 = ~n10284 & n10286;
  assign n10288 = ~n10079 & n10287;
  assign n10289 = ~n10110 & n10288;
  assign n10290 = ~n10112 & ~n10289;
  assign n10291 = ~n10096 & ~n10100;
  assign n10292 = n10290 & ~n10291;
  assign n10293 = ~n10111 & n10292;
  assign n10294 = ~n9971 & n10293;
  assign n10295 = n9971 & ~n10293;
  assign n10296 = ~n10294 & ~n10295;
  assign n10297 = pi0534 & n10089;
  assign n10298 = ~n9981 & ~n10003;
  assign n10299 = ~n10024 & ~n10047;
  assign n10300 = ~n10067 & ~n10238;
  assign n10301 = ~n10226 & n10261;
  assign n10302 = ~n10225 & ~n10301;
  assign n10303 = n10300 & ~n10302;
  assign n10304 = ~n10067 & n10237;
  assign n10305 = ~n10303 & ~n10304;
  assign n10306 = pi0506 & n10251;
  assign n10307 = pi0507 & ~n10226;
  assign n10308 = ~n10306 & ~n10307;
  assign n10309 = n10224 & n10251;
  assign n10310 = n10308 & ~n10309;
  assign n10311 = n10136 & ~n10152;
  assign n10312 = ~pi0510 & ~n10118;
  assign n10313 = n10185 & ~n10312;
  assign n10314 = pi0510 & n10118;
  assign n10315 = ~n10313 & ~n10314;
  assign n10316 = n10135 & n10151;
  assign n10317 = pi0508 & pi0509;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = pi0508 & n10135;
  assign n10320 = n10318 & ~n10319;
  assign n10321 = pi0509 & n10151;
  assign n10322 = n10320 & ~n10321;
  assign n10323 = ~n10315 & ~n10322;
  assign n10324 = ~n10311 & ~n10323;
  assign n10325 = ~n10153 & n10324;
  assign n10326 = ~n10310 & ~n10325;
  assign n10327 = n10300 & n10326;
  assign n10328 = ~n10066 & ~n10327;
  assign n10329 = n10305 & n10328;
  assign n10330 = n10299 & ~n10329;
  assign n10331 = n10298 & n10330;
  assign n10332 = ~n9981 & n10002;
  assign n10333 = ~n10024 & n10046;
  assign n10334 = ~n10023 & ~n10333;
  assign n10335 = n10298 & ~n10334;
  assign n10336 = ~n10332 & ~n10335;
  assign n10337 = ~n10331 & n10336;
  assign n10338 = ~n9982 & n10337;
  assign n10339 = ~pi0534 & ~n10089;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = ~n10297 & ~n10340;
  assign n10342 = ~n10097 & ~n10341;
  assign n10343 = n10097 & n10341;
  assign n10344 = ~n10342 & ~n10343;
  assign n10345 = n10296 & ~n10344;
  assign n10346 = ~n10101 & ~n10291;
  assign n10347 = n10081 & ~n10288;
  assign n10348 = n10083 & n10108;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = ~n10083 & ~n10108;
  assign n10351 = ~n10349 & ~n10350;
  assign n10352 = ~n10346 & ~n10351;
  assign n10353 = n10346 & n10351;
  assign n10354 = ~n10352 & ~n10353;
  assign n10355 = ~n10296 & ~n10354;
  assign n10356 = ~n10345 & ~n10355;
  assign n10357 = ~pi0568 & ~n10356;
  assign n10358 = ~n9969 & ~n10341;
  assign n10359 = ~n9965 & ~n10358;
  assign n10360 = pi0568 & ~n10359;
  assign n10361 = ~pi0568 & n10359;
  assign n10362 = ~n10360 & ~n10361;
  assign n10363 = ~n10354 & n10362;
  assign n10364 = ~n10344 & ~n10362;
  assign n10365 = ~n10363 & ~n10364;
  assign n10366 = pi0568 & ~n10365;
  assign n10367 = ~n10357 & ~n10366;
  assign n10368 = pi0666 & ~n9951;
  assign n10369 = ~pi0753 & n10368;
  assign n10370 = pi0666 & n9961;
  assign n10371 = ~n10369 & ~n10370;
  assign n10372 = n10367 & n10371;
  assign n10373 = n9829 & ~n10372;
  assign n10374 = n9394 & n9395;
  assign n10375 = pi2435 & n10374;
  assign n10376 = n9411 & n9412;
  assign n10377 = pi2268 & n10376;
  assign n10378 = ~n10375 & ~n10377;
  assign n10379 = n9404 & n9405;
  assign n10380 = pi1983 & n10379;
  assign n10381 = n9372 & n9385;
  assign n10382 = pi2445 & n10381;
  assign n10383 = ~n10380 & ~n10382;
  assign n10384 = n10378 & n10383;
  assign n10385 = ~n9829 & ~n10384;
  assign n10386 = ~n10373 & ~n10385;
  assign n10387 = n9911 & ~n10386;
  assign po0215 = ~n9910 | n10387;
  assign n10389 = pi3871 & n9804;
  assign n10390 = pi3887 & n9774;
  assign n10391 = ~n10389 & ~n10390;
  assign n10392 = pi3855 & n9802;
  assign n10393 = pi3919 & n9781;
  assign n10394 = pi3903 & n9771;
  assign n10395 = ~n10393 & ~n10394;
  assign n10396 = pi3951 & n9791;
  assign n10397 = pi3935 & n9788;
  assign n10398 = ~n10396 & ~n10397;
  assign n10399 = n10395 & n10398;
  assign n10400 = ~n10392 & n10399;
  assign n10401 = n10391 & n10400;
  assign n10402 = pi3871 & n9799;
  assign n10403 = n10401 & ~n10402;
  assign n10404 = pi3983 & n9783;
  assign n10405 = pi3967 & n9793;
  assign n10406 = ~n10404 & ~n10405;
  assign n10407 = n10403 & n10406;
  assign n10408 = ~n9472 & ~n10407;
  assign n10409 = pi1331 & ~n9257;
  assign n10410 = ~pi3233 & ~pi3329;
  assign n10411 = pi3512 & ~n10410;
  assign n10412 = ~n10409 & ~n10411;
  assign n10413 = pi0593 & pi1359;
  assign n10414 = pi0381 & pi1057;
  assign n10415 = ~n10413 & ~n10414;
  assign n10416 = n10412 & n10415;
  assign n10417 = n9475 & ~n10416;
  assign n10418 = pi0120 & ~pi0979;
  assign n10419 = pi0117 & pi0979;
  assign n10420 = ~n10418 & ~n10419;
  assign n10421 = pi0720 & ~n10420;
  assign n10422 = pi0241 & ~pi0979;
  assign n10423 = pi0240 & pi0979;
  assign n10424 = ~n10422 & ~n10423;
  assign n10425 = pi0721 & ~n10424;
  assign n10426 = ~n10421 & ~n10425;
  assign n10427 = ~pi0979 & pi2641;
  assign n10428 = pi0979 & pi3174;
  assign n10429 = ~n10427 & ~n10428;
  assign n10430 = pi0765 & ~n10429;
  assign n10431 = ~pi0979 & pi2895;
  assign n10432 = pi0979 & pi3143;
  assign n10433 = ~n10431 & ~n10432;
  assign n10434 = pi0766 & ~n10433;
  assign n10435 = ~n10430 & ~n10434;
  assign n10436 = ~pi0979 & pi2614;
  assign n10437 = pi0979 & pi2608;
  assign n10438 = ~n10436 & ~n10437;
  assign n10439 = pi0763 & ~n10438;
  assign n10440 = ~pi0979 & pi2627;
  assign n10441 = pi0979 & pi2621;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = pi0764 & ~n10442;
  assign n10444 = ~n10439 & ~n10443;
  assign n10445 = n10435 & n10444;
  assign n10446 = ~n9499 & n10445;
  assign n10447 = n10426 & n10446;
  assign n10448 = n9486 & ~n10447;
  assign n10449 = ~n10417 & ~n10448;
  assign n10450 = ~pi0979 & pi2853;
  assign n10451 = pi0979 & pi2136;
  assign n10452 = ~n10450 & ~n10451;
  assign n10453 = pi0717 & ~n10452;
  assign n10454 = pi0184 & ~pi0979;
  assign n10455 = pi0183 & pi0979;
  assign n10456 = ~n10454 & ~n10455;
  assign n10457 = pi0716 & ~n10456;
  assign n10458 = pi0272 & ~pi0979;
  assign n10459 = pi0271 & pi0979;
  assign n10460 = ~n10458 & ~n10459;
  assign n10461 = pi0761 & ~n10460;
  assign n10462 = ~n10457 & ~n10461;
  assign n10463 = ~n9535 & n10462;
  assign n10464 = ~n9531 & n10463;
  assign n10465 = ~n10453 & n10464;
  assign n10466 = n9523 & ~n10465;
  assign n10467 = pi0979 & pi2173;
  assign n10468 = ~pi0979 & pi2803;
  assign n10469 = ~n10467 & ~n10468;
  assign n10470 = pi0836 & ~n10469;
  assign n10471 = ~pi0979 & pi2949;
  assign n10472 = pi0979 & pi2189;
  assign n10473 = ~n10471 & ~n10472;
  assign n10474 = pi0837 & ~n10473;
  assign n10475 = ~n10470 & ~n10474;
  assign n10476 = pi0979 & pi2155;
  assign n10477 = ~pi0979 & pi2927;
  assign n10478 = ~n10476 & ~n10477;
  assign n10479 = pi0767 & ~n10478;
  assign n10480 = ~pi0979 & pi2430;
  assign n10481 = pi0979 & pi1965;
  assign n10482 = ~n10480 & ~n10481;
  assign n10483 = pi0768 & ~n10482;
  assign n10484 = ~n10479 & ~n10483;
  assign n10485 = pi0179 & ~pi0979;
  assign n10486 = pi0164 & pi0979;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = pi0838 & ~n10487;
  assign n10489 = n10484 & ~n10488;
  assign n10490 = n10475 & n10489;
  assign n10491 = n9549 & ~n10490;
  assign n10492 = ~n10466 & ~n10491;
  assign n10493 = pi1340 & pi2288;
  assign n10494 = pi1341 & pi2122;
  assign n10495 = ~n10493 & ~n10494;
  assign n10496 = pi1342 & pi2310;
  assign n10497 = n10495 & ~n10496;
  assign n10498 = pi1055 & pi2725;
  assign n10499 = n10497 & ~n10498;
  assign n10500 = pi1343 & pi2324;
  assign n10501 = pi1054 & pi2717;
  assign n10502 = ~n10500 & ~n10501;
  assign n10503 = pi1349 & pi2735;
  assign n10504 = pi1056 & pi2543;
  assign n10505 = ~n10503 & ~n10504;
  assign n10506 = pi1354 & pi2533;
  assign n10507 = n10505 & ~n10506;
  assign n10508 = pi1357 & pi2467;
  assign n10509 = n10507 & ~n10508;
  assign n10510 = pi1355 & pi2525;
  assign n10511 = pi1356 & pi2755;
  assign n10512 = ~n10510 & ~n10511;
  assign n10513 = n10509 & n10512;
  assign n10514 = n10502 & n10513;
  assign n10515 = n10499 & n10514;
  assign n10516 = n9736 & ~n10515;
  assign n10517 = pi1600 & pi2211;
  assign n10518 = pi1337 & pi2225;
  assign n10519 = ~n10517 & ~n10518;
  assign n10520 = pi1338 & pi2239;
  assign n10521 = n10519 & ~n10520;
  assign n10522 = pi1346 & pi2671;
  assign n10523 = n10521 & ~n10522;
  assign n10524 = pi1339 & pi2253;
  assign n10525 = pi1345 & pi2657;
  assign n10526 = ~n10524 & ~n10525;
  assign n10527 = pi1351 & pi2269;
  assign n10528 = pi1352 & pi2446;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = pi1353 & pi1984;
  assign n10531 = n10529 & ~n10530;
  assign n10532 = pi1350 & pi2436;
  assign n10533 = n10531 & ~n10532;
  assign n10534 = pi1347 & pi2685;
  assign n10535 = pi1348 & pi2695;
  assign n10536 = ~n10534 & ~n10535;
  assign n10537 = n10533 & n10536;
  assign n10538 = n10526 & n10537;
  assign n10539 = n10523 & n10538;
  assign n10540 = n9577 & ~n10539;
  assign n10541 = ~n10516 & ~n10540;
  assign n10542 = pi0189 & pi1336;
  assign n10543 = pi1333 & pi1744;
  assign n10544 = ~n10542 & ~n10543;
  assign n10545 = pi1332 & pi2579;
  assign n10546 = pi1335 & pi2594;
  assign n10547 = ~n10545 & ~n10546;
  assign n10548 = n10544 & n10547;
  assign n10549 = n9726 & ~n10548;
  assign n10550 = pi0961 & n9614;
  assign n10551 = pi2053 & n9618;
  assign n10552 = ~n10550 & ~n10551;
  assign n10553 = pi0972 & n9687;
  assign n10554 = pi1909 & n9691;
  assign n10555 = ~n10553 & ~n10554;
  assign n10556 = n10552 & n10555;
  assign n10557 = pi0796 & n9607;
  assign n10558 = pi1844 & n10557;
  assign n10559 = pi1837 & n9698;
  assign n10560 = ~n10558 & ~n10559;
  assign n10561 = pi0889 & n9715;
  assign n10562 = pi1874 & n9718;
  assign n10563 = ~n10561 & ~n10562;
  assign n10564 = pi0890 & n9702;
  assign n10565 = pi1842 & n10564;
  assign n10566 = pi0897 & n9707;
  assign n10567 = ~n10565 & ~n10566;
  assign n10568 = n10563 & n10567;
  assign n10569 = n10560 & n10568;
  assign n10570 = n10556 & n10569;
  assign n10571 = pi1762 & n9657;
  assign n10572 = pi1750 & n9659;
  assign n10573 = ~n10571 & ~n10572;
  assign n10574 = pi2102 & n9628;
  assign n10575 = pi1019 & n9631;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = pi2111 & n9622;
  assign n10578 = n10576 & ~n10577;
  assign n10579 = n10573 & n10578;
  assign n10580 = n10570 & n10579;
  assign n10581 = pi1880 & n9679;
  assign n10582 = pi0303 & n9682;
  assign n10583 = ~n10581 & ~n10582;
  assign n10584 = pi0779 & n9670;
  assign n10585 = pi0688 & n9676;
  assign n10586 = ~n10584 & ~n10585;
  assign n10587 = pi0819 & n9710;
  assign n10588 = pi1783 & n9712;
  assign n10589 = ~n10587 & ~n10588;
  assign n10590 = n10586 & n10589;
  assign n10591 = pi2989 & n9647;
  assign n10592 = pi0724 & n9654;
  assign n10593 = ~n10591 & ~n10592;
  assign n10594 = n10590 & n10593;
  assign n10595 = n10583 & n10594;
  assign n10596 = n10580 & n10595;
  assign n10597 = pi1934 & ~n10596;
  assign n10598 = ~n10549 & ~n10597;
  assign n10599 = n10541 & n10598;
  assign n10600 = n10492 & n10599;
  assign n10601 = n10449 & n10600;
  assign n10602 = pi3296 & po3871;
  assign n10603 = n10601 & ~n10602;
  assign n10604 = ~pi1787 & ~n10603;
  assign n10605 = pi1787 & pi2833;
  assign n10606 = ~n10604 & ~n10605;
  assign n10607 = n9472 & ~n10606;
  assign n10608 = ~n10408 & ~n10607;
  assign n10609 = n9464 & ~n10608;
  assign n10610 = pi1984 & n9832;
  assign n10611 = pi2446 & n9834;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = pi2436 & n9837;
  assign n10614 = pi2269 & n9839;
  assign n10615 = ~n10613 & ~n10614;
  assign n10616 = n10612 & n10615;
  assign n10617 = n9831 & ~n10616;
  assign n10618 = ~n9464 & n10617;
  assign n10619 = ~n10609 & ~n10618;
  assign n10620 = ~n9464 & ~n9829;
  assign n10621 = n9830 & n10620;
  assign n10622 = pi2557 & po3871;
  assign n10623 = pi0819 & n9853;
  assign n10624 = ~n10622 & ~n10623;
  assign n10625 = pi2529 & ~n9903;
  assign n10626 = n10624 & ~n10625;
  assign n10627 = ~n9850 & ~n10626;
  assign n10628 = pi0779 & n9850;
  assign n10629 = ~n10627 & ~n10628;
  assign n10630 = n10621 & ~n10629;
  assign n10631 = n10619 & ~n10630;
  assign n10632 = n10105 & ~n10338;
  assign n10633 = ~n10105 & n10338;
  assign n10634 = ~n10632 & ~n10633;
  assign n10635 = n10296 & ~n10634;
  assign n10636 = ~n10083 & n10108;
  assign n10637 = n10083 & ~n10108;
  assign n10638 = ~n10636 & ~n10637;
  assign n10639 = ~n10347 & n10638;
  assign n10640 = n10347 & ~n10638;
  assign n10641 = ~n10639 & ~n10640;
  assign n10642 = ~n10296 & ~n10641;
  assign n10643 = ~n10635 & ~n10642;
  assign n10644 = ~pi0568 & ~n10643;
  assign n10645 = n10362 & ~n10641;
  assign n10646 = ~n10362 & ~n10634;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = pi0568 & ~n10647;
  assign n10649 = ~n10644 & ~n10648;
  assign n10650 = pi0643 & n10084;
  assign n10651 = pi0643 & n10087;
  assign n10652 = ~n10650 & ~n10651;
  assign n10653 = n10649 & n10652;
  assign n10654 = n9829 & ~n10653;
  assign n10655 = pi2436 & n10374;
  assign n10656 = pi2269 & n10376;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = pi1984 & n10379;
  assign n10659 = pi2446 & n10381;
  assign n10660 = ~n10658 & ~n10659;
  assign n10661 = n10657 & n10660;
  assign n10662 = ~n9829 & ~n10661;
  assign n10663 = ~n10654 & ~n10662;
  assign n10664 = n9911 & ~n10663;
  assign po0214 = ~n10631 | n10664;
  assign n10666 = ~pi3680 & ~po0214;
  assign n10667 = po0215 & ~n10666;
  assign n10668 = ~n8567 & n8589;
  assign n10669 = pi2493 & n8577;
  assign n10670 = pi2404 & ~n8577;
  assign n10671 = ~n10669 & ~n10670;
  assign n10672 = ~n10668 & ~n10671;
  assign n10673 = pi1450 & n10668;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = n10667 & n10674;
  assign n10676 = pi2405 & ~n8577;
  assign n10677 = pi2494 & n8577;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = ~n10668 & ~n10678;
  assign n10680 = pi1451 & n10668;
  assign n10681 = ~n10679 & ~n10680;
  assign n10682 = pi2500 & n8577;
  assign n10683 = pi2409 & ~n8577;
  assign n10684 = ~n10682 & ~n10683;
  assign n10685 = ~n10668 & ~n10684;
  assign n10686 = pi1459 & n10668;
  assign n10687 = ~n10685 & ~n10686;
  assign n10688 = pi2501 & n8577;
  assign n10689 = pi2473 & ~n8577;
  assign n10690 = ~n10688 & ~n10689;
  assign n10691 = ~n10668 & ~n10690;
  assign n10692 = pi1460 & n10668;
  assign n10693 = ~n10691 & ~n10692;
  assign n10694 = n10687 & n10693;
  assign n10695 = n10681 & n10694;
  assign n10696 = n10675 & n10695;
  assign po0044 = ~n9357 & n10696;
  assign n10698 = ~n10681 & n10694;
  assign n10699 = n10675 & n10698;
  assign po0045 = ~n9357 & n10699;
  assign n10701 = n10667 & ~n10674;
  assign n10702 = n10695 & n10701;
  assign po0046 = ~n9357 & n10702;
  assign n10704 = n10698 & n10701;
  assign po0047 = ~n9357 & n10704;
  assign n10706 = n10667 & n10687;
  assign n10707 = n10681 & ~n10693;
  assign n10708 = n10706 & n10707;
  assign n10709 = n10674 & n10708;
  assign po0048 = ~n9357 & n10709;
  assign n10711 = ~n10681 & n10706;
  assign n10712 = ~n10693 & n10711;
  assign n10713 = n10674 & n10712;
  assign po0049 = ~n9357 & n10713;
  assign n10715 = ~n10674 & n10708;
  assign po0050 = ~n9357 & n10715;
  assign n10717 = ~n10674 & n10712;
  assign po0051 = ~n9357 & n10717;
  assign n10719 = ~n10696 & ~n10699;
  assign n10720 = ~n10702 & n10719;
  assign n10721 = ~n10709 & n10720;
  assign n10722 = ~n10704 & n10721;
  assign n10723 = ~n10713 & n10722;
  assign n10724 = ~n10715 & ~n10717;
  assign n10725 = n10723 & n10724;
  assign n10726 = ~pi3426 & ~n8561;
  assign n10727 = ~po3871 & ~n10726;
  assign n10728 = ~n9356 & ~n10727;
  assign n10729 = ~n8567 & ~n8604;
  assign n10730 = ~n10728 & ~n10729;
  assign po0052 = n10725 | n10730;
  assign n10732 = pi3378 & n9352;
  assign n10733 = pi1037 & n9640;
  assign n10734 = pi1013 & n9634;
  assign n10735 = pi1029 & n10734;
  assign n10736 = pi1038 & n10735;
  assign n10737 = pi1028 & n10736;
  assign n10738 = n10733 & n10737;
  assign n10739 = pi2789 & ~n10738;
  assign n10740 = ~pi0692 & n10739;
  assign n10741 = ~po3841 & n10740;
  assign n10742 = ~n9352 & n10741;
  assign n10743 = ~n10732 & ~n10742;
  assign n10744 = ~pi3426 & n10740;
  assign n10745 = ~n8561 & ~n10744;
  assign n10746 = ~pi0403 & pi0416;
  assign n10747 = ~pi0417 & n10746;
  assign n10748 = pi3055 & ~pi3641;
  assign n10749 = n10747 & ~n10748;
  assign n10750 = ~pi0419 & n10749;
  assign n10751 = pi0403 & pi0417;
  assign n10752 = ~pi0416 & n10751;
  assign n10753 = ~pi0418 & n10752;
  assign n10754 = ~n10750 & ~n10753;
  assign n10755 = pi0405 & ~pi0420;
  assign n10756 = ~pi0419 & n10755;
  assign n10757 = pi0418 & n10756;
  assign n10758 = ~pi0421 & n10757;
  assign n10759 = n8609 & n10758;
  assign n10760 = ~pi0422 & n10759;
  assign n10761 = ~n8615 & ~n10760;
  assign n10762 = n10754 & n10761;
  assign n10763 = ~po3841 & ~n10762;
  assign n10764 = n9345 & n10763;
  assign n10765 = n10745 & n10764;
  assign n10766 = pi3257 & n8561;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = pi1422 & pi2515;
  assign n10769 = n8589 & n10768;
  assign n10770 = ~n8580 & n8581;
  assign n10771 = pi2048 & ~pi2986;
  assign n10772 = pi3099 & ~n10771;
  assign n10773 = n10770 & n10772;
  assign n10774 = n8577 & n10773;
  assign n10775 = ~n10769 & ~n10774;
  assign n10776 = ~n8568 & n10775;
  assign n10777 = ~n9420 & n10776;
  assign n10778 = ~pi2048 & ~pi2986;
  assign n10779 = ~pi3099 & ~n10778;
  assign n10780 = n10770 & n10779;
  assign n10781 = n8577 & n10780;
  assign n10782 = pi1422 & pi2769;
  assign n10783 = n8589 & n10782;
  assign n10784 = ~n9419 & ~n10783;
  assign n10785 = ~n9422 & n10784;
  assign n10786 = ~n10781 & n10785;
  assign n10787 = n10777 & n10786;
  assign n10788 = ~n8567 & ~n10787;
  assign n10789 = n10767 & ~n10788;
  assign n10790 = n10743 & n10789;
  assign n10791 = ~pi0405 & n10759;
  assign n10792 = ~n8615 & ~n10791;
  assign n10793 = pi0416 & pi0417;
  assign n10794 = ~pi0418 & n10793;
  assign n10795 = n10792 & ~n10794;
  assign n10796 = ~n9424 & ~n9460;
  assign n10797 = ~n9415 & n9424;
  assign n10798 = ~n10796 & ~n10797;
  assign n10799 = n10795 & n10798;
  assign n10800 = ~pi0418 & n10749;
  assign n10801 = n10799 & ~n10800;
  assign n10802 = ~pi0417 & ~pi0418;
  assign n10803 = n10746 & n10802;
  assign n10804 = ~n10748 & n10803;
  assign n10805 = n10795 & ~n10804;
  assign n10806 = ~n9361 & n10805;
  assign n10807 = pi0405 & n10759;
  assign n10808 = pi0418 & n10793;
  assign n10809 = ~n10807 & ~n10808;
  assign n10810 = pi0418 & n10747;
  assign n10811 = ~n10748 & n10810;
  assign n10812 = n10809 & ~n10811;
  assign n10813 = n10805 & n10812;
  assign n10814 = ~n10806 & ~n10813;
  assign n10815 = ~n10801 & n10814;
  assign n10816 = ~po3841 & n10745;
  assign n10817 = pi3436 & ~pi3451;
  assign n10818 = n9387 & n10817;
  assign n10819 = pi2488 & ~pi3426;
  assign n10820 = n9360 & n10819;
  assign n10821 = pi3398 & n10820;
  assign n10822 = pi3392 & n10821;
  assign n10823 = ~pi0996 & ~n10822;
  assign n10824 = n9365 & ~n10823;
  assign n10825 = ~n10818 & ~n10824;
  assign n10826 = pi0414 & pi0415;
  assign n10827 = ~n10825 & n10826;
  assign n10828 = ~pi3398 & n9360;
  assign n10829 = n10819 & n10828;
  assign n10830 = ~pi3392 & n10829;
  assign n10831 = ~pi0999 & ~n10830;
  assign n10832 = n9365 & ~n10831;
  assign n10833 = ~pi3436 & ~pi3451;
  assign n10834 = n9363 & n10833;
  assign n10835 = ~n10832 & ~n10834;
  assign n10836 = ~pi0414 & ~pi0415;
  assign n10837 = ~n10835 & n10836;
  assign n10838 = ~n10827 & ~n10837;
  assign n10839 = pi3392 & n10829;
  assign n10840 = ~pi0998 & ~n10839;
  assign n10841 = n9365 & ~n10840;
  assign n10842 = n9363 & n10817;
  assign n10843 = ~n10841 & ~n10842;
  assign n10844 = ~pi0414 & pi0415;
  assign n10845 = ~n10843 & n10844;
  assign n10846 = n9387 & n10833;
  assign n10847 = ~pi3392 & n10821;
  assign n10848 = ~pi0997 & ~n10847;
  assign n10849 = n9365 & ~n10848;
  assign n10850 = ~n10846 & ~n10849;
  assign n10851 = pi0414 & ~pi0415;
  assign n10852 = ~n10850 & n10851;
  assign n10853 = ~n10845 & ~n10852;
  assign n10854 = n10838 & n10853;
  assign n10855 = n9424 & ~n10854;
  assign n10856 = n9440 & n9447;
  assign n10857 = ~n9433 & n10856;
  assign n10858 = ~n10843 & n10857;
  assign n10859 = n9433 & n10856;
  assign n10860 = ~n10835 & n10859;
  assign n10861 = ~n10858 & ~n10860;
  assign n10862 = ~n9440 & n9447;
  assign n10863 = ~n9433 & n10862;
  assign n10864 = ~n10825 & n10863;
  assign n10865 = n9433 & n10862;
  assign n10866 = ~n10850 & n10865;
  assign n10867 = ~n10864 & ~n10866;
  assign n10868 = n10861 & n10867;
  assign n10869 = ~n9424 & ~n10868;
  assign n10870 = ~n10855 & ~n10869;
  assign n10871 = n10798 & n10870;
  assign n10872 = n10816 & ~n10871;
  assign n10873 = ~pi2488 & n9360;
  assign n10874 = ~n10805 & ~n10873;
  assign n10875 = pi0830 & n10874;
  assign n10876 = n10872 & ~n10875;
  assign n10877 = n10815 & n10876;
  assign n10878 = ~n9426 & ~n10877;
  assign n10879 = ~n10798 & n10870;
  assign n10880 = n10816 & n10879;
  assign n10881 = ~n10805 & n10880;
  assign n10882 = ~n9361 & ~n10798;
  assign n10883 = n10870 & n10882;
  assign n10884 = ~n10881 & ~n10883;
  assign n10885 = ~n10878 & n10884;
  assign n10886 = ~n10805 & n10816;
  assign n10887 = ~n9361 & ~n10886;
  assign n10888 = ~pi0830 & n10886;
  assign n10889 = ~n10887 & ~n10888;
  assign n10890 = n10870 & ~n10889;
  assign n10891 = n9426 & n10870;
  assign n10892 = n10798 & n10891;
  assign n10893 = ~n10890 & ~n10892;
  assign n10894 = pi0830 & n10873;
  assign n10895 = ~n10805 & n10894;
  assign n10896 = ~n10870 & n10895;
  assign n10897 = ~n10801 & ~n10896;
  assign n10898 = n10816 & n10897;
  assign n10899 = ~n10806 & n10898;
  assign n10900 = ~n10813 & n10899;
  assign n10901 = ~n9426 & ~n10900;
  assign n10902 = n10893 & ~n10901;
  assign n10903 = n9426 & ~n10873;
  assign n10904 = ~n10870 & n10903;
  assign n10905 = ~n10870 & ~n10873;
  assign n10906 = ~pi0830 & n10905;
  assign n10907 = ~n10880 & ~n10906;
  assign n10908 = ~n10805 & ~n10907;
  assign n10909 = ~n10904 & ~n10908;
  assign n10910 = n10872 & ~n10895;
  assign n10911 = ~n10801 & ~n10813;
  assign n10912 = n10910 & n10911;
  assign n10913 = ~n9426 & ~n10912;
  assign n10914 = n10909 & ~n10913;
  assign n10915 = pi3859 & n9804;
  assign n10916 = pi3875 & n9774;
  assign n10917 = ~n10915 & ~n10916;
  assign n10918 = pi3843 & n9802;
  assign n10919 = pi3891 & n9771;
  assign n10920 = pi3955 & n9793;
  assign n10921 = ~n10919 & ~n10920;
  assign n10922 = pi3939 & n9791;
  assign n10923 = pi3923 & n9788;
  assign n10924 = ~n10922 & ~n10923;
  assign n10925 = n10921 & n10924;
  assign n10926 = ~n10918 & n10925;
  assign n10927 = n10917 & n10926;
  assign n10928 = pi3859 & n9799;
  assign n10929 = n10927 & ~n10928;
  assign n10930 = pi3907 & n9781;
  assign n10931 = pi3971 & n9783;
  assign n10932 = ~n10930 & ~n10931;
  assign n10933 = n10929 & n10932;
  assign n10934 = ~n9472 & ~n10933;
  assign n10935 = pi0393 & pi1057;
  assign n10936 = pi1059 & pi2981;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = pi1053 & pi2408;
  assign n10939 = n10937 & ~n10938;
  assign n10940 = pi0979 & pi1344;
  assign n10941 = n10939 & ~n10940;
  assign n10942 = pi1047 & pi1334;
  assign n10943 = pi0980 & pi1358;
  assign n10944 = ~n10942 & ~n10943;
  assign n10945 = pi1331 & ~n9028;
  assign n10946 = pi1058 & pi3361;
  assign n10947 = ~n10945 & ~n10946;
  assign n10948 = pi0585 & pi1359;
  assign n10949 = n10947 & ~n10948;
  assign n10950 = n10944 & n10949;
  assign n10951 = n10941 & n10950;
  assign n10952 = pi3520 & ~n10410;
  assign n10953 = n10951 & ~n10952;
  assign n10954 = n9475 & ~n10953;
  assign n10955 = ~pi0979 & pi3084;
  assign n10956 = pi0979 & pi3159;
  assign n10957 = ~n10955 & ~n10956;
  assign n10958 = pi0763 & ~n10957;
  assign n10959 = ~pi0979 & pi2879;
  assign n10960 = pi0979 & pi3166;
  assign n10961 = ~n10959 & ~n10960;
  assign n10962 = pi0764 & ~n10961;
  assign n10963 = ~n10958 & ~n10962;
  assign n10964 = pi0088 & ~pi0979;
  assign n10965 = pi0086 & pi0979;
  assign n10966 = ~n10964 & ~n10965;
  assign n10967 = pi0720 & ~n10966;
  assign n10968 = pi0751 & ~pi0979;
  assign n10969 = pi0750 & pi0979;
  assign n10970 = ~n10968 & ~n10969;
  assign n10971 = pi0721 & ~n10970;
  assign n10972 = ~n10967 & ~n10971;
  assign n10973 = pi0050 & ~pi0979;
  assign n10974 = pi0049 & pi0979;
  assign n10975 = ~n10973 & ~n10974;
  assign n10976 = pi0719 & ~n10975;
  assign n10977 = ~pi0979 & pi2537;
  assign n10978 = pi0979 & pi3127;
  assign n10979 = ~n10977 & ~n10978;
  assign n10980 = pi0765 & ~n10979;
  assign n10981 = ~pi0979 & pi2897;
  assign n10982 = pi0979 & pi3202;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = pi0766 & ~n10983;
  assign n10985 = ~n10980 & ~n10984;
  assign n10986 = ~n10976 & n10985;
  assign n10987 = n10972 & n10986;
  assign n10988 = n10963 & n10987;
  assign n10989 = n9486 & ~n10988;
  assign n10990 = ~n10954 & ~n10989;
  assign n10991 = pi0979 & pi2176;
  assign n10992 = ~pi0979 & pi2938;
  assign n10993 = ~n10991 & ~n10992;
  assign n10994 = pi0836 & ~n10993;
  assign n10995 = ~pi0979 & pi2950;
  assign n10996 = pi0979 & pi2192;
  assign n10997 = ~n10995 & ~n10996;
  assign n10998 = pi0837 & ~n10997;
  assign n10999 = ~n10994 & ~n10998;
  assign n11000 = ~pi0979 & pi2929;
  assign n11001 = pi0979 & pi2158;
  assign n11002 = ~n11000 & ~n11001;
  assign n11003 = pi0767 & ~n11002;
  assign n11004 = pi0144 & ~pi0979;
  assign n11005 = pi0129 & pi0979;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = pi0768 & ~n11006;
  assign n11008 = ~n11003 & ~n11007;
  assign n11009 = pi0182 & ~pi0979;
  assign n11010 = pi0174 & pi0979;
  assign n11011 = ~n11009 & ~n11010;
  assign n11012 = pi0838 & ~n11011;
  assign n11013 = pi0149 & pi1360;
  assign n11014 = ~n11012 & ~n11013;
  assign n11015 = n11008 & n11014;
  assign n11016 = n10999 & n11015;
  assign n11017 = n9549 & ~n11016;
  assign n11018 = pi0266 & ~pi0979;
  assign n11019 = pi0262 & pi0979;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = pi0716 & ~n11020;
  assign n11022 = pi0333 & ~pi0979;
  assign n11023 = pi0332 & pi0979;
  assign n11024 = ~n11022 & ~n11023;
  assign n11025 = pi0718 & ~n11024;
  assign n11026 = ~n11021 & ~n11025;
  assign n11027 = pi0979 & pi2139;
  assign n11028 = ~pi0979 & pi2856;
  assign n11029 = ~n11027 & ~n11028;
  assign n11030 = pi0717 & ~n11029;
  assign n11031 = pi0208 & ~pi0979;
  assign n11032 = pi0205 & pi0979;
  assign n11033 = ~n11031 & ~n11032;
  assign n11034 = pi1599 & ~n11033;
  assign n11035 = ~n11030 & ~n11034;
  assign n11036 = pi0311 & ~pi0979;
  assign n11037 = pi0309 & pi0979;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = pi0761 & ~n11038;
  assign n11040 = n11035 & ~n11039;
  assign n11041 = n11026 & n11040;
  assign n11042 = n9523 & ~n11041;
  assign n11043 = ~n11017 & ~n11042;
  assign n11044 = pi1339 & pi2256;
  assign n11045 = pi1345 & pi2660;
  assign n11046 = ~n11044 & ~n11045;
  assign n11047 = pi1346 & pi2674;
  assign n11048 = n11046 & ~n11047;
  assign n11049 = pi1338 & pi2242;
  assign n11050 = n11048 & ~n11049;
  assign n11051 = pi1600 & pi2214;
  assign n11052 = pi1337 & pi2228;
  assign n11053 = ~n11051 & ~n11052;
  assign n11054 = pi1347 & pi2603;
  assign n11055 = pi1348 & pi2562;
  assign n11056 = ~n11054 & ~n11055;
  assign n11057 = pi1350 & pi2437;
  assign n11058 = n11056 & ~n11057;
  assign n11059 = pi1353 & pi1985;
  assign n11060 = n11058 & ~n11059;
  assign n11061 = pi1351 & pi2270;
  assign n11062 = pi1352 & pi2447;
  assign n11063 = ~n11061 & ~n11062;
  assign n11064 = n11060 & n11063;
  assign n11065 = n11053 & n11064;
  assign n11066 = n11050 & n11065;
  assign n11067 = n9577 & ~n11066;
  assign n11068 = pi1349 & pi2552;
  assign n11069 = pi1056 & pi2542;
  assign n11070 = ~n11068 & ~n11069;
  assign n11071 = pi1354 & pi2964;
  assign n11072 = n11070 & ~n11071;
  assign n11073 = pi1357 & pi2470;
  assign n11074 = n11072 & ~n11073;
  assign n11075 = pi1355 & pi2524;
  assign n11076 = pi1356 & pi2968;
  assign n11077 = ~n11075 & ~n11076;
  assign n11078 = pi1340 & pi2291;
  assign n11079 = pi1341 & pi2302;
  assign n11080 = ~n11078 & ~n11079;
  assign n11081 = pi1342 & pi2313;
  assign n11082 = n11080 & ~n11081;
  assign n11083 = pi1055 & pi2727;
  assign n11084 = n11082 & ~n11083;
  assign n11085 = pi1343 & pi2327;
  assign n11086 = pi1054 & pi2532;
  assign n11087 = ~n11085 & ~n11086;
  assign n11088 = n11084 & n11087;
  assign n11089 = n11077 & n11088;
  assign n11090 = n11074 & n11089;
  assign n11091 = n9736 & ~n11090;
  assign n11092 = ~n11067 & ~n11091;
  assign n11093 = pi0479 & pi1336;
  assign n11094 = pi0128 & pi1333;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = pi1332 & pi2582;
  assign n11097 = pi1335 & pi2597;
  assign n11098 = ~n11096 & ~n11097;
  assign n11099 = n11095 & n11098;
  assign n11100 = n9726 & ~n11099;
  assign n11101 = n9624 & n9627;
  assign n11102 = pi1012 & n11101;
  assign n11103 = pi0741 & n9715;
  assign n11104 = n9626 & n9642;
  assign n11105 = pi1033 & pi1034;
  assign n11106 = n11104 & n11105;
  assign n11107 = pi1738 & n11106;
  assign n11108 = pi0748 & n9707;
  assign n11109 = ~n11107 & ~n11108;
  assign n11110 = pi0795 & n9614;
  assign n11111 = pi1907 & n9618;
  assign n11112 = ~n11110 & ~n11111;
  assign n11113 = pi0805 & n9687;
  assign n11114 = pi1447 & n9691;
  assign n11115 = ~n11113 & ~n11114;
  assign n11116 = pi0967 & n9607;
  assign n11117 = n11115 & ~n11116;
  assign n11118 = n11112 & n11117;
  assign n11119 = pi1839 & n9698;
  assign n11120 = n11118 & ~n11119;
  assign n11121 = pi1873 & n9718;
  assign n11122 = pi0953 & n9702;
  assign n11123 = ~n11121 & ~n11122;
  assign n11124 = n11120 & n11123;
  assign n11125 = n11109 & n11124;
  assign n11126 = ~n11103 & n11125;
  assign n11127 = pi2110 & n9628;
  assign n11128 = pi1103 & n9631;
  assign n11129 = ~n11127 & ~n11128;
  assign n11130 = pi1769 & n9657;
  assign n11131 = pi1760 & n9659;
  assign n11132 = ~n11130 & ~n11131;
  assign n11133 = n9621 & n9690;
  assign n11134 = pi1434 & n11133;
  assign n11135 = pi0849 & n9682;
  assign n11136 = ~n11134 & ~n11135;
  assign n11137 = pi1726 & n9679;
  assign n11138 = n11136 & ~n11137;
  assign n11139 = pi1933 & n9622;
  assign n11140 = n11138 & ~n11139;
  assign n11141 = n11132 & n11140;
  assign n11142 = n11129 & n11141;
  assign n11143 = pi1786 & n9712;
  assign n11144 = n11142 & ~n11143;
  assign n11145 = n9621 & n9717;
  assign n11146 = pi1461 & n11145;
  assign n11147 = pi0873 & n9710;
  assign n11148 = ~n11146 & ~n11147;
  assign n11149 = n11144 & n11148;
  assign n11150 = n11126 & n11149;
  assign n11151 = pi0749 & n9670;
  assign n11152 = pi2059 & n9676;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 = pi0787 & n9654;
  assign n11155 = n9624 & n9665;
  assign n11156 = n9641 & n11155;
  assign n11157 = n9636 & n11156;
  assign n11158 = pi2112 & n11157;
  assign n11159 = pi2502 & n11158;
  assign n11160 = ~n11154 & ~n11159;
  assign n11161 = pi2990 & n9647;
  assign n11162 = n11160 & ~n11161;
  assign n11163 = n11153 & n11162;
  assign n11164 = pi1033 & n9626;
  assign n11165 = n9643 & n11164;
  assign n11166 = pi1945 & n11165;
  assign n11167 = n11163 & ~n11166;
  assign n11168 = n11150 & n11167;
  assign n11169 = ~n11102 & n11168;
  assign n11170 = pi1934 & ~n11169;
  assign n11171 = ~n11100 & ~n11170;
  assign n11172 = n11092 & n11171;
  assign n11173 = n11043 & n11172;
  assign n11174 = n10990 & n11173;
  assign n11175 = pi3316 & po3871;
  assign n11176 = n11174 & ~n11175;
  assign n11177 = ~pi1787 & ~n11176;
  assign n11178 = pi1787 & pi2836;
  assign n11179 = ~n11177 & ~n11178;
  assign n11180 = n9472 & ~n11179;
  assign n11181 = ~n10934 & ~n11180;
  assign n11182 = ~n10914 & ~n11181;
  assign n11183 = ~n10902 & n11182;
  assign n11184 = n9426 & n10909;
  assign n11185 = n10909 & n10912;
  assign n11186 = ~n11184 & ~n11185;
  assign n11187 = ~n9424 & ~n9842;
  assign n11188 = n9424 & ~n10384;
  assign n11189 = ~n11187 & ~n11188;
  assign n11190 = n10843 & n10844;
  assign n11191 = pi2530 & n11190;
  assign n11192 = n10835 & n10836;
  assign n11193 = pi2410 & n11192;
  assign n11194 = ~n11191 & ~n11193;
  assign n11195 = n10850 & n10851;
  assign n11196 = pi2458 & n11195;
  assign n11197 = n10825 & n10826;
  assign n11198 = pi2748 & n11197;
  assign n11199 = ~n11196 & ~n11198;
  assign n11200 = n11194 & n11199;
  assign n11201 = n9424 & ~n11200;
  assign n11202 = n10835 & n10859;
  assign n11203 = pi2410 & n11202;
  assign n11204 = n10843 & n10857;
  assign n11205 = pi2530 & n11204;
  assign n11206 = ~n11203 & ~n11205;
  assign n11207 = n10825 & n10863;
  assign n11208 = pi2748 & n11207;
  assign n11209 = n10850 & n10865;
  assign n11210 = pi2458 & n11209;
  assign n11211 = ~n11208 & ~n11210;
  assign n11212 = n11206 & n11211;
  assign n11213 = ~n9424 & ~n11212;
  assign n11214 = ~n11201 & ~n11213;
  assign n11215 = n11189 & n11214;
  assign n11216 = ~n11186 & ~n11215;
  assign n11217 = ~n10902 & n11216;
  assign n11218 = ~n11183 & ~n11217;
  assign n11219 = n10885 & ~n11218;
  assign n11220 = pi0656 & pi0707;
  assign n11221 = ~pi0645 & ~pi0646;
  assign n11222 = ~pi0675 & n11221;
  assign n11223 = ~pi0676 & n11222;
  assign n11224 = pi0668 & ~n11223;
  assign n11225 = pi0676 & ~n11222;
  assign n11226 = ~n11224 & ~n11225;
  assign n11227 = pi0675 & ~n11221;
  assign n11228 = pi0645 & pi0646;
  assign n11229 = ~n11227 & ~n11228;
  assign n11230 = ~pi0673 & ~pi0674;
  assign n11231 = ~pi0668 & ~pi0676;
  assign n11232 = n11222 & n11231;
  assign n11233 = ~pi0644 & ~pi0669;
  assign n11234 = n11232 & n11233;
  assign n11235 = ~pi0670 & ~pi0671;
  assign n11236 = n11234 & n11235;
  assign n11237 = ~pi0657 & ~pi0672;
  assign n11238 = n11236 & n11237;
  assign n11239 = n11230 & n11238;
  assign n11240 = pi0656 & ~n11239;
  assign n11241 = ~n11230 & ~n11238;
  assign n11242 = pi0673 & pi0674;
  assign n11243 = ~n11241 & ~n11242;
  assign n11244 = ~pi0672 & n11236;
  assign n11245 = pi0657 & ~n11244;
  assign n11246 = ~pi0670 & n11234;
  assign n11247 = pi0671 & ~n11246;
  assign n11248 = pi0672 & ~n11236;
  assign n11249 = ~n11247 & ~n11248;
  assign n11250 = ~n11245 & n11249;
  assign n11251 = n11243 & n11250;
  assign n11252 = ~n11240 & n11251;
  assign n11253 = ~n11232 & ~n11233;
  assign n11254 = pi0670 & ~n11234;
  assign n11255 = ~n11253 & ~n11254;
  assign n11256 = pi0644 & pi0669;
  assign n11257 = n11255 & ~n11256;
  assign n11258 = n11252 & n11257;
  assign n11259 = n11229 & n11258;
  assign n11260 = n11226 & n11259;
  assign n11261 = n11220 & n11260;
  assign n11262 = ~pi0656 & ~pi0673;
  assign n11263 = ~pi0657 & ~pi0674;
  assign n11264 = n11262 & n11263;
  assign n11265 = ~pi0671 & ~pi0672;
  assign n11266 = ~pi0670 & n11265;
  assign n11267 = n11264 & n11266;
  assign n11268 = ~pi0644 & ~pi0668;
  assign n11269 = ~pi0676 & n11268;
  assign n11270 = n11267 & n11269;
  assign n11271 = n11222 & n11270;
  assign n11272 = ~pi0669 & n11271;
  assign n11273 = ~n11260 & ~n11272;
  assign n11274 = ~pi0656 & n11260;
  assign n11275 = ~n11273 & ~n11274;
  assign n11276 = pi0707 & ~n11275;
  assign n11277 = pi0521 & n11276;
  assign n11278 = ~pi0521 & ~n11276;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = ~pi0668 & n11223;
  assign n11281 = ~pi0669 & ~pi0670;
  assign n11282 = ~pi0644 & n11281;
  assign n11283 = ~pi0657 & n11265;
  assign n11284 = ~pi0674 & n11262;
  assign n11285 = n11283 & n11284;
  assign n11286 = n11282 & n11285;
  assign n11287 = n11280 & n11286;
  assign n11288 = n11260 & ~n11287;
  assign n11289 = ~pi0645 & ~n11260;
  assign n11290 = ~n11288 & ~n11289;
  assign n11291 = pi0680 & n11290;
  assign n11292 = pi0518 & n11291;
  assign n11293 = ~pi0518 & ~pi0645;
  assign n11294 = pi0518 & pi0645;
  assign n11295 = ~n11293 & ~n11294;
  assign n11296 = ~pi0518 & ~n11291;
  assign n11297 = ~n11295 & ~n11296;
  assign n11298 = ~n11292 & ~n11297;
  assign n11299 = ~pi0675 & ~pi0676;
  assign n11300 = ~pi0668 & n11299;
  assign n11301 = n11283 & n11300;
  assign n11302 = n11284 & n11301;
  assign n11303 = ~pi0646 & n11302;
  assign n11304 = n11282 & n11303;
  assign n11305 = n11260 & ~n11304;
  assign n11306 = n11221 & ~n11260;
  assign n11307 = ~n11305 & ~n11306;
  assign n11308 = pi0681 & n11307;
  assign n11309 = ~pi0518 & ~pi0646;
  assign n11310 = pi0518 & pi0646;
  assign n11311 = ~n11309 & ~n11310;
  assign n11312 = ~pi0589 & n11311;
  assign n11313 = n11308 & ~n11312;
  assign n11314 = pi0589 & ~n11311;
  assign n11315 = ~n11313 & ~n11314;
  assign n11316 = ~n11292 & ~n11296;
  assign n11317 = ~n11295 & ~n11316;
  assign n11318 = n11295 & n11316;
  assign n11319 = ~n11317 & ~n11318;
  assign n11320 = ~n11315 & ~n11319;
  assign n11321 = n11282 & n11302;
  assign n11322 = n11260 & ~n11321;
  assign n11323 = n11222 & ~n11260;
  assign n11324 = ~n11322 & ~n11323;
  assign n11325 = pi0682 & n11324;
  assign n11326 = pi0519 & n11325;
  assign n11327 = ~pi0518 & ~pi0675;
  assign n11328 = pi0518 & pi0675;
  assign n11329 = ~n11327 & ~n11328;
  assign n11330 = ~pi0519 & ~n11325;
  assign n11331 = ~n11329 & ~n11330;
  assign n11332 = ~n11326 & ~n11331;
  assign n11333 = pi0589 & n11308;
  assign n11334 = ~pi0589 & ~n11308;
  assign n11335 = ~n11333 & ~n11334;
  assign n11336 = ~n11311 & ~n11335;
  assign n11337 = n11311 & n11335;
  assign n11338 = ~n11336 & ~n11337;
  assign n11339 = n11332 & n11338;
  assign n11340 = ~n11319 & ~n11339;
  assign n11341 = ~n11315 & ~n11332;
  assign n11342 = ~n11340 & ~n11341;
  assign n11343 = ~n11315 & ~n11338;
  assign n11344 = n11342 & ~n11343;
  assign n11345 = ~pi0669 & n11235;
  assign n11346 = n11269 & n11345;
  assign n11347 = ~pi0672 & n11263;
  assign n11348 = n11346 & n11347;
  assign n11349 = n11262 & n11348;
  assign n11350 = n11260 & ~n11349;
  assign n11351 = n11223 & ~n11260;
  assign n11352 = ~n11350 & ~n11351;
  assign n11353 = pi0683 & n11352;
  assign n11354 = pi0520 & n11353;
  assign n11355 = ~pi0518 & ~pi0676;
  assign n11356 = pi0518 & pi0676;
  assign n11357 = ~n11355 & ~n11356;
  assign n11358 = ~pi0520 & ~n11353;
  assign n11359 = ~n11357 & ~n11358;
  assign n11360 = ~n11354 & ~n11359;
  assign n11361 = ~n11326 & ~n11330;
  assign n11362 = ~n11329 & ~n11361;
  assign n11363 = n11329 & n11361;
  assign n11364 = ~n11362 & ~n11363;
  assign n11365 = ~n11360 & ~n11364;
  assign n11366 = ~n11354 & ~n11358;
  assign n11367 = ~n11357 & ~n11366;
  assign n11368 = n11357 & n11366;
  assign n11369 = ~n11367 & ~n11368;
  assign n11370 = n11266 & n11268;
  assign n11371 = ~pi0669 & n11370;
  assign n11372 = n11264 & n11371;
  assign n11373 = n11260 & ~n11372;
  assign n11374 = n11232 & ~n11260;
  assign n11375 = ~n11373 & ~n11374;
  assign n11376 = pi0701 & n11375;
  assign n11377 = pi0511 & n11376;
  assign n11378 = ~pi0518 & ~pi0668;
  assign n11379 = pi0518 & pi0668;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = ~pi0511 & ~n11376;
  assign n11382 = ~n11380 & ~n11381;
  assign n11383 = ~n11377 & ~n11382;
  assign n11384 = n11369 & n11383;
  assign n11385 = ~n11360 & ~n11384;
  assign n11386 = ~n11377 & ~n11381;
  assign n11387 = ~n11380 & n11386;
  assign n11388 = n11380 & ~n11386;
  assign n11389 = ~n11387 & ~n11388;
  assign n11390 = pi0518 & pi0644;
  assign n11391 = ~pi0518 & ~pi0644;
  assign n11392 = ~n11390 & ~n11391;
  assign n11393 = n11264 & n11265;
  assign n11394 = n11282 & n11393;
  assign n11395 = n11260 & ~n11394;
  assign n11396 = n11221 & n11299;
  assign n11397 = n11268 & n11396;
  assign n11398 = ~n11260 & n11397;
  assign n11399 = ~n11395 & ~n11398;
  assign n11400 = pi0677 & n11399;
  assign n11401 = ~pi0512 & ~n11400;
  assign n11402 = ~n11392 & ~n11401;
  assign n11403 = pi0512 & n11400;
  assign n11404 = ~n11402 & ~n11403;
  assign n11405 = n11389 & ~n11404;
  assign n11406 = n11385 & n11405;
  assign n11407 = ~n11364 & ~n11384;
  assign n11408 = ~n11389 & n11404;
  assign n11409 = ~pi0512 & n11400;
  assign n11410 = pi0512 & ~n11400;
  assign n11411 = ~n11409 & ~n11410;
  assign n11412 = ~n11392 & n11411;
  assign n11413 = n11392 & ~n11411;
  assign n11414 = ~n11412 & ~n11413;
  assign n11415 = n11281 & n11393;
  assign n11416 = n11260 & ~n11415;
  assign n11417 = n11234 & ~n11260;
  assign n11418 = ~n11416 & ~n11417;
  assign n11419 = pi0702 & n11418;
  assign n11420 = pi0587 & n11419;
  assign n11421 = ~pi0587 & ~n11419;
  assign n11422 = ~pi0518 & ~pi0669;
  assign n11423 = pi0518 & pi0669;
  assign n11424 = ~n11422 & ~n11423;
  assign n11425 = ~n11421 & ~n11424;
  assign n11426 = ~n11420 & ~n11425;
  assign n11427 = ~n11414 & ~n11426;
  assign n11428 = ~n11408 & n11427;
  assign n11429 = n11407 & n11428;
  assign n11430 = ~n11406 & ~n11429;
  assign n11431 = ~n11369 & ~n11383;
  assign n11432 = n11360 & n11364;
  assign n11433 = n11431 & ~n11432;
  assign n11434 = n11405 & n11407;
  assign n11435 = n11385 & n11428;
  assign n11436 = ~n11434 & ~n11435;
  assign n11437 = ~n11433 & n11436;
  assign n11438 = n11430 & n11437;
  assign n11439 = ~n11365 & n11438;
  assign n11440 = ~n11344 & ~n11439;
  assign n11441 = ~n11320 & ~n11440;
  assign n11442 = n11315 & n11319;
  assign n11443 = ~n11332 & ~n11442;
  assign n11444 = ~n11338 & n11443;
  assign n11445 = n11260 & ~n11262;
  assign n11446 = ~pi0673 & n11222;
  assign n11447 = n11348 & n11446;
  assign n11448 = ~n11260 & n11447;
  assign n11449 = ~n11445 & ~n11448;
  assign n11450 = pi0679 & n11449;
  assign n11451 = ~pi0518 & ~pi0673;
  assign n11452 = pi0518 & pi0673;
  assign n11453 = ~n11451 & ~n11452;
  assign n11454 = ~pi0517 & n11453;
  assign n11455 = n11450 & ~n11454;
  assign n11456 = pi0517 & ~n11453;
  assign n11457 = ~n11455 & ~n11456;
  assign n11458 = ~pi0518 & ~pi0674;
  assign n11459 = pi0518 & pi0674;
  assign n11460 = ~n11458 & ~n11459;
  assign n11461 = ~pi0656 & n11230;
  assign n11462 = n11260 & ~n11461;
  assign n11463 = n11222 & n11347;
  assign n11464 = n11346 & n11463;
  assign n11465 = ~n11260 & n11464;
  assign n11466 = ~n11462 & ~n11465;
  assign n11467 = pi0706 & n11466;
  assign n11468 = ~pi0516 & ~n11467;
  assign n11469 = pi0516 & n11467;
  assign n11470 = ~n11468 & ~n11469;
  assign n11471 = ~n11460 & ~n11470;
  assign n11472 = n11460 & n11470;
  assign n11473 = ~n11471 & ~n11472;
  assign n11474 = ~n11457 & ~n11473;
  assign n11475 = ~pi0518 & ~pi0657;
  assign n11476 = pi0518 & pi0657;
  assign n11477 = ~n11475 & ~n11476;
  assign n11478 = n11260 & ~n11264;
  assign n11479 = n11221 & n11282;
  assign n11480 = n11301 & n11479;
  assign n11481 = ~n11260 & n11480;
  assign n11482 = ~n11478 & ~n11481;
  assign n11483 = pi0705 & n11482;
  assign n11484 = ~pi0588 & ~n11483;
  assign n11485 = pi0588 & n11483;
  assign n11486 = ~n11484 & ~n11485;
  assign n11487 = ~n11477 & ~n11486;
  assign n11488 = n11477 & n11486;
  assign n11489 = ~n11487 & ~n11488;
  assign n11490 = ~n11460 & ~n11468;
  assign n11491 = ~n11469 & ~n11490;
  assign n11492 = n11489 & n11491;
  assign n11493 = n11474 & ~n11492;
  assign n11494 = ~pi0518 & ~pi0656;
  assign n11495 = pi0518 & pi0656;
  assign n11496 = ~n11494 & ~n11495;
  assign n11497 = ~pi0521 & n11496;
  assign n11498 = n11276 & ~n11497;
  assign n11499 = pi0521 & ~n11496;
  assign n11500 = ~n11498 & ~n11499;
  assign n11501 = ~pi0517 & n11450;
  assign n11502 = pi0517 & ~n11450;
  assign n11503 = ~n11501 & ~n11502;
  assign n11504 = ~n11453 & ~n11503;
  assign n11505 = n11453 & n11503;
  assign n11506 = ~n11504 & ~n11505;
  assign n11507 = ~n11500 & n11506;
  assign n11508 = ~n11279 & ~n11496;
  assign n11509 = n11279 & n11496;
  assign n11510 = ~n11508 & ~n11509;
  assign n11511 = ~pi0518 & ~n11510;
  assign n11512 = n11500 & ~n11506;
  assign n11513 = n11511 & ~n11512;
  assign n11514 = ~n11507 & ~n11513;
  assign n11515 = ~n11473 & ~n11491;
  assign n11516 = ~n11457 & ~n11491;
  assign n11517 = n11457 & n11473;
  assign n11518 = ~n11489 & ~n11517;
  assign n11519 = ~n11516 & ~n11518;
  assign n11520 = ~n11515 & n11519;
  assign n11521 = ~n11514 & ~n11520;
  assign n11522 = ~n11489 & ~n11491;
  assign n11523 = ~n11521 & ~n11522;
  assign n11524 = ~n11493 & n11523;
  assign n11525 = ~n11420 & ~n11421;
  assign n11526 = ~n11424 & ~n11525;
  assign n11527 = n11424 & n11525;
  assign n11528 = ~n11526 & ~n11527;
  assign n11529 = n11235 & n11237;
  assign n11530 = n11461 & n11529;
  assign n11531 = n11260 & ~n11530;
  assign n11532 = n11281 & n11397;
  assign n11533 = ~n11260 & n11532;
  assign n11534 = ~n11531 & ~n11533;
  assign n11535 = pi0703 & n11534;
  assign n11536 = pi0513 & n11535;
  assign n11537 = ~pi0513 & ~n11535;
  assign n11538 = ~pi0518 & ~pi0670;
  assign n11539 = pi0518 & pi0670;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = ~n11537 & ~n11540;
  assign n11542 = ~n11536 & ~n11541;
  assign n11543 = n11528 & n11542;
  assign n11544 = ~n11536 & ~n11537;
  assign n11545 = ~n11540 & n11544;
  assign n11546 = n11540 & ~n11544;
  assign n11547 = ~n11545 & ~n11546;
  assign n11548 = n11260 & ~n11393;
  assign n11549 = n11345 & n11397;
  assign n11550 = ~n11260 & n11549;
  assign n11551 = ~n11548 & ~n11550;
  assign n11552 = pi0678 & n11551;
  assign n11553 = pi0514 & n11552;
  assign n11554 = ~pi0518 & ~pi0671;
  assign n11555 = pi0518 & pi0671;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = ~pi0514 & ~n11552;
  assign n11558 = ~n11556 & ~n11557;
  assign n11559 = ~n11553 & ~n11558;
  assign n11560 = ~n11547 & n11559;
  assign n11561 = ~n11543 & ~n11560;
  assign n11562 = ~pi0518 & ~pi0672;
  assign n11563 = pi0518 & pi0672;
  assign n11564 = ~n11562 & ~n11563;
  assign n11565 = n11237 & n11284;
  assign n11566 = n11260 & ~n11565;
  assign n11567 = n11371 & n11396;
  assign n11568 = ~n11260 & n11567;
  assign n11569 = ~n11566 & ~n11568;
  assign n11570 = pi0704 & n11569;
  assign n11571 = ~pi0515 & n11570;
  assign n11572 = pi0515 & ~n11570;
  assign n11573 = ~n11571 & ~n11572;
  assign n11574 = ~n11564 & n11573;
  assign n11575 = n11564 & ~n11573;
  assign n11576 = ~n11574 & ~n11575;
  assign n11577 = ~n11477 & ~n11484;
  assign n11578 = ~n11485 & ~n11577;
  assign n11579 = n11576 & n11578;
  assign n11580 = ~pi0515 & ~n11570;
  assign n11581 = ~n11564 & ~n11580;
  assign n11582 = pi0515 & n11570;
  assign n11583 = ~n11581 & ~n11582;
  assign n11584 = ~n11553 & ~n11557;
  assign n11585 = ~n11556 & ~n11584;
  assign n11586 = n11556 & n11584;
  assign n11587 = ~n11585 & ~n11586;
  assign n11588 = n11583 & n11587;
  assign n11589 = ~n11579 & ~n11588;
  assign n11590 = n11561 & n11589;
  assign n11591 = ~n11524 & n11590;
  assign n11592 = ~n11576 & ~n11578;
  assign n11593 = n11583 & ~n11592;
  assign n11594 = ~n11587 & ~n11593;
  assign n11595 = ~n11576 & ~n11583;
  assign n11596 = ~n11578 & n11595;
  assign n11597 = ~n11594 & ~n11596;
  assign n11598 = n11561 & ~n11597;
  assign n11599 = ~n11528 & ~n11542;
  assign n11600 = ~n11598 & ~n11599;
  assign n11601 = n11547 & ~n11559;
  assign n11602 = ~n11543 & n11601;
  assign n11603 = n11600 & ~n11602;
  assign n11604 = ~n11591 & n11603;
  assign n11605 = n11414 & n11426;
  assign n11606 = ~n11408 & ~n11605;
  assign n11607 = ~n11604 & n11606;
  assign n11608 = ~n11385 & ~n11407;
  assign n11609 = n11607 & ~n11608;
  assign n11610 = ~n11344 & n11609;
  assign n11611 = ~n11444 & ~n11610;
  assign n11612 = n11441 & n11611;
  assign n11613 = ~n11298 & n11612;
  assign n11614 = n11298 & ~n11612;
  assign n11615 = ~n11613 & ~n11614;
  assign n11616 = ~n11279 & n11615;
  assign n11617 = pi0518 & n11510;
  assign n11618 = ~n11511 & ~n11617;
  assign n11619 = ~n11615 & ~n11618;
  assign n11620 = ~n11616 & ~n11619;
  assign n11621 = ~pi0518 & ~n11620;
  assign n11622 = ~n11330 & ~n11358;
  assign n11623 = ~n11421 & n11536;
  assign n11624 = ~n11421 & ~n11537;
  assign n11625 = ~n11557 & n11582;
  assign n11626 = ~n11553 & ~n11625;
  assign n11627 = n11624 & ~n11626;
  assign n11628 = ~n11623 & ~n11627;
  assign n11629 = n11469 & ~n11484;
  assign n11630 = ~pi0517 & ~n11450;
  assign n11631 = n11277 & ~n11630;
  assign n11632 = pi0517 & n11450;
  assign n11633 = ~n11631 & ~n11632;
  assign n11634 = n11467 & n11483;
  assign n11635 = pi0516 & pi0588;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = pi0516 & n11483;
  assign n11638 = n11636 & ~n11637;
  assign n11639 = pi0588 & n11467;
  assign n11640 = n11638 & ~n11639;
  assign n11641 = ~n11633 & ~n11640;
  assign n11642 = ~n11629 & ~n11641;
  assign n11643 = ~n11485 & n11642;
  assign n11644 = ~n11557 & ~n11580;
  assign n11645 = n11624 & n11644;
  assign n11646 = ~n11643 & n11645;
  assign n11647 = n11628 & ~n11646;
  assign n11648 = ~n11420 & n11647;
  assign n11649 = ~n11381 & ~n11401;
  assign n11650 = ~n11648 & n11649;
  assign n11651 = n11622 & n11650;
  assign n11652 = ~n11330 & n11354;
  assign n11653 = ~n11381 & n11403;
  assign n11654 = ~n11377 & ~n11653;
  assign n11655 = n11622 & ~n11654;
  assign n11656 = ~n11652 & ~n11655;
  assign n11657 = ~n11651 & n11656;
  assign n11658 = ~n11326 & n11657;
  assign n11659 = ~n11334 & ~n11658;
  assign n11660 = ~n11333 & ~n11659;
  assign n11661 = ~n11296 & ~n11660;
  assign n11662 = ~n11292 & ~n11661;
  assign n11663 = pi0518 & ~n11662;
  assign n11664 = ~pi0518 & n11662;
  assign n11665 = ~n11663 & ~n11664;
  assign n11666 = ~n11618 & n11665;
  assign n11667 = ~n11279 & ~n11665;
  assign n11668 = ~n11666 & ~n11667;
  assign n11669 = pi0518 & ~n11668;
  assign n11670 = ~n11621 & ~n11669;
  assign n11671 = pi0707 & ~n11260;
  assign n11672 = n11272 & n11671;
  assign n11673 = ~n11670 & ~n11672;
  assign n11674 = ~n11261 & n11673;
  assign n11675 = ~n11186 & ~n11674;
  assign n11676 = pi2524 & n11195;
  assign n11677 = pi2968 & n11190;
  assign n11678 = ~n11676 & ~n11677;
  assign n11679 = pi2470 & n11192;
  assign n11680 = pi2964 & n11197;
  assign n11681 = ~n11679 & ~n11680;
  assign n11682 = n11678 & n11681;
  assign n11683 = n9424 & ~n11682;
  assign n11684 = pi2964 & n11207;
  assign n11685 = pi2524 & n11209;
  assign n11686 = ~n11684 & ~n11685;
  assign n11687 = pi2470 & n11202;
  assign n11688 = pi2968 & n11204;
  assign n11689 = ~n11687 & ~n11688;
  assign n11690 = n11686 & n11689;
  assign n11691 = ~n9424 & ~n11690;
  assign n11692 = ~n11683 & ~n11691;
  assign n11693 = n11186 & ~n11692;
  assign n11694 = ~n11675 & ~n11693;
  assign n11695 = n10902 & ~n11694;
  assign n11696 = ~n10892 & ~n10901;
  assign n11697 = ~n10890 & n11696;
  assign n11698 = ~n10372 & ~n11186;
  assign n11699 = ~n10774 & ~n10781;
  assign n11700 = ~n8567 & ~n11699;
  assign n11701 = ~n10812 & n10816;
  assign n11702 = ~n11189 & n11701;
  assign n11703 = ~n8561 & n10744;
  assign n11704 = ~po3841 & n11703;
  assign n11705 = n9897 & ~n11704;
  assign n11706 = ~po3848 & n11705;
  assign n11707 = pi1035 & ~n11706;
  assign n11708 = ~n8565 & n8589;
  assign n11709 = pi1422 & n11708;
  assign n11710 = pi0909 & n11709;
  assign n11711 = ~n9851 & ~n11710;
  assign n11712 = ~n11707 & n11711;
  assign n11713 = ~n11702 & n11712;
  assign n11714 = n10752 & n10816;
  assign n11715 = pi0421 & n11714;
  assign n11716 = n10886 & ~n11214;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = n11713 & n11717;
  assign n11719 = ~n11700 & ~n11718;
  assign n11720 = pi0752 & n11700;
  assign n11721 = ~n11719 & ~n11720;
  assign n11722 = ~n10914 & ~n11721;
  assign n11723 = ~n11698 & ~n11722;
  assign n11724 = ~n11697 & ~n11723;
  assign n11725 = ~n11695 & ~n11724;
  assign n11726 = ~n10885 & ~n11725;
  assign n11727 = n9825 & ~n11186;
  assign n11728 = pi0680 & n11288;
  assign n11729 = ~n11320 & ~n11442;
  assign n11730 = n11439 & ~n11609;
  assign n11731 = ~n11339 & ~n11730;
  assign n11732 = ~n11332 & ~n11338;
  assign n11733 = ~n11731 & ~n11732;
  assign n11734 = ~n11729 & ~n11733;
  assign n11735 = n11729 & n11733;
  assign n11736 = ~n11734 & ~n11735;
  assign n11737 = n11665 & ~n11736;
  assign n11738 = ~n11316 & ~n11660;
  assign n11739 = n11316 & n11660;
  assign n11740 = ~n11738 & ~n11739;
  assign n11741 = ~n11665 & ~n11740;
  assign n11742 = ~n11737 & ~n11741;
  assign n11743 = pi0518 & ~n11742;
  assign n11744 = n11615 & ~n11740;
  assign n11745 = ~n11615 & ~n11736;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = ~pi0518 & ~n11746;
  assign n11748 = ~n11743 & ~n11747;
  assign n11749 = ~n11728 & n11748;
  assign n11750 = ~pi0645 & pi0680;
  assign n11751 = ~n11260 & n11750;
  assign n11752 = n11749 & ~n11751;
  assign n11753 = n11186 & n11752;
  assign n11754 = ~n11727 & ~n11753;
  assign n11755 = n10885 & n11697;
  assign n11756 = n11754 & n11755;
  assign n11757 = ~n11726 & ~n11756;
  assign po0229 = n11219 | ~n11757;
  assign n11759 = ~n10608 & n10914;
  assign n11760 = n11335 & ~n11658;
  assign n11761 = ~n11335 & n11658;
  assign n11762 = ~n11760 & ~n11761;
  assign n11763 = n11615 & ~n11762;
  assign n11764 = ~n11339 & ~n11732;
  assign n11765 = ~n11730 & n11764;
  assign n11766 = n11730 & ~n11764;
  assign n11767 = ~n11765 & ~n11766;
  assign n11768 = ~n11615 & ~n11767;
  assign n11769 = ~n11763 & ~n11768;
  assign n11770 = ~pi0518 & ~n11769;
  assign n11771 = n11665 & ~n11767;
  assign n11772 = ~n11665 & ~n11762;
  assign n11773 = ~n11771 & ~n11772;
  assign n11774 = pi0518 & ~n11773;
  assign n11775 = ~n11770 & ~n11774;
  assign n11776 = pi0681 & ~n11304;
  assign n11777 = n11260 & n11776;
  assign n11778 = ~n11775 & ~n11777;
  assign n11779 = pi0681 & n11221;
  assign n11780 = ~n11260 & n11779;
  assign n11781 = n11778 & ~n11780;
  assign n11782 = ~n10914 & ~n11781;
  assign n11783 = ~n11759 & ~n11782;
  assign n11784 = n11755 & ~n11783;
  assign n11785 = ~n10902 & ~n11186;
  assign n11786 = ~n9424 & ~n10616;
  assign n11787 = n9424 & ~n10661;
  assign n11788 = ~n11786 & ~n11787;
  assign n11789 = pi2525 & n11195;
  assign n11790 = pi2755 & n11190;
  assign n11791 = ~n11789 & ~n11790;
  assign n11792 = pi2467 & n11192;
  assign n11793 = pi2533 & n11197;
  assign n11794 = ~n11792 & ~n11793;
  assign n11795 = n11791 & n11794;
  assign n11796 = n9424 & ~n11795;
  assign n11797 = pi2755 & n11204;
  assign n11798 = pi2525 & n11209;
  assign n11799 = ~n11797 & ~n11798;
  assign n11800 = pi2533 & n11207;
  assign n11801 = pi2467 & n11202;
  assign n11802 = ~n11800 & ~n11801;
  assign n11803 = n11799 & n11802;
  assign n11804 = ~n9424 & ~n11803;
  assign n11805 = ~n11796 & ~n11804;
  assign n11806 = n11788 & n11805;
  assign n11807 = n11785 & ~n11806;
  assign n11808 = pi0979 & pi2185;
  assign n11809 = ~pi0979 & pi2783;
  assign n11810 = ~n11808 & ~n11809;
  assign n11811 = pi0837 & ~n11810;
  assign n11812 = ~pi0979 & pi2935;
  assign n11813 = pi0979 & pi2169;
  assign n11814 = ~n11812 & ~n11813;
  assign n11815 = pi0836 & ~n11814;
  assign n11816 = ~n11811 & ~n11815;
  assign n11817 = pi0176 & ~pi0979;
  assign n11818 = pi0161 & pi0979;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = pi0838 & ~n11819;
  assign n11821 = pi0134 & pi1360;
  assign n11822 = ~n11820 & ~n11821;
  assign n11823 = pi0979 & pi2151;
  assign n11824 = ~pi0979 & pi2923;
  assign n11825 = ~n11823 & ~n11824;
  assign n11826 = pi0767 & ~n11825;
  assign n11827 = ~pi0979 & pi2159;
  assign n11828 = pi0979 & pi1790;
  assign n11829 = ~n11827 & ~n11828;
  assign n11830 = pi0768 & ~n11829;
  assign n11831 = ~n11826 & ~n11830;
  assign n11832 = n11822 & n11831;
  assign n11833 = n11816 & n11832;
  assign n11834 = n9549 & ~n11833;
  assign n11835 = pi0292 & ~pi0979;
  assign n11836 = pi0289 & pi0979;
  assign n11837 = ~n11835 & ~n11836;
  assign n11838 = pi0761 & ~n11837;
  assign n11839 = pi0395 & ~pi0979;
  assign n11840 = pi0394 & pi0979;
  assign n11841 = ~n11839 & ~n11840;
  assign n11842 = pi0718 & ~n11841;
  assign n11843 = ~n11838 & ~n11842;
  assign n11844 = pi0979 & pi2132;
  assign n11845 = ~pi0979 & pi2849;
  assign n11846 = ~n11844 & ~n11845;
  assign n11847 = pi0717 & ~n11846;
  assign n11848 = pi0206 & ~pi0979;
  assign n11849 = pi0202 & pi0979;
  assign n11850 = ~n11848 & ~n11849;
  assign n11851 = pi1599 & ~n11850;
  assign n11852 = ~n11847 & ~n11851;
  assign n11853 = pi0307 & ~pi0979;
  assign n11854 = pi0305 & pi0979;
  assign n11855 = ~n11853 & ~n11854;
  assign n11856 = pi0716 & ~n11855;
  assign n11857 = n11852 & ~n11856;
  assign n11858 = n11843 & n11857;
  assign n11859 = n9523 & ~n11858;
  assign n11860 = ~n11834 & ~n11859;
  assign n11861 = pi0370 & pi1336;
  assign n11862 = pi0073 & pi1333;
  assign n11863 = ~n11861 & ~n11862;
  assign n11864 = pi1332 & pi2575;
  assign n11865 = pi1335 & pi2590;
  assign n11866 = ~n11864 & ~n11865;
  assign n11867 = n11863 & n11866;
  assign n11868 = n9726 & ~n11867;
  assign n11869 = pi2986 & n9647;
  assign n11870 = pi0733 & n9654;
  assign n11871 = ~n11869 & ~n11870;
  assign n11872 = pi0778 & n9670;
  assign n11873 = pi2061 & n9676;
  assign n11874 = ~n11872 & ~n11873;
  assign n11875 = pi2499 & n11158;
  assign n11876 = n11874 & ~n11875;
  assign n11877 = n11871 & n11876;
  assign n11878 = pi1944 & n11165;
  assign n11879 = n11877 & ~n11878;
  assign n11880 = pi1433 & n11133;
  assign n11881 = pi0699 & n9682;
  assign n11882 = ~n11880 & ~n11881;
  assign n11883 = pi1721 & n9679;
  assign n11884 = n11882 & ~n11883;
  assign n11885 = pi1927 & n9622;
  assign n11886 = n11884 & ~n11885;
  assign n11887 = pi0739 & n9715;
  assign n11888 = pi1735 & n11106;
  assign n11889 = pi0747 & n9707;
  assign n11890 = ~n11888 & ~n11889;
  assign n11891 = pi1853 & n9698;
  assign n11892 = pi1862 & n9718;
  assign n11893 = pi0952 & n9702;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = ~n11891 & n11894;
  assign n11896 = n11890 & n11895;
  assign n11897 = ~n11887 & n11896;
  assign n11898 = pi0804 & n9687;
  assign n11899 = pi1444 & n9691;
  assign n11900 = ~n11898 & ~n11899;
  assign n11901 = pi0793 & n9614;
  assign n11902 = pi2052 & n9618;
  assign n11903 = ~n11901 & ~n11902;
  assign n11904 = pi0966 & n9607;
  assign n11905 = n11903 & ~n11904;
  assign n11906 = n11900 & n11905;
  assign n11907 = n11897 & n11906;
  assign n11908 = pi2108 & n9628;
  assign n11909 = pi1757 & n9659;
  assign n11910 = ~n11908 & ~n11909;
  assign n11911 = pi1023 & n9631;
  assign n11912 = pi1767 & n9657;
  assign n11913 = ~n11911 & ~n11912;
  assign n11914 = n11910 & n11913;
  assign n11915 = n11907 & n11914;
  assign n11916 = n11886 & n11915;
  assign n11917 = pi1780 & n9712;
  assign n11918 = n11916 & ~n11917;
  assign n11919 = pi1458 & n11145;
  assign n11920 = pi0908 & n9710;
  assign n11921 = ~n11919 & ~n11920;
  assign n11922 = n11918 & n11921;
  assign n11923 = ~n11102 & n11922;
  assign n11924 = n11879 & n11923;
  assign n11925 = pi1934 & ~n11924;
  assign n11926 = ~n11868 & ~n11925;
  assign n11927 = pi0210 & ~pi0979;
  assign n11928 = pi0209 & pi0979;
  assign n11929 = ~n11927 & ~n11928;
  assign n11930 = pi0720 & ~n11929;
  assign n11931 = pi0584 & ~pi0979;
  assign n11932 = pi0583 & pi0979;
  assign n11933 = ~n11931 & ~n11932;
  assign n11934 = pi0721 & ~n11933;
  assign n11935 = ~n11930 & ~n11934;
  assign n11936 = ~pi0979 & pi2781;
  assign n11937 = pi0979 & pi3157;
  assign n11938 = ~n11936 & ~n11937;
  assign n11939 = pi0763 & ~n11938;
  assign n11940 = ~pi0979 & pi2876;
  assign n11941 = pi0979 & pi3165;
  assign n11942 = ~n11940 & ~n11941;
  assign n11943 = pi0764 & ~n11942;
  assign n11944 = ~n11939 & ~n11943;
  assign n11945 = pi0047 & ~pi0979;
  assign n11946 = pi0046 & pi0979;
  assign n11947 = ~n11945 & ~n11946;
  assign n11948 = pi0719 & ~n11947;
  assign n11949 = ~pi0979 & pi2637;
  assign n11950 = pi0979 & pi3128;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = pi0765 & ~n11951;
  assign n11953 = ~pi0979 & pi2893;
  assign n11954 = pi0979 & pi3123;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = pi0766 & ~n11955;
  assign n11957 = ~n11952 & ~n11956;
  assign n11958 = ~n11948 & n11957;
  assign n11959 = n11944 & n11958;
  assign n11960 = n11935 & n11959;
  assign n11961 = n9486 & ~n11960;
  assign n11962 = n11926 & ~n11961;
  assign n11963 = n11860 & n11962;
  assign n11964 = pi1334 & pi2766;
  assign n11965 = pi0830 & pi1344;
  assign n11966 = ~n11964 & ~n11965;
  assign n11967 = pi1331 & ~n8802;
  assign n11968 = pi1058 & pi3360;
  assign n11969 = ~n11967 & ~n11968;
  assign n11970 = pi0632 & pi1359;
  assign n11971 = n11969 & ~n11970;
  assign n11972 = pi3511 & ~n10410;
  assign n11973 = n11971 & ~n11972;
  assign n11974 = pi0390 & pi1057;
  assign n11975 = pi1059 & pi2980;
  assign n11976 = ~n11974 & ~n11975;
  assign n11977 = pi1053 & pi2400;
  assign n11978 = n11976 & ~n11977;
  assign n11979 = pi0919 & pi1358;
  assign n11980 = n11978 & ~n11979;
  assign n11981 = n11973 & n11980;
  assign n11982 = n11966 & n11981;
  assign n11983 = n9475 & ~n11982;
  assign n11984 = n11963 & ~n11983;
  assign n11985 = pi1340 & pi2068;
  assign n11986 = pi1341 & pi2299;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = pi1342 & pi2308;
  assign n11989 = n11987 & ~n11988;
  assign n11990 = pi1055 & pi2773;
  assign n11991 = n11989 & ~n11990;
  assign n11992 = pi1343 & pi2322;
  assign n11993 = pi1054 & pi2715;
  assign n11994 = ~n11992 & ~n11993;
  assign n11995 = pi1349 & pi2734;
  assign n11996 = pi1056 & pi2743;
  assign n11997 = ~n11995 & ~n11996;
  assign n11998 = pi1354 & pi2747;
  assign n11999 = n11997 & ~n11998;
  assign n12000 = pi1357 & pi2466;
  assign n12001 = n11999 & ~n12000;
  assign n12002 = pi1355 & pi2457;
  assign n12003 = pi1356 & pi2754;
  assign n12004 = ~n12002 & ~n12003;
  assign n12005 = n12001 & n12004;
  assign n12006 = n11994 & n12005;
  assign n12007 = n11991 & n12006;
  assign n12008 = n9736 & ~n12007;
  assign n12009 = pi1351 & pi2267;
  assign n12010 = pi1352 & pi2444;
  assign n12011 = ~n12009 & ~n12010;
  assign n12012 = pi1353 & pi1982;
  assign n12013 = n12011 & ~n12012;
  assign n12014 = pi1350 & pi2434;
  assign n12015 = n12013 & ~n12014;
  assign n12016 = pi1347 & pi2683;
  assign n12017 = pi1348 & pi2693;
  assign n12018 = ~n12016 & ~n12017;
  assign n12019 = pi1600 & pi2209;
  assign n12020 = pi1337 & pi2223;
  assign n12021 = ~n12019 & ~n12020;
  assign n12022 = pi1338 & pi2237;
  assign n12023 = n12021 & ~n12022;
  assign n12024 = pi1346 & pi2669;
  assign n12025 = n12023 & ~n12024;
  assign n12026 = pi1339 & pi2251;
  assign n12027 = pi1345 & pi2655;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = n12025 & n12028;
  assign n12030 = n12018 & n12029;
  assign n12031 = n12015 & n12030;
  assign n12032 = n9577 & ~n12031;
  assign n12033 = ~n12008 & ~n12032;
  assign n12034 = n11984 & n12033;
  assign n12035 = pi3312 & po3871;
  assign n12036 = n12034 & ~n12035;
  assign n12037 = ~pi1787 & ~n12036;
  assign n12038 = pi1787 & pi2831;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = n9472 & ~n12039;
  assign n12041 = pi3860 & n9804;
  assign n12042 = pi3876 & n9774;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = pi3844 & n9802;
  assign n12045 = pi3972 & n9783;
  assign n12046 = pi3892 & n9771;
  assign n12047 = ~n12045 & ~n12046;
  assign n12048 = pi3940 & n9791;
  assign n12049 = pi3924 & n9788;
  assign n12050 = ~n12048 & ~n12049;
  assign n12051 = n12047 & n12050;
  assign n12052 = ~n12044 & n12051;
  assign n12053 = n12043 & n12052;
  assign n12054 = pi3860 & n9799;
  assign n12055 = n12053 & ~n12054;
  assign n12056 = pi3908 & n9781;
  assign n12057 = pi3956 & n9793;
  assign n12058 = ~n12056 & ~n12057;
  assign n12059 = n12055 & n12058;
  assign n12060 = ~n9472 & ~n12059;
  assign n12061 = ~n12040 & ~n12060;
  assign n12062 = ~n10914 & ~n12061;
  assign n12063 = ~n11697 & n12062;
  assign n12064 = ~n11807 & ~n12063;
  assign n12065 = n10885 & ~n12064;
  assign n12066 = ~n10653 & ~n11186;
  assign n12067 = n10886 & ~n11805;
  assign n12068 = pi0819 & n11709;
  assign n12069 = ~n10622 & ~n12068;
  assign n12070 = pi0405 & n11714;
  assign n12071 = n12069 & ~n12070;
  assign n12072 = n11701 & ~n11788;
  assign n12073 = pi1036 & ~n11706;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = n12071 & n12074;
  assign n12076 = ~n11700 & n12075;
  assign n12077 = ~n12067 & n12076;
  assign n12078 = ~pi0779 & n11700;
  assign n12079 = ~n12077 & ~n12078;
  assign n12080 = ~n10914 & n12079;
  assign n12081 = ~n12066 & ~n12080;
  assign n12082 = ~n10902 & ~n12081;
  assign n12083 = n11277 & n11503;
  assign n12084 = ~n11277 & ~n11503;
  assign n12085 = ~n12083 & ~n12084;
  assign n12086 = n11615 & ~n12085;
  assign n12087 = ~n11500 & ~n11506;
  assign n12088 = n11500 & n11506;
  assign n12089 = ~n12087 & ~n12088;
  assign n12090 = n11511 & n12089;
  assign n12091 = ~n11511 & ~n12089;
  assign n12092 = ~n12090 & ~n12091;
  assign n12093 = ~n11615 & ~n12092;
  assign n12094 = ~n12086 & ~n12093;
  assign n12095 = ~pi0518 & ~n12094;
  assign n12096 = n11665 & ~n12092;
  assign n12097 = ~n11665 & ~n12085;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = pi0518 & ~n12098;
  assign n12100 = ~n12095 & ~n12099;
  assign n12101 = pi0679 & ~n11262;
  assign n12102 = n11260 & n12101;
  assign n12103 = n12100 & ~n12102;
  assign n12104 = pi0679 & n11447;
  assign n12105 = ~n11260 & n12104;
  assign n12106 = n12103 & ~n12105;
  assign n12107 = ~n11186 & n12106;
  assign n12108 = pi2457 & n11195;
  assign n12109 = pi2747 & n11197;
  assign n12110 = ~n12108 & ~n12109;
  assign n12111 = pi2754 & n11190;
  assign n12112 = pi2466 & n11192;
  assign n12113 = ~n12111 & ~n12112;
  assign n12114 = n12110 & n12113;
  assign n12115 = n9424 & ~n12114;
  assign n12116 = pi2747 & n11207;
  assign n12117 = pi2754 & n11204;
  assign n12118 = ~n12116 & ~n12117;
  assign n12119 = pi2466 & n11202;
  assign n12120 = pi2457 & n11209;
  assign n12121 = ~n12119 & ~n12120;
  assign n12122 = n12118 & n12121;
  assign n12123 = ~n9424 & ~n12122;
  assign n12124 = ~n12115 & ~n12123;
  assign n12125 = n11186 & n12124;
  assign n12126 = ~n12107 & ~n12125;
  assign n12127 = n10902 & n12126;
  assign n12128 = ~n12082 & ~n12127;
  assign n12129 = ~n10885 & ~n12128;
  assign n12130 = ~n12065 & ~n12129;
  assign po0228 = n11784 | ~n12130;
  assign n12132 = pi2452 & n11195;
  assign n12133 = pi2413 & n11192;
  assign n12134 = ~n12132 & ~n12133;
  assign n12135 = pi2965 & n11190;
  assign n12136 = pi2960 & n11197;
  assign n12137 = ~n12135 & ~n12136;
  assign n12138 = n12134 & n12137;
  assign n12139 = n9424 & ~n12138;
  assign n12140 = pi2413 & n11202;
  assign n12141 = pi2452 & n11209;
  assign n12142 = ~n12140 & ~n12141;
  assign n12143 = pi2960 & n11207;
  assign n12144 = pi2965 & n11204;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = n12142 & n12145;
  assign n12147 = ~n9424 & ~n12146;
  assign n12148 = ~n12139 & ~n12147;
  assign n12149 = pi2257 & n9837;
  assign n12150 = pi2271 & n9834;
  assign n12151 = ~n12149 & ~n12150;
  assign n12152 = pi2261 & n9839;
  assign n12153 = pi1976 & n9832;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = n12151 & n12154;
  assign n12156 = ~n9424 & ~n12155;
  assign n12157 = pi2257 & n10374;
  assign n12158 = pi1976 & n10379;
  assign n12159 = ~n12157 & ~n12158;
  assign n12160 = pi2261 & n10376;
  assign n12161 = pi2271 & n10381;
  assign n12162 = ~n12160 & ~n12161;
  assign n12163 = n12159 & n12162;
  assign n12164 = n9424 & ~n12163;
  assign n12165 = ~n12156 & ~n12164;
  assign n12166 = n12148 & n12165;
  assign n12167 = n11785 & ~n12166;
  assign n12168 = pi3863 & n9804;
  assign n12169 = pi3879 & n9774;
  assign n12170 = ~n12168 & ~n12169;
  assign n12171 = pi3847 & n9802;
  assign n12172 = pi3911 & n9781;
  assign n12173 = pi3895 & n9771;
  assign n12174 = ~n12172 & ~n12173;
  assign n12175 = pi3943 & n9791;
  assign n12176 = pi3927 & n9788;
  assign n12177 = ~n12175 & ~n12176;
  assign n12178 = n12174 & n12177;
  assign n12179 = ~n12171 & n12178;
  assign n12180 = n12170 & n12179;
  assign n12181 = pi3863 & n9799;
  assign n12182 = n12180 & ~n12181;
  assign n12183 = pi3975 & n9783;
  assign n12184 = pi3959 & n9793;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186 = n12182 & n12185;
  assign n12187 = ~n9472 & ~n12186;
  assign n12188 = pi0387 & pi1057;
  assign n12189 = pi1053 & pi2405;
  assign n12190 = ~n12188 & ~n12189;
  assign n12191 = pi0917 & pi1358;
  assign n12192 = n12190 & ~n12191;
  assign n12193 = pi1334 & pi2380;
  assign n12194 = pi0868 & pi1344;
  assign n12195 = ~n12193 & ~n12194;
  assign n12196 = pi1331 & ~n8950;
  assign n12197 = pi1058 & pi3293;
  assign n12198 = ~n12196 & ~n12197;
  assign n12199 = pi0591 & pi1359;
  assign n12200 = n12198 & ~n12199;
  assign n12201 = n12195 & n12200;
  assign n12202 = n12192 & n12201;
  assign n12203 = pi3509 & ~n10410;
  assign n12204 = n12202 & ~n12203;
  assign n12205 = n9475 & ~n12204;
  assign n12206 = pi0495 & ~pi0979;
  assign n12207 = pi0494 & pi0979;
  assign n12208 = ~n12206 & ~n12207;
  assign n12209 = pi0718 & ~n12208;
  assign n12210 = ~pi0979 & pi2846;
  assign n12211 = pi0979 & pi2129;
  assign n12212 = ~n12210 & ~n12211;
  assign n12213 = pi0717 & ~n12212;
  assign n12214 = ~n12209 & ~n12213;
  assign n12215 = pi0270 & ~pi0979;
  assign n12216 = pi0269 & pi0979;
  assign n12217 = ~n12215 & ~n12216;
  assign n12218 = pi0716 & ~n12217;
  assign n12219 = pi0319 & ~pi0979;
  assign n12220 = pi0317 & pi0979;
  assign n12221 = ~n12219 & ~n12220;
  assign n12222 = pi0761 & ~n12221;
  assign n12223 = ~n12218 & ~n12222;
  assign n12224 = n12214 & n12223;
  assign n12225 = ~n9535 & n12224;
  assign n12226 = n9523 & ~n12225;
  assign n12227 = ~n12205 & ~n12226;
  assign n12228 = pi0979 & pi2166;
  assign n12229 = ~pi0979 & pi2933;
  assign n12230 = ~n12228 & ~n12229;
  assign n12231 = pi0836 & ~n12230;
  assign n12232 = ~pi0979 & pi2943;
  assign n12233 = pi0979 & pi2182;
  assign n12234 = ~n12232 & ~n12233;
  assign n12235 = pi0837 & ~n12234;
  assign n12236 = ~n12231 & ~n12235;
  assign n12237 = pi0979 & pi2148;
  assign n12238 = ~pi0979 & pi2920;
  assign n12239 = ~n12237 & ~n12238;
  assign n12240 = pi0767 & ~n12239;
  assign n12241 = ~pi0979 & pi2425;
  assign n12242 = pi0979 & pi1960;
  assign n12243 = ~n12241 & ~n12242;
  assign n12244 = pi0768 & ~n12243;
  assign n12245 = ~n12240 & ~n12244;
  assign n12246 = pi0172 & ~pi0979;
  assign n12247 = pi0158 & pi0979;
  assign n12248 = ~n12246 & ~n12247;
  assign n12249 = pi0838 & ~n12248;
  assign n12250 = pi0659 & pi1360;
  assign n12251 = ~n12249 & ~n12250;
  assign n12252 = n12245 & n12251;
  assign n12253 = n12236 & n12252;
  assign n12254 = n9549 & ~n12253;
  assign n12255 = pi0065 & ~pi0979;
  assign n12256 = pi0063 & pi0979;
  assign n12257 = ~n12255 & ~n12256;
  assign n12258 = pi0719 & ~n12257;
  assign n12259 = ~pi0979 & pi2635;
  assign n12260 = pi0979 & pi3132;
  assign n12261 = ~n12259 & ~n12260;
  assign n12262 = pi0765 & ~n12261;
  assign n12263 = ~pi0979 & pi3059;
  assign n12264 = pi0979 & pi3180;
  assign n12265 = ~n12263 & ~n12264;
  assign n12266 = pi0766 & ~n12265;
  assign n12267 = ~n12262 & ~n12266;
  assign n12268 = pi0186 & ~pi0979;
  assign n12269 = pi0185 & pi0979;
  assign n12270 = ~n12268 & ~n12269;
  assign n12271 = pi0720 & ~n12270;
  assign n12272 = pi0345 & ~pi0979;
  assign n12273 = pi0344 & pi0979;
  assign n12274 = ~n12272 & ~n12273;
  assign n12275 = pi0721 & ~n12274;
  assign n12276 = ~n12271 & ~n12275;
  assign n12277 = ~pi0979 & pi2782;
  assign n12278 = pi0979 & pi3154;
  assign n12279 = ~n12277 & ~n12278;
  assign n12280 = pi0763 & ~n12279;
  assign n12281 = ~pi0979 & pi2873;
  assign n12282 = pi0979 & pi3201;
  assign n12283 = ~n12281 & ~n12282;
  assign n12284 = pi0764 & ~n12283;
  assign n12285 = ~n12280 & ~n12284;
  assign n12286 = n12276 & n12285;
  assign n12287 = n12267 & n12286;
  assign n12288 = ~n12258 & n12287;
  assign n12289 = n9486 & ~n12288;
  assign n12290 = ~n12254 & ~n12289;
  assign n12291 = pi1343 & pi2319;
  assign n12292 = pi1054 & pi2712;
  assign n12293 = ~n12291 & ~n12292;
  assign n12294 = pi1055 & pi2722;
  assign n12295 = n12293 & ~n12294;
  assign n12296 = pi1342 & pi2087;
  assign n12297 = n12295 & ~n12296;
  assign n12298 = pi1340 & pi2284;
  assign n12299 = pi1341 & pi2296;
  assign n12300 = ~n12298 & ~n12299;
  assign n12301 = pi1355 & pi2455;
  assign n12302 = pi1356 & pi2966;
  assign n12303 = ~n12301 & ~n12302;
  assign n12304 = pi1357 & pi2464;
  assign n12305 = n12303 & ~n12304;
  assign n12306 = pi1354 & pi2963;
  assign n12307 = n12305 & ~n12306;
  assign n12308 = pi1349 & pi2732;
  assign n12309 = pi1056 & pi2546;
  assign n12310 = ~n12308 & ~n12309;
  assign n12311 = n12307 & n12310;
  assign n12312 = n12300 & n12311;
  assign n12313 = n12297 & n12312;
  assign n12314 = n9736 & ~n12313;
  assign n12315 = pi1347 & pi2680;
  assign n12316 = pi1348 & pi2690;
  assign n12317 = ~n12315 & ~n12316;
  assign n12318 = pi1350 & pi2259;
  assign n12319 = n12317 & ~n12318;
  assign n12320 = pi1353 & pi1979;
  assign n12321 = n12319 & ~n12320;
  assign n12322 = pi1351 & pi2264;
  assign n12323 = pi1352 & pi2273;
  assign n12324 = ~n12322 & ~n12323;
  assign n12325 = pi1600 & pi2206;
  assign n12326 = pi1337 & pi2220;
  assign n12327 = ~n12325 & ~n12326;
  assign n12328 = pi1338 & pi2234;
  assign n12329 = n12327 & ~n12328;
  assign n12330 = pi1346 & pi2666;
  assign n12331 = n12329 & ~n12330;
  assign n12332 = pi1339 & pi2248;
  assign n12333 = pi1345 & pi2652;
  assign n12334 = ~n12332 & ~n12333;
  assign n12335 = n12331 & n12334;
  assign n12336 = n12324 & n12335;
  assign n12337 = n12321 & n12336;
  assign n12338 = n9577 & ~n12337;
  assign n12339 = ~n12314 & ~n12338;
  assign n12340 = pi0329 & pi1336;
  assign n12341 = pi0330 & pi1333;
  assign n12342 = ~n12340 & ~n12341;
  assign n12343 = pi1332 & pi2572;
  assign n12344 = pi1335 & pi2587;
  assign n12345 = ~n12343 & ~n12344;
  assign n12346 = n12342 & n12345;
  assign n12347 = n9726 & ~n12346;
  assign n12348 = pi0883 & n9715;
  assign n12349 = pi1886 & n9718;
  assign n12350 = ~n12348 & ~n12349;
  assign n12351 = pi1732 & n11106;
  assign n12352 = pi0745 & n9707;
  assign n12353 = ~n12351 & ~n12352;
  assign n12354 = pi0951 & n9702;
  assign n12355 = n12353 & ~n12354;
  assign n12356 = n12350 & n12355;
  assign n12357 = pi1833 & n9698;
  assign n12358 = n12356 & ~n12357;
  assign n12359 = pi1017 & n9614;
  assign n12360 = pi1900 & n9618;
  assign n12361 = ~n12359 & ~n12360;
  assign n12362 = pi0900 & n9607;
  assign n12363 = n12361 & ~n12362;
  assign n12364 = pi0850 & n9687;
  assign n12365 = pi1441 & n9691;
  assign n12366 = ~n12364 & ~n12365;
  assign n12367 = n12363 & n12366;
  assign n12368 = pi0782 & n9654;
  assign n12369 = pi2513 & n11158;
  assign n12370 = ~n12368 & ~n12369;
  assign n12371 = pi0775 & n9670;
  assign n12372 = pi1467 & n9676;
  assign n12373 = ~n12371 & ~n12372;
  assign n12374 = pi2505 & n9647;
  assign n12375 = n12373 & ~n12374;
  assign n12376 = n12370 & n12375;
  assign n12377 = pi1941 & n11165;
  assign n12378 = n12376 & ~n12377;
  assign n12379 = pi2106 & n9628;
  assign n12380 = pi1100 & n9631;
  assign n12381 = ~n12379 & ~n12380;
  assign n12382 = pi1765 & n9657;
  assign n12383 = pi1754 & n9659;
  assign n12384 = ~n12382 & ~n12383;
  assign n12385 = n12381 & n12384;
  assign n12386 = pi1430 & n11133;
  assign n12387 = pi0863 & n9682;
  assign n12388 = ~n12386 & ~n12387;
  assign n12389 = pi1718 & n9679;
  assign n12390 = n12388 & ~n12389;
  assign n12391 = pi1924 & n9622;
  assign n12392 = n12390 & ~n12391;
  assign n12393 = n12385 & n12392;
  assign n12394 = ~n11102 & n12393;
  assign n12395 = n12378 & n12394;
  assign n12396 = pi1777 & n9712;
  assign n12397 = n12395 & ~n12396;
  assign n12398 = pi1455 & n11145;
  assign n12399 = pi0906 & n9710;
  assign n12400 = ~n12398 & ~n12399;
  assign n12401 = n12397 & n12400;
  assign n12402 = n12367 & n12401;
  assign n12403 = n12358 & n12402;
  assign n12404 = pi1934 & ~n12403;
  assign n12405 = ~n12347 & ~n12404;
  assign n12406 = n12339 & n12405;
  assign n12407 = n12290 & n12406;
  assign n12408 = n12227 & n12407;
  assign n12409 = pi3310 & po3871;
  assign n12410 = n12408 & ~n12409;
  assign n12411 = ~pi1787 & ~n12410;
  assign n12412 = pi1787 & pi2828;
  assign n12413 = ~n12411 & ~n12412;
  assign n12414 = n9472 & ~n12413;
  assign n12415 = ~n12187 & ~n12414;
  assign n12416 = ~n10914 & ~n12415;
  assign n12417 = ~n10902 & n12416;
  assign n12418 = ~n12167 & ~n12417;
  assign n12419 = n10885 & ~n12418;
  assign n12420 = ~n10047 & ~n10329;
  assign n12421 = ~n10046 & ~n12420;
  assign n12422 = n10034 & n12421;
  assign n12423 = ~n10034 & ~n12421;
  assign n12424 = ~n12422 & ~n12423;
  assign n12425 = n10296 & ~n12424;
  assign n12426 = ~n10284 & ~n10285;
  assign n12427 = ~n10073 & ~n12426;
  assign n12428 = n10037 & ~n10052;
  assign n12429 = ~n10037 & n10052;
  assign n12430 = ~n12428 & ~n12429;
  assign n12431 = n12427 & ~n12430;
  assign n12432 = ~n12427 & n12430;
  assign n12433 = ~n12431 & ~n12432;
  assign n12434 = ~n10296 & ~n12433;
  assign n12435 = ~n12425 & ~n12434;
  assign n12436 = ~pi0568 & ~n12435;
  assign n12437 = n10362 & ~n12433;
  assign n12438 = ~n10362 & ~n12424;
  assign n12439 = ~n12437 & ~n12438;
  assign n12440 = pi0568 & ~n12439;
  assign n12441 = ~n12436 & ~n12440;
  assign n12442 = pi0660 & n10020;
  assign n12443 = pi0660 & n10019;
  assign n12444 = ~n12442 & ~n12443;
  assign n12445 = n12441 & n12444;
  assign n12446 = ~n11186 & ~n12445;
  assign n12447 = pi1028 & ~n11706;
  assign n12448 = pi0902 & n11709;
  assign n12449 = n11701 & ~n12165;
  assign n12450 = ~n12448 & ~n12449;
  assign n12451 = ~n12447 & n12450;
  assign n12452 = n10886 & ~n12148;
  assign n12453 = pi2448 & po3871;
  assign n12454 = pi0424 & n11714;
  assign n12455 = ~n12453 & ~n12454;
  assign n12456 = ~n12452 & n12455;
  assign n12457 = n12451 & n12456;
  assign n12458 = ~n11700 & ~n12457;
  assign n12459 = pi0845 & n11700;
  assign n12460 = ~n12458 & ~n12459;
  assign n12461 = ~n10914 & ~n12460;
  assign n12462 = ~n12446 & ~n12461;
  assign n12463 = ~n10902 & ~n12462;
  assign n12464 = ~n11573 & n11643;
  assign n12465 = n11573 & ~n11643;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = n11615 & ~n12466;
  assign n12468 = ~n11576 & n11578;
  assign n12469 = n11576 & ~n11578;
  assign n12470 = ~n12468 & ~n12469;
  assign n12471 = n11524 & ~n12470;
  assign n12472 = ~n11524 & n12470;
  assign n12473 = ~n12471 & ~n12472;
  assign n12474 = ~n11615 & ~n12473;
  assign n12475 = ~n12467 & ~n12474;
  assign n12476 = ~pi0518 & ~n12475;
  assign n12477 = n11665 & ~n12473;
  assign n12478 = ~n11665 & ~n12466;
  assign n12479 = ~n12477 & ~n12478;
  assign n12480 = pi0518 & ~n12479;
  assign n12481 = ~n12476 & ~n12480;
  assign n12482 = pi0704 & n11566;
  assign n12483 = pi0704 & n11568;
  assign n12484 = ~n12482 & ~n12483;
  assign n12485 = n12481 & n12484;
  assign n12486 = ~n11186 & n12485;
  assign n12487 = pi2966 & n11190;
  assign n12488 = pi2963 & n11197;
  assign n12489 = ~n12487 & ~n12488;
  assign n12490 = pi2455 & n11195;
  assign n12491 = pi2464 & n11192;
  assign n12492 = ~n12490 & ~n12491;
  assign n12493 = n12489 & n12492;
  assign n12494 = n9424 & ~n12493;
  assign n12495 = pi2963 & n11207;
  assign n12496 = pi2464 & n11202;
  assign n12497 = ~n12495 & ~n12496;
  assign n12498 = pi2966 & n11204;
  assign n12499 = pi2455 & n11209;
  assign n12500 = ~n12498 & ~n12499;
  assign n12501 = n12497 & n12500;
  assign n12502 = ~n9424 & ~n12501;
  assign n12503 = ~n12494 & ~n12502;
  assign n12504 = n11186 & n12503;
  assign n12505 = ~n12486 & ~n12504;
  assign n12506 = n10902 & n12505;
  assign n12507 = ~n12463 & ~n12506;
  assign n12508 = ~n10885 & ~n12507;
  assign n12509 = pi1787 & pi3149;
  assign n12510 = ~pi0979 & pi2841;
  assign n12511 = pi0979 & pi2124;
  assign n12512 = ~n12510 & ~n12511;
  assign n12513 = pi0717 & ~n12512;
  assign n12514 = pi0198 & ~pi0979;
  assign n12515 = pi0197 & pi0979;
  assign n12516 = ~n12514 & ~n12515;
  assign n12517 = pi0716 & ~n12516;
  assign n12518 = pi0252 & ~pi0979;
  assign n12519 = pi0249 & pi0979;
  assign n12520 = ~n12518 & ~n12519;
  assign n12521 = pi0761 & ~n12520;
  assign n12522 = ~n12517 & ~n12521;
  assign n12523 = ~n9535 & n12522;
  assign n12524 = ~n9531 & n12523;
  assign n12525 = ~n12513 & n12524;
  assign n12526 = n9523 & ~n12525;
  assign n12527 = pi0979 & pi2177;
  assign n12528 = ~pi0979 & pi2939;
  assign n12529 = ~n12527 & ~n12528;
  assign n12530 = pi0837 & ~n12529;
  assign n12531 = ~pi0979 & pi2931;
  assign n12532 = pi0979 & pi2161;
  assign n12533 = ~n12531 & ~n12532;
  assign n12534 = pi0836 & ~n12533;
  assign n12535 = ~n12530 & ~n12534;
  assign n12536 = pi0979 & pi2144;
  assign n12537 = ~pi0979 & pi2916;
  assign n12538 = ~n12536 & ~n12537;
  assign n12539 = pi0767 & ~n12538;
  assign n12540 = ~pi0979 & pi2420;
  assign n12541 = pi0979 & pi1955;
  assign n12542 = ~n12540 & ~n12541;
  assign n12543 = pi0768 & ~n12542;
  assign n12544 = ~n12539 & ~n12543;
  assign n12545 = pi0167 & ~pi0979;
  assign n12546 = pi0153 & pi0979;
  assign n12547 = ~n12545 & ~n12546;
  assign n12548 = pi0838 & ~n12547;
  assign n12549 = n12544 & ~n12548;
  assign n12550 = n12535 & n12549;
  assign n12551 = n9549 & ~n12550;
  assign n12552 = ~n12526 & ~n12551;
  assign n12553 = pi1333 & pi1742;
  assign n12554 = pi1335 & pi2583;
  assign n12555 = ~n12553 & ~n12554;
  assign n12556 = pi1332 & pi2768;
  assign n12557 = pi0237 & pi1336;
  assign n12558 = ~n12556 & ~n12557;
  assign n12559 = n12555 & n12558;
  assign n12560 = n9726 & ~n12559;
  assign n12561 = pi1846 & n10564;
  assign n12562 = pi0738 & n9715;
  assign n12563 = pi1952 & n9718;
  assign n12564 = ~n12562 & ~n12563;
  assign n12565 = ~n12561 & n12564;
  assign n12566 = pi1727 & n11106;
  assign n12567 = pi0869 & n9707;
  assign n12568 = ~n12566 & ~n12567;
  assign n12569 = pi0977 & n9687;
  assign n12570 = pi1436 & n9691;
  assign n12571 = ~n12569 & ~n12570;
  assign n12572 = pi0792 & n9614;
  assign n12573 = pi2057 & n9618;
  assign n12574 = ~n12572 & ~n12573;
  assign n12575 = pi1849 & n10557;
  assign n12576 = n12574 & ~n12575;
  assign n12577 = n12571 & n12576;
  assign n12578 = pi1828 & n9698;
  assign n12579 = n12577 & ~n12578;
  assign n12580 = ~n11102 & n12579;
  assign n12581 = n12568 & n12580;
  assign n12582 = n12565 & n12581;
  assign n12583 = pi1772 & n9712;
  assign n12584 = n12582 & ~n12583;
  assign n12585 = pi1450 & n11145;
  assign n12586 = pi0902 & n9710;
  assign n12587 = ~n12585 & ~n12586;
  assign n12588 = pi0723 & n9654;
  assign n12589 = pi2493 & n11158;
  assign n12590 = ~n12588 & ~n12589;
  assign n12591 = pi0845 & n9670;
  assign n12592 = pi1066 & n9676;
  assign n12593 = ~n12591 & ~n12592;
  assign n12594 = pi3107 & n9647;
  assign n12595 = n12593 & ~n12594;
  assign n12596 = n12590 & n12595;
  assign n12597 = pi1918 & n9622;
  assign n12598 = n12596 & ~n12597;
  assign n12599 = pi1877 & n9679;
  assign n12600 = pi0398 & n9682;
  assign n12601 = ~n12599 & ~n12600;
  assign n12602 = n12598 & n12601;
  assign n12603 = n12587 & n12602;
  assign n12604 = n12584 & n12603;
  assign n12605 = pi1934 & ~n12604;
  assign n12606 = ~n12560 & ~n12605;
  assign n12607 = pi0137 & ~pi0979;
  assign n12608 = pi0135 & pi0979;
  assign n12609 = ~n12607 & ~n12608;
  assign n12610 = pi0720 & ~n12609;
  assign n12611 = pi0268 & ~pi0979;
  assign n12612 = pi0267 & pi0979;
  assign n12613 = ~n12611 & ~n12612;
  assign n12614 = pi0721 & ~n12613;
  assign n12615 = ~n12610 & ~n12614;
  assign n12616 = ~pi0979 & pi2630;
  assign n12617 = pi0979 & pi3167;
  assign n12618 = ~n12616 & ~n12617;
  assign n12619 = pi0765 & ~n12618;
  assign n12620 = ~pi0979 & pi2888;
  assign n12621 = pi0979 & pi3126;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = pi0766 & ~n12622;
  assign n12624 = ~n12619 & ~n12623;
  assign n12625 = ~pi0979 & pi2611;
  assign n12626 = pi0979 & pi2605;
  assign n12627 = ~n12625 & ~n12626;
  assign n12628 = pi0763 & ~n12627;
  assign n12629 = ~pi0979 & pi2624;
  assign n12630 = pi0979 & pi2618;
  assign n12631 = ~n12629 & ~n12630;
  assign n12632 = pi0764 & ~n12631;
  assign n12633 = ~n12628 & ~n12632;
  assign n12634 = n12624 & n12633;
  assign n12635 = ~n9499 & n12634;
  assign n12636 = n12615 & n12635;
  assign n12637 = n9486 & ~n12636;
  assign n12638 = n12606 & ~n12637;
  assign n12639 = n12552 & n12638;
  assign n12640 = pi1331 & ~n9105;
  assign n12641 = pi0590 & pi1359;
  assign n12642 = ~n12640 & ~n12641;
  assign n12643 = pi0912 & pi1358;
  assign n12644 = pi0382 & pi1057;
  assign n12645 = ~n12643 & ~n12644;
  assign n12646 = pi3514 & ~n10410;
  assign n12647 = n12645 & ~n12646;
  assign n12648 = n12642 & n12647;
  assign n12649 = n9475 & ~n12648;
  assign n12650 = n12639 & ~n12649;
  assign n12651 = pi1340 & pi2279;
  assign n12652 = pi1341 & pi2292;
  assign n12653 = ~n12651 & ~n12652;
  assign n12654 = pi1342 & pi2303;
  assign n12655 = n12653 & ~n12654;
  assign n12656 = pi1055 & pi2719;
  assign n12657 = n12655 & ~n12656;
  assign n12658 = pi1343 & pi2314;
  assign n12659 = pi1054 & pi2708;
  assign n12660 = ~n12658 & ~n12659;
  assign n12661 = pi1349 & pi2728;
  assign n12662 = pi1056 & pi2738;
  assign n12663 = ~n12661 & ~n12662;
  assign n12664 = pi1354 & pi2960;
  assign n12665 = n12663 & ~n12664;
  assign n12666 = pi1357 & pi2413;
  assign n12667 = n12665 & ~n12666;
  assign n12668 = pi1355 & pi2452;
  assign n12669 = pi1356 & pi2965;
  assign n12670 = ~n12668 & ~n12669;
  assign n12671 = n12667 & n12670;
  assign n12672 = n12660 & n12671;
  assign n12673 = n12657 & n12672;
  assign n12674 = n9736 & ~n12673;
  assign n12675 = pi1347 & pi2675;
  assign n12676 = pi1348 & pi2602;
  assign n12677 = ~n12675 & ~n12676;
  assign n12678 = pi1350 & pi2257;
  assign n12679 = n12677 & ~n12678;
  assign n12680 = pi1353 & pi1976;
  assign n12681 = n12679 & ~n12680;
  assign n12682 = pi1351 & pi2261;
  assign n12683 = pi1352 & pi2271;
  assign n12684 = ~n12682 & ~n12683;
  assign n12685 = pi1339 & pi2243;
  assign n12686 = pi1345 & pi2550;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = pi1346 & pi2661;
  assign n12689 = n12687 & ~n12688;
  assign n12690 = pi1338 & pi2229;
  assign n12691 = n12689 & ~n12690;
  assign n12692 = pi1600 & pi2201;
  assign n12693 = pi1337 & pi2215;
  assign n12694 = ~n12692 & ~n12693;
  assign n12695 = n12691 & n12694;
  assign n12696 = n12684 & n12695;
  assign n12697 = n12681 & n12696;
  assign n12698 = n9577 & ~n12697;
  assign n12699 = ~n12674 & ~n12698;
  assign n12700 = n12650 & n12699;
  assign n12701 = pi3306 & po3871;
  assign n12702 = n12700 & ~n12701;
  assign n12703 = ~pi1787 & ~n12702;
  assign n12704 = ~n12509 & ~n12703;
  assign n12705 = n9472 & ~n12704;
  assign n12706 = pi3868 & n9804;
  assign n12707 = pi3884 & n9774;
  assign n12708 = ~n12706 & ~n12707;
  assign n12709 = pi3852 & n9802;
  assign n12710 = pi3900 & n9771;
  assign n12711 = pi3964 & n9793;
  assign n12712 = ~n12710 & ~n12711;
  assign n12713 = pi3948 & n9791;
  assign n12714 = pi3932 & n9788;
  assign n12715 = ~n12713 & ~n12714;
  assign n12716 = n12712 & n12715;
  assign n12717 = ~n12709 & n12716;
  assign n12718 = n12708 & n12717;
  assign n12719 = pi3868 & n9799;
  assign n12720 = n12718 & ~n12719;
  assign n12721 = pi3916 & n9781;
  assign n12722 = pi3980 & n9783;
  assign n12723 = ~n12721 & ~n12722;
  assign n12724 = n12720 & n12723;
  assign n12725 = ~n9472 & ~n12724;
  assign n12726 = ~n12705 & ~n12725;
  assign n12727 = n10914 & ~n12726;
  assign n12728 = ~n11401 & ~n11648;
  assign n12729 = ~n11403 & ~n12728;
  assign n12730 = n11386 & n12729;
  assign n12731 = ~n11386 & ~n12729;
  assign n12732 = ~n12730 & ~n12731;
  assign n12733 = n11615 & ~n12732;
  assign n12734 = ~n11405 & ~n11408;
  assign n12735 = ~n11604 & ~n11605;
  assign n12736 = ~n11427 & ~n12735;
  assign n12737 = ~n12734 & ~n12736;
  assign n12738 = n12734 & n12736;
  assign n12739 = ~n12737 & ~n12738;
  assign n12740 = ~n11615 & ~n12739;
  assign n12741 = ~n12733 & ~n12740;
  assign n12742 = ~pi0518 & ~n12741;
  assign n12743 = n11665 & ~n12739;
  assign n12744 = ~n11665 & ~n12732;
  assign n12745 = ~n12743 & ~n12744;
  assign n12746 = pi0518 & ~n12745;
  assign n12747 = ~n12742 & ~n12746;
  assign n12748 = pi0701 & n11373;
  assign n12749 = pi0701 & n11374;
  assign n12750 = ~n12748 & ~n12749;
  assign n12751 = n12747 & n12750;
  assign n12752 = ~n10914 & ~n12751;
  assign n12753 = ~n12727 & ~n12752;
  assign n12754 = n11755 & ~n12753;
  assign n12755 = ~n12508 & ~n12754;
  assign po0225 = n12419 | ~n12755;
  assign n12757 = n10302 & ~n10326;
  assign n12758 = ~n10238 & ~n12757;
  assign n12759 = ~n10237 & ~n12758;
  assign n12760 = n10233 & n12759;
  assign n12761 = ~n10233 & ~n12759;
  assign n12762 = ~n12760 & ~n12761;
  assign n12763 = n10296 & ~n12762;
  assign n12764 = ~n10203 & n10270;
  assign n12765 = n10277 & ~n12764;
  assign n12766 = ~n10232 & ~n12765;
  assign n12767 = ~n10281 & ~n12766;
  assign n12768 = n10236 & ~n10240;
  assign n12769 = ~n10236 & n10240;
  assign n12770 = ~n12768 & ~n12769;
  assign n12771 = ~n12767 & n12770;
  assign n12772 = n12767 & ~n12770;
  assign n12773 = ~n12771 & ~n12772;
  assign n12774 = ~n10296 & ~n12773;
  assign n12775 = ~n12763 & ~n12774;
  assign n12776 = ~pi0568 & ~n12775;
  assign n12777 = n10362 & ~n12773;
  assign n12778 = ~n10362 & ~n12762;
  assign n12779 = ~n12777 & ~n12778;
  assign n12780 = pi0568 & ~n12779;
  assign n12781 = ~n12776 & ~n12780;
  assign n12782 = pi0755 & n10063;
  assign n12783 = pi0755 & n10062;
  assign n12784 = ~n12782 & ~n12783;
  assign n12785 = n12781 & n12784;
  assign n12786 = n10914 & ~n12785;
  assign n12787 = pi2699 & n9837;
  assign n12788 = pi2702 & n9834;
  assign n12789 = ~n12787 & ~n12788;
  assign n12790 = pi2439 & n9839;
  assign n12791 = pi2276 & n9832;
  assign n12792 = ~n12790 & ~n12791;
  assign n12793 = n12789 & n12792;
  assign n12794 = ~n9424 & ~n12793;
  assign n12795 = pi2439 & n10376;
  assign n12796 = pi2702 & n10381;
  assign n12797 = ~n12795 & ~n12796;
  assign n12798 = pi2699 & n10374;
  assign n12799 = pi2276 & n10379;
  assign n12800 = ~n12798 & ~n12799;
  assign n12801 = n12797 & n12800;
  assign n12802 = n9424 & ~n12801;
  assign n12803 = ~n12794 & ~n12802;
  assign n12804 = n11701 & ~n12803;
  assign n12805 = pi2449 & po3871;
  assign n12806 = pi0876 & n11709;
  assign n12807 = pi1030 & ~n11706;
  assign n12808 = pi0425 & n11714;
  assign n12809 = ~n12807 & ~n12808;
  assign n12810 = ~n12806 & n12809;
  assign n12811 = ~n12805 & n12810;
  assign n12812 = ~n11700 & n12811;
  assign n12813 = pi2461 & n11192;
  assign n12814 = pi2961 & n11197;
  assign n12815 = ~n12813 & ~n12814;
  assign n12816 = pi2453 & n11195;
  assign n12817 = pi3096 & n11190;
  assign n12818 = ~n12816 & ~n12817;
  assign n12819 = n12815 & n12818;
  assign n12820 = n9424 & ~n12819;
  assign n12821 = pi2961 & n11207;
  assign n12822 = pi2461 & n11202;
  assign n12823 = ~n12821 & ~n12822;
  assign n12824 = pi3096 & n11204;
  assign n12825 = pi2453 & n11209;
  assign n12826 = ~n12824 & ~n12825;
  assign n12827 = n12823 & n12826;
  assign n12828 = ~n9424 & ~n12827;
  assign n12829 = ~n12820 & ~n12828;
  assign n12830 = n10886 & ~n12829;
  assign n12831 = n12812 & ~n12830;
  assign n12832 = ~n12804 & n12831;
  assign n12833 = ~pi0861 & n11700;
  assign n12834 = ~n12832 & ~n12833;
  assign n12835 = n11186 & n12834;
  assign n12836 = ~n12786 & ~n12835;
  assign n12837 = ~n10902 & ~n12836;
  assign n12838 = pi0703 & ~n11530;
  assign n12839 = n11260 & n12838;
  assign n12840 = pi0703 & n11533;
  assign n12841 = ~n11643 & n11644;
  assign n12842 = n11626 & ~n12841;
  assign n12843 = ~n11544 & ~n12842;
  assign n12844 = n11544 & n12842;
  assign n12845 = ~n12843 & ~n12844;
  assign n12846 = n11615 & ~n12845;
  assign n12847 = ~n11560 & ~n11601;
  assign n12848 = ~n11524 & n11589;
  assign n12849 = n11597 & ~n12848;
  assign n12850 = ~n12847 & ~n12849;
  assign n12851 = n12847 & n12849;
  assign n12852 = ~n12850 & ~n12851;
  assign n12853 = ~n11615 & ~n12852;
  assign n12854 = ~n12846 & ~n12853;
  assign n12855 = ~pi0518 & ~n12854;
  assign n12856 = n11665 & ~n12852;
  assign n12857 = ~n11665 & ~n12845;
  assign n12858 = ~n12856 & ~n12857;
  assign n12859 = pi0518 & ~n12858;
  assign n12860 = ~n12855 & ~n12859;
  assign n12861 = ~n12840 & n12860;
  assign n12862 = ~n12839 & n12861;
  assign n12863 = n10914 & n12862;
  assign n12864 = pi2462 & n11192;
  assign n12865 = pi2962 & n11197;
  assign n12866 = ~n12864 & ~n12865;
  assign n12867 = pi2454 & n11195;
  assign n12868 = pi3093 & n11190;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = n12866 & n12869;
  assign n12871 = n9424 & ~n12870;
  assign n12872 = pi2462 & n11202;
  assign n12873 = pi3093 & n11204;
  assign n12874 = ~n12872 & ~n12873;
  assign n12875 = pi2962 & n11207;
  assign n12876 = pi2454 & n11209;
  assign n12877 = ~n12875 & ~n12876;
  assign n12878 = n12874 & n12877;
  assign n12879 = ~n9424 & ~n12878;
  assign n12880 = ~n12871 & ~n12879;
  assign n12881 = ~n10914 & n12880;
  assign n12882 = ~n12863 & ~n12881;
  assign n12883 = n10902 & n12882;
  assign n12884 = ~n12837 & ~n12883;
  assign n12885 = ~n10885 & ~n12884;
  assign n12886 = pi3866 & n9804;
  assign n12887 = pi3882 & n9774;
  assign n12888 = ~n12886 & ~n12887;
  assign n12889 = pi3850 & n9802;
  assign n12890 = pi3914 & n9781;
  assign n12891 = pi3898 & n9771;
  assign n12892 = ~n12890 & ~n12891;
  assign n12893 = pi3946 & n9791;
  assign n12894 = pi3930 & n9788;
  assign n12895 = ~n12893 & ~n12894;
  assign n12896 = n12892 & n12895;
  assign n12897 = ~n12889 & n12896;
  assign n12898 = n12888 & n12897;
  assign n12899 = pi3866 & n9799;
  assign n12900 = n12898 & ~n12899;
  assign n12901 = pi3978 & n9783;
  assign n12902 = pi3962 & n9793;
  assign n12903 = ~n12901 & ~n12902;
  assign n12904 = n12900 & n12903;
  assign n12905 = ~n9472 & ~n12904;
  assign n12906 = pi1331 & ~n8913;
  assign n12907 = pi0571 & pi1359;
  assign n12908 = ~n12906 & ~n12907;
  assign n12909 = pi3516 & ~n10410;
  assign n12910 = pi1334 & pi3285;
  assign n12911 = pi0914 & pi1358;
  assign n12912 = ~n12910 & ~n12911;
  assign n12913 = pi1053 & pi2409;
  assign n12914 = pi0384 & pi1057;
  assign n12915 = ~n12913 & ~n12914;
  assign n12916 = n12912 & n12915;
  assign n12917 = ~n12909 & n12916;
  assign n12918 = n12908 & n12917;
  assign n12919 = n9475 & ~n12918;
  assign n12920 = ~pi0979 & pi2862;
  assign n12921 = pi0979 & pi3151;
  assign n12922 = ~n12920 & ~n12921;
  assign n12923 = pi0763 & ~n12922;
  assign n12924 = ~pi0979 & pi2870;
  assign n12925 = pi0979 & pi3160;
  assign n12926 = ~n12924 & ~n12925;
  assign n12927 = pi0764 & ~n12926;
  assign n12928 = ~n12923 & ~n12927;
  assign n12929 = ~pi0979 & pi2632;
  assign n12930 = pi0979 & pi3169;
  assign n12931 = ~n12929 & ~n12930;
  assign n12932 = pi0765 & ~n12931;
  assign n12933 = ~pi0979 & pi3075;
  assign n12934 = pi0979 & pi3125;
  assign n12935 = ~n12933 & ~n12934;
  assign n12936 = pi0766 & ~n12935;
  assign n12937 = ~n12932 & ~n12936;
  assign n12938 = pi0138 & ~pi0979;
  assign n12939 = pi0136 & pi0979;
  assign n12940 = ~n12938 & ~n12939;
  assign n12941 = pi0720 & ~n12940;
  assign n12942 = pi0313 & ~pi0979;
  assign n12943 = pi0312 & pi0979;
  assign n12944 = ~n12942 & ~n12943;
  assign n12945 = pi0721 & ~n12944;
  assign n12946 = ~n12941 & ~n12945;
  assign n12947 = n12937 & n12946;
  assign n12948 = ~n9499 & n12947;
  assign n12949 = n12928 & n12948;
  assign n12950 = n9486 & ~n12949;
  assign n12951 = ~n12919 & ~n12950;
  assign n12952 = ~pi0979 & pi2843;
  assign n12953 = pi0979 & pi2126;
  assign n12954 = ~n12952 & ~n12953;
  assign n12955 = pi0717 & ~n12954;
  assign n12956 = pi0280 & ~pi0979;
  assign n12957 = pi0279 & pi0979;
  assign n12958 = ~n12956 & ~n12957;
  assign n12959 = pi0716 & ~n12958;
  assign n12960 = pi0253 & ~pi0979;
  assign n12961 = pi0250 & pi0979;
  assign n12962 = ~n12960 & ~n12961;
  assign n12963 = pi0761 & ~n12962;
  assign n12964 = ~n12959 & ~n12963;
  assign n12965 = ~n9535 & n12964;
  assign n12966 = ~n9531 & n12965;
  assign n12967 = ~n12955 & n12966;
  assign n12968 = n9523 & ~n12967;
  assign n12969 = pi0979 & pi2163;
  assign n12970 = ~pi0979 & pi2932;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = pi0836 & ~n12971;
  assign n12973 = ~pi0979 & pi2784;
  assign n12974 = pi0979 & pi2179;
  assign n12975 = ~n12973 & ~n12974;
  assign n12976 = pi0837 & ~n12975;
  assign n12977 = ~n12972 & ~n12976;
  assign n12978 = pi0979 & pi2146;
  assign n12979 = ~pi0979 & pi2918;
  assign n12980 = ~n12978 & ~n12979;
  assign n12981 = pi0767 & ~n12980;
  assign n12982 = ~pi0979 & pi2422;
  assign n12983 = pi0979 & pi1957;
  assign n12984 = ~n12982 & ~n12983;
  assign n12985 = pi0768 & ~n12984;
  assign n12986 = ~n12981 & ~n12985;
  assign n12987 = pi0169 & ~pi0979;
  assign n12988 = pi0155 & pi0979;
  assign n12989 = ~n12987 & ~n12988;
  assign n12990 = pi0838 & ~n12989;
  assign n12991 = pi0586 & pi1360;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = n12986 & n12992;
  assign n12994 = n12977 & n12993;
  assign n12995 = n9549 & ~n12994;
  assign n12996 = ~n12968 & ~n12995;
  assign n12997 = pi1343 & pi2316;
  assign n12998 = pi1054 & pi2710;
  assign n12999 = ~n12997 & ~n12998;
  assign n13000 = pi1055 & pi2531;
  assign n13001 = n12999 & ~n13000;
  assign n13002 = pi1342 & pi2304;
  assign n13003 = n13001 & ~n13002;
  assign n13004 = pi1340 & pi2281;
  assign n13005 = pi1341 & pi2293;
  assign n13006 = ~n13004 & ~n13005;
  assign n13007 = pi1349 & pi2729;
  assign n13008 = pi1056 & pi2548;
  assign n13009 = ~n13007 & ~n13008;
  assign n13010 = pi1354 & pi2961;
  assign n13011 = n13009 & ~n13010;
  assign n13012 = pi1357 & pi2461;
  assign n13013 = n13011 & ~n13012;
  assign n13014 = pi1355 & pi2453;
  assign n13015 = pi1356 & pi3096;
  assign n13016 = ~n13014 & ~n13015;
  assign n13017 = n13013 & n13016;
  assign n13018 = n13006 & n13017;
  assign n13019 = n13003 & n13018;
  assign n13020 = n9736 & ~n13019;
  assign n13021 = pi1351 & pi2439;
  assign n13022 = pi1352 & pi2702;
  assign n13023 = ~n13021 & ~n13022;
  assign n13024 = pi1353 & pi2276;
  assign n13025 = n13023 & ~n13024;
  assign n13026 = pi1350 & pi2699;
  assign n13027 = n13025 & ~n13026;
  assign n13028 = pi1347 & pi2677;
  assign n13029 = pi1348 & pi2688;
  assign n13030 = ~n13028 & ~n13029;
  assign n13031 = pi1600 & pi2203;
  assign n13032 = pi1337 & pi2217;
  assign n13033 = ~n13031 & ~n13032;
  assign n13034 = pi1338 & pi2231;
  assign n13035 = n13033 & ~n13034;
  assign n13036 = pi1346 & pi2663;
  assign n13037 = n13035 & ~n13036;
  assign n13038 = pi1339 & pi2245;
  assign n13039 = pi1345 & pi2649;
  assign n13040 = ~n13038 & ~n13039;
  assign n13041 = n13037 & n13040;
  assign n13042 = n13030 & n13041;
  assign n13043 = n13027 & n13042;
  assign n13044 = n9577 & ~n13043;
  assign n13045 = ~n13020 & ~n13044;
  assign n13046 = pi0247 & pi1336;
  assign n13047 = pi1333 & pi1867;
  assign n13048 = ~n13046 & ~n13047;
  assign n13049 = pi1332 & pi2569;
  assign n13050 = pi1335 & pi2585;
  assign n13051 = ~n13049 & ~n13050;
  assign n13052 = n13048 & n13051;
  assign n13053 = n9726 & ~n13052;
  assign n13054 = pi0956 & n9614;
  assign n13055 = pi2055 & n9618;
  assign n13056 = ~n13054 & ~n13055;
  assign n13057 = pi0800 & n9687;
  assign n13058 = pi1438 & n9691;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = pi0963 & n9607;
  assign n13061 = n13059 & ~n13060;
  assign n13062 = n13056 & n13061;
  assign n13063 = pi1830 & n9698;
  assign n13064 = n13062 & ~n13063;
  assign n13065 = pi0880 & n9715;
  assign n13066 = pi1884 & n9718;
  assign n13067 = ~n13065 & ~n13066;
  assign n13068 = pi0948 & n9702;
  assign n13069 = n13067 & ~n13068;
  assign n13070 = pi1729 & n11106;
  assign n13071 = pi0742 & n9707;
  assign n13072 = ~n13070 & ~n13071;
  assign n13073 = n13069 & n13072;
  assign n13074 = pi0769 & n9654;
  assign n13075 = pi2495 & n11158;
  assign n13076 = ~n13074 & ~n13075;
  assign n13077 = pi0861 & n9670;
  assign n13078 = pi1602 & n9676;
  assign n13079 = ~n13077 & ~n13078;
  assign n13080 = pi2503 & n9647;
  assign n13081 = n13079 & ~n13080;
  assign n13082 = n13076 & n13081;
  assign n13083 = pi1938 & n11165;
  assign n13084 = n13082 & ~n13083;
  assign n13085 = pi2103 & n9628;
  assign n13086 = pi1020 & n9631;
  assign n13087 = ~n13085 & ~n13086;
  assign n13088 = pi1857 & n9657;
  assign n13089 = pi1751 & n9659;
  assign n13090 = ~n13088 & ~n13089;
  assign n13091 = n13087 & n13090;
  assign n13092 = pi1427 & n11133;
  assign n13093 = pi0496 & n9682;
  assign n13094 = ~n13092 & ~n13093;
  assign n13095 = pi1706 & n9679;
  assign n13096 = n13094 & ~n13095;
  assign n13097 = pi1921 & n9622;
  assign n13098 = n13096 & ~n13097;
  assign n13099 = n13091 & n13098;
  assign n13100 = ~n11102 & n13099;
  assign n13101 = n13084 & n13100;
  assign n13102 = pi1774 & n9712;
  assign n13103 = n13101 & ~n13102;
  assign n13104 = pi1452 & n11145;
  assign n13105 = pi0876 & n9710;
  assign n13106 = ~n13104 & ~n13105;
  assign n13107 = n13103 & n13106;
  assign n13108 = n13073 & n13107;
  assign n13109 = n13064 & n13108;
  assign n13110 = pi1934 & ~n13109;
  assign n13111 = ~n13053 & ~n13110;
  assign n13112 = n13045 & n13111;
  assign n13113 = n12996 & n13112;
  assign n13114 = n12951 & n13113;
  assign n13115 = pi3308 & po3871;
  assign n13116 = n13114 & ~n13115;
  assign n13117 = ~pi1787 & ~n13116;
  assign n13118 = pi1787 & pi2826;
  assign n13119 = ~n13117 & ~n13118;
  assign n13120 = n9472 & ~n13119;
  assign n13121 = ~n12905 & ~n13120;
  assign n13122 = n10914 & n13121;
  assign n13123 = ~n11537 & ~n12842;
  assign n13124 = ~n11536 & ~n13123;
  assign n13125 = n11525 & n13124;
  assign n13126 = ~n11525 & ~n13124;
  assign n13127 = ~n13125 & ~n13126;
  assign n13128 = n11615 & ~n13127;
  assign n13129 = n11528 & ~n11542;
  assign n13130 = ~n11528 & n11542;
  assign n13131 = ~n13129 & ~n13130;
  assign n13132 = ~n11560 & ~n12849;
  assign n13133 = ~n11601 & ~n13132;
  assign n13134 = ~n13131 & n13133;
  assign n13135 = n13131 & ~n13133;
  assign n13136 = ~n13134 & ~n13135;
  assign n13137 = ~n11615 & ~n13136;
  assign n13138 = ~n13128 & ~n13137;
  assign n13139 = ~pi0518 & ~n13138;
  assign n13140 = n11665 & ~n13136;
  assign n13141 = ~n11665 & ~n13127;
  assign n13142 = ~n13140 & ~n13141;
  assign n13143 = pi0518 & ~n13142;
  assign n13144 = ~n13139 & ~n13143;
  assign n13145 = pi0702 & n11416;
  assign n13146 = pi0702 & ~n11260;
  assign n13147 = n11234 & n13146;
  assign n13148 = ~n13145 & ~n13147;
  assign n13149 = n13144 & n13148;
  assign n13150 = ~n10914 & n13149;
  assign n13151 = ~n13122 & ~n13150;
  assign n13152 = n11755 & n13151;
  assign n13153 = pi0979 & pi2164;
  assign n13154 = ~pi0979 & pi2808;
  assign n13155 = ~n13153 & ~n13154;
  assign n13156 = pi0836 & ~n13155;
  assign n13157 = ~pi0979 & pi2941;
  assign n13158 = pi0979 & pi2180;
  assign n13159 = ~n13157 & ~n13158;
  assign n13160 = pi0837 & ~n13159;
  assign n13161 = ~n13156 & ~n13160;
  assign n13162 = pi0979 & pi2147;
  assign n13163 = ~pi0979 & pi2919;
  assign n13164 = ~n13162 & ~n13163;
  assign n13165 = pi0767 & ~n13164;
  assign n13166 = ~pi0979 & pi2423;
  assign n13167 = pi0979 & pi1958;
  assign n13168 = ~n13166 & ~n13167;
  assign n13169 = pi0768 & ~n13168;
  assign n13170 = ~n13165 & ~n13169;
  assign n13171 = pi0170 & ~pi0979;
  assign n13172 = pi0156 & pi0979;
  assign n13173 = ~n13171 & ~n13172;
  assign n13174 = pi0838 & ~n13173;
  assign n13175 = pi1360 & ~pi3633;
  assign n13176 = ~n13174 & ~n13175;
  assign n13177 = n13170 & n13176;
  assign n13178 = n13161 & n13177;
  assign n13179 = n9549 & ~n13178;
  assign n13180 = pi0054 & ~pi0979;
  assign n13181 = pi0052 & pi0979;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = pi0719 & ~n13182;
  assign n13184 = ~pi0979 & pi2633;
  assign n13185 = pi0979 & pi3133;
  assign n13186 = ~n13184 & ~n13185;
  assign n13187 = pi0765 & ~n13186;
  assign n13188 = ~pi0979 & pi2890;
  assign n13189 = pi0979 & pi3178;
  assign n13190 = ~n13188 & ~n13189;
  assign n13191 = pi0766 & ~n13190;
  assign n13192 = ~n13187 & ~n13191;
  assign n13193 = ~pi0979 & pi2863;
  assign n13194 = pi0979 & pi3152;
  assign n13195 = ~n13193 & ~n13194;
  assign n13196 = pi0763 & ~n13195;
  assign n13197 = ~pi0979 & pi2871;
  assign n13198 = pi0979 & pi3161;
  assign n13199 = ~n13197 & ~n13198;
  assign n13200 = pi0764 & ~n13199;
  assign n13201 = ~n13196 & ~n13200;
  assign n13202 = pi0131 & ~pi0979;
  assign n13203 = pi0130 & pi0979;
  assign n13204 = ~n13202 & ~n13203;
  assign n13205 = pi0720 & ~n13204;
  assign n13206 = pi0328 & ~pi0979;
  assign n13207 = pi0327 & pi0979;
  assign n13208 = ~n13206 & ~n13207;
  assign n13209 = pi0721 & ~n13208;
  assign n13210 = ~n13205 & ~n13209;
  assign n13211 = n13201 & n13210;
  assign n13212 = n13192 & n13211;
  assign n13213 = ~n13183 & n13212;
  assign n13214 = n9486 & ~n13213;
  assign n13215 = ~n13179 & ~n13214;
  assign n13216 = pi0248 & pi1336;
  assign n13217 = pi0368 & pi1333;
  assign n13218 = ~n13216 & ~n13217;
  assign n13219 = pi1332 & pi2570;
  assign n13220 = pi1335 & pi2586;
  assign n13221 = ~n13219 & ~n13220;
  assign n13222 = n13218 & n13221;
  assign n13223 = n9726 & ~n13222;
  assign n13224 = pi0954 & n9614;
  assign n13225 = pi1899 & n9618;
  assign n13226 = ~n13224 & ~n13225;
  assign n13227 = pi0801 & n9687;
  assign n13228 = pi1439 & n9691;
  assign n13229 = ~n13227 & ~n13228;
  assign n13230 = pi0964 & n9607;
  assign n13231 = n13229 & ~n13230;
  assign n13232 = n13226 & n13231;
  assign n13233 = pi1831 & n9698;
  assign n13234 = n13232 & ~n13233;
  assign n13235 = pi0881 & n9715;
  assign n13236 = pi1885 & n9718;
  assign n13237 = ~n13235 & ~n13236;
  assign n13238 = pi0949 & n9702;
  assign n13239 = n13237 & ~n13238;
  assign n13240 = pi1730 & n11106;
  assign n13241 = pi0743 & n9707;
  assign n13242 = ~n13240 & ~n13241;
  assign n13243 = n13239 & n13242;
  assign n13244 = pi0770 & n9654;
  assign n13245 = pi2496 & n11158;
  assign n13246 = ~n13244 & ~n13245;
  assign n13247 = pi0773 & n9670;
  assign n13248 = pi1474 & n9676;
  assign n13249 = ~n13247 & ~n13248;
  assign n13250 = pi2504 & n9647;
  assign n13251 = n13249 & ~n13250;
  assign n13252 = n13246 & n13251;
  assign n13253 = pi1939 & n11165;
  assign n13254 = n13252 & ~n13253;
  assign n13255 = pi2104 & n9628;
  assign n13256 = pi1099 & n9631;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = pi1763 & n9657;
  assign n13259 = pi1752 & n9659;
  assign n13260 = ~n13258 & ~n13259;
  assign n13261 = n13257 & n13260;
  assign n13262 = pi1428 & n11133;
  assign n13263 = pi0577 & n9682;
  assign n13264 = ~n13262 & ~n13263;
  assign n13265 = pi1716 & n9679;
  assign n13266 = n13264 & ~n13265;
  assign n13267 = pi1922 & n9622;
  assign n13268 = n13266 & ~n13267;
  assign n13269 = n13261 & n13268;
  assign n13270 = ~n11102 & n13269;
  assign n13271 = n13254 & n13270;
  assign n13272 = pi1775 & n9712;
  assign n13273 = n13271 & ~n13272;
  assign n13274 = pi1453 & n11145;
  assign n13275 = pi0904 & n9710;
  assign n13276 = ~n13274 & ~n13275;
  assign n13277 = n13273 & n13276;
  assign n13278 = n13243 & n13277;
  assign n13279 = n13234 & n13278;
  assign n13280 = pi1934 & ~n13279;
  assign n13281 = ~n13223 & ~n13280;
  assign n13282 = pi0487 & ~pi0979;
  assign n13283 = pi0484 & pi0979;
  assign n13284 = ~n13282 & ~n13283;
  assign n13285 = pi0718 & ~n13284;
  assign n13286 = ~pi0979 & pi2844;
  assign n13287 = pi0979 & pi2127;
  assign n13288 = ~n13286 & ~n13287;
  assign n13289 = pi0717 & ~n13288;
  assign n13290 = ~n13285 & ~n13289;
  assign n13291 = pi0264 & ~pi0979;
  assign n13292 = pi0260 & pi0979;
  assign n13293 = ~n13291 & ~n13292;
  assign n13294 = pi0716 & ~n13293;
  assign n13295 = pi0290 & ~pi0979;
  assign n13296 = pi0287 & pi0979;
  assign n13297 = ~n13295 & ~n13296;
  assign n13298 = pi0761 & ~n13297;
  assign n13299 = ~n13294 & ~n13298;
  assign n13300 = n13290 & n13299;
  assign n13301 = ~n9535 & n13300;
  assign n13302 = n9523 & ~n13301;
  assign n13303 = n13281 & ~n13302;
  assign n13304 = n13215 & n13303;
  assign n13305 = pi0385 & pi1057;
  assign n13306 = pi1053 & pi2473;
  assign n13307 = ~n13305 & ~n13306;
  assign n13308 = pi0915 & pi1358;
  assign n13309 = n13307 & ~n13308;
  assign n13310 = pi1334 & pi2767;
  assign n13311 = pi0826 & pi1344;
  assign n13312 = ~n13310 & ~n13311;
  assign n13313 = pi3517 & ~n10410;
  assign n13314 = pi1331 & ~n8987;
  assign n13315 = pi0572 & pi1359;
  assign n13316 = ~n13314 & ~n13315;
  assign n13317 = ~n13313 & n13316;
  assign n13318 = n13312 & n13317;
  assign n13319 = n13309 & n13318;
  assign n13320 = n9475 & ~n13319;
  assign n13321 = n13304 & ~n13320;
  assign n13322 = pi1355 & pi2454;
  assign n13323 = pi1356 & pi3093;
  assign n13324 = ~n13322 & ~n13323;
  assign n13325 = pi1357 & pi2462;
  assign n13326 = n13324 & ~n13325;
  assign n13327 = pi1354 & pi2962;
  assign n13328 = n13326 & ~n13327;
  assign n13329 = pi1349 & pi2730;
  assign n13330 = pi1056 & pi2740;
  assign n13331 = ~n13329 & ~n13330;
  assign n13332 = pi1340 & pi2282;
  assign n13333 = pi1341 & pi2294;
  assign n13334 = ~n13332 & ~n13333;
  assign n13335 = pi1342 & pi2305;
  assign n13336 = n13334 & ~n13335;
  assign n13337 = pi1055 & pi2528;
  assign n13338 = n13336 & ~n13337;
  assign n13339 = pi1343 & pi2317;
  assign n13340 = pi1054 & pi2711;
  assign n13341 = ~n13339 & ~n13340;
  assign n13342 = n13338 & n13341;
  assign n13343 = n13331 & n13342;
  assign n13344 = n13328 & n13343;
  assign n13345 = n9736 & ~n13344;
  assign n13346 = pi1600 & pi2204;
  assign n13347 = pi1337 & pi2218;
  assign n13348 = ~n13346 & ~n13347;
  assign n13349 = pi1338 & pi2232;
  assign n13350 = n13348 & ~n13349;
  assign n13351 = pi1346 & pi2664;
  assign n13352 = n13350 & ~n13351;
  assign n13353 = pi1339 & pi2246;
  assign n13354 = pi1345 & pi2650;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = pi1351 & pi2262;
  assign n13357 = pi1352 & pi2272;
  assign n13358 = ~n13356 & ~n13357;
  assign n13359 = pi1353 & pi1977;
  assign n13360 = n13358 & ~n13359;
  assign n13361 = pi1350 & pi2258;
  assign n13362 = n13360 & ~n13361;
  assign n13363 = pi1347 & pi2678;
  assign n13364 = pi1348 & pi2563;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = n13362 & n13365;
  assign n13367 = n13355 & n13366;
  assign n13368 = n13352 & n13367;
  assign n13369 = n9577 & ~n13368;
  assign n13370 = ~n13345 & ~n13369;
  assign n13371 = n13321 & n13370;
  assign n13372 = pi3298 & po3871;
  assign n13373 = n13371 & ~n13372;
  assign n13374 = ~pi1787 & ~n13373;
  assign n13375 = pi1787 & pi2819;
  assign n13376 = ~n13374 & ~n13375;
  assign n13377 = n9472 & ~n13376;
  assign n13378 = pi3865 & n9804;
  assign n13379 = pi3881 & n9774;
  assign n13380 = ~n13378 & ~n13379;
  assign n13381 = pi3849 & n9802;
  assign n13382 = pi3913 & n9781;
  assign n13383 = pi3897 & n9771;
  assign n13384 = ~n13382 & ~n13383;
  assign n13385 = pi3945 & n9791;
  assign n13386 = pi3929 & n9788;
  assign n13387 = ~n13385 & ~n13386;
  assign n13388 = n13384 & n13387;
  assign n13389 = ~n13381 & n13388;
  assign n13390 = n13380 & n13389;
  assign n13391 = pi3865 & n9799;
  assign n13392 = n13390 & ~n13391;
  assign n13393 = pi3977 & n9783;
  assign n13394 = pi3961 & n9793;
  assign n13395 = ~n13393 & ~n13394;
  assign n13396 = n13392 & n13395;
  assign n13397 = ~n9472 & ~n13396;
  assign n13398 = ~n13377 & ~n13397;
  assign n13399 = n11186 & ~n13398;
  assign n13400 = ~n10902 & n13399;
  assign n13401 = n12803 & n12829;
  assign n13402 = ~n11697 & ~n13401;
  assign n13403 = ~n11186 & n13402;
  assign n13404 = ~n13400 & ~n13403;
  assign n13405 = n10885 & ~n13404;
  assign n13406 = ~n13152 & ~n13405;
  assign po0223 = n12885 | ~n13406;
  assign n13408 = n11186 & ~n13121;
  assign n13409 = ~n10902 & n13408;
  assign n13410 = pi2258 & n9837;
  assign n13411 = pi2272 & n9834;
  assign n13412 = ~n13410 & ~n13411;
  assign n13413 = pi2262 & n9839;
  assign n13414 = pi1977 & n9832;
  assign n13415 = ~n13413 & ~n13414;
  assign n13416 = n13412 & n13415;
  assign n13417 = ~n9424 & ~n13416;
  assign n13418 = pi2258 & n10374;
  assign n13419 = pi2272 & n10381;
  assign n13420 = ~n13418 & ~n13419;
  assign n13421 = pi2262 & n10376;
  assign n13422 = pi1977 & n10379;
  assign n13423 = ~n13421 & ~n13422;
  assign n13424 = n13420 & n13423;
  assign n13425 = n9424 & ~n13424;
  assign n13426 = ~n13417 & ~n13425;
  assign n13427 = n12880 & n13426;
  assign n13428 = ~n11697 & ~n13427;
  assign n13429 = ~n11186 & n13428;
  assign n13430 = ~n13409 & ~n13429;
  assign n13431 = n10885 & ~n13430;
  assign n13432 = n10216 & ~n12757;
  assign n13433 = ~n10216 & n12757;
  assign n13434 = ~n13432 & ~n13433;
  assign n13435 = n10296 & ~n13434;
  assign n13436 = ~n10232 & ~n10281;
  assign n13437 = ~n12765 & ~n13436;
  assign n13438 = n12765 & n13436;
  assign n13439 = ~n13437 & ~n13438;
  assign n13440 = ~n10296 & ~n13439;
  assign n13441 = ~n13435 & ~n13440;
  assign n13442 = ~pi0568 & ~n13441;
  assign n13443 = n10362 & ~n13439;
  assign n13444 = ~n10362 & ~n13434;
  assign n13445 = ~n13443 & ~n13444;
  assign n13446 = pi0568 & ~n13445;
  assign n13447 = ~n13442 & ~n13446;
  assign n13448 = pi0642 & n10209;
  assign n13449 = pi0642 & n10211;
  assign n13450 = ~n13448 & ~n13449;
  assign n13451 = n13447 & n13450;
  assign n13452 = ~n11186 & ~n13451;
  assign n13453 = n11701 & ~n13426;
  assign n13454 = pi1031 & ~n11706;
  assign n13455 = pi0904 & n11709;
  assign n13456 = pi2450 & po3871;
  assign n13457 = ~n13455 & ~n13456;
  assign n13458 = pi0426 & n11714;
  assign n13459 = n13457 & ~n13458;
  assign n13460 = ~n13454 & n13459;
  assign n13461 = ~n11700 & n13460;
  assign n13462 = n10886 & ~n12880;
  assign n13463 = n13461 & ~n13462;
  assign n13464 = ~n13453 & n13463;
  assign n13465 = ~pi0773 & n11700;
  assign n13466 = ~n13464 & ~n13465;
  assign n13467 = ~n10914 & n13466;
  assign n13468 = ~n13452 & ~n13467;
  assign n13469 = ~n11697 & ~n13468;
  assign n13470 = ~n11186 & ~n13149;
  assign n13471 = n11186 & ~n12829;
  assign n13472 = ~n13470 & ~n13471;
  assign n13473 = n10902 & ~n13472;
  assign n13474 = ~n13469 & ~n13473;
  assign n13475 = ~n10885 & ~n13474;
  assign n13476 = n10914 & n13398;
  assign n13477 = ~n10914 & n12862;
  assign n13478 = ~n13476 & ~n13477;
  assign n13479 = n11755 & n13478;
  assign n13480 = ~n13475 & ~n13479;
  assign po0222 = n13431 | ~n13480;
  assign n13482 = po0223 & po0222;
  assign n13483 = po0229 & n13482;
  assign n13484 = pi3867 & n9804;
  assign n13485 = pi3883 & n9774;
  assign n13486 = ~n13484 & ~n13485;
  assign n13487 = pi3851 & n9802;
  assign n13488 = pi3915 & n9781;
  assign n13489 = pi3899 & n9771;
  assign n13490 = ~n13488 & ~n13489;
  assign n13491 = pi3947 & n9791;
  assign n13492 = pi3931 & n9788;
  assign n13493 = ~n13491 & ~n13492;
  assign n13494 = n13490 & n13493;
  assign n13495 = ~n13487 & n13494;
  assign n13496 = n13486 & n13495;
  assign n13497 = pi3867 & n9799;
  assign n13498 = n13496 & ~n13497;
  assign n13499 = pi3979 & n9783;
  assign n13500 = pi3963 & n9793;
  assign n13501 = ~n13499 & ~n13500;
  assign n13502 = n13498 & n13501;
  assign n13503 = ~n9472 & ~n13502;
  assign n13504 = pi0913 & pi1358;
  assign n13505 = pi0383 & pi1057;
  assign n13506 = ~n13504 & ~n13505;
  assign n13507 = pi3518 & ~n10410;
  assign n13508 = pi1331 & ~n9142;
  assign n13509 = pi0602 & pi1359;
  assign n13510 = ~n13508 & ~n13509;
  assign n13511 = ~n13507 & n13510;
  assign n13512 = n13506 & n13511;
  assign n13513 = n9475 & ~n13512;
  assign n13514 = ~pi0979 & pi2612;
  assign n13515 = pi0979 & pi2606;
  assign n13516 = ~n13514 & ~n13515;
  assign n13517 = pi0763 & ~n13516;
  assign n13518 = ~pi0979 & pi2625;
  assign n13519 = pi0979 & pi2619;
  assign n13520 = ~n13518 & ~n13519;
  assign n13521 = pi0764 & ~n13520;
  assign n13522 = ~n13517 & ~n13521;
  assign n13523 = ~pi0979 & pi2631;
  assign n13524 = pi0979 & pi3168;
  assign n13525 = ~n13523 & ~n13524;
  assign n13526 = pi0765 & ~n13525;
  assign n13527 = ~pi0979 & pi2889;
  assign n13528 = pi0979 & pi3177;
  assign n13529 = ~n13527 & ~n13528;
  assign n13530 = pi0766 & ~n13529;
  assign n13531 = ~n13526 & ~n13530;
  assign n13532 = pi0146 & ~pi0979;
  assign n13533 = pi0145 & pi0979;
  assign n13534 = ~n13532 & ~n13533;
  assign n13535 = pi0720 & ~n13534;
  assign n13536 = pi0294 & ~pi0979;
  assign n13537 = pi0293 & pi0979;
  assign n13538 = ~n13536 & ~n13537;
  assign n13539 = pi0721 & ~n13538;
  assign n13540 = ~n13535 & ~n13539;
  assign n13541 = n13531 & n13540;
  assign n13542 = ~n9499 & n13541;
  assign n13543 = n13522 & n13542;
  assign n13544 = n9486 & ~n13543;
  assign n13545 = ~n13513 & ~n13544;
  assign n13546 = ~pi0979 & pi2842;
  assign n13547 = pi0979 & pi2125;
  assign n13548 = ~n13546 & ~n13547;
  assign n13549 = pi0717 & ~n13548;
  assign n13550 = pi0239 & ~pi0979;
  assign n13551 = pi0238 & pi0979;
  assign n13552 = ~n13550 & ~n13551;
  assign n13553 = pi0716 & ~n13552;
  assign n13554 = pi0236 & ~pi0979;
  assign n13555 = pi0235 & pi0979;
  assign n13556 = ~n13554 & ~n13555;
  assign n13557 = pi0761 & ~n13556;
  assign n13558 = ~n13553 & ~n13557;
  assign n13559 = ~n9535 & n13558;
  assign n13560 = ~n9531 & n13559;
  assign n13561 = ~n13549 & n13560;
  assign n13562 = n9523 & ~n13561;
  assign n13563 = pi0979 & pi2162;
  assign n13564 = ~pi0979 & pi2809;
  assign n13565 = ~n13563 & ~n13564;
  assign n13566 = pi0836 & ~n13565;
  assign n13567 = ~pi0979 & pi2940;
  assign n13568 = pi0979 & pi2178;
  assign n13569 = ~n13567 & ~n13568;
  assign n13570 = pi0837 & ~n13569;
  assign n13571 = ~n13566 & ~n13570;
  assign n13572 = pi0979 & pi2145;
  assign n13573 = ~pi0979 & pi2917;
  assign n13574 = ~n13572 & ~n13573;
  assign n13575 = pi0767 & ~n13574;
  assign n13576 = ~pi0979 & pi2421;
  assign n13577 = pi0979 & pi1956;
  assign n13578 = ~n13576 & ~n13577;
  assign n13579 = pi0768 & ~n13578;
  assign n13580 = ~n13575 & ~n13579;
  assign n13581 = pi0168 & ~pi0979;
  assign n13582 = pi0154 & pi0979;
  assign n13583 = ~n13581 & ~n13582;
  assign n13584 = pi0838 & ~n13583;
  assign n13585 = n13580 & ~n13584;
  assign n13586 = n13571 & n13585;
  assign n13587 = n9549 & ~n13586;
  assign n13588 = ~n13562 & ~n13587;
  assign n13589 = pi1347 & pi2676;
  assign n13590 = pi1348 & pi2687;
  assign n13591 = ~n13589 & ~n13590;
  assign n13592 = pi1350 & pi2698;
  assign n13593 = n13591 & ~n13592;
  assign n13594 = pi1353 & pi2275;
  assign n13595 = n13593 & ~n13594;
  assign n13596 = pi1351 & pi2438;
  assign n13597 = pi1352 & pi2701;
  assign n13598 = ~n13596 & ~n13597;
  assign n13599 = pi1600 & pi2202;
  assign n13600 = pi1337 & pi2216;
  assign n13601 = ~n13599 & ~n13600;
  assign n13602 = pi1338 & pi2230;
  assign n13603 = n13601 & ~n13602;
  assign n13604 = pi1346 & pi2662;
  assign n13605 = n13603 & ~n13604;
  assign n13606 = pi1339 & pi2244;
  assign n13607 = pi1345 & pi2648;
  assign n13608 = ~n13606 & ~n13607;
  assign n13609 = n13605 & n13608;
  assign n13610 = n13598 & n13609;
  assign n13611 = n13595 & n13610;
  assign n13612 = n9577 & ~n13611;
  assign n13613 = pi1355 & pi2520;
  assign n13614 = pi1356 & pi2752;
  assign n13615 = ~n13613 & ~n13614;
  assign n13616 = pi1357 & pi2412;
  assign n13617 = n13615 & ~n13616;
  assign n13618 = pi1354 & pi2535;
  assign n13619 = n13617 & ~n13618;
  assign n13620 = pi1349 & pi2566;
  assign n13621 = pi1056 & pi2739;
  assign n13622 = ~n13620 & ~n13621;
  assign n13623 = pi1343 & pi2315;
  assign n13624 = pi1054 & pi2709;
  assign n13625 = ~n13623 & ~n13624;
  assign n13626 = pi1055 & pi2720;
  assign n13627 = n13625 & ~n13626;
  assign n13628 = pi1342 & pi2089;
  assign n13629 = n13627 & ~n13628;
  assign n13630 = pi1340 & pi2280;
  assign n13631 = pi1341 & pi2067;
  assign n13632 = ~n13630 & ~n13631;
  assign n13633 = n13629 & n13632;
  assign n13634 = n13622 & n13633;
  assign n13635 = n13619 & n13634;
  assign n13636 = n9736 & ~n13635;
  assign n13637 = ~n13612 & ~n13636;
  assign n13638 = pi0232 & pi1336;
  assign n13639 = pi1333 & pi1741;
  assign n13640 = ~n13638 & ~n13639;
  assign n13641 = pi1332 & pi2568;
  assign n13642 = pi1335 & pi2584;
  assign n13643 = ~n13641 & ~n13642;
  assign n13644 = n13640 & n13643;
  assign n13645 = n9726 & ~n13644;
  assign n13646 = pi1848 & n10557;
  assign n13647 = pi0941 & n9614;
  assign n13648 = pi1898 & n9618;
  assign n13649 = ~n13647 & ~n13648;
  assign n13650 = ~n13646 & n13649;
  assign n13651 = pi0968 & n9687;
  assign n13652 = pi1437 & n9691;
  assign n13653 = ~n13651 & ~n13652;
  assign n13654 = pi0790 & n9715;
  assign n13655 = pi1883 & n9718;
  assign n13656 = ~n13654 & ~n13655;
  assign n13657 = pi1728 & n11106;
  assign n13658 = pi0894 & n9707;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = pi1847 & n10564;
  assign n13661 = n13659 & ~n13660;
  assign n13662 = n13656 & n13661;
  assign n13663 = pi1829 & n9698;
  assign n13664 = n13662 & ~n13663;
  assign n13665 = ~n11102 & n13664;
  assign n13666 = n13653 & n13665;
  assign n13667 = n13650 & n13666;
  assign n13668 = pi1773 & n9712;
  assign n13669 = n13667 & ~n13668;
  assign n13670 = pi1451 & n11145;
  assign n13671 = pi0903 & n9710;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = pi0732 & n9654;
  assign n13674 = pi3101 & n9647;
  assign n13675 = ~n13673 & ~n13674;
  assign n13676 = pi0862 & n9670;
  assign n13677 = pi0928 & n9676;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = pi2494 & n11158;
  assign n13680 = n13678 & ~n13679;
  assign n13681 = n13675 & n13680;
  assign n13682 = pi1919 & n9622;
  assign n13683 = n13681 & ~n13682;
  assign n13684 = pi1878 & n9679;
  assign n13685 = pi0458 & n9682;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = n13683 & n13686;
  assign n13688 = n13672 & n13687;
  assign n13689 = n13669 & n13688;
  assign n13690 = pi1934 & ~n13689;
  assign n13691 = ~n13645 & ~n13690;
  assign n13692 = n13637 & n13691;
  assign n13693 = n13588 & n13692;
  assign n13694 = n13545 & n13693;
  assign n13695 = pi3307 & po3871;
  assign n13696 = n13694 & ~n13695;
  assign n13697 = ~pi1787 & ~n13696;
  assign n13698 = pi1787 & pi3150;
  assign n13699 = ~n13697 & ~n13698;
  assign n13700 = n9472 & ~n13699;
  assign n13701 = ~n13503 & ~n13700;
  assign n13702 = ~n10914 & ~n13701;
  assign n13703 = ~n11697 & n13702;
  assign n13704 = pi2753 & n11190;
  assign n13705 = pi2746 & n11197;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = pi2527 & n11195;
  assign n13708 = pi2463 & n11192;
  assign n13709 = ~n13707 & ~n13708;
  assign n13710 = n13706 & n13709;
  assign n13711 = n9424 & ~n13710;
  assign n13712 = pi2753 & n11204;
  assign n13713 = pi2527 & n11209;
  assign n13714 = ~n13712 & ~n13713;
  assign n13715 = pi2746 & n11207;
  assign n13716 = pi2463 & n11202;
  assign n13717 = ~n13715 & ~n13716;
  assign n13718 = n13714 & n13717;
  assign n13719 = ~n9424 & ~n13718;
  assign n13720 = ~n13711 & ~n13719;
  assign n13721 = pi1978 & n9832;
  assign n13722 = pi2442 & n9834;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = pi2432 & n9837;
  assign n13725 = pi2263 & n9839;
  assign n13726 = ~n13724 & ~n13725;
  assign n13727 = n13723 & n13726;
  assign n13728 = ~n9424 & ~n13727;
  assign n13729 = pi2432 & n10374;
  assign n13730 = pi2442 & n10381;
  assign n13731 = ~n13729 & ~n13730;
  assign n13732 = pi2263 & n10376;
  assign n13733 = pi1978 & n10379;
  assign n13734 = ~n13732 & ~n13733;
  assign n13735 = n13731 & n13734;
  assign n13736 = n9424 & ~n13735;
  assign n13737 = ~n13728 & ~n13736;
  assign n13738 = n13720 & n13737;
  assign n13739 = ~n11697 & ~n13738;
  assign n13740 = ~n11186 & n13739;
  assign n13741 = ~n13703 & ~n13740;
  assign n13742 = n10885 & ~n13741;
  assign n13743 = pi3864 & n9804;
  assign n13744 = pi3880 & n9774;
  assign n13745 = ~n13743 & ~n13744;
  assign n13746 = pi3848 & n9802;
  assign n13747 = pi3912 & n9781;
  assign n13748 = pi3896 & n9771;
  assign n13749 = ~n13747 & ~n13748;
  assign n13750 = pi3944 & n9791;
  assign n13751 = pi3928 & n9788;
  assign n13752 = ~n13750 & ~n13751;
  assign n13753 = n13749 & n13752;
  assign n13754 = ~n13746 & n13753;
  assign n13755 = n13745 & n13754;
  assign n13756 = pi3864 & n9799;
  assign n13757 = n13755 & ~n13756;
  assign n13758 = pi3976 & n9783;
  assign n13759 = pi3960 & n9793;
  assign n13760 = ~n13758 & ~n13759;
  assign n13761 = n13757 & n13760;
  assign n13762 = ~n9472 & ~n13761;
  assign n13763 = pi0916 & pi1358;
  assign n13764 = pi0386 & pi1057;
  assign n13765 = pi1053 & pi2404;
  assign n13766 = ~n13764 & ~n13765;
  assign n13767 = pi1331 & ~n8876;
  assign n13768 = pi0578 & pi1359;
  assign n13769 = ~n13767 & ~n13768;
  assign n13770 = pi1334 & pi2379;
  assign n13771 = pi0827 & pi1344;
  assign n13772 = ~n13770 & ~n13771;
  assign n13773 = n13769 & n13772;
  assign n13774 = n13766 & n13773;
  assign n13775 = ~n13763 & n13774;
  assign n13776 = pi3508 & ~n10410;
  assign n13777 = n13775 & ~n13776;
  assign n13778 = n9475 & ~n13777;
  assign n13779 = pi0488 & ~pi0979;
  assign n13780 = pi0485 & pi0979;
  assign n13781 = ~n13779 & ~n13780;
  assign n13782 = pi0718 & ~n13781;
  assign n13783 = ~pi0979 & pi2845;
  assign n13784 = pi0979 & pi2128;
  assign n13785 = ~n13783 & ~n13784;
  assign n13786 = pi0717 & ~n13785;
  assign n13787 = ~n13782 & ~n13786;
  assign n13788 = pi0263 & ~pi0979;
  assign n13789 = pi0259 & pi0979;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = pi0716 & ~n13790;
  assign n13792 = pi0291 & ~pi0979;
  assign n13793 = pi0288 & pi0979;
  assign n13794 = ~n13792 & ~n13793;
  assign n13795 = pi0761 & ~n13794;
  assign n13796 = ~n13791 & ~n13795;
  assign n13797 = n13787 & n13796;
  assign n13798 = ~n9535 & n13797;
  assign n13799 = n9523 & ~n13798;
  assign n13800 = ~n13778 & ~n13799;
  assign n13801 = pi0979 & pi2165;
  assign n13802 = ~pi0979 & pi2807;
  assign n13803 = ~n13801 & ~n13802;
  assign n13804 = pi0836 & ~n13803;
  assign n13805 = ~pi0979 & pi2942;
  assign n13806 = pi0979 & pi2181;
  assign n13807 = ~n13805 & ~n13806;
  assign n13808 = pi0837 & ~n13807;
  assign n13809 = ~n13804 & ~n13808;
  assign n13810 = pi0979 & pi2085;
  assign n13811 = ~pi0979 & pi2787;
  assign n13812 = ~n13810 & ~n13811;
  assign n13813 = pi0767 & ~n13812;
  assign n13814 = ~pi0979 & pi2424;
  assign n13815 = pi0979 & pi1959;
  assign n13816 = ~n13814 & ~n13815;
  assign n13817 = pi0768 & ~n13816;
  assign n13818 = ~n13813 & ~n13817;
  assign n13819 = pi0171 & ~pi0979;
  assign n13820 = pi0157 & pi0979;
  assign n13821 = ~n13819 & ~n13820;
  assign n13822 = pi0838 & ~n13821;
  assign n13823 = pi0143 & pi1360;
  assign n13824 = ~n13822 & ~n13823;
  assign n13825 = n13818 & n13824;
  assign n13826 = n13809 & n13825;
  assign n13827 = n9549 & ~n13826;
  assign n13828 = ~pi0979 & pi2864;
  assign n13829 = pi0979 & pi3153;
  assign n13830 = ~n13828 & ~n13829;
  assign n13831 = pi0763 & ~n13830;
  assign n13832 = ~pi0979 & pi2872;
  assign n13833 = pi0979 & pi3162;
  assign n13834 = ~n13832 & ~n13833;
  assign n13835 = pi0764 & ~n13834;
  assign n13836 = ~n13831 & ~n13835;
  assign n13837 = pi0191 & ~pi0979;
  assign n13838 = pi0190 & pi0979;
  assign n13839 = ~n13837 & ~n13838;
  assign n13840 = pi0720 & ~n13839;
  assign n13841 = pi0335 & ~pi0979;
  assign n13842 = pi0334 & pi0979;
  assign n13843 = ~n13841 & ~n13842;
  assign n13844 = pi0721 & ~n13843;
  assign n13845 = ~n13840 & ~n13844;
  assign n13846 = pi0064 & ~pi0979;
  assign n13847 = pi0062 & pi0979;
  assign n13848 = ~n13846 & ~n13847;
  assign n13849 = pi0719 & ~n13848;
  assign n13850 = ~pi0979 & pi2634;
  assign n13851 = pi0979 & pi3134;
  assign n13852 = ~n13850 & ~n13851;
  assign n13853 = pi0765 & ~n13852;
  assign n13854 = ~pi0979 & pi3074;
  assign n13855 = pi0979 & pi3179;
  assign n13856 = ~n13854 & ~n13855;
  assign n13857 = pi0766 & ~n13856;
  assign n13858 = ~n13853 & ~n13857;
  assign n13859 = ~n13849 & n13858;
  assign n13860 = n13845 & n13859;
  assign n13861 = n13836 & n13860;
  assign n13862 = n9486 & ~n13861;
  assign n13863 = ~n13827 & ~n13862;
  assign n13864 = pi1340 & pi2283;
  assign n13865 = pi1341 & pi2295;
  assign n13866 = ~n13864 & ~n13865;
  assign n13867 = pi1342 & pi2084;
  assign n13868 = n13866 & ~n13867;
  assign n13869 = pi1055 & pi2721;
  assign n13870 = n13868 & ~n13869;
  assign n13871 = pi1343 & pi2318;
  assign n13872 = pi1054 & pi2536;
  assign n13873 = ~n13871 & ~n13872;
  assign n13874 = pi1355 & pi2527;
  assign n13875 = pi1356 & pi2753;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = pi1357 & pi2463;
  assign n13878 = n13876 & ~n13877;
  assign n13879 = pi1354 & pi2746;
  assign n13880 = n13878 & ~n13879;
  assign n13881 = pi1349 & pi2731;
  assign n13882 = pi1056 & pi2741;
  assign n13883 = ~n13881 & ~n13882;
  assign n13884 = n13880 & n13883;
  assign n13885 = n13873 & n13884;
  assign n13886 = n13870 & n13885;
  assign n13887 = n9736 & ~n13886;
  assign n13888 = pi1339 & pi2247;
  assign n13889 = pi1345 & pi2651;
  assign n13890 = ~n13888 & ~n13889;
  assign n13891 = pi1346 & pi2665;
  assign n13892 = n13890 & ~n13891;
  assign n13893 = pi1338 & pi2233;
  assign n13894 = n13892 & ~n13893;
  assign n13895 = pi1600 & pi2205;
  assign n13896 = pi1337 & pi2219;
  assign n13897 = ~n13895 & ~n13896;
  assign n13898 = pi1347 & pi2679;
  assign n13899 = pi1348 & pi2689;
  assign n13900 = ~n13898 & ~n13899;
  assign n13901 = pi1350 & pi2432;
  assign n13902 = n13900 & ~n13901;
  assign n13903 = pi1353 & pi1978;
  assign n13904 = n13902 & ~n13903;
  assign n13905 = pi1351 & pi2263;
  assign n13906 = pi1352 & pi2442;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = n13904 & n13907;
  assign n13909 = n13897 & n13908;
  assign n13910 = n13894 & n13909;
  assign n13911 = n9577 & ~n13910;
  assign n13912 = ~n13887 & ~n13911;
  assign n13913 = pi0278 & pi1336;
  assign n13914 = pi0314 & pi1333;
  assign n13915 = ~n13913 & ~n13914;
  assign n13916 = pi1332 & pi2571;
  assign n13917 = pi1335 & pi2764;
  assign n13918 = ~n13916 & ~n13917;
  assign n13919 = n13915 & n13918;
  assign n13920 = n9726 & ~n13919;
  assign n13921 = pi0882 & n9715;
  assign n13922 = pi1920 & n9718;
  assign n13923 = ~n13921 & ~n13922;
  assign n13924 = pi1731 & n11106;
  assign n13925 = pi0744 & n9707;
  assign n13926 = ~n13924 & ~n13925;
  assign n13927 = pi0950 & n9702;
  assign n13928 = n13926 & ~n13927;
  assign n13929 = n13923 & n13928;
  assign n13930 = pi1832 & n9698;
  assign n13931 = n13929 & ~n13930;
  assign n13932 = pi0955 & n9614;
  assign n13933 = pi2054 & n9618;
  assign n13934 = ~n13932 & ~n13933;
  assign n13935 = pi0965 & n9607;
  assign n13936 = n13934 & ~n13935;
  assign n13937 = pi0802 & n9687;
  assign n13938 = pi1440 & n9691;
  assign n13939 = ~n13937 & ~n13938;
  assign n13940 = n13936 & n13939;
  assign n13941 = pi0774 & n9670;
  assign n13942 = pi1603 & n9676;
  assign n13943 = ~n13941 & ~n13942;
  assign n13944 = pi0771 & n9654;
  assign n13945 = pi2497 & n11158;
  assign n13946 = ~n13944 & ~n13945;
  assign n13947 = pi2522 & n9647;
  assign n13948 = n13946 & ~n13947;
  assign n13949 = n13943 & n13948;
  assign n13950 = pi1940 & n11165;
  assign n13951 = n13949 & ~n13950;
  assign n13952 = pi2105 & n9628;
  assign n13953 = pi1021 & n9631;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = pi1764 & n9657;
  assign n13956 = pi1753 & n9659;
  assign n13957 = ~n13955 & ~n13956;
  assign n13958 = n13954 & n13957;
  assign n13959 = pi1429 & n11133;
  assign n13960 = pi0653 & n9682;
  assign n13961 = ~n13959 & ~n13960;
  assign n13962 = pi1717 & n9679;
  assign n13963 = n13961 & ~n13962;
  assign n13964 = pi1923 & n9622;
  assign n13965 = n13963 & ~n13964;
  assign n13966 = n13958 & n13965;
  assign n13967 = ~n11102 & n13966;
  assign n13968 = n13951 & n13967;
  assign n13969 = pi1776 & n9712;
  assign n13970 = n13968 & ~n13969;
  assign n13971 = pi1454 & n11145;
  assign n13972 = pi0905 & n9710;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = n13970 & n13973;
  assign n13975 = n13940 & n13974;
  assign n13976 = n13931 & n13975;
  assign n13977 = pi1934 & ~n13976;
  assign n13978 = ~n13920 & ~n13977;
  assign n13979 = n13912 & n13978;
  assign n13980 = n13863 & n13979;
  assign n13981 = n13800 & n13980;
  assign n13982 = pi3309 & po3871;
  assign n13983 = n13981 & ~n13982;
  assign n13984 = ~pi1787 & ~n13983;
  assign n13985 = pi1787 & pi2827;
  assign n13986 = ~n13984 & ~n13985;
  assign n13987 = n9472 & ~n13986;
  assign n13988 = ~n13762 & ~n13987;
  assign n13989 = ~n11186 & n13988;
  assign n13990 = pi0678 & ~n11393;
  assign n13991 = n11260 & n13990;
  assign n13992 = pi0678 & n11550;
  assign n13993 = ~n11580 & ~n11643;
  assign n13994 = ~n11582 & ~n13993;
  assign n13995 = n11584 & n13994;
  assign n13996 = ~n11584 & ~n13994;
  assign n13997 = ~n13995 & ~n13996;
  assign n13998 = n11615 & ~n13997;
  assign n13999 = ~n11524 & ~n11579;
  assign n14000 = ~n11592 & ~n13999;
  assign n14001 = ~n11583 & n11587;
  assign n14002 = n11583 & ~n11587;
  assign n14003 = ~n14001 & ~n14002;
  assign n14004 = n14000 & ~n14003;
  assign n14005 = ~n14000 & n14003;
  assign n14006 = ~n14004 & ~n14005;
  assign n14007 = ~n11615 & ~n14006;
  assign n14008 = ~n13998 & ~n14007;
  assign n14009 = ~pi0518 & ~n14008;
  assign n14010 = n11665 & ~n14006;
  assign n14011 = ~n11665 & ~n13997;
  assign n14012 = ~n14010 & ~n14011;
  assign n14013 = pi0518 & ~n14012;
  assign n14014 = ~n14009 & ~n14013;
  assign n14015 = ~n13992 & n14014;
  assign n14016 = ~n13991 & n14015;
  assign n14017 = n11186 & n14016;
  assign n14018 = ~n13989 & ~n14017;
  assign n14019 = n11755 & n14018;
  assign n14020 = ~n10262 & ~n10325;
  assign n14021 = ~n10261 & ~n14020;
  assign n14022 = n10265 & n14021;
  assign n14023 = ~n10265 & ~n14021;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = n10296 & ~n14024;
  assign n14026 = ~n10203 & ~n10260;
  assign n14027 = ~n10273 & ~n14026;
  assign n14028 = ~n10264 & n10268;
  assign n14029 = n10264 & ~n10268;
  assign n14030 = ~n14028 & ~n14029;
  assign n14031 = n14027 & ~n14030;
  assign n14032 = ~n14027 & n14030;
  assign n14033 = ~n14031 & ~n14032;
  assign n14034 = ~n10296 & ~n14033;
  assign n14035 = ~n14025 & ~n14034;
  assign n14036 = ~pi0568 & ~n14035;
  assign n14037 = n10362 & ~n14033;
  assign n14038 = ~n10362 & ~n14024;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = pi0568 & ~n14039;
  assign n14041 = ~n14036 & ~n14040;
  assign n14042 = pi0661 & n10222;
  assign n14043 = pi0661 & n9951;
  assign n14044 = ~n10038 & n14043;
  assign n14045 = ~n14042 & ~n14044;
  assign n14046 = n14041 & n14045;
  assign n14047 = n10914 & ~n14046;
  assign n14048 = n11701 & ~n13737;
  assign n14049 = pi1013 & ~n11706;
  assign n14050 = pi0905 & n11709;
  assign n14051 = pi2451 & po3871;
  assign n14052 = ~n14050 & ~n14051;
  assign n14053 = pi0409 & n11714;
  assign n14054 = n14052 & ~n14053;
  assign n14055 = ~n14049 & n14054;
  assign n14056 = ~n11700 & n14055;
  assign n14057 = n10886 & ~n13720;
  assign n14058 = n14056 & ~n14057;
  assign n14059 = ~n14048 & n14058;
  assign n14060 = ~pi0774 & n11700;
  assign n14061 = ~n14059 & ~n14060;
  assign n14062 = n11186 & n14061;
  assign n14063 = ~n14047 & ~n14062;
  assign n14064 = ~n10902 & ~n14063;
  assign n14065 = pi0677 & ~n11394;
  assign n14066 = n11260 & n14065;
  assign n14067 = pi0677 & n11398;
  assign n14068 = ~n11411 & n11648;
  assign n14069 = n11411 & ~n11648;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071 = n11615 & ~n14070;
  assign n14072 = ~n11414 & n11426;
  assign n14073 = n11414 & ~n11426;
  assign n14074 = ~n14072 & ~n14073;
  assign n14075 = n11604 & ~n14074;
  assign n14076 = ~n11604 & n14074;
  assign n14077 = ~n14075 & ~n14076;
  assign n14078 = ~n11615 & ~n14077;
  assign n14079 = ~n14071 & ~n14078;
  assign n14080 = ~pi0518 & ~n14079;
  assign n14081 = n11665 & ~n14077;
  assign n14082 = ~n11665 & ~n14070;
  assign n14083 = ~n14081 & ~n14082;
  assign n14084 = pi0518 & ~n14083;
  assign n14085 = ~n14080 & ~n14084;
  assign n14086 = ~n14067 & n14085;
  assign n14087 = ~n14066 & n14086;
  assign n14088 = n10914 & n14087;
  assign n14089 = pi2520 & n11195;
  assign n14090 = pi2535 & n11197;
  assign n14091 = ~n14089 & ~n14090;
  assign n14092 = pi2752 & n11190;
  assign n14093 = pi2412 & n11192;
  assign n14094 = ~n14092 & ~n14093;
  assign n14095 = n14091 & n14094;
  assign n14096 = n9424 & ~n14095;
  assign n14097 = pi2535 & n11207;
  assign n14098 = pi2520 & n11209;
  assign n14099 = ~n14097 & ~n14098;
  assign n14100 = pi2412 & n11202;
  assign n14101 = pi2752 & n11204;
  assign n14102 = ~n14100 & ~n14101;
  assign n14103 = n14099 & n14102;
  assign n14104 = ~n9424 & ~n14103;
  assign n14105 = ~n14096 & ~n14104;
  assign n14106 = ~n10914 & n14105;
  assign n14107 = ~n14088 & ~n14106;
  assign n14108 = n11697 & n14107;
  assign n14109 = ~n14064 & ~n14108;
  assign n14110 = ~n10885 & ~n14109;
  assign n14111 = ~n14019 & ~n14110;
  assign po0221 = n13742 | ~n14111;
  assign n14113 = ~n10057 & n10329;
  assign n14114 = n10057 & ~n10329;
  assign n14115 = ~n14113 & ~n14114;
  assign n14116 = n10296 & ~n14115;
  assign n14117 = ~n10060 & n10072;
  assign n14118 = n10060 & ~n10072;
  assign n14119 = ~n14117 & ~n14118;
  assign n14120 = n10284 & ~n14119;
  assign n14121 = ~n10284 & n14119;
  assign n14122 = ~n14120 & ~n14121;
  assign n14123 = ~n10296 & ~n14122;
  assign n14124 = ~n14116 & ~n14123;
  assign n14125 = ~pi0568 & ~n14124;
  assign n14126 = n10362 & ~n14122;
  assign n14127 = ~n10362 & ~n14115;
  assign n14128 = ~n14126 & ~n14127;
  assign n14129 = pi0568 & ~n14128;
  assign n14130 = ~n14125 & ~n14129;
  assign n14131 = pi0754 & n10043;
  assign n14132 = pi0754 & n10040;
  assign n14133 = ~n14131 & ~n14132;
  assign n14134 = n14130 & n14133;
  assign n14135 = n10914 & ~n14134;
  assign n14136 = pi1029 & ~n11706;
  assign n14137 = pi0903 & n11709;
  assign n14138 = pi2438 & n9839;
  assign n14139 = pi2701 & n9834;
  assign n14140 = ~n14138 & ~n14139;
  assign n14141 = pi2698 & n9837;
  assign n14142 = pi2275 & n9832;
  assign n14143 = ~n14141 & ~n14142;
  assign n14144 = n14140 & n14143;
  assign n14145 = ~n9424 & ~n14144;
  assign n14146 = pi2438 & n10376;
  assign n14147 = pi2701 & n10381;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = pi2698 & n10374;
  assign n14150 = pi2275 & n10379;
  assign n14151 = ~n14149 & ~n14150;
  assign n14152 = n14148 & n14151;
  assign n14153 = n9424 & ~n14152;
  assign n14154 = ~n14145 & ~n14153;
  assign n14155 = n11701 & ~n14154;
  assign n14156 = ~n14137 & ~n14155;
  assign n14157 = ~n14136 & n14156;
  assign n14158 = pi2415 & po3871;
  assign n14159 = n10886 & ~n14105;
  assign n14160 = pi0406 & n11714;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = ~n14158 & n14161;
  assign n14163 = n14157 & n14162;
  assign n14164 = ~n11700 & ~n14163;
  assign n14165 = pi0862 & n11700;
  assign n14166 = ~n14164 & ~n14165;
  assign n14167 = n11186 & ~n14166;
  assign n14168 = ~n14135 & ~n14167;
  assign n14169 = ~n10902 & ~n14168;
  assign n14170 = n10914 & n14016;
  assign n14171 = ~n10914 & n13720;
  assign n14172 = ~n14170 & ~n14171;
  assign n14173 = n11697 & n14172;
  assign n14174 = ~n14169 & ~n14173;
  assign n14175 = ~n10885 & ~n14174;
  assign n14176 = n10914 & n13701;
  assign n14177 = ~n10914 & n14087;
  assign n14178 = ~n14176 & ~n14177;
  assign n14179 = n11755 & n14178;
  assign n14180 = n11186 & ~n13988;
  assign n14181 = ~n10902 & n14180;
  assign n14182 = n14105 & n14154;
  assign n14183 = ~n11697 & ~n14182;
  assign n14184 = ~n11186 & n14183;
  assign n14185 = ~n14181 & ~n14184;
  assign n14186 = n10885 & ~n14185;
  assign n14187 = ~n14179 & ~n14186;
  assign po0224 = n14175 | ~n14187;
  assign n14189 = pi3869 & n9804;
  assign n14190 = pi3885 & n9774;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = pi3853 & n9802;
  assign n14193 = pi3981 & n9783;
  assign n14194 = pi3901 & n9771;
  assign n14195 = ~n14193 & ~n14194;
  assign n14196 = pi3949 & n9791;
  assign n14197 = pi3933 & n9788;
  assign n14198 = ~n14196 & ~n14197;
  assign n14199 = n14195 & n14198;
  assign n14200 = ~n14192 & n14199;
  assign n14201 = n14191 & n14200;
  assign n14202 = pi3869 & n9799;
  assign n14203 = n14201 & ~n14202;
  assign n14204 = pi3917 & n9781;
  assign n14205 = pi3965 & n9793;
  assign n14206 = ~n14204 & ~n14205;
  assign n14207 = n14203 & n14206;
  assign n14208 = ~n9472 & ~n14207;
  assign n14209 = pi1331 & ~n9179;
  assign n14210 = pi3504 & ~n10410;
  assign n14211 = ~n14209 & ~n14210;
  assign n14212 = pi0594 & pi1359;
  assign n14213 = pi0392 & pi1057;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = n14211 & n14214;
  assign n14216 = n9475 & ~n14215;
  assign n14217 = pi0069 & ~pi0979;
  assign n14218 = pi0068 & pi0979;
  assign n14219 = ~n14217 & ~n14218;
  assign n14220 = pi0720 & ~n14219;
  assign n14221 = pi0258 & ~pi0979;
  assign n14222 = pi0256 & pi0979;
  assign n14223 = ~n14221 & ~n14222;
  assign n14224 = pi0721 & ~n14223;
  assign n14225 = ~n14220 & ~n14224;
  assign n14226 = ~pi0979 & pi2642;
  assign n14227 = pi0979 & pi3176;
  assign n14228 = ~n14226 & ~n14227;
  assign n14229 = pi0765 & ~n14228;
  assign n14230 = ~pi0979 & pi2840;
  assign n14231 = pi0979 & pi3185;
  assign n14232 = ~n14230 & ~n14231;
  assign n14233 = pi0766 & ~n14232;
  assign n14234 = ~n14229 & ~n14233;
  assign n14235 = ~pi0979 & pi2617;
  assign n14236 = pi0979 & pi2610;
  assign n14237 = ~n14235 & ~n14236;
  assign n14238 = pi0763 & ~n14237;
  assign n14239 = ~pi0979 & pi2629;
  assign n14240 = pi0979 & pi2623;
  assign n14241 = ~n14239 & ~n14240;
  assign n14242 = pi0764 & ~n14241;
  assign n14243 = ~n14238 & ~n14242;
  assign n14244 = n14234 & n14243;
  assign n14245 = ~n9499 & n14244;
  assign n14246 = n14225 & n14245;
  assign n14247 = n9486 & ~n14246;
  assign n14248 = ~n14216 & ~n14247;
  assign n14249 = ~pi0979 & pi2855;
  assign n14250 = pi0979 & pi2138;
  assign n14251 = ~n14249 & ~n14250;
  assign n14252 = pi0717 & ~n14251;
  assign n14253 = pi0227 & ~pi0979;
  assign n14254 = pi0226 & pi0979;
  assign n14255 = ~n14253 & ~n14254;
  assign n14256 = pi0716 & ~n14255;
  assign n14257 = pi0284 & ~pi0979;
  assign n14258 = pi0282 & pi0979;
  assign n14259 = ~n14257 & ~n14258;
  assign n14260 = pi0761 & ~n14259;
  assign n14261 = ~n14256 & ~n14260;
  assign n14262 = ~n9535 & n14261;
  assign n14263 = ~n9531 & n14262;
  assign n14264 = ~n14252 & n14263;
  assign n14265 = n9523 & ~n14264;
  assign n14266 = pi0979 & pi2175;
  assign n14267 = ~pi0979 & pi2937;
  assign n14268 = ~n14266 & ~n14267;
  assign n14269 = pi0836 & ~n14268;
  assign n14270 = ~pi0979 & pi3113;
  assign n14271 = pi0979 & pi2191;
  assign n14272 = ~n14270 & ~n14271;
  assign n14273 = pi0837 & ~n14272;
  assign n14274 = ~n14269 & ~n14273;
  assign n14275 = ~pi0979 & pi2431;
  assign n14276 = pi0979 & pi1967;
  assign n14277 = ~n14275 & ~n14276;
  assign n14278 = pi0768 & ~n14277;
  assign n14279 = ~pi0979 & pi2928;
  assign n14280 = pi0979 & pi2157;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = pi0767 & ~n14281;
  assign n14283 = ~n14278 & ~n14282;
  assign n14284 = pi0181 & ~pi0979;
  assign n14285 = pi0166 & pi0979;
  assign n14286 = ~n14284 & ~n14285;
  assign n14287 = pi0838 & ~n14286;
  assign n14288 = n14283 & ~n14287;
  assign n14289 = n14274 & n14288;
  assign n14290 = n9549 & ~n14289;
  assign n14291 = ~n14265 & ~n14290;
  assign n14292 = pi1343 & pi2326;
  assign n14293 = pi1054 & pi2718;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = pi1055 & pi2726;
  assign n14296 = n14294 & ~n14295;
  assign n14297 = pi1342 & pi2312;
  assign n14298 = n14296 & ~n14297;
  assign n14299 = pi1340 & pi2290;
  assign n14300 = pi1341 & pi2301;
  assign n14301 = ~n14299 & ~n14300;
  assign n14302 = pi1355 & pi2460;
  assign n14303 = pi1356 & pi2756;
  assign n14304 = ~n14302 & ~n14303;
  assign n14305 = pi1357 & pi2469;
  assign n14306 = n14304 & ~n14305;
  assign n14307 = pi1354 & pi2750;
  assign n14308 = n14306 & ~n14307;
  assign n14309 = pi1349 & pi2737;
  assign n14310 = pi1056 & pi2745;
  assign n14311 = ~n14309 & ~n14310;
  assign n14312 = n14308 & n14311;
  assign n14313 = n14301 & n14312;
  assign n14314 = n14298 & n14313;
  assign n14315 = n9736 & ~n14314;
  assign n14316 = pi1339 & pi2255;
  assign n14317 = pi1345 & pi2659;
  assign n14318 = ~n14316 & ~n14317;
  assign n14319 = pi1346 & pi2673;
  assign n14320 = n14318 & ~n14319;
  assign n14321 = pi1338 & pi2241;
  assign n14322 = n14320 & ~n14321;
  assign n14323 = pi1600 & pi2213;
  assign n14324 = pi1337 & pi2227;
  assign n14325 = ~n14323 & ~n14324;
  assign n14326 = pi1351 & pi2441;
  assign n14327 = pi1352 & pi2751;
  assign n14328 = ~n14326 & ~n14327;
  assign n14329 = pi1353 & pi2278;
  assign n14330 = n14328 & ~n14329;
  assign n14331 = pi1350 & pi2700;
  assign n14332 = n14330 & ~n14331;
  assign n14333 = pi1347 & pi2686;
  assign n14334 = pi1348 & pi2697;
  assign n14335 = ~n14333 & ~n14334;
  assign n14336 = n14332 & n14335;
  assign n14337 = n14325 & n14336;
  assign n14338 = n14322 & n14337;
  assign n14339 = n9577 & ~n14338;
  assign n14340 = ~n14315 & ~n14339;
  assign n14341 = pi1333 & pi1745;
  assign n14342 = pi0225 & pi1336;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = pi1332 & pi2581;
  assign n14345 = pi1335 & pi2596;
  assign n14346 = ~n14344 & ~n14345;
  assign n14347 = n14343 & n14346;
  assign n14348 = n9726 & ~n14347;
  assign n14349 = pi1629 & n10557;
  assign n14350 = pi0794 & n9614;
  assign n14351 = pi2051 & n9618;
  assign n14352 = ~n14350 & ~n14351;
  assign n14353 = pi0740 & n9715;
  assign n14354 = pi1891 & n9718;
  assign n14355 = ~n14353 & ~n14354;
  assign n14356 = pi1737 & n11106;
  assign n14357 = pi0871 & n9707;
  assign n14358 = ~n14356 & ~n14357;
  assign n14359 = pi1702 & n10564;
  assign n14360 = n14358 & ~n14359;
  assign n14361 = n14355 & n14360;
  assign n14362 = pi1705 & n9698;
  assign n14363 = n14361 & ~n14362;
  assign n14364 = pi0978 & n9687;
  assign n14365 = pi1446 & n9691;
  assign n14366 = ~n14364 & ~n14365;
  assign n14367 = n14363 & n14366;
  assign n14368 = n14352 & n14367;
  assign n14369 = ~n14349 & n14368;
  assign n14370 = pi1785 & n9712;
  assign n14371 = n14369 & ~n14370;
  assign n14372 = pi1460 & n11145;
  assign n14373 = pi0910 & n9710;
  assign n14374 = ~n14372 & ~n14373;
  assign n14375 = pi0781 & n9670;
  assign n14376 = pi1090 & n9676;
  assign n14377 = ~n14375 & ~n14376;
  assign n14378 = pi0726 & n9654;
  assign n14379 = pi2501 & n11158;
  assign n14380 = ~n14378 & ~n14379;
  assign n14381 = pi3063 & n9647;
  assign n14382 = n14380 & ~n14381;
  assign n14383 = n14377 & n14382;
  assign n14384 = pi1932 & n9622;
  assign n14385 = n14383 & ~n14384;
  assign n14386 = pi1725 & n9679;
  assign n14387 = pi0367 & n9682;
  assign n14388 = ~n14386 & ~n14387;
  assign n14389 = n14385 & n14388;
  assign n14390 = n14374 & n14389;
  assign n14391 = n14371 & n14390;
  assign n14392 = pi1934 & ~n14391;
  assign n14393 = ~n14348 & ~n14392;
  assign n14394 = n14340 & n14393;
  assign n14395 = n14291 & n14394;
  assign n14396 = n14248 & n14395;
  assign n14397 = pi3315 & po3871;
  assign n14398 = n14396 & ~n14397;
  assign n14399 = ~pi1787 & ~n14398;
  assign n14400 = pi1787 & pi2835;
  assign n14401 = ~n14399 & ~n14400;
  assign n14402 = n9472 & ~n14401;
  assign n14403 = ~n14208 & ~n14402;
  assign n14404 = n10914 & ~n14403;
  assign n14405 = ~n11650 & n11654;
  assign n14406 = ~n11366 & ~n14405;
  assign n14407 = n11366 & n14405;
  assign n14408 = ~n14406 & ~n14407;
  assign n14409 = n11615 & ~n14408;
  assign n14410 = ~n11369 & n11383;
  assign n14411 = n11369 & ~n11383;
  assign n14412 = ~n14410 & ~n14411;
  assign n14413 = ~n11428 & ~n11607;
  assign n14414 = ~n11405 & n14413;
  assign n14415 = ~n14412 & n14414;
  assign n14416 = n14412 & ~n14414;
  assign n14417 = ~n14415 & ~n14416;
  assign n14418 = ~n11615 & ~n14417;
  assign n14419 = ~n14409 & ~n14418;
  assign n14420 = ~pi0518 & ~n14419;
  assign n14421 = n11665 & ~n14417;
  assign n14422 = ~n11665 & ~n14408;
  assign n14423 = ~n14421 & ~n14422;
  assign n14424 = pi0518 & ~n14423;
  assign n14425 = ~n14420 & ~n14424;
  assign n14426 = pi0683 & n11350;
  assign n14427 = pi0683 & ~n11260;
  assign n14428 = n11223 & n14427;
  assign n14429 = ~n14426 & ~n14428;
  assign n14430 = n14425 & n14429;
  assign n14431 = ~n10914 & ~n14430;
  assign n14432 = ~n14404 & ~n14431;
  assign n14433 = n11755 & ~n14432;
  assign n14434 = ~n10330 & n10334;
  assign n14435 = n10010 & n14434;
  assign n14436 = ~n10010 & ~n14434;
  assign n14437 = ~n14435 & ~n14436;
  assign n14438 = n10296 & ~n14437;
  assign n14439 = n10075 & ~n10287;
  assign n14440 = ~n10013 & n10029;
  assign n14441 = n10013 & ~n10029;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = ~n14439 & n14442;
  assign n14444 = n14439 & ~n14442;
  assign n14445 = ~n14443 & ~n14444;
  assign n14446 = ~n10296 & ~n14445;
  assign n14447 = ~n14438 & ~n14446;
  assign n14448 = ~pi0568 & ~n14447;
  assign n14449 = n10362 & ~n14445;
  assign n14450 = ~n10362 & ~n14437;
  assign n14451 = ~n14449 & ~n14450;
  assign n14452 = pi0568 & ~n14451;
  assign n14453 = ~n14448 & ~n14452;
  assign n14454 = pi0757 & n9998;
  assign n14455 = pi0757 & ~n9951;
  assign n14456 = n9917 & n14455;
  assign n14457 = ~n14454 & ~n14456;
  assign n14458 = n14453 & n14457;
  assign n14459 = n10914 & ~n14458;
  assign n14460 = ~pi0781 & n11700;
  assign n14461 = pi1038 & ~n11706;
  assign n14462 = pi0910 & n11709;
  assign n14463 = pi2707 & po3871;
  assign n14464 = ~n14462 & ~n14463;
  assign n14465 = pi0423 & n11714;
  assign n14466 = n14464 & ~n14465;
  assign n14467 = ~n14461 & n14466;
  assign n14468 = ~n11700 & n14467;
  assign n14469 = pi2756 & n11190;
  assign n14470 = pi2469 & n11192;
  assign n14471 = ~n14469 & ~n14470;
  assign n14472 = pi2460 & n11195;
  assign n14473 = pi2750 & n11197;
  assign n14474 = ~n14472 & ~n14473;
  assign n14475 = n14471 & n14474;
  assign n14476 = n9424 & ~n14475;
  assign n14477 = pi2750 & n11207;
  assign n14478 = pi2756 & n11204;
  assign n14479 = ~n14477 & ~n14478;
  assign n14480 = pi2469 & n11202;
  assign n14481 = pi2460 & n11209;
  assign n14482 = ~n14480 & ~n14481;
  assign n14483 = n14479 & n14482;
  assign n14484 = ~n9424 & ~n14483;
  assign n14485 = ~n14476 & ~n14484;
  assign n14486 = n10886 & ~n14485;
  assign n14487 = n14468 & ~n14486;
  assign n14488 = pi2700 & n9837;
  assign n14489 = pi2751 & n9834;
  assign n14490 = ~n14488 & ~n14489;
  assign n14491 = pi2441 & n9839;
  assign n14492 = pi2278 & n9832;
  assign n14493 = ~n14491 & ~n14492;
  assign n14494 = n14490 & n14493;
  assign n14495 = ~n9424 & ~n14494;
  assign n14496 = pi2441 & n10376;
  assign n14497 = pi2751 & n10381;
  assign n14498 = ~n14496 & ~n14497;
  assign n14499 = pi2700 & n10374;
  assign n14500 = pi2278 & n10379;
  assign n14501 = ~n14499 & ~n14500;
  assign n14502 = n14498 & n14501;
  assign n14503 = n9424 & ~n14502;
  assign n14504 = ~n14495 & ~n14503;
  assign n14505 = n11701 & ~n14504;
  assign n14506 = n14487 & ~n14505;
  assign n14507 = ~n14460 & ~n14506;
  assign n14508 = n11186 & n14507;
  assign n14509 = ~n14459 & ~n14508;
  assign n14510 = ~n10902 & ~n14509;
  assign n14511 = ~n11468 & ~n11633;
  assign n14512 = ~n11469 & ~n14511;
  assign n14513 = n11486 & ~n14512;
  assign n14514 = ~n11486 & n14512;
  assign n14515 = ~n14513 & ~n14514;
  assign n14516 = n11615 & ~n14515;
  assign n14517 = ~n11514 & ~n11517;
  assign n14518 = ~n11474 & ~n14517;
  assign n14519 = n11489 & ~n11491;
  assign n14520 = ~n11489 & n11491;
  assign n14521 = ~n14519 & ~n14520;
  assign n14522 = n14518 & n14521;
  assign n14523 = ~n14518 & ~n14521;
  assign n14524 = ~n14522 & ~n14523;
  assign n14525 = ~n11615 & ~n14524;
  assign n14526 = ~n14516 & ~n14525;
  assign n14527 = ~pi0518 & ~n14526;
  assign n14528 = n11665 & ~n14524;
  assign n14529 = ~n11665 & ~n14515;
  assign n14530 = ~n14528 & ~n14529;
  assign n14531 = pi0518 & ~n14530;
  assign n14532 = ~n14527 & ~n14531;
  assign n14533 = pi0705 & n11260;
  assign n14534 = ~n11264 & n14533;
  assign n14535 = pi0705 & n11481;
  assign n14536 = ~n14534 & ~n14535;
  assign n14537 = ~n14532 & n14536;
  assign n14538 = n10914 & n14537;
  assign n14539 = pi2456 & n11195;
  assign n14540 = pi2465 & n11192;
  assign n14541 = ~n14539 & ~n14540;
  assign n14542 = pi2810 & n11190;
  assign n14543 = pi2780 & n11197;
  assign n14544 = ~n14542 & ~n14543;
  assign n14545 = n14541 & n14544;
  assign n14546 = n9424 & ~n14545;
  assign n14547 = pi2780 & n11207;
  assign n14548 = pi2810 & n11204;
  assign n14549 = ~n14547 & ~n14548;
  assign n14550 = pi2465 & n11202;
  assign n14551 = pi2456 & n11209;
  assign n14552 = ~n14550 & ~n14551;
  assign n14553 = n14549 & n14552;
  assign n14554 = ~n9424 & ~n14553;
  assign n14555 = ~n14546 & ~n14554;
  assign n14556 = ~n10914 & n14555;
  assign n14557 = ~n14538 & ~n14556;
  assign n14558 = n11697 & n14557;
  assign n14559 = ~n14510 & ~n14558;
  assign n14560 = ~n10885 & ~n14559;
  assign n14561 = n14485 & n14504;
  assign n14562 = n11785 & ~n14561;
  assign n14563 = pi3862 & n9804;
  assign n14564 = pi3878 & n9774;
  assign n14565 = ~n14563 & ~n14564;
  assign n14566 = pi3846 & n9802;
  assign n14567 = pi3910 & n9781;
  assign n14568 = pi3894 & n9771;
  assign n14569 = ~n14567 & ~n14568;
  assign n14570 = pi3942 & n9791;
  assign n14571 = pi3926 & n9788;
  assign n14572 = ~n14570 & ~n14571;
  assign n14573 = n14569 & n14572;
  assign n14574 = ~n14566 & n14573;
  assign n14575 = n14565 & n14574;
  assign n14576 = pi3862 & n9799;
  assign n14577 = n14575 & ~n14576;
  assign n14578 = pi3974 & n9783;
  assign n14579 = pi3958 & n9793;
  assign n14580 = ~n14578 & ~n14579;
  assign n14581 = n14577 & n14580;
  assign n14582 = ~n9472 & ~n14581;
  assign n14583 = pi1334 & pi3204;
  assign n14584 = pi0828 & pi1344;
  assign n14585 = ~n14583 & ~n14584;
  assign n14586 = pi0708 & pi1358;
  assign n14587 = n14585 & ~n14586;
  assign n14588 = pi1053 & pi2472;
  assign n14589 = n14587 & ~n14588;
  assign n14590 = pi1059 & pi2978;
  assign n14591 = pi0388 & pi1057;
  assign n14592 = ~n14590 & ~n14591;
  assign n14593 = pi1331 & ~n8839;
  assign n14594 = pi1058 & pi3407;
  assign n14595 = ~n14593 & ~n14594;
  assign n14596 = pi0603 & pi1359;
  assign n14597 = n14595 & ~n14596;
  assign n14598 = n14592 & n14597;
  assign n14599 = n14589 & n14598;
  assign n14600 = pi3521 & ~n10410;
  assign n14601 = n14599 & ~n14600;
  assign n14602 = n9475 & ~n14601;
  assign n14603 = pi0306 & ~pi0979;
  assign n14604 = pi0304 & pi0979;
  assign n14605 = ~n14603 & ~n14604;
  assign n14606 = pi0716 & ~n14605;
  assign n14607 = pi0324 & ~pi0979;
  assign n14608 = pi0323 & pi0979;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = pi0761 & ~n14609;
  assign n14611 = ~n14606 & ~n14610;
  assign n14612 = pi0979 & pi2130;
  assign n14613 = ~pi0979 & pi2847;
  assign n14614 = ~n14612 & ~n14613;
  assign n14615 = pi0717 & ~n14614;
  assign n14616 = pi0204 & ~pi0979;
  assign n14617 = pi0200 & pi0979;
  assign n14618 = ~n14616 & ~n14617;
  assign n14619 = pi1599 & ~n14618;
  assign n14620 = ~n14615 & ~n14619;
  assign n14621 = pi0481 & ~pi0979;
  assign n14622 = pi0480 & pi0979;
  assign n14623 = ~n14621 & ~n14622;
  assign n14624 = pi0718 & ~n14623;
  assign n14625 = n14620 & ~n14624;
  assign n14626 = n14611 & n14625;
  assign n14627 = n9523 & ~n14626;
  assign n14628 = ~n14602 & ~n14627;
  assign n14629 = pi0979 & pi2167;
  assign n14630 = ~pi0979 & pi2793;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = pi0836 & ~n14631;
  assign n14633 = ~pi0979 & pi2944;
  assign n14634 = pi0979 & pi2183;
  assign n14635 = ~n14633 & ~n14634;
  assign n14636 = pi0837 & ~n14635;
  assign n14637 = ~n14632 & ~n14636;
  assign n14638 = pi0979 & pi2149;
  assign n14639 = ~pi0979 & pi2921;
  assign n14640 = ~n14638 & ~n14639;
  assign n14641 = pi0767 & ~n14640;
  assign n14642 = ~pi0979 & pi2426;
  assign n14643 = pi0979 & pi1961;
  assign n14644 = ~n14642 & ~n14643;
  assign n14645 = pi0768 & ~n14644;
  assign n14646 = ~n14641 & ~n14645;
  assign n14647 = pi0173 & ~pi0979;
  assign n14648 = pi0159 & pi0979;
  assign n14649 = ~n14647 & ~n14648;
  assign n14650 = pi0838 & ~n14649;
  assign n14651 = pi0196 & pi1360;
  assign n14652 = ~n14650 & ~n14651;
  assign n14653 = n14646 & n14652;
  assign n14654 = n14637 & n14653;
  assign n14655 = n9549 & ~n14654;
  assign n14656 = ~pi0979 & pi2865;
  assign n14657 = pi0979 & pi3155;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = pi0763 & ~n14658;
  assign n14660 = ~pi0979 & pi2874;
  assign n14661 = pi0979 & pi3163;
  assign n14662 = ~n14660 & ~n14661;
  assign n14663 = pi0764 & ~n14662;
  assign n14664 = ~n14659 & ~n14663;
  assign n14665 = ~pi0979 & pi2541;
  assign n14666 = pi0979 & pi3131;
  assign n14667 = ~n14665 & ~n14666;
  assign n14668 = pi0765 & ~n14667;
  assign n14669 = ~pi0979 & pi2891;
  assign n14670 = pi0979 & pi3181;
  assign n14671 = ~n14669 & ~n14670;
  assign n14672 = pi0766 & ~n14671;
  assign n14673 = ~n14668 & ~n14672;
  assign n14674 = pi0218 & ~pi0979;
  assign n14675 = pi0215 & pi0979;
  assign n14676 = ~n14674 & ~n14675;
  assign n14677 = pi0720 & ~n14676;
  assign n14678 = pi0397 & ~pi0979;
  assign n14679 = pi0396 & pi0979;
  assign n14680 = ~n14678 & ~n14679;
  assign n14681 = pi0721 & ~n14680;
  assign n14682 = ~n14677 & ~n14681;
  assign n14683 = pi0041 & ~pi0979;
  assign n14684 = pi0039 & pi0979;
  assign n14685 = ~n14683 & ~n14684;
  assign n14686 = pi0719 & ~n14685;
  assign n14687 = n14682 & ~n14686;
  assign n14688 = n14673 & n14687;
  assign n14689 = n14664 & n14688;
  assign n14690 = n9486 & ~n14689;
  assign n14691 = ~n14655 & ~n14690;
  assign n14692 = pi1355 & pi2456;
  assign n14693 = pi1356 & pi2810;
  assign n14694 = ~n14692 & ~n14693;
  assign n14695 = pi1357 & pi2465;
  assign n14696 = n14694 & ~n14695;
  assign n14697 = pi1354 & pi2780;
  assign n14698 = n14696 & ~n14697;
  assign n14699 = pi1349 & pi2733;
  assign n14700 = pi1056 & pi2742;
  assign n14701 = ~n14699 & ~n14700;
  assign n14702 = pi1343 & pi2320;
  assign n14703 = pi1054 & pi2713;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = pi1055 & pi2723;
  assign n14706 = n14704 & ~n14705;
  assign n14707 = pi1342 & pi2306;
  assign n14708 = n14706 & ~n14707;
  assign n14709 = pi1340 & pi2285;
  assign n14710 = pi1341 & pi2297;
  assign n14711 = ~n14709 & ~n14710;
  assign n14712 = n14708 & n14711;
  assign n14713 = n14701 & n14712;
  assign n14714 = n14698 & n14713;
  assign n14715 = n9736 & ~n14714;
  assign n14716 = pi1347 & pi2681;
  assign n14717 = pi1348 & pi2691;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = pi1350 & pi2260;
  assign n14720 = n14718 & ~n14719;
  assign n14721 = pi1346 & pi2667;
  assign n14722 = n14720 & ~n14721;
  assign n14723 = pi1339 & pi2249;
  assign n14724 = pi1345 & pi2653;
  assign n14725 = ~n14723 & ~n14724;
  assign n14726 = pi1600 & pi2207;
  assign n14727 = pi1337 & pi2221;
  assign n14728 = ~n14726 & ~n14727;
  assign n14729 = pi1338 & pi2235;
  assign n14730 = n14728 & ~n14729;
  assign n14731 = pi1353 & pi1980;
  assign n14732 = n14730 & ~n14731;
  assign n14733 = pi1351 & pi2265;
  assign n14734 = pi1352 & pi2443;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = n14732 & n14735;
  assign n14737 = n14725 & n14736;
  assign n14738 = n14722 & n14737;
  assign n14739 = n9577 & ~n14738;
  assign n14740 = ~n14715 & ~n14739;
  assign n14741 = pi0331 & pi1336;
  assign n14742 = pi0072 & pi1333;
  assign n14743 = ~n14741 & ~n14742;
  assign n14744 = pi1332 & pi2573;
  assign n14745 = pi1335 & pi2588;
  assign n14746 = ~n14744 & ~n14745;
  assign n14747 = n14743 & n14746;
  assign n14748 = n9726 & ~n14747;
  assign n14749 = pi0884 & n9715;
  assign n14750 = pi1887 & n9718;
  assign n14751 = ~n14749 & ~n14750;
  assign n14752 = pi1733 & n11106;
  assign n14753 = pi0746 & n9707;
  assign n14754 = ~n14752 & ~n14753;
  assign n14755 = pi0891 & n9702;
  assign n14756 = n14754 & ~n14755;
  assign n14757 = n14751 & n14756;
  assign n14758 = pi1852 & n9698;
  assign n14759 = n14757 & ~n14758;
  assign n14760 = pi0957 & n9614;
  assign n14761 = pi1901 & n9618;
  assign n14762 = ~n14760 & ~n14761;
  assign n14763 = pi0797 & n9607;
  assign n14764 = n14762 & ~n14763;
  assign n14765 = pi0803 & n9687;
  assign n14766 = pi1442 & n9691;
  assign n14767 = ~n14765 & ~n14766;
  assign n14768 = n14764 & n14767;
  assign n14769 = pi0772 & n9654;
  assign n14770 = pi2498 & n11158;
  assign n14771 = ~n14769 & ~n14770;
  assign n14772 = pi0776 & n9670;
  assign n14773 = pi1841 & n9676;
  assign n14774 = ~n14772 & ~n14773;
  assign n14775 = pi3100 & n9647;
  assign n14776 = n14774 & ~n14775;
  assign n14777 = n14771 & n14776;
  assign n14778 = pi1942 & n11165;
  assign n14779 = n14777 & ~n14778;
  assign n14780 = pi2107 & n9628;
  assign n14781 = pi1022 & n9631;
  assign n14782 = ~n14780 & ~n14781;
  assign n14783 = pi1858 & n9657;
  assign n14784 = pi1755 & n9659;
  assign n14785 = ~n14783 & ~n14784;
  assign n14786 = n14782 & n14785;
  assign n14787 = pi1431 & n11133;
  assign n14788 = pi0822 & n9682;
  assign n14789 = ~n14787 & ~n14788;
  assign n14790 = pi1719 & n9679;
  assign n14791 = n14789 & ~n14790;
  assign n14792 = pi1925 & n9622;
  assign n14793 = n14791 & ~n14792;
  assign n14794 = n14786 & n14793;
  assign n14795 = ~n11102 & n14794;
  assign n14796 = n14779 & n14795;
  assign n14797 = pi1778 & n9712;
  assign n14798 = n14796 & ~n14797;
  assign n14799 = pi1456 & n11145;
  assign n14800 = pi0874 & n9710;
  assign n14801 = ~n14799 & ~n14800;
  assign n14802 = n14798 & n14801;
  assign n14803 = n14768 & n14802;
  assign n14804 = n14759 & n14803;
  assign n14805 = pi1934 & ~n14804;
  assign n14806 = ~n14748 & ~n14805;
  assign n14807 = n14740 & n14806;
  assign n14808 = n14691 & n14807;
  assign n14809 = n14628 & n14808;
  assign n14810 = pi3311 & po3871;
  assign n14811 = n14809 & ~n14810;
  assign n14812 = ~pi1787 & ~n14811;
  assign n14813 = pi1787 & pi2829;
  assign n14814 = ~n14812 & ~n14813;
  assign n14815 = n9472 & ~n14814;
  assign n14816 = ~n14582 & ~n14815;
  assign n14817 = ~n10914 & ~n14816;
  assign n14818 = ~n11697 & n14817;
  assign n14819 = ~n14562 & ~n14818;
  assign n14820 = n10885 & ~n14819;
  assign n14821 = ~n14560 & ~n14820;
  assign po0226 = n14433 | ~n14821;
  assign n14823 = po0224 & po0226;
  assign n14824 = po0221 & n14823;
  assign n14825 = n13483 & n14824;
  assign n14826 = pi2544 & n11190;
  assign n14827 = pi2468 & n11192;
  assign n14828 = ~n14826 & ~n14827;
  assign n14829 = pi2459 & n11195;
  assign n14830 = pi2749 & n11197;
  assign n14831 = ~n14829 & ~n14830;
  assign n14832 = n14828 & n14831;
  assign n14833 = n9424 & ~n14832;
  assign n14834 = pi2749 & n11207;
  assign n14835 = pi2544 & n11204;
  assign n14836 = ~n14834 & ~n14835;
  assign n14837 = pi2468 & n11202;
  assign n14838 = pi2459 & n11209;
  assign n14839 = ~n14837 & ~n14838;
  assign n14840 = n14836 & n14839;
  assign n14841 = ~n9424 & ~n14840;
  assign n14842 = ~n14833 & ~n14841;
  assign n14843 = pi2539 & n9837;
  assign n14844 = pi2440 & n9839;
  assign n14845 = ~n14843 & ~n14844;
  assign n14846 = pi2277 & n9832;
  assign n14847 = pi2703 & n9834;
  assign n14848 = ~n14846 & ~n14847;
  assign n14849 = n14845 & n14848;
  assign n14850 = ~n9424 & ~n14849;
  assign n14851 = pi2539 & n10374;
  assign n14852 = pi2440 & n10376;
  assign n14853 = ~n14851 & ~n14852;
  assign n14854 = pi2277 & n10379;
  assign n14855 = pi2703 & n10381;
  assign n14856 = ~n14854 & ~n14855;
  assign n14857 = n14853 & n14856;
  assign n14858 = n9424 & ~n14857;
  assign n14859 = ~n14850 & ~n14858;
  assign n14860 = n14842 & n14859;
  assign n14861 = n11785 & ~n14860;
  assign n14862 = pi0979 & pi2168;
  assign n14863 = ~pi0979 & pi2934;
  assign n14864 = ~n14862 & ~n14863;
  assign n14865 = pi0836 & ~n14864;
  assign n14866 = ~pi0979 & pi2945;
  assign n14867 = pi0979 & pi2184;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = pi0837 & ~n14868;
  assign n14870 = ~n14865 & ~n14869;
  assign n14871 = pi0979 & pi2150;
  assign n14872 = ~pi0979 & pi2922;
  assign n14873 = ~n14871 & ~n14872;
  assign n14874 = pi0767 & ~n14873;
  assign n14875 = ~pi0979 & pi2427;
  assign n14876 = pi0979 & pi1962;
  assign n14877 = ~n14875 & ~n14876;
  assign n14878 = pi0768 & ~n14877;
  assign n14879 = ~n14874 & ~n14878;
  assign n14880 = pi0175 & ~pi0979;
  assign n14881 = pi0160 & pi0979;
  assign n14882 = ~n14880 & ~n14881;
  assign n14883 = pi0838 & ~n14882;
  assign n14884 = pi0152 & pi1360;
  assign n14885 = ~n14883 & ~n14884;
  assign n14886 = n14879 & n14885;
  assign n14887 = n14870 & n14886;
  assign n14888 = n9549 & ~n14887;
  assign n14889 = pi0042 & ~pi0979;
  assign n14890 = pi0040 & pi0979;
  assign n14891 = ~n14889 & ~n14890;
  assign n14892 = pi0719 & ~n14891;
  assign n14893 = ~pi0979 & pi2636;
  assign n14894 = pi0979 & pi3170;
  assign n14895 = ~n14893 & ~n14894;
  assign n14896 = pi0765 & ~n14895;
  assign n14897 = ~pi0979 & pi2892;
  assign n14898 = pi0979 & pi3122;
  assign n14899 = ~n14897 & ~n14898;
  assign n14900 = pi0766 & ~n14899;
  assign n14901 = ~n14896 & ~n14900;
  assign n14902 = ~pi0979 & pi2866;
  assign n14903 = pi0979 & pi3156;
  assign n14904 = ~n14902 & ~n14903;
  assign n14905 = pi0763 & ~n14904;
  assign n14906 = ~pi0979 & pi2875;
  assign n14907 = pi0979 & pi3164;
  assign n14908 = ~n14906 & ~n14907;
  assign n14909 = pi0764 & ~n14908;
  assign n14910 = ~n14905 & ~n14909;
  assign n14911 = pi0217 & ~pi0979;
  assign n14912 = pi0216 & pi0979;
  assign n14913 = ~n14911 & ~n14912;
  assign n14914 = pi0720 & ~n14913;
  assign n14915 = pi0490 & ~pi0979;
  assign n14916 = pi0489 & pi0979;
  assign n14917 = ~n14915 & ~n14916;
  assign n14918 = pi0721 & ~n14917;
  assign n14919 = ~n14914 & ~n14918;
  assign n14920 = n14910 & n14919;
  assign n14921 = n14901 & n14920;
  assign n14922 = ~n14892 & n14921;
  assign n14923 = n9486 & ~n14922;
  assign n14924 = ~n14888 & ~n14923;
  assign n14925 = pi0350 & pi1336;
  assign n14926 = pi0127 & pi1333;
  assign n14927 = ~n14925 & ~n14926;
  assign n14928 = pi1332 & pi2574;
  assign n14929 = pi1335 & pi2589;
  assign n14930 = ~n14928 & ~n14929;
  assign n14931 = n14927 & n14930;
  assign n14932 = n9726 & ~n14931;
  assign n14933 = pi0885 & n9715;
  assign n14934 = pi1888 & n9718;
  assign n14935 = ~n14933 & ~n14934;
  assign n14936 = pi1734 & n11106;
  assign n14937 = pi0737 & n9707;
  assign n14938 = ~n14936 & ~n14937;
  assign n14939 = pi0892 & n9702;
  assign n14940 = n14938 & ~n14939;
  assign n14941 = n14935 & n14940;
  assign n14942 = pi1834 & n9698;
  assign n14943 = n14941 & ~n14942;
  assign n14944 = pi1009 & n9614;
  assign n14945 = pi1902 & n9618;
  assign n14946 = ~n14944 & ~n14945;
  assign n14947 = pi0798 & n9607;
  assign n14948 = n14946 & ~n14947;
  assign n14949 = pi0846 & n9687;
  assign n14950 = pi1443 & n9691;
  assign n14951 = ~n14949 & ~n14950;
  assign n14952 = n14948 & n14951;
  assign n14953 = pi0786 & n9654;
  assign n14954 = pi2512 & n11158;
  assign n14955 = ~n14953 & ~n14954;
  assign n14956 = pi0777 & n9670;
  assign n14957 = pi2058 & n9676;
  assign n14958 = ~n14956 & ~n14957;
  assign n14959 = pi3099 & n9647;
  assign n14960 = n14958 & ~n14959;
  assign n14961 = n14955 & n14960;
  assign n14962 = pi1943 & n11165;
  assign n14963 = n14961 & ~n14962;
  assign n14964 = pi2141 & n9628;
  assign n14965 = pi1101 & n9631;
  assign n14966 = ~n14964 & ~n14965;
  assign n14967 = pi1766 & n9657;
  assign n14968 = pi1756 & n9659;
  assign n14969 = ~n14967 & ~n14968;
  assign n14970 = n14966 & n14969;
  assign n14971 = pi1432 & n11133;
  assign n14972 = pi0728 & n9682;
  assign n14973 = ~n14971 & ~n14972;
  assign n14974 = pi1720 & n9679;
  assign n14975 = n14973 & ~n14974;
  assign n14976 = pi1926 & n9622;
  assign n14977 = n14975 & ~n14976;
  assign n14978 = n14970 & n14977;
  assign n14979 = ~n11102 & n14978;
  assign n14980 = n14963 & n14979;
  assign n14981 = pi1779 & n9712;
  assign n14982 = n14980 & ~n14981;
  assign n14983 = pi1457 & n11145;
  assign n14984 = pi0907 & n9710;
  assign n14985 = ~n14983 & ~n14984;
  assign n14986 = n14982 & n14985;
  assign n14987 = n14952 & n14986;
  assign n14988 = n14943 & n14987;
  assign n14989 = pi1934 & ~n14988;
  assign n14990 = ~n14932 & ~n14989;
  assign n14991 = pi0316 & ~pi0979;
  assign n14992 = pi0315 & pi0979;
  assign n14993 = ~n14991 & ~n14992;
  assign n14994 = pi0716 & ~n14993;
  assign n14995 = pi0300 & ~pi0979;
  assign n14996 = pi0299 & pi0979;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = pi0761 & ~n14997;
  assign n14999 = ~n14994 & ~n14998;
  assign n15000 = pi0979 & pi2131;
  assign n15001 = ~pi0979 & pi2848;
  assign n15002 = ~n15000 & ~n15001;
  assign n15003 = pi0717 & ~n15002;
  assign n15004 = pi0207 & ~pi0979;
  assign n15005 = pi0201 & pi0979;
  assign n15006 = ~n15004 & ~n15005;
  assign n15007 = pi1599 & ~n15006;
  assign n15008 = ~n15003 & ~n15007;
  assign n15009 = pi0400 & ~pi0979;
  assign n15010 = pi0399 & pi0979;
  assign n15011 = ~n15009 & ~n15010;
  assign n15012 = pi0718 & ~n15011;
  assign n15013 = n15008 & ~n15012;
  assign n15014 = n14999 & n15013;
  assign n15015 = n9523 & ~n15014;
  assign n15016 = n14990 & ~n15015;
  assign n15017 = n14924 & n15016;
  assign n15018 = pi0685 & pi1334;
  assign n15019 = pi0829 & pi1344;
  assign n15020 = ~n15018 & ~n15019;
  assign n15021 = pi1331 & ~n9065;
  assign n15022 = pi1058 & pi3328;
  assign n15023 = ~n15021 & ~n15022;
  assign n15024 = pi0592 & pi1359;
  assign n15025 = n15023 & ~n15024;
  assign n15026 = pi3510 & ~n10410;
  assign n15027 = n15025 & ~n15026;
  assign n15028 = pi1059 & pi2979;
  assign n15029 = pi0389 & pi1057;
  assign n15030 = ~n15028 & ~n15029;
  assign n15031 = pi1053 & pi2514;
  assign n15032 = n15030 & ~n15031;
  assign n15033 = pi0918 & pi1358;
  assign n15034 = n15032 & ~n15033;
  assign n15035 = n15027 & n15034;
  assign n15036 = n15020 & n15035;
  assign n15037 = n9475 & ~n15036;
  assign n15038 = n15017 & ~n15037;
  assign n15039 = pi1349 & pi2560;
  assign n15040 = pi1056 & pi2547;
  assign n15041 = ~n15039 & ~n15040;
  assign n15042 = pi1354 & pi2776;
  assign n15043 = n15041 & ~n15042;
  assign n15044 = pi1357 & pi2411;
  assign n15045 = n15043 & ~n15044;
  assign n15046 = pi1355 & pi2526;
  assign n15047 = pi1356 & pi2967;
  assign n15048 = ~n15046 & ~n15047;
  assign n15049 = pi1343 & pi2321;
  assign n15050 = pi1054 & pi2714;
  assign n15051 = ~n15049 & ~n15050;
  assign n15052 = pi1055 & pi2724;
  assign n15053 = n15051 & ~n15052;
  assign n15054 = pi1342 & pi2307;
  assign n15055 = n15053 & ~n15054;
  assign n15056 = pi1340 & pi2286;
  assign n15057 = pi1341 & pi2298;
  assign n15058 = ~n15056 & ~n15057;
  assign n15059 = n15055 & n15058;
  assign n15060 = n15048 & n15059;
  assign n15061 = n15045 & n15060;
  assign n15062 = n9736 & ~n15061;
  assign n15063 = pi1339 & pi2250;
  assign n15064 = pi1345 & pi2654;
  assign n15065 = ~n15063 & ~n15064;
  assign n15066 = pi1346 & pi2668;
  assign n15067 = n15065 & ~n15066;
  assign n15068 = pi1338 & pi2236;
  assign n15069 = n15067 & ~n15068;
  assign n15070 = pi1600 & pi2208;
  assign n15071 = pi1337 & pi2222;
  assign n15072 = ~n15070 & ~n15071;
  assign n15073 = pi1351 & pi2266;
  assign n15074 = pi1352 & pi2274;
  assign n15075 = ~n15073 & ~n15074;
  assign n15076 = pi1353 & pi1981;
  assign n15077 = n15075 & ~n15076;
  assign n15078 = pi1350 & pi2433;
  assign n15079 = n15077 & ~n15078;
  assign n15080 = pi1347 & pi2682;
  assign n15081 = pi1348 & pi2692;
  assign n15082 = ~n15080 & ~n15081;
  assign n15083 = n15079 & n15082;
  assign n15084 = n15072 & n15083;
  assign n15085 = n15069 & n15084;
  assign n15086 = n9577 & ~n15085;
  assign n15087 = ~n15062 & ~n15086;
  assign n15088 = n15038 & n15087;
  assign n15089 = pi3297 & po3871;
  assign n15090 = n15088 & ~n15089;
  assign n15091 = ~pi1787 & ~n15090;
  assign n15092 = pi1787 & pi2830;
  assign n15093 = ~n15091 & ~n15092;
  assign n15094 = n9472 & ~n15093;
  assign n15095 = pi3861 & n9804;
  assign n15096 = pi3877 & n9774;
  assign n15097 = ~n15095 & ~n15096;
  assign n15098 = pi3845 & n9802;
  assign n15099 = pi3893 & n9771;
  assign n15100 = pi3957 & n9793;
  assign n15101 = ~n15099 & ~n15100;
  assign n15102 = pi3941 & n9791;
  assign n15103 = pi3925 & n9788;
  assign n15104 = ~n15102 & ~n15103;
  assign n15105 = n15101 & n15104;
  assign n15106 = ~n15098 & n15105;
  assign n15107 = n15097 & n15106;
  assign n15108 = pi3861 & n9799;
  assign n15109 = n15107 & ~n15108;
  assign n15110 = pi3909 & n9781;
  assign n15111 = pi3973 & n9783;
  assign n15112 = ~n15110 & ~n15111;
  assign n15113 = n15109 & n15112;
  assign n15114 = ~n9472 & ~n15113;
  assign n15115 = ~n15094 & ~n15114;
  assign n15116 = n11186 & ~n15115;
  assign n15117 = ~n10902 & n15116;
  assign n15118 = ~n14861 & ~n15117;
  assign n15119 = n10885 & ~n15118;
  assign n15120 = ~n10076 & ~n14439;
  assign n15121 = ~n10030 & ~n15120;
  assign n15122 = n9989 & ~n10008;
  assign n15123 = ~n9989 & n10008;
  assign n15124 = ~n15122 & ~n15123;
  assign n15125 = n15121 & n15124;
  assign n15126 = ~n15121 & ~n15124;
  assign n15127 = ~n15125 & ~n15126;
  assign n15128 = n10362 & ~n15127;
  assign n15129 = ~n10003 & ~n14434;
  assign n15130 = ~n10002 & ~n15129;
  assign n15131 = n9983 & ~n15130;
  assign n15132 = ~n9983 & n15130;
  assign n15133 = ~n15131 & ~n15132;
  assign n15134 = ~n10362 & ~n15133;
  assign n15135 = ~n15128 & ~n15134;
  assign n15136 = pi0568 & ~n15135;
  assign n15137 = n10296 & ~n15133;
  assign n15138 = ~n10296 & ~n15127;
  assign n15139 = ~n15137 & ~n15138;
  assign n15140 = ~pi0568 & ~n15139;
  assign n15141 = ~n15136 & ~n15140;
  assign n15142 = pi0756 & n9977;
  assign n15143 = pi0756 & ~n9951;
  assign n15144 = n9916 & n15143;
  assign n15145 = ~n15142 & ~n15144;
  assign n15146 = ~n15141 & n15145;
  assign n15147 = n10914 & ~n15146;
  assign n15148 = ~pi0780 & n11700;
  assign n15149 = n10886 & ~n14842;
  assign n15150 = pi2706 & po3871;
  assign n15151 = pi0820 & n11709;
  assign n15152 = pi1037 & ~n11706;
  assign n15153 = pi0422 & n11714;
  assign n15154 = ~n15152 & ~n15153;
  assign n15155 = ~n15151 & n15154;
  assign n15156 = ~n15150 & n15155;
  assign n15157 = ~n11700 & n15156;
  assign n15158 = n11701 & ~n14859;
  assign n15159 = n15157 & ~n15158;
  assign n15160 = ~n15149 & n15159;
  assign n15161 = ~n15148 & ~n15160;
  assign n15162 = ~n10914 & n15161;
  assign n15163 = ~n15147 & ~n15162;
  assign n15164 = ~n10902 & ~n15163;
  assign n15165 = ~n11470 & ~n11633;
  assign n15166 = n11470 & n11633;
  assign n15167 = ~n15165 & ~n15166;
  assign n15168 = n11615 & ~n15167;
  assign n15169 = ~n11457 & n11473;
  assign n15170 = n11457 & ~n11473;
  assign n15171 = ~n15169 & ~n15170;
  assign n15172 = ~n11514 & n15171;
  assign n15173 = n11514 & ~n15171;
  assign n15174 = ~n15172 & ~n15173;
  assign n15175 = ~n11615 & ~n15174;
  assign n15176 = ~n15168 & ~n15175;
  assign n15177 = ~pi0518 & ~n15176;
  assign n15178 = n11665 & ~n15174;
  assign n15179 = ~n11665 & ~n15167;
  assign n15180 = ~n15178 & ~n15179;
  assign n15181 = pi0518 & ~n15180;
  assign n15182 = ~n15177 & ~n15181;
  assign n15183 = pi0706 & n11260;
  assign n15184 = ~n11461 & n15183;
  assign n15185 = pi0706 & n11465;
  assign n15186 = ~n15184 & ~n15185;
  assign n15187 = n15182 & n15186;
  assign n15188 = ~n11186 & n15187;
  assign n15189 = pi2967 & n11190;
  assign n15190 = pi2411 & n11192;
  assign n15191 = ~n15189 & ~n15190;
  assign n15192 = pi2526 & n11195;
  assign n15193 = pi2776 & n11197;
  assign n15194 = ~n15192 & ~n15193;
  assign n15195 = n15191 & n15194;
  assign n15196 = n9424 & ~n15195;
  assign n15197 = pi2776 & n11207;
  assign n15198 = pi2967 & n11204;
  assign n15199 = ~n15197 & ~n15198;
  assign n15200 = pi2411 & n11202;
  assign n15201 = pi2526 & n11209;
  assign n15202 = ~n15200 & ~n15201;
  assign n15203 = n15199 & n15202;
  assign n15204 = ~n9424 & ~n15203;
  assign n15205 = ~n15196 & ~n15204;
  assign n15206 = n11186 & n15205;
  assign n15207 = ~n15188 & ~n15206;
  assign n15208 = n10902 & n15207;
  assign n15209 = ~n15164 & ~n15208;
  assign n15210 = ~n10885 & ~n15209;
  assign n15211 = pi3870 & n9804;
  assign n15212 = pi3886 & n9774;
  assign n15213 = ~n15211 & ~n15212;
  assign n15214 = pi3854 & n9802;
  assign n15215 = pi3918 & n9781;
  assign n15216 = pi3902 & n9771;
  assign n15217 = ~n15215 & ~n15216;
  assign n15218 = pi3950 & n9791;
  assign n15219 = pi3934 & n9788;
  assign n15220 = ~n15218 & ~n15219;
  assign n15221 = n15217 & n15220;
  assign n15222 = ~n15214 & n15221;
  assign n15223 = n15213 & n15222;
  assign n15224 = pi3870 & n9799;
  assign n15225 = n15223 & ~n15224;
  assign n15226 = pi3982 & n9783;
  assign n15227 = pi3966 & n9793;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = n15225 & n15228;
  assign n15230 = ~n9472 & ~n15229;
  assign n15231 = pi1331 & ~n9216;
  assign n15232 = pi3513 & ~n10410;
  assign n15233 = ~n15231 & ~n15232;
  assign n15234 = pi0595 & pi1359;
  assign n15235 = pi0391 & pi1057;
  assign n15236 = ~n15234 & ~n15235;
  assign n15237 = n15233 & n15236;
  assign n15238 = n9475 & ~n15237;
  assign n15239 = ~pi0979 & pi2616;
  assign n15240 = pi0979 & pi2609;
  assign n15241 = ~n15239 & ~n15240;
  assign n15242 = pi0763 & ~n15241;
  assign n15243 = ~pi0979 & pi2628;
  assign n15244 = pi0979 & pi2622;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = pi0764 & ~n15245;
  assign n15247 = ~n15242 & ~n15246;
  assign n15248 = ~pi0979 & pi2538;
  assign n15249 = pi0979 & pi3175;
  assign n15250 = ~n15248 & ~n15249;
  assign n15251 = pi0765 & ~n15250;
  assign n15252 = ~pi0979 & pi2896;
  assign n15253 = pi0979 & pi3184;
  assign n15254 = ~n15252 & ~n15253;
  assign n15255 = pi0766 & ~n15254;
  assign n15256 = ~n15251 & ~n15255;
  assign n15257 = pi0087 & ~pi0979;
  assign n15258 = pi0085 & pi0979;
  assign n15259 = ~n15257 & ~n15258;
  assign n15260 = pi0720 & ~n15259;
  assign n15261 = pi0257 & ~pi0979;
  assign n15262 = pi0255 & pi0979;
  assign n15263 = ~n15261 & ~n15262;
  assign n15264 = pi0721 & ~n15263;
  assign n15265 = ~n15260 & ~n15264;
  assign n15266 = n15256 & n15265;
  assign n15267 = ~n9499 & n15266;
  assign n15268 = n15247 & n15267;
  assign n15269 = n9486 & ~n15268;
  assign n15270 = ~n15238 & ~n15269;
  assign n15271 = ~pi0979 & pi2854;
  assign n15272 = pi0979 & pi2137;
  assign n15273 = ~n15271 & ~n15272;
  assign n15274 = pi0717 & ~n15273;
  assign n15275 = pi0234 & ~pi0979;
  assign n15276 = pi0233 & pi0979;
  assign n15277 = ~n15275 & ~n15276;
  assign n15278 = pi0716 & ~n15277;
  assign n15279 = pi0283 & ~pi0979;
  assign n15280 = pi0281 & pi0979;
  assign n15281 = ~n15279 & ~n15280;
  assign n15282 = pi0761 & ~n15281;
  assign n15283 = ~n15278 & ~n15282;
  assign n15284 = ~n9535 & n15283;
  assign n15285 = ~n9531 & n15284;
  assign n15286 = ~n15274 & n15285;
  assign n15287 = n9523 & ~n15286;
  assign n15288 = pi0979 & pi2156;
  assign n15289 = ~pi0979 & pi2778;
  assign n15290 = ~n15288 & ~n15289;
  assign n15291 = pi0767 & ~n15290;
  assign n15292 = ~pi0979 & pi2511;
  assign n15293 = pi0979 & pi1966;
  assign n15294 = ~n15292 & ~n15293;
  assign n15295 = pi0768 & ~n15294;
  assign n15296 = ~n15291 & ~n15295;
  assign n15297 = pi0979 & pi2174;
  assign n15298 = ~pi0979 & pi2801;
  assign n15299 = ~n15297 & ~n15298;
  assign n15300 = pi0836 & ~n15299;
  assign n15301 = ~pi0979 & pi3079;
  assign n15302 = pi0979 & pi2190;
  assign n15303 = ~n15301 & ~n15302;
  assign n15304 = pi0837 & ~n15303;
  assign n15305 = ~n15300 & ~n15304;
  assign n15306 = pi0180 & ~pi0979;
  assign n15307 = pi0165 & pi0979;
  assign n15308 = ~n15306 & ~n15307;
  assign n15309 = pi0838 & ~n15308;
  assign n15310 = n15305 & ~n15309;
  assign n15311 = n15296 & n15310;
  assign n15312 = n9549 & ~n15311;
  assign n15313 = ~n15287 & ~n15312;
  assign n15314 = pi1600 & pi2212;
  assign n15315 = pi1337 & pi2226;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = pi1338 & pi2240;
  assign n15318 = n15316 & ~n15317;
  assign n15319 = pi1346 & pi2672;
  assign n15320 = n15318 & ~n15319;
  assign n15321 = pi1339 & pi2254;
  assign n15322 = pi1345 & pi2658;
  assign n15323 = ~n15321 & ~n15322;
  assign n15324 = pi1347 & pi2615;
  assign n15325 = pi1348 & pi2696;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = pi1350 & pi2539;
  assign n15328 = n15326 & ~n15327;
  assign n15329 = pi1353 & pi2277;
  assign n15330 = n15328 & ~n15329;
  assign n15331 = pi1351 & pi2440;
  assign n15332 = pi1352 & pi2703;
  assign n15333 = ~n15331 & ~n15332;
  assign n15334 = n15330 & n15333;
  assign n15335 = n15323 & n15334;
  assign n15336 = n15320 & n15335;
  assign n15337 = n9577 & ~n15336;
  assign n15338 = pi1349 & pi2736;
  assign n15339 = pi1056 & pi2545;
  assign n15340 = ~n15338 & ~n15339;
  assign n15341 = pi1354 & pi2749;
  assign n15342 = n15340 & ~n15341;
  assign n15343 = pi1357 & pi2468;
  assign n15344 = n15342 & ~n15343;
  assign n15345 = pi1355 & pi2459;
  assign n15346 = pi1356 & pi2544;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = pi1340 & pi2289;
  assign n15349 = pi1341 & pi2088;
  assign n15350 = ~n15348 & ~n15349;
  assign n15351 = pi1342 & pi2311;
  assign n15352 = n15350 & ~n15351;
  assign n15353 = pi1055 & pi2565;
  assign n15354 = n15352 & ~n15353;
  assign n15355 = pi1343 & pi2325;
  assign n15356 = pi1054 & pi2534;
  assign n15357 = ~n15355 & ~n15356;
  assign n15358 = n15354 & n15357;
  assign n15359 = n15347 & n15358;
  assign n15360 = n15344 & n15359;
  assign n15361 = n9736 & ~n15360;
  assign n15362 = ~n15337 & ~n15361;
  assign n15363 = pi0224 & pi1336;
  assign n15364 = pi1333 & pi1714;
  assign n15365 = ~n15363 & ~n15364;
  assign n15366 = pi1332 & pi2580;
  assign n15367 = pi1335 & pi2595;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = n15365 & n15368;
  assign n15370 = n9726 & ~n15369;
  assign n15371 = pi1687 & n10557;
  assign n15372 = pi0971 & n9687;
  assign n15373 = pi1445 & n9691;
  assign n15374 = ~n15372 & ~n15373;
  assign n15375 = ~n15371 & n15374;
  assign n15376 = pi0899 & n9614;
  assign n15377 = pi1906 & n9618;
  assign n15378 = ~n15376 & ~n15377;
  assign n15379 = pi1736 & n11106;
  assign n15380 = pi0872 & n9707;
  assign n15381 = ~n15379 & ~n15380;
  assign n15382 = pi0791 & n9715;
  assign n15383 = pi1892 & n9718;
  assign n15384 = ~n15382 & ~n15383;
  assign n15385 = pi1684 & n10564;
  assign n15386 = n15384 & ~n15385;
  assign n15387 = n15381 & n15386;
  assign n15388 = pi1838 & n9698;
  assign n15389 = n15387 & ~n15388;
  assign n15390 = ~n11102 & n15389;
  assign n15391 = n15378 & n15390;
  assign n15392 = n15375 & n15391;
  assign n15393 = pi1784 & n9712;
  assign n15394 = n15392 & ~n15393;
  assign n15395 = pi1459 & n11145;
  assign n15396 = pi0820 & n9710;
  assign n15397 = ~n15395 & ~n15396;
  assign n15398 = pi3091 & n9647;
  assign n15399 = pi0725 & n9654;
  assign n15400 = ~n15398 & ~n15399;
  assign n15401 = pi0780 & n9670;
  assign n15402 = pi0930 & n9676;
  assign n15403 = ~n15401 & ~n15402;
  assign n15404 = pi2500 & n11158;
  assign n15405 = n15403 & ~n15404;
  assign n15406 = n15400 & n15405;
  assign n15407 = pi1931 & n9622;
  assign n15408 = n15406 & ~n15407;
  assign n15409 = pi1724 & n9679;
  assign n15410 = pi0336 & n9682;
  assign n15411 = ~n15409 & ~n15410;
  assign n15412 = n15408 & n15411;
  assign n15413 = n15397 & n15412;
  assign n15414 = n15394 & n15413;
  assign n15415 = pi1934 & ~n15414;
  assign n15416 = ~n15370 & ~n15415;
  assign n15417 = n15362 & n15416;
  assign n15418 = n15313 & n15417;
  assign n15419 = n15270 & n15418;
  assign n15420 = pi3295 & po3871;
  assign n15421 = n15419 & ~n15420;
  assign n15422 = ~pi1787 & ~n15421;
  assign n15423 = pi1787 & pi2834;
  assign n15424 = ~n15422 & ~n15423;
  assign n15425 = n9472 & ~n15424;
  assign n15426 = ~n15230 & ~n15425;
  assign n15427 = n10914 & ~n15426;
  assign n15428 = ~n11360 & n11364;
  assign n15429 = n11360 & ~n11364;
  assign n15430 = ~n15428 & ~n15429;
  assign n15431 = ~n11384 & ~n14414;
  assign n15432 = ~n11431 & ~n15431;
  assign n15433 = ~n15430 & ~n15432;
  assign n15434 = n15430 & n15432;
  assign n15435 = ~n15433 & ~n15434;
  assign n15436 = n11665 & ~n15435;
  assign n15437 = ~n11358 & ~n14405;
  assign n15438 = ~n11354 & ~n15437;
  assign n15439 = n11361 & ~n15438;
  assign n15440 = ~n11361 & n15438;
  assign n15441 = ~n15439 & ~n15440;
  assign n15442 = ~n11665 & ~n15441;
  assign n15443 = ~n15436 & ~n15442;
  assign n15444 = pi0518 & ~n15443;
  assign n15445 = n11615 & ~n15441;
  assign n15446 = ~n11615 & ~n15435;
  assign n15447 = ~n15445 & ~n15446;
  assign n15448 = ~pi0518 & ~n15447;
  assign n15449 = ~n15444 & ~n15448;
  assign n15450 = pi0682 & n11322;
  assign n15451 = pi0682 & ~n11260;
  assign n15452 = n11222 & n15451;
  assign n15453 = ~n15450 & ~n15452;
  assign n15454 = ~n15449 & n15453;
  assign n15455 = ~n10914 & ~n15454;
  assign n15456 = ~n15427 & ~n15455;
  assign n15457 = n11755 & ~n15456;
  assign n15458 = ~n15210 & ~n15457;
  assign po0227 = n15119 | ~n15458;
  assign n15460 = n14825 & po0227;
  assign n15461 = po0225 & n15460;
  assign n15462 = po0228 & n15461;
  assign n15463 = po0229 & ~n15462;
  assign po0061 = ~n10790 & n15463;
  assign n15465 = pi2497 & n8577;
  assign n15466 = pi2980 & ~n8577;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = ~n10668 & ~n15467;
  assign n15469 = pi1454 & n10668;
  assign n15470 = ~n15468 & ~n15469;
  assign n15471 = ~n11219 & ~n11756;
  assign n15472 = n15470 & n15471;
  assign n15473 = ~n11726 & n15472;
  assign n15474 = pi2513 & n8577;
  assign n15475 = pi2981 & ~n8577;
  assign n15476 = ~n15474 & ~n15475;
  assign n15477 = ~n10668 & ~n15476;
  assign n15478 = pi1455 & n10668;
  assign n15479 = ~n15477 & ~n15478;
  assign n15480 = pi2496 & n8577;
  assign n15481 = pi2979 & ~n8577;
  assign n15482 = ~n15480 & ~n15481;
  assign n15483 = ~n10668 & ~n15482;
  assign n15484 = pi1453 & n10668;
  assign n15485 = ~n15483 & ~n15484;
  assign n15486 = pi2495 & n8577;
  assign n15487 = pi2978 & ~n8577;
  assign n15488 = ~n15486 & ~n15487;
  assign n15489 = ~n10668 & ~n15488;
  assign n15490 = pi1452 & n10668;
  assign n15491 = ~n15489 & ~n15490;
  assign n15492 = n15485 & n15491;
  assign n15493 = n15479 & n15492;
  assign n15494 = n15473 & n15493;
  assign po0062 = ~n10790 & n15494;
  assign n15496 = ~n15479 & n15492;
  assign n15497 = n15473 & n15496;
  assign po0063 = ~n10790 & n15497;
  assign n15499 = ~n11756 & ~n15470;
  assign n15500 = ~n11726 & n15499;
  assign n15501 = ~n11219 & n15500;
  assign n15502 = n15493 & n15501;
  assign po0064 = ~n10790 & n15502;
  assign n15504 = n15496 & n15501;
  assign po0065 = ~n10790 & n15504;
  assign n15506 = ~n15485 & n15491;
  assign n15507 = n15479 & n15506;
  assign n15508 = n15473 & n15507;
  assign po0066 = ~n10790 & n15508;
  assign n15510 = ~n15479 & n15506;
  assign n15511 = n15473 & n15510;
  assign po0067 = ~n10790 & n15511;
  assign n15513 = n15501 & n15507;
  assign po0068 = ~n10790 & n15513;
  assign n15515 = n15501 & n15510;
  assign po0069 = ~n10790 & n15515;
  assign n15517 = ~n9365 & ~po3871;
  assign n15518 = ~n10743 & ~n15517;
  assign n15519 = ~n8567 & ~n10786;
  assign n15520 = ~n15518 & ~n15519;
  assign n15521 = ~n11784 & ~n12129;
  assign n15522 = ~n12065 & n15521;
  assign n15523 = n15461 & ~n15522;
  assign n15524 = po0229 & ~n15523;
  assign n15525 = ~n15494 & ~n15497;
  assign n15526 = ~n15524 & n15525;
  assign n15527 = ~n15502 & ~n15504;
  assign n15528 = ~n15515 & n15527;
  assign n15529 = ~n15513 & n15528;
  assign n15530 = ~n15508 & n15529;
  assign n15531 = ~n15511 & n15530;
  assign n15532 = n15526 & n15531;
  assign po0070 = n15520 | n15532;
  assign n15534 = pi3236 & pi3547;
  assign n15535 = pi0684 & pi3528;
  assign n15536 = ~n15534 & ~n15535;
  assign n15537 = pi3362 & ~n9873;
  assign n15538 = pi3505 & ~pi3515;
  assign n15539 = pi0684 & n15538;
  assign n15540 = ~n15537 & ~n15539;
  assign po3948 = ~n15536 | ~n15540;
  assign n15542 = ~pi3548 & ~n15538;
  assign n15543 = pi0404 & ~n15542;
  assign po3850 = ~pi0684 & n15543;
  assign po3627 = ~po3948 & ~po3850;
  assign n15546 = ~po3831 & po3627;
  assign n15547 = ~pi3551 & n15546;
  assign n15548 = ~po3841 & ~n15547;
  assign n15549 = pi3055 & n10747;
  assign n15550 = ~pi3641 & n15549;
  assign n15551 = n15548 & ~n15550;
  assign n15552 = ~pi3390 & n15551;
  assign n15553 = ~pi0684 & n9873;
  assign n15554 = pi2489 & ~n8670;
  assign n15555 = n9266 & ~n15554;
  assign n15556 = n8698 & n15555;
  assign n15557 = ~n9342 & ~n15556;
  assign n15558 = ~n15554 & n15557;
  assign n15559 = ~pi3481 & ~n15558;
  assign n15560 = pi0540 & ~n15555;
  assign n15561 = n15559 & ~n15560;
  assign n15562 = n15553 & ~n15561;
  assign n15563 = pi3401 & pi3422;
  assign n15564 = pi3400 & pi3403;
  assign n15565 = pi3402 & n15564;
  assign n15566 = pi3404 & n15565;
  assign n15567 = pi3414 & n15566;
  assign n15568 = pi3413 & n15567;
  assign n15569 = pi3405 & n15568;
  assign n15570 = pi3406 & pi3411;
  assign n15571 = n15569 & n15570;
  assign n15572 = n15563 & n15571;
  assign n15573 = pi3421 & n15572;
  assign n15574 = pi3420 & n15573;
  assign n15575 = pi3430 & n15574;
  assign n15576 = ~pi3430 & ~n15574;
  assign n15577 = ~n15575 & ~n15576;
  assign n15578 = n15562 & n15577;
  assign n15579 = pi3236 & n15553;
  assign n15580 = pi0814 & n15579;
  assign n15581 = ~n15578 & ~n15580;
  assign n15582 = ~pi0684 & ~pi3236;
  assign n15583 = ~pi3481 & n9342;
  assign n15584 = ~pi0540 & n15583;
  assign n15585 = n15582 & n15584;
  assign n15586 = n15553 & n15585;
  assign n15587 = pi3641 & n9373;
  assign n15588 = n9374 & n10755;
  assign n15589 = n15587 & n15588;
  assign n15590 = pi2193 & n15589;
  assign n15591 = n15586 & n15590;
  assign n15592 = ~pi1713 & pi1798;
  assign n15593 = pi1800 & n15592;
  assign n15594 = pi1713 & pi1798;
  assign n15595 = pi1799 & n15594;
  assign n15596 = ~n15593 & ~n15595;
  assign n15597 = pi1713 & ~pi1798;
  assign n15598 = pi1996 & n15597;
  assign n15599 = ~pi1713 & ~pi1798;
  assign n15600 = pi2008 & n15599;
  assign n15601 = ~n15598 & ~n15600;
  assign n15602 = n15596 & n15601;
  assign n15603 = ~pi3437 & n15602;
  assign n15604 = pi3437 & ~n15602;
  assign n15605 = ~n15603 & ~n15604;
  assign n15606 = pi2071 & n15597;
  assign n15607 = pi1999 & n15592;
  assign n15608 = ~n15606 & ~n15607;
  assign n15609 = pi2361 & n15599;
  assign n15610 = pi1988 & n15594;
  assign n15611 = ~n15609 & ~n15610;
  assign n15612 = n15608 & n15611;
  assign n15613 = ~pi3433 & n15612;
  assign n15614 = pi3433 & ~n15612;
  assign n15615 = ~n15613 & ~n15614;
  assign n15616 = pi1997 & n15597;
  assign n15617 = pi2000 & n15592;
  assign n15618 = ~n15616 & ~n15617;
  assign n15619 = pi2009 & n15599;
  assign n15620 = pi1989 & n15594;
  assign n15621 = ~n15619 & ~n15620;
  assign n15622 = n15618 & n15621;
  assign n15623 = ~pi3460 & n15622;
  assign n15624 = pi3460 & ~n15622;
  assign n15625 = ~n15623 & ~n15624;
  assign n15626 = pi2337 & n15597;
  assign n15627 = pi2352 & n15592;
  assign n15628 = ~n15626 & ~n15627;
  assign n15629 = pi2360 & n15599;
  assign n15630 = pi1986 & n15594;
  assign n15631 = ~n15629 & ~n15630;
  assign n15632 = n15628 & n15631;
  assign n15633 = ~pi3457 & n15632;
  assign n15634 = pi3457 & ~n15632;
  assign n15635 = ~n15633 & ~n15634;
  assign n15636 = ~n15625 & ~n15635;
  assign n15637 = ~n15615 & n15636;
  assign n15638 = ~n15605 & n15637;
  assign n15639 = pi2371 & n15599;
  assign n15640 = pi2333 & n15594;
  assign n15641 = ~n15639 & ~n15640;
  assign n15642 = pi2349 & n15597;
  assign n15643 = pi2007 & n15592;
  assign n15644 = ~n15642 & ~n15643;
  assign n15645 = n15641 & n15644;
  assign n15646 = ~pi3454 & n15645;
  assign n15647 = pi3454 & ~n15645;
  assign n15648 = ~n15646 & ~n15647;
  assign n15649 = pi2073 & n15597;
  assign n15650 = pi1998 & n15592;
  assign n15651 = ~n15649 & ~n15650;
  assign n15652 = pi2389 & n15599;
  assign n15653 = pi2075 & n15594;
  assign n15654 = ~n15652 & ~n15653;
  assign n15655 = n15651 & n15654;
  assign n15656 = ~pi3434 & n15655;
  assign n15657 = pi3434 & ~n15655;
  assign n15658 = ~n15656 & ~n15657;
  assign n15659 = pi2350 & n15597;
  assign n15660 = pi2388 & n15592;
  assign n15661 = ~n15659 & ~n15660;
  assign n15662 = pi2372 & n15599;
  assign n15663 = pi2334 & n15594;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = n15661 & n15664;
  assign n15666 = ~pi3455 & n15665;
  assign n15667 = pi3455 & ~n15665;
  assign n15668 = ~n15666 & ~n15667;
  assign n15669 = pi2336 & n15597;
  assign n15670 = pi2351 & n15592;
  assign n15671 = ~n15669 & ~n15670;
  assign n15672 = pi2359 & n15599;
  assign n15673 = pi1987 & n15594;
  assign n15674 = ~n15672 & ~n15673;
  assign n15675 = n15671 & n15674;
  assign n15676 = ~pi3456 & n15675;
  assign n15677 = pi3456 & ~n15675;
  assign n15678 = ~n15676 & ~n15677;
  assign n15679 = ~n15668 & ~n15678;
  assign n15680 = ~n15658 & n15679;
  assign n15681 = ~n15648 & n15680;
  assign n15682 = n15638 & n15681;
  assign n15683 = pi2342 & n15597;
  assign n15684 = pi2355 & n15592;
  assign n15685 = ~n15683 & ~n15684;
  assign n15686 = pi2072 & n15599;
  assign n15687 = pi2074 & n15594;
  assign n15688 = ~n15686 & ~n15687;
  assign n15689 = n15685 & n15688;
  assign n15690 = ~pi2408 & n15689;
  assign n15691 = pi2408 & ~n15689;
  assign n15692 = ~n15690 & ~n15691;
  assign n15693 = pi2341 & n15597;
  assign n15694 = pi2391 & n15592;
  assign n15695 = ~n15693 & ~n15694;
  assign n15696 = pi2365 & n15599;
  assign n15697 = pi1992 & n15594;
  assign n15698 = ~n15696 & ~n15697;
  assign n15699 = n15695 & n15698;
  assign n15700 = ~pi2400 & n15699;
  assign n15701 = pi2400 & ~n15699;
  assign n15702 = ~n15700 & ~n15701;
  assign n15703 = pi2344 & n15597;
  assign n15704 = pi2356 & n15592;
  assign n15705 = ~n15703 & ~n15704;
  assign n15706 = pi2367 & n15599;
  assign n15707 = pi1994 & n15594;
  assign n15708 = ~n15706 & ~n15707;
  assign n15709 = n15705 & n15708;
  assign n15710 = ~pi3450 & n15709;
  assign n15711 = pi3450 & ~n15709;
  assign n15712 = ~n15710 & ~n15711;
  assign n15713 = pi2366 & n15599;
  assign n15714 = pi1993 & n15594;
  assign n15715 = ~n15713 & ~n15714;
  assign n15716 = pi2343 & n15597;
  assign n15717 = pi2003 & n15592;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = n15715 & n15718;
  assign n15720 = ~pi3458 & n15719;
  assign n15721 = pi3458 & ~n15719;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = ~n15712 & ~n15722;
  assign n15724 = ~n15702 & n15723;
  assign n15725 = ~n15692 & n15724;
  assign n15726 = pi2069 & n15599;
  assign n15727 = pi1995 & n15594;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = pi2345 & n15597;
  assign n15730 = pi2004 & n15592;
  assign n15731 = ~n15729 & ~n15730;
  assign n15732 = n15728 & n15731;
  assign n15733 = ~pi3478 & n15732;
  assign n15734 = pi3478 & ~n15732;
  assign n15735 = ~n15733 & ~n15734;
  assign n15736 = pi2348 & n15597;
  assign n15737 = pi2006 & n15592;
  assign n15738 = ~n15736 & ~n15737;
  assign n15739 = pi2370 & n15599;
  assign n15740 = pi2332 & n15594;
  assign n15741 = ~n15739 & ~n15740;
  assign n15742 = n15738 & n15741;
  assign n15743 = ~pi3453 & n15742;
  assign n15744 = pi3453 & ~n15742;
  assign n15745 = ~n15743 & ~n15744;
  assign n15746 = pi2347 & n15597;
  assign n15747 = pi2357 & n15592;
  assign n15748 = ~n15746 & ~n15747;
  assign n15749 = pi2369 & n15599;
  assign n15750 = pi2331 & n15594;
  assign n15751 = ~n15749 & ~n15750;
  assign n15752 = n15748 & n15751;
  assign n15753 = ~pi3432 & n15752;
  assign n15754 = pi3432 & ~n15752;
  assign n15755 = ~n15753 & ~n15754;
  assign n15756 = pi2346 & n15597;
  assign n15757 = pi2005 & n15592;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = pi2368 & n15599;
  assign n15760 = pi2330 & n15594;
  assign n15761 = ~n15759 & ~n15760;
  assign n15762 = n15758 & n15761;
  assign n15763 = ~pi3459 & n15762;
  assign n15764 = pi3459 & ~n15762;
  assign n15765 = ~n15763 & ~n15764;
  assign n15766 = ~n15755 & ~n15765;
  assign n15767 = ~n15745 & n15766;
  assign n15768 = ~n15735 & n15767;
  assign n15769 = n15725 & n15768;
  assign n15770 = pi2339 & n15597;
  assign n15771 = pi2002 & n15592;
  assign n15772 = ~n15770 & ~n15771;
  assign n15773 = pi2363 & n15599;
  assign n15774 = pi1991 & n15594;
  assign n15775 = ~n15773 & ~n15774;
  assign n15776 = n15772 & n15775;
  assign n15777 = pi2514 & n15776;
  assign n15778 = ~pi2514 & ~n15776;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = ~pi1797 & n15779;
  assign n15781 = pi2070 & n15597;
  assign n15782 = pi2390 & n15592;
  assign n15783 = ~n15781 & ~n15782;
  assign n15784 = pi2076 & n15599;
  assign n15785 = pi2077 & n15594;
  assign n15786 = ~n15784 & ~n15785;
  assign n15787 = n15783 & n15786;
  assign n15788 = ~pi2472 & n15787;
  assign n15789 = pi2472 & ~n15787;
  assign n15790 = ~n15788 & ~n15789;
  assign n15791 = n15780 & ~n15790;
  assign n15792 = n15769 & n15791;
  assign n15793 = n15682 & n15792;
  assign n15794 = n15591 & n15793;
  assign n15795 = ~n8712 & ~n8734;
  assign n15796 = ~pi0976 & ~n15795;
  assign n15797 = pi1044 & ~n8742;
  assign n15798 = ~n8743 & ~n15797;
  assign n15799 = pi1043 & ~n8734;
  assign n15800 = ~n8742 & ~n15799;
  assign n15801 = ~n15798 & n15800;
  assign n15802 = n15796 & n15801;
  assign n15803 = pi1297 & n15802;
  assign n15804 = pi0976 & ~n15795;
  assign n15805 = ~n15798 & ~n15800;
  assign n15806 = n15804 & n15805;
  assign n15807 = pi1255 & n15806;
  assign n15808 = ~n15803 & ~n15807;
  assign n15809 = pi0976 & n15795;
  assign n15810 = n15805 & n15809;
  assign n15811 = pi1283 & n15810;
  assign n15812 = n15801 & n15809;
  assign n15813 = pi1129 & n15812;
  assign n15814 = ~n15811 & ~n15813;
  assign n15815 = n15798 & n15800;
  assign n15816 = ~pi0976 & n15795;
  assign n15817 = n15815 & n15816;
  assign n15818 = pi1227 & n15817;
  assign n15819 = n15796 & n15815;
  assign n15820 = pi1199 & n15819;
  assign n15821 = ~n15818 & ~n15820;
  assign n15822 = n15798 & ~n15800;
  assign n15823 = n15816 & n15822;
  assign n15824 = pi1171 & n15823;
  assign n15825 = n15804 & n15815;
  assign n15826 = pi1213 & n15825;
  assign n15827 = ~n15824 & ~n15826;
  assign n15828 = n15821 & n15827;
  assign n15829 = n15814 & n15828;
  assign n15830 = n15808 & n15829;
  assign n15831 = n15796 & n15822;
  assign n15832 = pi1143 & n15831;
  assign n15833 = n15804 & n15822;
  assign n15834 = pi1157 & n15833;
  assign n15835 = ~n15832 & ~n15834;
  assign n15836 = n15805 & n15816;
  assign n15837 = pi1269 & n15836;
  assign n15838 = n15796 & n15805;
  assign n15839 = pi1241 & n15838;
  assign n15840 = ~n15837 & ~n15839;
  assign n15841 = n15809 & n15815;
  assign n15842 = pi1325 & n15841;
  assign n15843 = n15809 & n15822;
  assign n15844 = pi1185 & n15843;
  assign n15845 = ~n15842 & ~n15844;
  assign n15846 = n15801 & n15816;
  assign n15847 = pi1115 & n15846;
  assign n15848 = n15801 & n15804;
  assign n15849 = pi1311 & n15848;
  assign n15850 = ~n15847 & ~n15849;
  assign n15851 = n15845 & n15850;
  assign n15852 = n15840 & n15851;
  assign n15853 = n15835 & n15852;
  assign n15854 = n15830 & n15853;
  assign n15855 = n15794 & ~n15854;
  assign n15856 = n15585 & n15793;
  assign n15857 = ~n15590 & n15856;
  assign n15858 = n8698 & ~n9342;
  assign n15859 = n15555 & n15858;
  assign n15860 = ~n15554 & n15859;
  assign n15861 = pi0540 & n15556;
  assign n15862 = ~n15860 & ~n15861;
  assign n15863 = ~n15857 & n15862;
  assign n15864 = ~pi0008 & ~pi3459;
  assign n15865 = pi0008 & pi3459;
  assign n15866 = ~n15864 & ~n15865;
  assign n15867 = ~pi0010 & ~pi3450;
  assign n15868 = pi0010 & pi3450;
  assign n15869 = ~n15867 & ~n15868;
  assign n15870 = pi0007 & pi3432;
  assign n15871 = ~pi0007 & ~pi3432;
  assign n15872 = ~n15870 & ~n15871;
  assign n15873 = pi3352 & pi3457;
  assign n15874 = pi3331 & pi3433;
  assign n15875 = n15873 & n15874;
  assign n15876 = ~pi3331 & ~pi3433;
  assign n15877 = ~pi3352 & ~pi3457;
  assign n15878 = n15876 & n15877;
  assign n15879 = ~n15875 & ~n15878;
  assign n15880 = n15874 & n15877;
  assign n15881 = n15879 & ~n15880;
  assign n15882 = n15873 & n15876;
  assign n15883 = n15881 & ~n15882;
  assign n15884 = ~pi3347 & ~pi3437;
  assign n15885 = pi3347 & pi3437;
  assign n15886 = ~n15884 & ~n15885;
  assign n15887 = pi3332 & pi3460;
  assign n15888 = ~n15886 & n15887;
  assign n15889 = ~pi3332 & ~pi3460;
  assign n15890 = pi3347 & n15889;
  assign n15891 = pi3437 & n15890;
  assign n15892 = ~n15888 & ~n15891;
  assign n15893 = n15884 & n15889;
  assign n15894 = n15892 & ~n15893;
  assign n15895 = ~pi3354 & ~pi3456;
  assign n15896 = pi3354 & pi3456;
  assign n15897 = ~n15895 & ~n15896;
  assign n15898 = pi3423 & ~n15897;
  assign n15899 = ~n15894 & n15898;
  assign n15900 = ~n15883 & n15899;
  assign n15901 = pi1930 & ~n15900;
  assign n15902 = ~pi0004 & ~pi3455;
  assign n15903 = pi0004 & pi3455;
  assign n15904 = ~n15902 & ~n15903;
  assign n15905 = n15901 & ~n15904;
  assign n15906 = ~pi0011 & ~pi3458;
  assign n15907 = pi0011 & pi3458;
  assign n15908 = ~n15906 & ~n15907;
  assign n15909 = ~pi0003 & ~pi3434;
  assign n15910 = pi0003 & pi3434;
  assign n15911 = ~n15909 & ~n15910;
  assign n15912 = ~n15908 & ~n15911;
  assign n15913 = n15905 & n15912;
  assign n15914 = ~pi0005 & ~pi3454;
  assign n15915 = pi0005 & pi3454;
  assign n15916 = ~n15914 & ~n15915;
  assign n15917 = ~pi0006 & ~pi3453;
  assign n15918 = pi0006 & pi3453;
  assign n15919 = ~n15917 & ~n15918;
  assign n15920 = ~n15916 & ~n15919;
  assign n15921 = n15913 & n15920;
  assign n15922 = pi0002 & n15921;
  assign n15923 = ~n15872 & n15922;
  assign n15924 = ~pi0009 & ~pi3478;
  assign n15925 = pi0009 & pi3478;
  assign n15926 = ~n15924 & ~n15925;
  assign n15927 = n15923 & ~n15926;
  assign n15928 = ~n15869 & n15927;
  assign n15929 = ~n15866 & n15928;
  assign n15930 = pi3355 & ~n15901;
  assign n15931 = pi0000 & n15901;
  assign n15932 = ~n15930 & ~n15931;
  assign n15933 = pi3353 & ~n15901;
  assign n15934 = pi0001 & n15901;
  assign n15935 = ~n15933 & ~n15934;
  assign n15936 = n15932 & n15935;
  assign n15937 = n15929 & ~n15936;
  assign n15938 = n15585 & n15937;
  assign n15939 = n15863 & ~n15938;
  assign n15940 = n15553 & ~n15939;
  assign n15941 = ~n8765 & n15940;
  assign n15942 = ~n15855 & ~n15941;
  assign n15943 = n15553 & n15554;
  assign n15944 = ~n9342 & n15943;
  assign n15945 = pi2763 & ~n8670;
  assign n15946 = pi2375 & n15945;
  assign n15947 = ~n8765 & ~n15945;
  assign n15948 = ~n15946 & ~n15947;
  assign n15949 = n15944 & ~n15948;
  assign n15950 = pi0013 & n15901;
  assign n15951 = ~n15933 & ~n15950;
  assign n15952 = pi0012 & n15901;
  assign n15953 = ~n15930 & ~n15952;
  assign n15954 = n15951 & n15953;
  assign n15955 = ~pi0032 & ~pi3453;
  assign n15956 = pi0032 & pi3453;
  assign n15957 = ~n15955 & ~n15956;
  assign n15958 = ~pi0033 & ~pi3432;
  assign n15959 = pi0033 & pi3432;
  assign n15960 = ~n15958 & ~n15959;
  assign n15961 = pi0036 & pi3450;
  assign n15962 = ~pi0036 & ~pi3450;
  assign n15963 = ~n15961 & ~n15962;
  assign n15964 = ~pi0037 & ~pi3458;
  assign n15965 = pi0037 & pi3458;
  assign n15966 = ~n15964 & ~n15965;
  assign n15967 = n15901 & ~n15966;
  assign n15968 = ~pi0029 & ~pi3434;
  assign n15969 = pi0029 & pi3434;
  assign n15970 = ~n15968 & ~n15969;
  assign n15971 = ~pi0030 & ~pi3455;
  assign n15972 = pi0030 & pi3455;
  assign n15973 = ~n15971 & ~n15972;
  assign n15974 = ~n15970 & ~n15973;
  assign n15975 = n15967 & n15974;
  assign n15976 = ~pi0034 & ~pi3459;
  assign n15977 = pi0034 & pi3459;
  assign n15978 = ~n15976 & ~n15977;
  assign n15979 = ~pi0035 & ~pi3478;
  assign n15980 = pi0035 & pi3478;
  assign n15981 = ~n15979 & ~n15980;
  assign n15982 = ~n15978 & ~n15981;
  assign n15983 = n15975 & n15982;
  assign n15984 = pi0028 & n15983;
  assign n15985 = ~n15963 & n15984;
  assign n15986 = ~pi0031 & ~pi3454;
  assign n15987 = pi0031 & pi3454;
  assign n15988 = ~n15986 & ~n15987;
  assign n15989 = n15985 & ~n15988;
  assign n15990 = ~n15960 & n15989;
  assign n15991 = ~n15957 & n15990;
  assign n15992 = ~n15954 & n15991;
  assign n15993 = n15586 & n15992;
  assign n15994 = pi0027 & n15993;
  assign n15995 = ~n15949 & ~n15994;
  assign n15996 = ~pi3236 & ~pi3481;
  assign n15997 = n9342 & ~n15992;
  assign n15998 = ~n15793 & n15997;
  assign n15999 = n15996 & n15998;
  assign n16000 = ~n8698 & n15555;
  assign n16001 = pi0540 & ~n16000;
  assign n16002 = n15999 & ~n16001;
  assign n16003 = ~n15937 & n16002;
  assign n16004 = ~pi3589 & n16003;
  assign n16005 = ~pi0684 & n8563;
  assign n16006 = n16004 & n16005;
  assign n16007 = pi3432 & pi3450;
  assign n16008 = pi3434 & pi3455;
  assign n16009 = pi3437 & pi3460;
  assign n16010 = pi3433 & pi3457;
  assign n16011 = pi3456 & n16010;
  assign n16012 = n16009 & n16011;
  assign n16013 = pi3453 & pi3454;
  assign n16014 = n16012 & n16013;
  assign n16015 = n16008 & n16014;
  assign n16016 = pi3478 & n16015;
  assign n16017 = pi3459 & n16016;
  assign n16018 = n16007 & n16017;
  assign n16019 = pi3458 & n16018;
  assign n16020 = ~pi3458 & ~n16018;
  assign n16021 = ~n16019 & ~n16020;
  assign n16022 = n16006 & n16021;
  assign n16023 = n15995 & ~n16022;
  assign n16024 = n15942 & n16023;
  assign n16025 = n15581 & n16024;
  assign n16026 = n15552 & ~n16025;
  assign n16027 = pi0909 & n8589;
  assign n16028 = po3841 & n16027;
  assign n16029 = ~n8589 & po3841;
  assign n16030 = pi0752 & n8577;
  assign n16031 = n16029 & n16030;
  assign n16032 = ~n16028 & ~n16031;
  assign n16033 = ~n15552 & ~n16032;
  assign n16034 = ~po3841 & ~n15552;
  assign n16035 = ~pi3390 & ~n15550;
  assign n16036 = pi3519 & n8561;
  assign n16037 = pi0421 & ~n8561;
  assign po3845 = n16036 | n16037;
  assign n16039 = ~n16035 & po3845;
  assign n16040 = pi3458 & n16035;
  assign n16041 = ~n16039 & ~n16040;
  assign n16042 = n16034 & ~n16041;
  assign n16043 = ~n16033 & ~n16042;
  assign po0243 = n16026 | ~n16043;
  assign n16045 = pi3433 & n16009;
  assign n16046 = pi3457 & n16045;
  assign n16047 = n16008 & n16046;
  assign n16048 = pi3456 & n16047;
  assign n16049 = pi3454 & n16048;
  assign n16050 = pi3478 & n16049;
  assign n16051 = pi3459 & n16050;
  assign n16052 = pi3453 & n16051;
  assign n16053 = pi3432 & n16052;
  assign n16054 = ~pi3450 & ~n16053;
  assign n16055 = pi3450 & n16053;
  assign n16056 = ~n16054 & ~n16055;
  assign n16057 = n16006 & n16056;
  assign n16058 = pi1298 & n15802;
  assign n16059 = pi1256 & n15806;
  assign n16060 = ~n16058 & ~n16059;
  assign n16061 = pi1284 & n15810;
  assign n16062 = pi1130 & n15812;
  assign n16063 = ~n16061 & ~n16062;
  assign n16064 = pi1228 & n15817;
  assign n16065 = pi1200 & n15819;
  assign n16066 = ~n16064 & ~n16065;
  assign n16067 = pi1172 & n15823;
  assign n16068 = pi1214 & n15825;
  assign n16069 = ~n16067 & ~n16068;
  assign n16070 = n16066 & n16069;
  assign n16071 = n16063 & n16070;
  assign n16072 = n16060 & n16071;
  assign n16073 = pi1270 & n15836;
  assign n16074 = pi1242 & n15838;
  assign n16075 = ~n16073 & ~n16074;
  assign n16076 = pi1116 & n15846;
  assign n16077 = pi1312 & n15848;
  assign n16078 = ~n16076 & ~n16077;
  assign n16079 = pi1144 & n15831;
  assign n16080 = pi1158 & n15833;
  assign n16081 = ~n16079 & ~n16080;
  assign n16082 = pi1326 & n15841;
  assign n16083 = pi1186 & n15843;
  assign n16084 = ~n16082 & ~n16083;
  assign n16085 = n16081 & n16084;
  assign n16086 = n16078 & n16085;
  assign n16087 = n16075 & n16086;
  assign n16088 = n16072 & n16087;
  assign n16089 = n15794 & ~n16088;
  assign n16090 = ~n9257 & n15940;
  assign n16091 = ~n16089 & ~n16090;
  assign n16092 = pi3406 & n15569;
  assign n16093 = n15563 & n16092;
  assign n16094 = pi3411 & n16093;
  assign n16095 = pi3420 & n16094;
  assign n16096 = ~pi3421 & ~n16095;
  assign n16097 = pi3421 & n16095;
  assign n16098 = ~n16096 & ~n16097;
  assign n16099 = n15562 & n16098;
  assign n16100 = pi0815 & n15579;
  assign n16101 = ~n16099 & ~n16100;
  assign n16102 = pi2376 & n15945;
  assign n16103 = ~n9257 & ~n15945;
  assign n16104 = ~n16102 & ~n16103;
  assign n16105 = n15944 & ~n16104;
  assign n16106 = pi0026 & n15993;
  assign n16107 = ~n16105 & ~n16106;
  assign n16108 = n16101 & n16107;
  assign n16109 = n16091 & n16108;
  assign n16110 = ~n16057 & n16109;
  assign n16111 = n15552 & ~n16110;
  assign n16112 = pi0819 & n8589;
  assign n16113 = n8577 & ~n8589;
  assign n16114 = pi0779 & n16113;
  assign n16115 = ~n16112 & ~n16114;
  assign n16116 = po3841 & ~n16115;
  assign n16117 = ~n15552 & n16116;
  assign n16118 = ~n16111 & ~n16117;
  assign n16119 = pi3450 & n16035;
  assign n16120 = pi3512 & n8561;
  assign n16121 = pi0405 & ~n8561;
  assign po3838 = n16120 | n16121;
  assign n16123 = ~n16035 & po3838;
  assign n16124 = ~n16119 & ~n16123;
  assign n16125 = n16034 & ~n16124;
  assign po0242 = ~n16118 | n16125;
  assign n16127 = pi3680 & po0242;
  assign n16128 = ~po0243 & ~n16127;
  assign n16129 = ~pi0404 & n15538;
  assign n16130 = ~pi0684 & pi3190;
  assign n16131 = n16129 & n16130;
  assign n16132 = pi3523 & n8551;
  assign n16133 = ~n16131 & ~n16132;
  assign n16134 = ~pi0404 & pi3190;
  assign n16135 = pi3547 & n16134;
  assign n16136 = ~pi0684 & n16135;
  assign po3849 = ~n16133 | n16136;
  assign n16138 = n8564 & n8626;
  assign n16139 = n15547 & n16138;
  assign n16140 = n9897 & n16139;
  assign n16141 = ~po3850 & n16140;
  assign n16142 = ~po3849 & n16141;
  assign n16143 = ~n8577 & ~n8589;
  assign po3893 = pi3586 & pi3591;
  assign n16145 = po3850 & ~po3893;
  assign n16146 = n16143 & n16145;
  assign n16147 = n16035 & po3849;
  assign n16148 = ~n16146 & ~n16147;
  assign n16149 = ~pi3682 & n16148;
  assign n16150 = ~n16142 & n16149;
  assign po0080 = n16128 & n16150;
  assign n16152 = pi2502 & n8577;
  assign n16153 = pi2408 & ~n8577;
  assign n16154 = ~n16152 & ~n16153;
  assign n16155 = ~n10668 & ~n16154;
  assign n16156 = pi1461 & n10668;
  assign n16157 = ~n16155 & ~n16156;
  assign n16158 = ~n16142 & n16157;
  assign n16159 = pi2499 & n8577;
  assign n16160 = pi2400 & ~n8577;
  assign n16161 = ~n16159 & ~n16160;
  assign n16162 = ~n10668 & ~n16161;
  assign n16163 = pi1458 & n10668;
  assign n16164 = ~n16162 & ~n16163;
  assign n16165 = pi2498 & n8577;
  assign n16166 = pi2472 & ~n8577;
  assign n16167 = ~n16165 & ~n16166;
  assign n16168 = ~n10668 & ~n16167;
  assign n16169 = pi1456 & n10668;
  assign n16170 = ~n16168 & ~n16169;
  assign n16171 = pi2512 & n8577;
  assign n16172 = pi2514 & ~n8577;
  assign n16173 = ~n16171 & ~n16172;
  assign n16174 = ~n10668 & ~n16173;
  assign n16175 = pi1457 & n10668;
  assign n16176 = ~n16174 & ~n16175;
  assign n16177 = n16170 & n16176;
  assign n16178 = n16149 & n16177;
  assign n16179 = ~po0243 & po0242;
  assign n16180 = pi3680 & n16179;
  assign n16181 = ~pi3680 & po0243;
  assign n16182 = ~po0242 & n16181;
  assign n16183 = ~n16180 & ~n16182;
  assign n16184 = n16178 & ~n16183;
  assign n16185 = n16164 & n16184;
  assign po0081 = n16158 & n16185;
  assign n16187 = ~n16142 & ~n16157;
  assign po0082 = n16185 & n16187;
  assign n16189 = ~n16142 & n16184;
  assign n16190 = n16157 & ~n16164;
  assign po0083 = n16189 & n16190;
  assign n16192 = ~n16157 & ~n16164;
  assign po0084 = n16189 & n16192;
  assign n16194 = n16164 & ~n16176;
  assign n16195 = n16157 & n16194;
  assign n16196 = n16150 & ~n16183;
  assign n16197 = n16170 & n16196;
  assign po0085 = n16195 & n16197;
  assign n16199 = ~n16157 & n16194;
  assign po0086 = n16197 & n16199;
  assign n16201 = ~n16164 & ~n16176;
  assign n16202 = n16157 & n16201;
  assign po0087 = n16197 & n16202;
  assign n16204 = ~n16157 & n16201;
  assign po0088 = n16197 & n16204;
  assign n16206 = pi0418 & ~n8561;
  assign n16207 = n15550 & n16206;
  assign n16208 = po3849 & ~n16207;
  assign n16209 = pi0752 & ~n8584;
  assign n16210 = n8581 & ~n16209;
  assign n16211 = n8580 & n16210;
  assign n16212 = pi1840 & n16211;
  assign n16213 = ~pi1861 & n16212;
  assign n16214 = ~pi3099 & n16213;
  assign n16215 = n8577 & n16214;
  assign n16216 = ~n8591 & n8602;
  assign n16217 = ~n16215 & ~n16216;
  assign n16218 = ~n8567 & ~n16217;
  assign n16219 = ~po3849 & ~n16218;
  assign po0089 = n16208 | n16219;
  assign n16221 = pi2059 & ~pi3626;
  assign n16222 = pi2540 & ~po0014;
  assign n16223 = pi1039 & ~po0015;
  assign n16224 = ~n16222 & ~n16223;
  assign n16225 = pi3350 & n8389;
  assign n16226 = pi3496 & n16225;
  assign n16227 = pi3350 & ~n8389;
  assign n16228 = pi0375 & n16227;
  assign n16229 = ~n16226 & ~n16228;
  assign n16230 = pi3520 & ~po0017;
  assign n16231 = n16229 & ~n16230;
  assign n16232 = n16224 & n16231;
  assign n16233 = pi3626 & ~n16232;
  assign po0099 = n16221 | n16233;
  assign n16235 = pi2061 & ~pi3626;
  assign n16236 = pi2549 & ~po0014;
  assign n16237 = pi1012 & ~po0015;
  assign n16238 = ~n16236 & ~n16237;
  assign n16239 = pi3497 & n16225;
  assign n16240 = pi0374 & n16227;
  assign n16241 = ~n16239 & ~n16240;
  assign n16242 = pi3511 & ~po0017;
  assign n16243 = n16241 & ~n16242;
  assign n16244 = n16238 & n16243;
  assign n16245 = pi3626 & ~n16244;
  assign po0100 = n16235 | n16245;
  assign n16247 = pi2058 & ~pi3626;
  assign n16248 = pi2646 & ~po0014;
  assign n16249 = pi1034 & ~po0015;
  assign n16250 = ~n16248 & ~n16249;
  assign n16251 = pi3495 & n16225;
  assign n16252 = pi0373 & n16227;
  assign n16253 = ~n16251 & ~n16252;
  assign n16254 = pi3510 & ~po0017;
  assign n16255 = n16253 & ~n16254;
  assign n16256 = n16250 & n16255;
  assign n16257 = pi3626 & ~n16256;
  assign po0101 = n16247 | n16257;
  assign n16259 = pi1841 & ~pi3626;
  assign n16260 = pi2551 & ~po0014;
  assign n16261 = pi1033 & ~po0015;
  assign n16262 = ~n16260 & ~n16261;
  assign n16263 = pi3500 & n16225;
  assign n16264 = pi0372 & n16227;
  assign n16265 = ~n16263 & ~n16264;
  assign n16266 = pi3521 & ~po0017;
  assign n16267 = n16265 & ~n16266;
  assign n16268 = n16262 & n16267;
  assign n16269 = pi3626 & ~n16268;
  assign po0102 = n16259 | n16269;
  assign n16271 = pi1467 & ~pi3626;
  assign n16272 = pi2553 & ~po0014;
  assign n16273 = pi1032 & ~po0015;
  assign n16274 = ~n16272 & ~n16273;
  assign n16275 = pi3499 & n16225;
  assign n16276 = pi0371 & n16227;
  assign n16277 = ~n16275 & ~n16276;
  assign n16278 = pi3509 & ~po0017;
  assign n16279 = n16277 & ~n16278;
  assign n16280 = n16274 & n16279;
  assign n16281 = pi3626 & ~n16280;
  assign po0103 = n16271 | n16281;
  assign n16283 = pi1603 & ~pi3626;
  assign n16284 = pi2645 & ~po0014;
  assign n16285 = pi1013 & ~po0015;
  assign n16286 = ~n16284 & ~n16285;
  assign n16287 = pi3503 & n16225;
  assign n16288 = pi0369 & n16227;
  assign n16289 = ~n16287 & ~n16288;
  assign n16290 = pi3508 & ~po0017;
  assign n16291 = n16289 & ~n16290;
  assign n16292 = n16286 & n16291;
  assign n16293 = pi3626 & ~n16292;
  assign po0104 = n16283 | n16293;
  assign n16295 = pi1474 & ~pi3626;
  assign n16296 = pi2797 & ~po0014;
  assign n16297 = pi1031 & ~po0015;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = pi3489 & n16225;
  assign n16300 = pi0380 & n16227;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = pi3517 & ~po0017;
  assign n16303 = n16301 & ~n16302;
  assign n16304 = n16298 & n16303;
  assign n16305 = pi3626 & ~n16304;
  assign po0105 = n16295 | n16305;
  assign n16307 = pi1602 & ~pi3626;
  assign n16308 = pi2644 & ~po0014;
  assign n16309 = pi1030 & ~po0015;
  assign n16310 = ~n16308 & ~n16309;
  assign n16311 = pi3492 & n16225;
  assign n16312 = pi0379 & n16227;
  assign n16313 = ~n16311 & ~n16312;
  assign n16314 = pi3516 & ~po0017;
  assign n16315 = n16313 & ~n16314;
  assign n16316 = n16310 & n16315;
  assign n16317 = pi3626 & ~n16316;
  assign po0106 = n16307 | n16317;
  assign n16319 = ~n16225 & ~n16227;
  assign n16320 = pi3501 & ~n16319;
  assign n16321 = pi2796 & ~po0014;
  assign n16322 = pi1029 & ~po0015;
  assign n16323 = ~n16321 & ~n16322;
  assign n16324 = ~n16320 & n16323;
  assign n16325 = pi3518 & ~po0017;
  assign n16326 = n16324 & ~n16325;
  assign n16327 = pi3626 & ~n16326;
  assign n16328 = pi0928 & ~pi3626;
  assign po0107 = n16327 | n16328;
  assign n16330 = pi3491 & ~n16319;
  assign n16331 = pi2794 & ~po0014;
  assign n16332 = pi1028 & ~po0015;
  assign n16333 = ~n16331 & ~n16332;
  assign n16334 = ~n16330 & n16333;
  assign n16335 = pi3514 & ~po0017;
  assign n16336 = n16334 & ~n16335;
  assign n16337 = pi3626 & ~n16336;
  assign n16338 = pi1066 & ~pi3626;
  assign po0108 = n16337 | n16338;
  assign n16340 = pi3494 & ~n16319;
  assign n16341 = pi2788 & ~po0014;
  assign n16342 = pi1038 & ~po0015;
  assign n16343 = ~n16341 & ~n16342;
  assign n16344 = ~n16340 & n16343;
  assign n16345 = pi3504 & ~po0017;
  assign n16346 = n16344 & ~n16345;
  assign n16347 = pi3626 & ~n16346;
  assign n16348 = pi1090 & ~pi3626;
  assign po0109 = n16347 | n16348;
  assign n16350 = pi1037 & ~po0015;
  assign n16351 = pi2953 & ~po0014;
  assign n16352 = pi3498 & ~n16319;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = ~n16350 & n16353;
  assign n16355 = pi3626 & ~n16354;
  assign n16356 = pi0930 & ~pi3626;
  assign po0110 = n16355 | n16356;
  assign n16358 = pi0688 & ~pi3626;
  assign n16359 = pi1036 & ~po0015;
  assign n16360 = ~pi2472 & po0243;
  assign n16361 = pi2408 & n16360;
  assign n16362 = ~pi2400 & ~po0242;
  assign n16363 = pi2514 & n16362;
  assign n16364 = n16361 & n16363;
  assign n16365 = ~pi2514 & n16362;
  assign n16366 = n16361 & n16365;
  assign n16367 = ~pi2514 & ~po0242;
  assign n16368 = pi2400 & n16367;
  assign n16369 = n16361 & n16368;
  assign n16370 = ~n16366 & ~n16369;
  assign n16371 = pi2400 & pi2514;
  assign n16372 = ~po0242 & ~n16371;
  assign n16373 = po0243 & n16372;
  assign n16374 = ~pi2472 & n16373;
  assign n16375 = pi3449 & ~n16374;
  assign n16376 = n16370 & ~n16375;
  assign n16377 = ~n16364 & n16376;
  assign n16378 = ~pi3680 & ~n16377;
  assign n16379 = ~pi2408 & ~po0243;
  assign n16380 = pi2400 & n16379;
  assign n16381 = ~pi2472 & po0242;
  assign n16382 = ~pi2514 & n16381;
  assign n16383 = n16380 & n16382;
  assign n16384 = ~pi2400 & n16379;
  assign n16385 = pi2514 & n16381;
  assign n16386 = n16384 & n16385;
  assign n16387 = ~n16383 & ~n16386;
  assign n16388 = pi3449 & n16382;
  assign n16389 = n16384 & n16388;
  assign n16390 = n16380 & n16385;
  assign n16391 = ~n16389 & ~n16390;
  assign n16392 = n16387 & n16391;
  assign n16393 = pi3680 & ~n16392;
  assign n16394 = ~n16378 & ~n16393;
  assign n16395 = n16227 & ~n16394;
  assign n16396 = n16225 & ~n16394;
  assign n16397 = pi2405 & ~pi3680;
  assign n16398 = pi2529 & pi3680;
  assign n16399 = ~n16397 & ~n16398;
  assign n16400 = ~po0014 & ~n16399;
  assign n16401 = ~n16396 & ~n16400;
  assign n16402 = ~n16395 & n16401;
  assign n16403 = ~n16359 & n16402;
  assign n16404 = pi3626 & ~n16403;
  assign po0111 = n16358 | n16404;
  assign n16406 = pi0929 & ~pi3626;
  assign n16407 = pi2404 & ~pi3680;
  assign n16408 = pi2405 & pi3680;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = ~po0014 & ~n16409;
  assign n16411 = pi2981 & ~po0015;
  assign n16412 = ~n16410 & ~n16411;
  assign n16413 = ~pi2408 & n16360;
  assign n16414 = n16363 & n16413;
  assign n16415 = n16365 & n16413;
  assign n16416 = ~n16366 & ~n16415;
  assign n16417 = ~n16364 & n16416;
  assign n16418 = ~n16414 & n16417;
  assign n16419 = ~pi3680 & ~n16418;
  assign n16420 = pi2408 & ~po0243;
  assign n16421 = ~pi2400 & n16420;
  assign n16422 = n16382 & n16421;
  assign n16423 = ~n16383 & ~n16422;
  assign n16424 = n16385 & n16421;
  assign n16425 = ~n16390 & ~n16424;
  assign n16426 = n16423 & n16425;
  assign n16427 = pi3680 & ~n16426;
  assign n16428 = ~n16419 & ~n16427;
  assign n16429 = ~n16319 & ~n16428;
  assign n16430 = n16412 & ~n16429;
  assign n16431 = pi3626 & ~n16430;
  assign po0112 = n16406 | n16431;
  assign n16433 = pi3101 & ~pi3626;
  assign n16434 = pi2980 & ~po0015;
  assign n16435 = n16368 & n16413;
  assign n16436 = ~n16364 & ~n16435;
  assign n16437 = ~n16369 & ~n16414;
  assign n16438 = n16436 & n16437;
  assign n16439 = ~pi3680 & ~n16438;
  assign n16440 = ~n16386 & ~n16424;
  assign n16441 = n16382 & n16420;
  assign n16442 = pi2400 & n16441;
  assign n16443 = ~n16390 & ~n16442;
  assign n16444 = n16440 & n16443;
  assign n16445 = pi3680 & ~n16444;
  assign n16446 = ~n16439 & ~n16445;
  assign n16447 = n16225 & ~n16446;
  assign n16448 = n16227 & ~n16446;
  assign n16449 = pi2473 & ~pi3680;
  assign n16450 = pi2404 & pi3680;
  assign n16451 = ~n16449 & ~n16450;
  assign n16452 = ~po0014 & ~n16451;
  assign n16453 = ~n16448 & ~n16452;
  assign n16454 = ~n16447 & n16453;
  assign n16455 = ~n16434 & n16454;
  assign n16456 = pi3626 & ~n16455;
  assign po0113 = n16433 | n16456;
  assign n16458 = pi0942 & n8405;
  assign n16459 = pi3624 & ~po0014;
  assign n16460 = po0017 & po0015;
  assign n16461 = pi3625 & ~n16460;
  assign n16462 = n16459 & ~n16461;
  assign n16463 = pi0574 & ~po3871;
  assign n16464 = ~n11016 & n16463;
  assign n16465 = pi0537 & ~po3871;
  assign n16466 = ~n11041 & n16465;
  assign n16467 = ~n16464 & ~n16466;
  assign n16468 = pi0523 & ~po3871;
  assign n16469 = ~n10988 & n16468;
  assign n16470 = n16467 & ~n16469;
  assign n16471 = ~pi2419 & ~n16470;
  assign n16472 = pi2121 & pi2419;
  assign n16473 = ~n16471 & ~n16472;
  assign n16474 = ~pi3366 & ~pi3383;
  assign n16475 = ~pi3369 & ~pi3384;
  assign n16476 = n16474 & n16475;
  assign n16477 = ~pi3379 & n16476;
  assign n16478 = ~pi3368 & ~pi3381;
  assign n16479 = ~pi3380 & n16478;
  assign n16480 = n16477 & n16479;
  assign n16481 = ~n16473 & n16480;
  assign n16482 = ~pi3380 & n16477;
  assign n16483 = pi3368 & ~pi3381;
  assign n16484 = n16482 & n16483;
  assign n16485 = ~pi3368 & n16482;
  assign n16486 = pi3381 & n16485;
  assign n16487 = ~n16484 & ~n16486;
  assign n16488 = pi3380 & n16478;
  assign n16489 = n16477 & n16488;
  assign n16490 = ~pi3379 & n16479;
  assign n16491 = ~pi3383 & n16490;
  assign n16492 = pi3366 & n16475;
  assign n16493 = n16491 & n16492;
  assign n16494 = pi3369 & n16491;
  assign n16495 = ~pi3366 & ~pi3384;
  assign n16496 = n16494 & n16495;
  assign n16497 = ~pi3369 & n16491;
  assign n16498 = ~pi3366 & pi3384;
  assign n16499 = n16497 & n16498;
  assign n16500 = n16475 & n16490;
  assign n16501 = ~pi3366 & pi3383;
  assign n16502 = n16500 & n16501;
  assign n16503 = pi3379 & n16479;
  assign n16504 = n16476 & n16503;
  assign n16505 = ~n16502 & ~n16504;
  assign n16506 = ~n16499 & n16505;
  assign n16507 = ~n16496 & n16506;
  assign n16508 = ~n16493 & n16507;
  assign n16509 = ~n16489 & n16508;
  assign n16510 = n16487 & n16509;
  assign n16511 = pi3715 & n16510;
  assign n16512 = pi3827 & n16504;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = pi3795 & n16486;
  assign n16515 = n16513 & ~n16514;
  assign n16516 = pi3747 & n16502;
  assign n16517 = n16515 & ~n16516;
  assign n16518 = pi3715 & n16499;
  assign n16519 = pi3731 & n16493;
  assign n16520 = ~n16518 & ~n16519;
  assign n16521 = pi3779 & n16484;
  assign n16522 = pi3811 & n16489;
  assign n16523 = ~n16521 & ~n16522;
  assign n16524 = pi3763 & n16496;
  assign n16525 = n16523 & ~n16524;
  assign n16526 = n16520 & n16525;
  assign n16527 = n16517 & n16526;
  assign n16528 = ~n16480 & ~n16527;
  assign n16529 = ~n16481 & ~n16528;
  assign n16530 = n16462 & ~n16529;
  assign n16531 = pi3625 & ~n16459;
  assign n16532 = ~n16460 & n16531;
  assign n16533 = ~n11181 & n16532;
  assign n16534 = ~n16530 & ~n16533;
  assign n16535 = ~n16462 & ~n16532;
  assign n16536 = pi0393 & n16535;
  assign n16537 = n16534 & ~n16536;
  assign n16538 = po0021 & ~n16537;
  assign po0114 = n16458 | n16538;
  assign n16540 = pi0927 & n8405;
  assign n16541 = ~n11833 & n16463;
  assign n16542 = ~n11858 & n16465;
  assign n16543 = ~n16541 & ~n16542;
  assign n16544 = ~n11960 & n16468;
  assign n16545 = n16543 & ~n16544;
  assign n16546 = ~pi2419 & ~n16545;
  assign n16547 = pi2120 & pi2419;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = n16480 & ~n16548;
  assign n16550 = pi3716 & n16510;
  assign n16551 = pi3828 & n16504;
  assign n16552 = ~n16550 & ~n16551;
  assign n16553 = pi3796 & n16486;
  assign n16554 = n16552 & ~n16553;
  assign n16555 = pi3748 & n16502;
  assign n16556 = n16554 & ~n16555;
  assign n16557 = pi3716 & n16499;
  assign n16558 = pi3732 & n16493;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = pi3780 & n16484;
  assign n16561 = pi3812 & n16489;
  assign n16562 = ~n16560 & ~n16561;
  assign n16563 = pi3764 & n16496;
  assign n16564 = n16562 & ~n16563;
  assign n16565 = n16559 & n16564;
  assign n16566 = n16556 & n16565;
  assign n16567 = ~n16480 & ~n16566;
  assign n16568 = ~n16549 & ~n16567;
  assign n16569 = n16462 & ~n16568;
  assign n16570 = ~n12061 & n16532;
  assign n16571 = ~n16569 & ~n16570;
  assign n16572 = pi0390 & n16535;
  assign n16573 = n16571 & ~n16572;
  assign n16574 = po0021 & ~n16573;
  assign po0115 = n16540 | n16574;
  assign n16576 = pi0926 & n8405;
  assign n16577 = ~n14887 & n16463;
  assign n16578 = ~n14922 & n16468;
  assign n16579 = ~n16577 & ~n16578;
  assign n16580 = ~n15014 & n16465;
  assign n16581 = n16579 & ~n16580;
  assign n16582 = ~pi2419 & ~n16581;
  assign n16583 = pi2119 & pi2419;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = n16480 & ~n16584;
  assign n16586 = pi3717 & n16510;
  assign n16587 = pi3829 & n16504;
  assign n16588 = ~n16586 & ~n16587;
  assign n16589 = pi3797 & n16486;
  assign n16590 = n16588 & ~n16589;
  assign n16591 = pi3749 & n16502;
  assign n16592 = n16590 & ~n16591;
  assign n16593 = pi3717 & n16499;
  assign n16594 = pi3733 & n16493;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = pi3765 & n16496;
  assign n16597 = pi3781 & n16484;
  assign n16598 = ~n16596 & ~n16597;
  assign n16599 = pi3813 & n16489;
  assign n16600 = n16598 & ~n16599;
  assign n16601 = n16595 & n16600;
  assign n16602 = n16592 & n16601;
  assign n16603 = ~n16480 & ~n16602;
  assign n16604 = ~n16585 & ~n16603;
  assign n16605 = n16462 & ~n16604;
  assign n16606 = ~n15115 & n16532;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = pi0389 & n16535;
  assign n16609 = n16607 & ~n16608;
  assign n16610 = po0021 & ~n16609;
  assign po0116 = n16576 | n16610;
  assign n16612 = pi0925 & n8405;
  assign n16613 = ~n14654 & n16463;
  assign n16614 = ~n14626 & n16465;
  assign n16615 = ~n16613 & ~n16614;
  assign n16616 = ~n14689 & n16468;
  assign n16617 = n16615 & ~n16616;
  assign n16618 = ~pi2419 & ~n16617;
  assign n16619 = pi2118 & pi2419;
  assign n16620 = ~n16618 & ~n16619;
  assign n16621 = n16480 & ~n16620;
  assign n16622 = pi3718 & n16510;
  assign n16623 = pi3830 & n16504;
  assign n16624 = ~n16622 & ~n16623;
  assign n16625 = pi3798 & n16486;
  assign n16626 = n16624 & ~n16625;
  assign n16627 = pi3750 & n16502;
  assign n16628 = n16626 & ~n16627;
  assign n16629 = pi3718 & n16499;
  assign n16630 = pi3734 & n16493;
  assign n16631 = ~n16629 & ~n16630;
  assign n16632 = pi3782 & n16484;
  assign n16633 = pi3814 & n16489;
  assign n16634 = ~n16632 & ~n16633;
  assign n16635 = pi3766 & n16496;
  assign n16636 = n16634 & ~n16635;
  assign n16637 = n16631 & n16636;
  assign n16638 = n16628 & n16637;
  assign n16639 = ~n16480 & ~n16638;
  assign n16640 = ~n16621 & ~n16639;
  assign n16641 = n16462 & ~n16640;
  assign n16642 = ~n14816 & n16532;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = pi0388 & n16535;
  assign n16645 = n16643 & ~n16644;
  assign n16646 = po0021 & ~n16645;
  assign po0117 = n16612 | n16646;
  assign n16648 = pi0943 & n8405;
  assign n16649 = ~n12225 & n16465;
  assign n16650 = ~n12253 & n16463;
  assign n16651 = ~n16649 & ~n16650;
  assign n16652 = ~n12288 & n16468;
  assign n16653 = n16651 & ~n16652;
  assign n16654 = ~pi2419 & ~n16653;
  assign n16655 = pi2117 & pi2419;
  assign n16656 = ~n16654 & ~n16655;
  assign n16657 = n16480 & ~n16656;
  assign n16658 = pi3719 & n16510;
  assign n16659 = pi3831 & n16504;
  assign n16660 = ~n16658 & ~n16659;
  assign n16661 = pi3799 & n16486;
  assign n16662 = n16660 & ~n16661;
  assign n16663 = pi3751 & n16502;
  assign n16664 = n16662 & ~n16663;
  assign n16665 = pi3719 & n16499;
  assign n16666 = pi3735 & n16493;
  assign n16667 = ~n16665 & ~n16666;
  assign n16668 = pi3783 & n16484;
  assign n16669 = pi3815 & n16489;
  assign n16670 = ~n16668 & ~n16669;
  assign n16671 = pi3767 & n16496;
  assign n16672 = n16670 & ~n16671;
  assign n16673 = n16667 & n16672;
  assign n16674 = n16664 & n16673;
  assign n16675 = ~n16480 & ~n16674;
  assign n16676 = ~n16657 & ~n16675;
  assign n16677 = n16462 & ~n16676;
  assign n16678 = ~n12415 & n16532;
  assign n16679 = ~n16677 & ~n16678;
  assign n16680 = pi0387 & n16535;
  assign n16681 = n16679 & ~n16680;
  assign n16682 = po0021 & ~n16681;
  assign po0118 = n16648 | n16682;
  assign n16684 = pi0924 & n8405;
  assign n16685 = ~n13798 & n16465;
  assign n16686 = ~n13826 & n16463;
  assign n16687 = ~n16685 & ~n16686;
  assign n16688 = ~n13861 & n16468;
  assign n16689 = n16687 & ~n16688;
  assign n16690 = ~pi2419 & ~n16689;
  assign n16691 = pi2078 & pi2419;
  assign n16692 = ~n16690 & ~n16691;
  assign n16693 = n16480 & ~n16692;
  assign n16694 = pi3720 & n16510;
  assign n16695 = pi3832 & n16504;
  assign n16696 = ~n16694 & ~n16695;
  assign n16697 = pi3800 & n16486;
  assign n16698 = n16696 & ~n16697;
  assign n16699 = pi3752 & n16502;
  assign n16700 = n16698 & ~n16699;
  assign n16701 = pi3720 & n16499;
  assign n16702 = pi3736 & n16493;
  assign n16703 = ~n16701 & ~n16702;
  assign n16704 = pi3784 & n16484;
  assign n16705 = pi3816 & n16489;
  assign n16706 = ~n16704 & ~n16705;
  assign n16707 = pi3768 & n16496;
  assign n16708 = n16706 & ~n16707;
  assign n16709 = n16703 & n16708;
  assign n16710 = n16700 & n16709;
  assign n16711 = ~n16480 & ~n16710;
  assign n16712 = ~n16693 & ~n16711;
  assign n16713 = n16462 & ~n16712;
  assign n16714 = ~n13988 & n16532;
  assign n16715 = ~n16713 & ~n16714;
  assign n16716 = pi0386 & n16535;
  assign n16717 = n16715 & ~n16716;
  assign n16718 = po0021 & ~n16717;
  assign po0119 = n16684 | n16718;
  assign n16720 = pi0923 & n8405;
  assign n16721 = ~n13301 & n16465;
  assign n16722 = ~n13178 & n16463;
  assign n16723 = ~n16721 & ~n16722;
  assign n16724 = ~n13213 & n16468;
  assign n16725 = n16723 & ~n16724;
  assign n16726 = ~pi2419 & ~n16725;
  assign n16727 = pi2116 & pi2419;
  assign n16728 = ~n16726 & ~n16727;
  assign n16729 = n16480 & ~n16728;
  assign n16730 = pi3721 & n16510;
  assign n16731 = pi3833 & n16504;
  assign n16732 = ~n16730 & ~n16731;
  assign n16733 = pi3801 & n16486;
  assign n16734 = n16732 & ~n16733;
  assign n16735 = pi3753 & n16502;
  assign n16736 = n16734 & ~n16735;
  assign n16737 = pi3721 & n16499;
  assign n16738 = pi3737 & n16493;
  assign n16739 = ~n16737 & ~n16738;
  assign n16740 = pi3785 & n16484;
  assign n16741 = pi3817 & n16489;
  assign n16742 = ~n16740 & ~n16741;
  assign n16743 = pi3769 & n16496;
  assign n16744 = n16742 & ~n16743;
  assign n16745 = n16739 & n16744;
  assign n16746 = n16736 & n16745;
  assign n16747 = ~n16480 & ~n16746;
  assign n16748 = ~n16729 & ~n16747;
  assign n16749 = n16462 & ~n16748;
  assign n16750 = ~n13398 & n16532;
  assign n16751 = ~n16749 & ~n16750;
  assign n16752 = pi0385 & n16535;
  assign n16753 = n16751 & ~n16752;
  assign n16754 = po0021 & ~n16753;
  assign po0120 = n16720 | n16754;
  assign n16756 = pi0922 & n8405;
  assign n16757 = ~n12967 & n16465;
  assign n16758 = ~n12994 & n16463;
  assign n16759 = ~n16757 & ~n16758;
  assign n16760 = ~n12949 & n16468;
  assign n16761 = n16759 & ~n16760;
  assign n16762 = ~pi2419 & ~n16761;
  assign n16763 = pi2115 & pi2419;
  assign n16764 = ~n16762 & ~n16763;
  assign n16765 = n16480 & ~n16764;
  assign n16766 = pi3722 & n16510;
  assign n16767 = pi3834 & n16504;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = pi3802 & n16486;
  assign n16770 = n16768 & ~n16769;
  assign n16771 = pi3754 & n16502;
  assign n16772 = n16770 & ~n16771;
  assign n16773 = pi3722 & n16499;
  assign n16774 = pi3738 & n16493;
  assign n16775 = ~n16773 & ~n16774;
  assign n16776 = pi3786 & n16484;
  assign n16777 = pi3818 & n16489;
  assign n16778 = ~n16776 & ~n16777;
  assign n16779 = pi3770 & n16496;
  assign n16780 = n16778 & ~n16779;
  assign n16781 = n16775 & n16780;
  assign n16782 = n16772 & n16781;
  assign n16783 = ~n16480 & ~n16782;
  assign n16784 = ~n16765 & ~n16783;
  assign n16785 = n16462 & ~n16784;
  assign n16786 = ~n13121 & n16532;
  assign n16787 = ~n16785 & ~n16786;
  assign n16788 = pi0384 & n16535;
  assign n16789 = n16787 & ~n16788;
  assign n16790 = po0021 & ~n16789;
  assign po0121 = n16756 | n16790;
  assign n16792 = ~n13561 & n16465;
  assign n16793 = ~n13543 & n16468;
  assign n16794 = ~n16792 & ~n16793;
  assign n16795 = ~n13586 & n16463;
  assign n16796 = n16794 & ~n16795;
  assign n16797 = ~pi2419 & ~n16796;
  assign n16798 = pi2414 & pi2419;
  assign n16799 = ~n16797 & ~n16798;
  assign n16800 = n16480 & ~n16799;
  assign n16801 = pi3723 & n16510;
  assign n16802 = pi3835 & n16504;
  assign n16803 = ~n16801 & ~n16802;
  assign n16804 = pi3803 & n16486;
  assign n16805 = n16803 & ~n16804;
  assign n16806 = pi3755 & n16502;
  assign n16807 = n16805 & ~n16806;
  assign n16808 = pi3723 & n16499;
  assign n16809 = pi3739 & n16493;
  assign n16810 = ~n16808 & ~n16809;
  assign n16811 = pi3787 & n16484;
  assign n16812 = pi3819 & n16489;
  assign n16813 = ~n16811 & ~n16812;
  assign n16814 = pi3771 & n16496;
  assign n16815 = n16813 & ~n16814;
  assign n16816 = n16810 & n16815;
  assign n16817 = n16807 & n16816;
  assign n16818 = ~n16480 & ~n16817;
  assign n16819 = ~n16800 & ~n16818;
  assign n16820 = n16462 & ~n16819;
  assign n16821 = ~n13701 & n16532;
  assign n16822 = ~n16820 & ~n16821;
  assign n16823 = pi0383 & n16535;
  assign n16824 = n16822 & ~n16823;
  assign n16825 = po0021 & ~n16824;
  assign n16826 = pi3107 & ~pi3626;
  assign po0122 = n16825 | n16826;
  assign n16828 = ~n12525 & n16465;
  assign n16829 = ~n12636 & n16468;
  assign n16830 = ~n16828 & ~n16829;
  assign n16831 = ~n12550 & n16463;
  assign n16832 = n16830 & ~n16831;
  assign n16833 = ~pi2419 & ~n16832;
  assign n16834 = pi2418 & pi2419;
  assign n16835 = ~n16833 & ~n16834;
  assign n16836 = n16480 & ~n16835;
  assign n16837 = pi3724 & n16510;
  assign n16838 = pi3836 & n16504;
  assign n16839 = ~n16837 & ~n16838;
  assign n16840 = pi3804 & n16486;
  assign n16841 = n16839 & ~n16840;
  assign n16842 = pi3756 & n16502;
  assign n16843 = n16841 & ~n16842;
  assign n16844 = pi3724 & n16499;
  assign n16845 = pi3740 & n16493;
  assign n16846 = ~n16844 & ~n16845;
  assign n16847 = pi3772 & n16496;
  assign n16848 = pi3820 & n16489;
  assign n16849 = ~n16847 & ~n16848;
  assign n16850 = pi3788 & n16484;
  assign n16851 = n16849 & ~n16850;
  assign n16852 = n16846 & n16851;
  assign n16853 = n16843 & n16852;
  assign n16854 = ~n16480 & ~n16853;
  assign n16855 = ~n16836 & ~n16854;
  assign n16856 = n16462 & ~n16855;
  assign n16857 = ~n12726 & n16532;
  assign n16858 = ~n16856 & ~n16857;
  assign n16859 = pi0382 & n16535;
  assign n16860 = n16858 & ~n16859;
  assign n16861 = po0021 & ~n16860;
  assign n16862 = pi3063 & ~pi3626;
  assign po0123 = n16861 | n16862;
  assign n16864 = ~n14264 & n16465;
  assign n16865 = ~n14246 & n16468;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = ~n14289 & n16463;
  assign n16868 = n16866 & ~n16867;
  assign n16869 = ~pi2419 & ~n16868;
  assign n16870 = pi1951 & pi2419;
  assign n16871 = ~n16869 & ~n16870;
  assign n16872 = n16480 & ~n16871;
  assign n16873 = pi3725 & n16510;
  assign n16874 = pi3837 & n16504;
  assign n16875 = ~n16873 & ~n16874;
  assign n16876 = pi3805 & n16486;
  assign n16877 = n16875 & ~n16876;
  assign n16878 = pi3757 & n16502;
  assign n16879 = n16877 & ~n16878;
  assign n16880 = pi3725 & n16499;
  assign n16881 = pi3741 & n16493;
  assign n16882 = ~n16880 & ~n16881;
  assign n16883 = pi3773 & n16496;
  assign n16884 = pi3821 & n16489;
  assign n16885 = ~n16883 & ~n16884;
  assign n16886 = pi3789 & n16484;
  assign n16887 = n16885 & ~n16886;
  assign n16888 = n16882 & n16887;
  assign n16889 = n16879 & n16888;
  assign n16890 = ~n16480 & ~n16889;
  assign n16891 = ~n16872 & ~n16890;
  assign n16892 = n16462 & ~n16891;
  assign n16893 = ~n14403 & n16532;
  assign n16894 = ~n16892 & ~n16893;
  assign n16895 = pi0392 & n16535;
  assign n16896 = n16894 & ~n16895;
  assign n16897 = po0021 & ~n16896;
  assign n16898 = pi3091 & ~pi3626;
  assign po0124 = n16897 | n16898;
  assign n16900 = ~n15286 & n16465;
  assign n16901 = ~n15268 & n16468;
  assign n16902 = ~n16900 & ~n16901;
  assign n16903 = ~n15311 & n16463;
  assign n16904 = n16902 & ~n16903;
  assign n16905 = ~pi2419 & ~n16904;
  assign n16906 = pi1950 & pi2419;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = n16480 & ~n16907;
  assign n16909 = pi3726 & n16510;
  assign n16910 = pi3838 & n16504;
  assign n16911 = ~n16909 & ~n16910;
  assign n16912 = pi3806 & n16486;
  assign n16913 = n16911 & ~n16912;
  assign n16914 = pi3758 & n16502;
  assign n16915 = n16913 & ~n16914;
  assign n16916 = pi3726 & n16499;
  assign n16917 = pi3742 & n16493;
  assign n16918 = ~n16916 & ~n16917;
  assign n16919 = pi3774 & n16496;
  assign n16920 = pi3790 & n16484;
  assign n16921 = ~n16919 & ~n16920;
  assign n16922 = pi3822 & n16489;
  assign n16923 = n16921 & ~n16922;
  assign n16924 = n16918 & n16923;
  assign n16925 = n16915 & n16924;
  assign n16926 = ~n16480 & ~n16925;
  assign n16927 = ~n16908 & ~n16926;
  assign n16928 = n16462 & ~n16927;
  assign n16929 = ~n15426 & n16532;
  assign n16930 = ~n16928 & ~n16929;
  assign n16931 = pi0391 & n16535;
  assign n16932 = n16930 & ~n16931;
  assign n16933 = po0021 & ~n16932;
  assign n16934 = pi2989 & ~pi3626;
  assign po0125 = n16933 | n16934;
  assign n16936 = ~n10465 & n16465;
  assign n16937 = ~n10447 & n16468;
  assign n16938 = ~n16936 & ~n16937;
  assign n16939 = ~n10490 & n16463;
  assign n16940 = n16938 & ~n16939;
  assign n16941 = ~pi2419 & ~n16940;
  assign n16942 = pi1949 & pi2419;
  assign n16943 = ~n16941 & ~n16942;
  assign n16944 = n16480 & ~n16943;
  assign n16945 = pi3727 & n16510;
  assign n16946 = pi3839 & n16504;
  assign n16947 = ~n16945 & ~n16946;
  assign n16948 = pi3807 & n16486;
  assign n16949 = n16947 & ~n16948;
  assign n16950 = pi3759 & n16502;
  assign n16951 = n16949 & ~n16950;
  assign n16952 = pi3727 & n16499;
  assign n16953 = pi3743 & n16493;
  assign n16954 = ~n16952 & ~n16953;
  assign n16955 = pi3775 & n16496;
  assign n16956 = pi3791 & n16484;
  assign n16957 = ~n16955 & ~n16956;
  assign n16958 = pi3823 & n16489;
  assign n16959 = n16957 & ~n16958;
  assign n16960 = n16954 & n16959;
  assign n16961 = n16951 & n16960;
  assign n16962 = ~n16480 & ~n16961;
  assign n16963 = ~n16944 & ~n16962;
  assign n16964 = n16462 & ~n16963;
  assign n16965 = ~n10608 & n16532;
  assign n16966 = ~n16964 & ~n16965;
  assign n16967 = pi0381 & n16535;
  assign n16968 = n16966 & ~n16967;
  assign n16969 = po0021 & ~n16968;
  assign n16970 = pi2988 & ~pi3626;
  assign po0126 = n16969 | n16970;
  assign n16972 = ~n9547 & n16465;
  assign n16973 = ~n9520 & n16468;
  assign n16974 = ~n16972 & ~n16973;
  assign n16975 = ~n9573 & n16463;
  assign n16976 = n16974 & ~n16975;
  assign n16977 = ~pi2419 & ~n16976;
  assign n16978 = pi1948 & pi2419;
  assign n16979 = ~n16977 & ~n16978;
  assign n16980 = n16480 & ~n16979;
  assign n16981 = pi3728 & n16510;
  assign n16982 = pi3840 & n16504;
  assign n16983 = ~n16981 & ~n16982;
  assign n16984 = pi3808 & n16486;
  assign n16985 = n16983 & ~n16984;
  assign n16986 = pi3760 & n16502;
  assign n16987 = n16985 & ~n16986;
  assign n16988 = pi3728 & n16499;
  assign n16989 = pi3744 & n16493;
  assign n16990 = ~n16988 & ~n16989;
  assign n16991 = pi3792 & n16484;
  assign n16992 = pi3824 & n16489;
  assign n16993 = ~n16991 & ~n16992;
  assign n16994 = pi3776 & n16496;
  assign n16995 = n16993 & ~n16994;
  assign n16996 = n16990 & n16995;
  assign n16997 = n16987 & n16996;
  assign n16998 = ~n16480 & ~n16997;
  assign n16999 = ~n16980 & ~n16998;
  assign n17000 = n16462 & ~n16999;
  assign n17001 = ~n9825 & n16532;
  assign n17002 = ~n17000 & ~n17001;
  assign n17003 = pi0378 & n16535;
  assign n17004 = n17002 & ~n17003;
  assign n17005 = po0021 & ~n17004;
  assign n17006 = pi2987 & ~pi3626;
  assign po0127 = n17005 | n17006;
  assign n17008 = ~pi0979 & pi2851;
  assign n17009 = pi0979 & pi2134;
  assign n17010 = ~n17008 & ~n17009;
  assign n17011 = pi0717 & ~n17010;
  assign n17012 = pi0298 & ~pi0979;
  assign n17013 = pi0297 & pi0979;
  assign n17014 = ~n17012 & ~n17013;
  assign n17015 = pi0716 & ~n17014;
  assign n17016 = pi0320 & ~pi0979;
  assign n17017 = pi0318 & pi0979;
  assign n17018 = ~n17016 & ~n17017;
  assign n17019 = pi0761 & ~n17018;
  assign n17020 = ~n17015 & ~n17019;
  assign n17021 = ~n9535 & n17020;
  assign n17022 = ~n9531 & n17021;
  assign n17023 = ~n17011 & n17022;
  assign n17024 = n16465 & ~n17023;
  assign n17025 = pi0979 & pi2153;
  assign n17026 = ~pi0979 & pi2925;
  assign n17027 = ~n17025 & ~n17026;
  assign n17028 = pi0767 & ~n17027;
  assign n17029 = ~pi0979 & pi2160;
  assign n17030 = pi0979 & pi1791;
  assign n17031 = ~n17029 & ~n17030;
  assign n17032 = pi0768 & ~n17031;
  assign n17033 = ~n17028 & ~n17032;
  assign n17034 = pi0979 & pi2171;
  assign n17035 = ~pi0979 & pi2804;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = pi0836 & ~n17036;
  assign n17038 = ~pi0979 & pi2947;
  assign n17039 = pi0979 & pi2187;
  assign n17040 = ~n17038 & ~n17039;
  assign n17041 = pi0837 & ~n17040;
  assign n17042 = ~n17037 & ~n17041;
  assign n17043 = pi0177 & ~pi0979;
  assign n17044 = pi0162 & pi0979;
  assign n17045 = ~n17043 & ~n17044;
  assign n17046 = pi0838 & ~n17045;
  assign n17047 = n17042 & ~n17046;
  assign n17048 = n17033 & n17047;
  assign n17049 = n16463 & ~n17048;
  assign n17050 = ~n17024 & ~n17049;
  assign n17051 = ~pi0979 & pi2868;
  assign n17052 = pi0979 & pi2861;
  assign n17053 = ~n17051 & ~n17052;
  assign n17054 = pi0763 & ~n17053;
  assign n17055 = ~pi0979 & pi2878;
  assign n17056 = pi0979 & pi2869;
  assign n17057 = ~n17055 & ~n17056;
  assign n17058 = pi0764 & ~n17057;
  assign n17059 = ~n17054 & ~n17058;
  assign n17060 = ~pi0979 & pi2639;
  assign n17061 = pi0979 & pi3172;
  assign n17062 = ~n17060 & ~n17061;
  assign n17063 = pi0765 & ~n17062;
  assign n17064 = ~pi0979 & pi2914;
  assign n17065 = pi0979 & pi3183;
  assign n17066 = ~n17064 & ~n17065;
  assign n17067 = pi0766 & ~n17066;
  assign n17068 = ~n17063 & ~n17067;
  assign n17069 = pi0119 & ~pi0979;
  assign n17070 = pi0115 & pi0979;
  assign n17071 = ~n17069 & ~n17070;
  assign n17072 = pi0720 & ~n17071;
  assign n17073 = pi0212 & ~pi0979;
  assign n17074 = pi0211 & pi0979;
  assign n17075 = ~n17073 & ~n17074;
  assign n17076 = pi0721 & ~n17075;
  assign n17077 = ~n17072 & ~n17076;
  assign n17078 = n17068 & n17077;
  assign n17079 = ~n9499 & n17078;
  assign n17080 = n17059 & n17079;
  assign n17081 = n16468 & ~n17080;
  assign n17082 = n17050 & ~n17081;
  assign n17083 = ~pi2419 & ~n17082;
  assign n17084 = pi1947 & pi2419;
  assign n17085 = ~n17083 & ~n17084;
  assign n17086 = n16480 & ~n17085;
  assign n17087 = pi3729 & n16510;
  assign n17088 = pi3841 & n16504;
  assign n17089 = ~n17087 & ~n17088;
  assign n17090 = pi3809 & n16486;
  assign n17091 = n17089 & ~n17090;
  assign n17092 = pi3761 & n16502;
  assign n17093 = n17091 & ~n17092;
  assign n17094 = pi3729 & n16499;
  assign n17095 = pi3745 & n16493;
  assign n17096 = ~n17094 & ~n17095;
  assign n17097 = pi3793 & n16484;
  assign n17098 = pi3825 & n16489;
  assign n17099 = ~n17097 & ~n17098;
  assign n17100 = pi3777 & n16496;
  assign n17101 = n17099 & ~n17100;
  assign n17102 = n17096 & n17101;
  assign n17103 = n17093 & n17102;
  assign n17104 = ~n16480 & ~n17103;
  assign n17105 = ~n17086 & ~n17104;
  assign n17106 = n16462 & ~n17105;
  assign n17107 = n9486 & ~n17080;
  assign n17108 = n9523 & ~n17023;
  assign n17109 = n9549 & ~n17048;
  assign n17110 = ~n17108 & ~n17109;
  assign n17111 = pi3233 & pi3396;
  assign n17112 = pi0377 & pi1057;
  assign n17113 = ~n17111 & ~n17112;
  assign n17114 = n9475 & ~n17113;
  assign n17115 = pi0607 & pi1336;
  assign n17116 = pi1333 & pi1866;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = pi1332 & pi2577;
  assign n17119 = pi1335 & pi2592;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = n17117 & n17120;
  assign n17122 = n9726 & ~n17121;
  assign n17123 = pi2123 & n9628;
  assign n17124 = pi1102 & n9631;
  assign n17125 = ~n17123 & ~n17124;
  assign n17126 = pi1929 & n9622;
  assign n17127 = n17125 & ~n17126;
  assign n17128 = pi1854 & n9657;
  assign n17129 = pi1759 & n9659;
  assign n17130 = ~n17128 & ~n17129;
  assign n17131 = pi1422 & n9710;
  assign n17132 = pi1781 & n9712;
  assign n17133 = ~n17131 & ~n17132;
  assign n17134 = pi3680 & n11102;
  assign n17135 = pi2987 & n9647;
  assign n17136 = ~n17134 & ~n17135;
  assign n17137 = n17133 & n17136;
  assign n17138 = pi0896 & n9707;
  assign n17139 = pi0887 & n9715;
  assign n17140 = pi1869 & n9718;
  assign n17141 = ~n17139 & ~n17140;
  assign n17142 = pi0959 & n9614;
  assign n17143 = pi1904 & n9618;
  assign n17144 = ~n17142 & ~n17143;
  assign n17145 = pi0970 & n9687;
  assign n17146 = pi1917 & n9691;
  assign n17147 = ~n17145 & ~n17146;
  assign n17148 = n17144 & n17147;
  assign n17149 = ~n10557 & n17148;
  assign n17150 = pi1792 & n9698;
  assign n17151 = n17149 & ~n17150;
  assign n17152 = ~n10564 & n17151;
  assign n17153 = n17141 & n17152;
  assign n17154 = ~n17138 & n17153;
  assign n17155 = n17137 & n17154;
  assign n17156 = pi1723 & n9679;
  assign n17157 = pi0246 & n9682;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = n17155 & n17158;
  assign n17160 = n17130 & n17159;
  assign n17161 = n17127 & n17160;
  assign n17162 = pi1934 & ~n17161;
  assign n17163 = ~n17122 & ~n17162;
  assign n17164 = ~n17114 & n17163;
  assign n17165 = n17110 & n17164;
  assign n17166 = ~n17107 & n17165;
  assign n17167 = n9577 & ~n9594;
  assign n17168 = n9736 & ~n9753;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = n9475 & n9479;
  assign n17171 = n17169 & ~n17170;
  assign n17172 = n17166 & n17171;
  assign n17173 = pi3314 & po3871;
  assign n17174 = n17172 & ~n17173;
  assign n17175 = ~pi1787 & ~n17174;
  assign n17176 = pi1787 & pi2832;
  assign n17177 = ~n17175 & ~n17176;
  assign n17178 = n9472 & ~n17177;
  assign n17179 = pi3873 & n9804;
  assign n17180 = pi3889 & n9774;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = pi3857 & n9802;
  assign n17183 = pi3921 & n9781;
  assign n17184 = pi3905 & n9771;
  assign n17185 = ~n17183 & ~n17184;
  assign n17186 = pi3953 & n9791;
  assign n17187 = pi3937 & n9788;
  assign n17188 = ~n17186 & ~n17187;
  assign n17189 = n17185 & n17188;
  assign n17190 = ~n17182 & n17189;
  assign n17191 = n17181 & n17190;
  assign n17192 = pi3873 & n9799;
  assign n17193 = n17191 & ~n17192;
  assign n17194 = pi3985 & n9783;
  assign n17195 = pi3969 & n9793;
  assign n17196 = ~n17194 & ~n17195;
  assign n17197 = n17193 & n17196;
  assign n17198 = ~n9472 & ~n17197;
  assign n17199 = ~n17178 & ~n17198;
  assign n17200 = n16532 & ~n17199;
  assign n17201 = ~n17106 & ~n17200;
  assign n17202 = pi0377 & n16535;
  assign n17203 = n17201 & ~n17202;
  assign n17204 = po0021 & ~n17203;
  assign n17205 = pi3097 & ~pi3626;
  assign po0128 = n17204 | n17205;
  assign n17207 = pi3233 & pi3393;
  assign n17208 = n9475 & n17207;
  assign n17209 = n17169 & ~n17208;
  assign n17210 = ~n17170 & n17209;
  assign n17211 = ~pi0979 & pi2850;
  assign n17212 = pi0979 & pi2133;
  assign n17213 = ~n17211 & ~n17212;
  assign n17214 = pi0717 & ~n17213;
  assign n17215 = pi0286 & ~pi0979;
  assign n17216 = pi0285 & pi0979;
  assign n17217 = ~n17215 & ~n17216;
  assign n17218 = pi0716 & ~n17217;
  assign n17219 = pi0254 & ~pi0979;
  assign n17220 = pi0251 & pi0979;
  assign n17221 = ~n17219 & ~n17220;
  assign n17222 = pi0761 & ~n17221;
  assign n17223 = ~n17218 & ~n17222;
  assign n17224 = ~n9535 & n17223;
  assign n17225 = ~n9531 & n17224;
  assign n17226 = ~n17214 & n17225;
  assign n17227 = n9523 & ~n17226;
  assign n17228 = pi0979 & pi2152;
  assign n17229 = ~pi0979 & pi2924;
  assign n17230 = ~n17228 & ~n17229;
  assign n17231 = pi0767 & ~n17230;
  assign n17232 = ~pi0979 & pi2428;
  assign n17233 = pi0979 & pi1963;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = pi0768 & ~n17234;
  assign n17236 = ~n17231 & ~n17235;
  assign n17237 = pi0979 & pi2170;
  assign n17238 = ~pi0979 & pi2805;
  assign n17239 = ~n17237 & ~n17238;
  assign n17240 = pi0836 & ~n17239;
  assign n17241 = ~pi0979 & pi2946;
  assign n17242 = pi0979 & pi2186;
  assign n17243 = ~n17241 & ~n17242;
  assign n17244 = pi0837 & ~n17243;
  assign n17245 = ~n17240 & ~n17244;
  assign n17246 = pi0151 & ~pi0979;
  assign n17247 = pi0150 & pi0979;
  assign n17248 = ~n17246 & ~n17247;
  assign n17249 = pi0838 & ~n17248;
  assign n17250 = n17245 & ~n17249;
  assign n17251 = n17236 & n17250;
  assign n17252 = n9549 & ~n17251;
  assign n17253 = ~n17227 & ~n17252;
  assign n17254 = pi1057 & n9475;
  assign n17255 = pi0376 & n17254;
  assign n17256 = pi0605 & pi1336;
  assign n17257 = pi1335 & pi2591;
  assign n17258 = ~n17256 & ~n17257;
  assign n17259 = pi1332 & pi2576;
  assign n17260 = pi1333 & pi1897;
  assign n17261 = ~n17259 & ~n17260;
  assign n17262 = n17258 & n17261;
  assign n17263 = n9726 & ~n17262;
  assign n17264 = pi2109 & n9628;
  assign n17265 = pi1768 & n9657;
  assign n17266 = ~n17264 & ~n17265;
  assign n17267 = pi1426 & n11133;
  assign n17268 = pi0223 & n9682;
  assign n17269 = ~n17267 & ~n17268;
  assign n17270 = pi1722 & n9679;
  assign n17271 = n17269 & ~n17270;
  assign n17272 = pi1928 & n9622;
  assign n17273 = n17271 & ~n17272;
  assign n17274 = pi1024 & n9631;
  assign n17275 = pi1758 & n9659;
  assign n17276 = ~n17274 & ~n17275;
  assign n17277 = n17273 & n17276;
  assign n17278 = n17266 & n17277;
  assign n17279 = pi1934 & ~n17278;
  assign n17280 = ~n17263 & ~n17279;
  assign n17281 = pi2385 & n11102;
  assign n17282 = pi3097 & n9647;
  assign n17283 = ~n17281 & ~n17282;
  assign n17284 = pi1934 & ~n17283;
  assign n17285 = pi0895 & n9707;
  assign n17286 = pi0893 & n9702;
  assign n17287 = ~n17285 & ~n17286;
  assign n17288 = pi1835 & n9698;
  assign n17289 = n17287 & ~n17288;
  assign n17290 = pi0886 & n9715;
  assign n17291 = pi1889 & n9718;
  assign n17292 = ~n17290 & ~n17291;
  assign n17293 = pi0958 & n9614;
  assign n17294 = pi1903 & n9618;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = pi0799 & n9607;
  assign n17297 = n17295 & ~n17296;
  assign n17298 = pi0969 & n9687;
  assign n17299 = pi1908 & n9691;
  assign n17300 = ~n17298 & ~n17299;
  assign n17301 = n17297 & n17300;
  assign n17302 = n17292 & n17301;
  assign n17303 = n17289 & n17302;
  assign n17304 = pi1934 & ~n17303;
  assign n17305 = ~n17284 & ~n17304;
  assign n17306 = n17280 & n17305;
  assign n17307 = ~pi0979 & pi2867;
  assign n17308 = pi0979 & pi3158;
  assign n17309 = ~n17307 & ~n17308;
  assign n17310 = pi0763 & ~n17309;
  assign n17311 = ~pi0979 & pi2877;
  assign n17312 = pi0979 & pi3140;
  assign n17313 = ~n17311 & ~n17312;
  assign n17314 = pi0764 & ~n17313;
  assign n17315 = ~n17310 & ~n17314;
  assign n17316 = ~pi0979 & pi2638;
  assign n17317 = pi0979 & pi3171;
  assign n17318 = ~n17316 & ~n17317;
  assign n17319 = pi0765 & ~n17318;
  assign n17320 = ~pi0979 & pi2894;
  assign n17321 = pi0979 & pi3182;
  assign n17322 = ~n17320 & ~n17321;
  assign n17323 = pi0766 & ~n17322;
  assign n17324 = ~n17319 & ~n17323;
  assign n17325 = pi0059 & ~pi0979;
  assign n17326 = pi0058 & pi0979;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = pi0720 & ~n17327;
  assign n17329 = pi0193 & ~pi0979;
  assign n17330 = pi0192 & pi0979;
  assign n17331 = ~n17329 & ~n17330;
  assign n17332 = pi0721 & ~n17331;
  assign n17333 = ~n17328 & ~n17332;
  assign n17334 = n17324 & n17333;
  assign n17335 = ~n9499 & n17334;
  assign n17336 = n17315 & n17335;
  assign n17337 = n9486 & ~n17336;
  assign n17338 = n17306 & ~n17337;
  assign n17339 = ~n17255 & n17338;
  assign n17340 = n17253 & n17339;
  assign n17341 = n17210 & n17340;
  assign n17342 = pi3313 & po3871;
  assign n17343 = n17341 & ~n17342;
  assign n17344 = ~pi1787 & ~n17343;
  assign n17345 = pi1787 & pi2816;
  assign n17346 = ~n17344 & ~n17345;
  assign n17347 = n9472 & ~n17346;
  assign n17348 = pi3874 & n9804;
  assign n17349 = pi3890 & n9774;
  assign n17350 = ~n17348 & ~n17349;
  assign n17351 = pi3858 & n9802;
  assign n17352 = pi3922 & n9781;
  assign n17353 = pi3906 & n9771;
  assign n17354 = ~n17352 & ~n17353;
  assign n17355 = pi3954 & n9791;
  assign n17356 = pi3938 & n9788;
  assign n17357 = ~n17355 & ~n17356;
  assign n17358 = n17354 & n17357;
  assign n17359 = ~n17351 & n17358;
  assign n17360 = n17350 & n17359;
  assign n17361 = pi3874 & n9799;
  assign n17362 = n17360 & ~n17361;
  assign n17363 = pi3986 & n9783;
  assign n17364 = pi3970 & n9793;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = n17362 & n17365;
  assign n17367 = ~n9472 & ~n17366;
  assign n17368 = ~n17347 & ~n17367;
  assign n17369 = n16532 & ~n17368;
  assign n17370 = n16465 & ~n17226;
  assign n17371 = n16463 & ~n17251;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = n16468 & ~n17336;
  assign n17374 = n17372 & ~n17373;
  assign n17375 = ~pi2419 & ~n17374;
  assign n17376 = pi1946 & pi2419;
  assign n17377 = ~n17375 & ~n17376;
  assign n17378 = n16480 & ~n17377;
  assign n17379 = pi3730 & n16510;
  assign n17380 = pi3842 & n16504;
  assign n17381 = ~n17379 & ~n17380;
  assign n17382 = pi3810 & n16486;
  assign n17383 = n17381 & ~n17382;
  assign n17384 = pi3762 & n16502;
  assign n17385 = n17383 & ~n17384;
  assign n17386 = pi3730 & n16499;
  assign n17387 = pi3746 & n16493;
  assign n17388 = ~n17386 & ~n17387;
  assign n17389 = pi3794 & n16484;
  assign n17390 = pi3826 & n16489;
  assign n17391 = ~n17389 & ~n17390;
  assign n17392 = pi3778 & n16496;
  assign n17393 = n17391 & ~n17392;
  assign n17394 = n17388 & n17393;
  assign n17395 = n17385 & n17394;
  assign n17396 = ~n16480 & ~n17395;
  assign n17397 = ~n17378 & ~n17396;
  assign n17398 = n16462 & ~n17397;
  assign n17399 = ~n17369 & ~n17398;
  assign n17400 = pi0376 & n16535;
  assign po0129 = ~n17399 | n17400;
  assign n17402 = ~pi1422 & ~pi1856;
  assign n17403 = pi0366 & ~n17402;
  assign n17404 = pi0434 & n17402;
  assign n17405 = ~n17403 & ~n17404;
  assign po0130 = pi3641 & ~n17405;
  assign n17407 = pi0359 & ~n17402;
  assign n17408 = pi0433 & n17402;
  assign n17409 = ~n17407 & ~n17408;
  assign po0131 = pi3641 & ~n17409;
  assign n17411 = pi0432 & n17402;
  assign n17412 = pi0358 & ~n17402;
  assign n17413 = ~n17411 & ~n17412;
  assign po0132 = ~pi3641 | ~n17413;
  assign n17415 = pi0357 & ~n17402;
  assign n17416 = pi0431 & n17402;
  assign n17417 = ~n17415 & ~n17416;
  assign po0133 = pi3641 & ~n17417;
  assign n17419 = pi0356 & ~n17402;
  assign n17420 = pi0430 & n17402;
  assign n17421 = ~n17419 & ~n17420;
  assign po0134 = pi3641 & ~n17421;
  assign n17423 = pi0429 & n17402;
  assign n17424 = pi0355 & ~n17402;
  assign n17425 = ~n17423 & ~n17424;
  assign po0135 = ~pi3641 | ~n17425;
  assign n17427 = pi0354 & ~n17402;
  assign n17428 = pi0428 & n17402;
  assign n17429 = ~n17427 & ~n17428;
  assign po0136 = pi3641 & ~n17429;
  assign n17431 = pi0435 & n17402;
  assign n17432 = pi0353 & ~n17402;
  assign n17433 = ~n17431 & ~n17432;
  assign po0137 = ~pi3641 | ~n17433;
  assign n17435 = pi3641 & ~n17402;
  assign po0138 = pi0352 & n17435;
  assign po0139 = pi0351 & n17435;
  assign n17438 = pi0365 & ~n17402;
  assign po0140 = ~pi3641 | n17438;
  assign po0141 = pi0364 & n17435;
  assign po0142 = pi0363 & n17435;
  assign n17442 = pi0362 & ~n17402;
  assign po0143 = ~pi3641 | n17442;
  assign po0144 = pi0361 & n17435;
  assign n17445 = pi0360 & ~n17402;
  assign po0145 = ~pi3641 | n17445;
  assign n17447 = ~n8567 & n8603;
  assign n17448 = pi0366 & n17447;
  assign n17449 = ~n8567 & n8600;
  assign n17450 = pi1092 & n17449;
  assign n17451 = ~n11175 & n16470;
  assign n17452 = ~n17449 & ~n17451;
  assign n17453 = ~n17450 & ~n17452;
  assign n17454 = ~n17447 & ~n17453;
  assign po0146 = n17448 | n17454;
  assign n17456 = pi0359 & n17447;
  assign n17457 = ~pi1060 & n17449;
  assign n17458 = ~n12035 & ~n17449;
  assign n17459 = n16545 & n17458;
  assign n17460 = ~n17457 & ~n17459;
  assign n17461 = ~n17447 & n17460;
  assign po0147 = n17456 | n17461;
  assign n17463 = pi0358 & n17447;
  assign n17464 = pi1089 & n17449;
  assign n17465 = ~n15089 & n16581;
  assign n17466 = ~n17449 & ~n17465;
  assign n17467 = ~n17464 & ~n17466;
  assign n17468 = ~n17447 & ~n17467;
  assign po0148 = n17463 | n17468;
  assign n17470 = pi0357 & n17447;
  assign n17471 = ~pi1065 & n17449;
  assign n17472 = ~n14810 & ~n17449;
  assign n17473 = n16617 & n17472;
  assign n17474 = ~n17471 & ~n17473;
  assign n17475 = ~n17447 & n17474;
  assign po0149 = n17470 | n17475;
  assign n17477 = pi0356 & n17447;
  assign n17478 = pi1064 & n17449;
  assign n17479 = ~n12409 & n16653;
  assign n17480 = ~n17449 & ~n17479;
  assign n17481 = ~n17478 & ~n17480;
  assign n17482 = ~n17447 & ~n17481;
  assign po0150 = n17477 | n17482;
  assign n17484 = pi0355 & n17447;
  assign n17485 = pi1063 & n17449;
  assign n17486 = ~n13982 & n16689;
  assign n17487 = ~n17449 & ~n17486;
  assign n17488 = ~n17485 & ~n17487;
  assign n17489 = ~n17447 & ~n17488;
  assign po0151 = n17484 | n17489;
  assign n17491 = pi0354 & n17447;
  assign n17492 = ~pi1062 & n17449;
  assign n17493 = ~n13372 & ~n17449;
  assign n17494 = n16725 & n17493;
  assign n17495 = ~n17492 & ~n17494;
  assign n17496 = ~n17447 & n17495;
  assign po0152 = n17491 | n17496;
  assign n17498 = pi0353 & n17447;
  assign n17499 = ~pi1061 & n17449;
  assign n17500 = ~n13115 & ~n17449;
  assign n17501 = n16761 & n17500;
  assign n17502 = ~n17499 & ~n17501;
  assign n17503 = ~n17447 & n17502;
  assign po0153 = n17498 | n17503;
  assign n17505 = pi0352 & n17447;
  assign n17506 = ~pi3106 & n17449;
  assign n17507 = ~n13695 & ~n17449;
  assign n17508 = n16796 & n17507;
  assign n17509 = ~n17506 & ~n17508;
  assign n17510 = ~n17447 & n17509;
  assign po0154 = n17505 | n17510;
  assign n17512 = pi0351 & n17447;
  assign n17513 = ~pi3105 & n17449;
  assign n17514 = ~n12701 & ~n17449;
  assign n17515 = n16832 & n17514;
  assign n17516 = ~n17513 & ~n17515;
  assign n17517 = ~n17447 & n17516;
  assign po0155 = n17512 | n17517;
  assign n17519 = pi0365 & n17447;
  assign n17520 = pi3104 & n17449;
  assign n17521 = ~n14397 & n16868;
  assign n17522 = ~n17449 & ~n17521;
  assign n17523 = ~n17520 & ~n17522;
  assign n17524 = ~n17447 & ~n17523;
  assign po0156 = n17519 | n17524;
  assign n17526 = pi0364 & n17447;
  assign n17527 = pi2985 & n17449;
  assign n17528 = ~n15420 & n16904;
  assign n17529 = ~n17449 & ~n17528;
  assign n17530 = ~n17527 & ~n17529;
  assign n17531 = ~n17447 & ~n17530;
  assign po0157 = n17526 | n17531;
  assign n17533 = pi0363 & n17447;
  assign n17534 = pi3102 & n17449;
  assign n17535 = ~n10602 & n16940;
  assign n17536 = ~n17449 & ~n17535;
  assign n17537 = ~n17534 & ~n17536;
  assign n17538 = ~n17447 & ~n17537;
  assign po0158 = n17533 | n17538;
  assign n17540 = pi0362 & n17447;
  assign n17541 = pi3109 & n17449;
  assign n17542 = ~n9763 & n16976;
  assign n17543 = ~n17449 & ~n17542;
  assign n17544 = ~n17541 & ~n17543;
  assign n17545 = ~n17447 & ~n17544;
  assign po0159 = n17540 | n17545;
  assign n17547 = pi0361 & n17447;
  assign n17548 = ~pi3111 & n17449;
  assign n17549 = ~n17173 & ~n17449;
  assign n17550 = n17082 & n17549;
  assign n17551 = ~n17548 & ~n17550;
  assign n17552 = ~n17447 & n17551;
  assign po0160 = n17547 | n17552;
  assign n17554 = pi0360 & n17447;
  assign n17555 = pi3112 & n17449;
  assign n17556 = ~n17342 & n17374;
  assign n17557 = ~n17449 & ~n17556;
  assign n17558 = ~n17555 & ~n17557;
  assign n17559 = ~n17447 & ~n17558;
  assign po0161 = n17554 | n17559;
  assign n17561 = ~n8627 & n9422;
  assign n17562 = ~n8627 & n9419;
  assign n17563 = ~n8567 & n10781;
  assign n17564 = ~n8567 & n10783;
  assign n17565 = ~n17563 & ~n17564;
  assign n17566 = ~n17562 & n17565;
  assign n17567 = ~n17561 & n17566;
  assign n17568 = ~n11176 & n17567;
  assign n17569 = pi0844 & n17563;
  assign n17570 = pi0366 & n17564;
  assign n17571 = ~n17569 & ~n17570;
  assign n17572 = pi0479 & n17561;
  assign n17573 = pi2597 & n17562;
  assign n17574 = ~n17572 & ~n17573;
  assign n17575 = n17571 & n17574;
  assign n17576 = ~n17567 & ~n17575;
  assign po0162 = n17568 | n17576;
  assign n17578 = ~n12036 & n17567;
  assign n17579 = pi0843 & n17563;
  assign n17580 = pi0359 & n17564;
  assign n17581 = ~n17579 & ~n17580;
  assign n17582 = pi0370 & n17561;
  assign n17583 = pi2590 & n17562;
  assign n17584 = ~n17582 & ~n17583;
  assign n17585 = n17581 & n17584;
  assign n17586 = ~n17567 & ~n17585;
  assign po0163 = n17578 | n17586;
  assign n17588 = ~n15090 & n17567;
  assign n17589 = pi0842 & n17563;
  assign n17590 = pi0358 & n17564;
  assign n17591 = ~n17589 & ~n17590;
  assign n17592 = pi0350 & n17561;
  assign n17593 = pi2589 & n17562;
  assign n17594 = ~n17592 & ~n17593;
  assign n17595 = n17591 & n17594;
  assign n17596 = ~n17567 & ~n17595;
  assign po0164 = n17588 | n17596;
  assign n17598 = ~n14811 & n17567;
  assign n17599 = pi0864 & n17563;
  assign n17600 = pi0357 & n17564;
  assign n17601 = ~n17599 & ~n17600;
  assign n17602 = pi0331 & n17561;
  assign n17603 = pi2588 & n17562;
  assign n17604 = ~n17602 & ~n17603;
  assign n17605 = n17601 & n17604;
  assign n17606 = ~n17567 & ~n17605;
  assign po0165 = n17598 | n17606;
  assign n17608 = ~n12410 & n17567;
  assign n17609 = pi0841 & n17563;
  assign n17610 = pi0356 & n17564;
  assign n17611 = ~n17609 & ~n17610;
  assign n17612 = pi0329 & n17561;
  assign n17613 = pi2587 & n17562;
  assign n17614 = ~n17612 & ~n17613;
  assign n17615 = n17611 & n17614;
  assign n17616 = ~n17567 & ~n17615;
  assign po0166 = n17608 | n17616;
  assign n17618 = ~n13983 & n17567;
  assign n17619 = pi0865 & n17563;
  assign n17620 = pi0355 & n17564;
  assign n17621 = ~n17619 & ~n17620;
  assign n17622 = pi0278 & n17561;
  assign n17623 = pi2764 & n17562;
  assign n17624 = ~n17622 & ~n17623;
  assign n17625 = n17621 & n17624;
  assign n17626 = ~n17567 & ~n17625;
  assign po0167 = n17618 | n17626;
  assign n17628 = ~n13373 & n17567;
  assign n17629 = pi0840 & n17563;
  assign n17630 = pi0354 & n17564;
  assign n17631 = ~n17629 & ~n17630;
  assign n17632 = pi0248 & n17561;
  assign n17633 = pi2586 & n17562;
  assign n17634 = ~n17632 & ~n17633;
  assign n17635 = n17631 & n17634;
  assign n17636 = ~n17567 & ~n17635;
  assign po0168 = n17628 | n17636;
  assign n17638 = ~n13116 & n17567;
  assign n17639 = pi0839 & n17563;
  assign n17640 = pi0353 & n17564;
  assign n17641 = ~n17639 & ~n17640;
  assign n17642 = pi0247 & n17561;
  assign n17643 = pi2585 & n17562;
  assign n17644 = ~n17642 & ~n17643;
  assign n17645 = n17641 & n17644;
  assign n17646 = ~n17567 & ~n17645;
  assign po0169 = n17638 | n17646;
  assign n17648 = ~n13696 & n17567;
  assign n17649 = pi1092 & n17563;
  assign n17650 = pi0352 & n17564;
  assign n17651 = ~n17649 & ~n17650;
  assign n17652 = pi0232 & n17561;
  assign n17653 = pi2584 & n17562;
  assign n17654 = ~n17652 & ~n17653;
  assign n17655 = n17651 & n17654;
  assign n17656 = ~n17567 & ~n17655;
  assign po0170 = n17648 | n17656;
  assign n17658 = ~n12702 & n17567;
  assign n17659 = pi1060 & n17563;
  assign n17660 = pi0351 & n17564;
  assign n17661 = ~n17659 & ~n17660;
  assign n17662 = pi0237 & n17561;
  assign n17663 = pi2583 & n17562;
  assign n17664 = ~n17662 & ~n17663;
  assign n17665 = n17661 & n17664;
  assign n17666 = ~n17567 & ~n17665;
  assign po0171 = n17658 | n17666;
  assign n17668 = ~n14398 & n17567;
  assign n17669 = pi1089 & n17563;
  assign n17670 = pi0365 & n17564;
  assign n17671 = ~n17669 & ~n17670;
  assign n17672 = pi0225 & n17561;
  assign n17673 = pi2596 & n17562;
  assign n17674 = ~n17672 & ~n17673;
  assign n17675 = n17671 & n17674;
  assign n17676 = ~n17567 & ~n17675;
  assign po0172 = n17668 | n17676;
  assign n17678 = ~n15421 & n17567;
  assign n17679 = pi1065 & n17563;
  assign n17680 = pi0364 & n17564;
  assign n17681 = ~n17679 & ~n17680;
  assign n17682 = pi0224 & n17561;
  assign n17683 = pi2595 & n17562;
  assign n17684 = ~n17682 & ~n17683;
  assign n17685 = n17681 & n17684;
  assign n17686 = ~n17567 & ~n17685;
  assign po0173 = n17678 | n17686;
  assign n17688 = ~n10603 & n17567;
  assign n17689 = pi1064 & n17563;
  assign n17690 = pi0363 & n17564;
  assign n17691 = ~n17689 & ~n17690;
  assign n17692 = pi0189 & n17561;
  assign n17693 = pi2594 & n17562;
  assign n17694 = ~n17692 & ~n17693;
  assign n17695 = n17691 & n17694;
  assign n17696 = ~n17567 & ~n17695;
  assign po0174 = n17688 | n17696;
  assign n17698 = ~n9764 & n17567;
  assign n17699 = pi1063 & n17563;
  assign n17700 = pi0362 & n17564;
  assign n17701 = ~n17699 & ~n17700;
  assign n17702 = pi0606 & n17561;
  assign n17703 = pi2593 & n17562;
  assign n17704 = ~n17702 & ~n17703;
  assign n17705 = n17701 & n17704;
  assign n17706 = ~n17567 & ~n17705;
  assign po0175 = n17698 | n17706;
  assign n17708 = ~n17174 & n17567;
  assign n17709 = pi1062 & n17563;
  assign n17710 = pi0361 & n17564;
  assign n17711 = ~n17709 & ~n17710;
  assign n17712 = pi0607 & n17561;
  assign n17713 = pi2592 & n17562;
  assign n17714 = ~n17712 & ~n17713;
  assign n17715 = n17711 & n17714;
  assign n17716 = ~n17567 & ~n17715;
  assign po0176 = n17708 | n17716;
  assign n17718 = ~n17343 & n17567;
  assign n17719 = pi1061 & n17563;
  assign n17720 = pi0360 & n17564;
  assign n17721 = ~n17719 & ~n17720;
  assign n17722 = pi0605 & n17561;
  assign n17723 = pi2591 & n17562;
  assign n17724 = ~n17722 & ~n17723;
  assign n17725 = n17721 & n17724;
  assign n17726 = ~n17567 & ~n17725;
  assign po0177 = n17718 | n17726;
  assign n17728 = pi2437 & n10374;
  assign n17729 = pi1985 & n10379;
  assign n17730 = ~n17728 & ~n17729;
  assign n17731 = pi2270 & n10376;
  assign n17732 = pi2447 & n10381;
  assign n17733 = ~n17731 & ~n17732;
  assign n17734 = n17730 & n17733;
  assign n17735 = ~n9829 & ~n17734;
  assign n17736 = ~n10187 & n10296;
  assign n17737 = pi0568 & n10190;
  assign n17738 = ~n10191 & ~n17737;
  assign n17739 = ~n10296 & ~n17738;
  assign n17740 = ~n17736 & ~n17739;
  assign n17741 = ~pi0568 & ~n17740;
  assign n17742 = n10362 & ~n17738;
  assign n17743 = ~n10187 & ~n10362;
  assign n17744 = ~n17742 & ~n17743;
  assign n17745 = pi0568 & ~n17744;
  assign n17746 = ~n17741 & ~n17745;
  assign n17747 = pi0667 & n10166;
  assign n17748 = pi0667 & n9951;
  assign n17749 = pi0641 & n17748;
  assign n17750 = ~n17747 & ~n17749;
  assign n17751 = ~n17746 & n17750;
  assign n17752 = n9829 & ~n17751;
  assign n17753 = ~n17735 & ~n17752;
  assign n17754 = ~n9830 & ~n17753;
  assign n17755 = ~pi0749 & n9850;
  assign n17756 = pi2554 & po3871;
  assign n17757 = pi0873 & n9853;
  assign n17758 = ~n17756 & ~n17757;
  assign n17759 = pi2540 & ~n9903;
  assign n17760 = n17758 & ~n17759;
  assign n17761 = ~n9850 & n17760;
  assign n17762 = ~n17755 & ~n17761;
  assign n17763 = ~n9829 & n17762;
  assign n17764 = pi2437 & n9837;
  assign n17765 = pi2447 & n9834;
  assign n17766 = ~n17764 & ~n17765;
  assign n17767 = pi2270 & n9839;
  assign n17768 = pi1985 & n9832;
  assign n17769 = ~n17767 & ~n17768;
  assign n17770 = n17766 & n17769;
  assign n17771 = n9829 & ~n17770;
  assign n17772 = ~n17763 & ~n17771;
  assign n17773 = n9830 & ~n17772;
  assign n17774 = ~n17754 & ~n17773;
  assign n17775 = ~n9464 & ~n17774;
  assign n17776 = n9464 & ~n11181;
  assign po0202 = n17775 | n17776;
  assign n17778 = pi2434 & n10374;
  assign n17779 = pi2267 & n10376;
  assign n17780 = ~n17778 & ~n17779;
  assign n17781 = pi1982 & n10379;
  assign n17782 = pi2444 & n10381;
  assign n17783 = ~n17781 & ~n17782;
  assign n17784 = n17780 & n17783;
  assign n17785 = ~n9829 & ~n17784;
  assign n17786 = n10179 & n10185;
  assign n17787 = ~n10179 & ~n10185;
  assign n17788 = ~n17786 & ~n17787;
  assign n17789 = n10296 & ~n17788;
  assign n17790 = ~n10176 & ~n10182;
  assign n17791 = n10176 & n10182;
  assign n17792 = ~n17790 & ~n17791;
  assign n17793 = n10191 & n17792;
  assign n17794 = ~n10191 & ~n17792;
  assign n17795 = ~n17793 & ~n17794;
  assign n17796 = ~n10296 & ~n17795;
  assign n17797 = ~n17789 & ~n17796;
  assign n17798 = ~pi0568 & ~n17797;
  assign n17799 = n10362 & ~n17795;
  assign n17800 = ~n10362 & ~n17788;
  assign n17801 = ~n17799 & ~n17800;
  assign n17802 = pi0568 & ~n17801;
  assign n17803 = ~n17798 & ~n17802;
  assign n17804 = pi0665 & n10114;
  assign n17805 = ~n9951 & n17804;
  assign n17806 = n17803 & ~n17805;
  assign n17807 = pi0665 & ~n9956;
  assign n17808 = n9951 & n17807;
  assign n17809 = n17806 & ~n17808;
  assign n17810 = n9829 & ~n17809;
  assign n17811 = ~n17785 & ~n17810;
  assign n17812 = ~n9830 & ~n17811;
  assign n17813 = ~pi0778 & n9850;
  assign n17814 = pi2559 & po3871;
  assign n17815 = pi0908 & n9853;
  assign n17816 = ~n17814 & ~n17815;
  assign n17817 = pi2549 & ~n9903;
  assign n17818 = n17816 & ~n17817;
  assign n17819 = ~n9850 & n17818;
  assign n17820 = ~n17813 & ~n17819;
  assign n17821 = ~n9829 & n17820;
  assign n17822 = pi2434 & n9837;
  assign n17823 = pi1982 & n9832;
  assign n17824 = ~n17822 & ~n17823;
  assign n17825 = pi2267 & n9839;
  assign n17826 = pi2444 & n9834;
  assign n17827 = ~n17825 & ~n17826;
  assign n17828 = n17824 & n17827;
  assign n17829 = n9829 & ~n17828;
  assign n17830 = ~n17821 & ~n17829;
  assign n17831 = n9830 & ~n17830;
  assign n17832 = ~n17812 & ~n17831;
  assign n17833 = ~n9464 & ~n17832;
  assign n17834 = n9464 & ~n12061;
  assign po0203 = n17833 | n17834;
  assign n17836 = pi2266 & n10376;
  assign n17837 = pi2274 & n10381;
  assign n17838 = ~n17836 & ~n17837;
  assign n17839 = pi2433 & n10374;
  assign n17840 = pi1981 & n10379;
  assign n17841 = ~n17839 & ~n17840;
  assign n17842 = n17838 & n17841;
  assign n17843 = ~n9829 & ~n17842;
  assign n17844 = ~n10138 & ~n10315;
  assign n17845 = n10138 & n10315;
  assign n17846 = ~n17844 & ~n17845;
  assign n17847 = n10296 & ~n17846;
  assign n17848 = ~n10125 & ~n10141;
  assign n17849 = n10125 & n10141;
  assign n17850 = ~n17848 & ~n17849;
  assign n17851 = ~n10193 & n17850;
  assign n17852 = n10193 & ~n17850;
  assign n17853 = ~n17851 & ~n17852;
  assign n17854 = ~n10296 & ~n17853;
  assign n17855 = ~n17847 & ~n17854;
  assign n17856 = ~pi0568 & ~n17855;
  assign n17857 = n10362 & ~n17853;
  assign n17858 = ~n10362 & ~n17846;
  assign n17859 = ~n17857 & ~n17858;
  assign n17860 = pi0568 & ~n17859;
  assign n17861 = ~n17856 & ~n17860;
  assign n17862 = pi0664 & n10133;
  assign n17863 = pi0664 & n9951;
  assign n17864 = ~n10129 & n17863;
  assign n17865 = ~n17862 & ~n17864;
  assign n17866 = n17861 & n17865;
  assign n17867 = n9829 & ~n17866;
  assign n17868 = ~n17843 & ~n17867;
  assign n17869 = ~n9830 & ~n17868;
  assign n17870 = ~pi0777 & n9850;
  assign n17871 = pi2705 & po3871;
  assign n17872 = pi0907 & n9853;
  assign n17873 = ~n17871 & ~n17872;
  assign n17874 = pi2646 & ~n9903;
  assign n17875 = n17873 & ~n17874;
  assign n17876 = ~n9850 & n17875;
  assign n17877 = ~n17870 & ~n17876;
  assign n17878 = ~n9829 & n17877;
  assign n17879 = pi1981 & n9832;
  assign n17880 = pi2274 & n9834;
  assign n17881 = ~n17879 & ~n17880;
  assign n17882 = pi2433 & n9837;
  assign n17883 = pi2266 & n9839;
  assign n17884 = ~n17882 & ~n17883;
  assign n17885 = n17881 & n17884;
  assign n17886 = n9829 & ~n17885;
  assign n17887 = ~n17878 & ~n17886;
  assign n17888 = n9830 & ~n17887;
  assign n17889 = ~n17869 & ~n17888;
  assign n17890 = ~n9464 & ~n17889;
  assign n17891 = n9464 & ~n15115;
  assign po0204 = n17890 | n17891;
  assign n17893 = pi2260 & n10374;
  assign n17894 = pi2265 & n10376;
  assign n17895 = ~n17893 & ~n17894;
  assign n17896 = pi1980 & n10379;
  assign n17897 = pi2443 & n10381;
  assign n17898 = ~n17896 & ~n17897;
  assign n17899 = n17895 & n17898;
  assign n17900 = ~n9829 & ~n17899;
  assign n17901 = ~n10137 & ~n10315;
  assign n17902 = ~n10136 & ~n17901;
  assign n17903 = n10154 & ~n17902;
  assign n17904 = ~n10154 & n17902;
  assign n17905 = ~n17903 & ~n17904;
  assign n17906 = n10296 & ~n17905;
  assign n17907 = ~n10193 & ~n10196;
  assign n17908 = ~n10142 & ~n17907;
  assign n17909 = n10157 & ~n10159;
  assign n17910 = ~n10157 & n10159;
  assign n17911 = ~n17909 & ~n17910;
  assign n17912 = n17908 & n17911;
  assign n17913 = ~n17908 & ~n17911;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = ~n10296 & ~n17914;
  assign n17916 = ~n17906 & ~n17915;
  assign n17917 = ~pi0568 & ~n17916;
  assign n17918 = n10362 & ~n17914;
  assign n17919 = ~n10362 & ~n17905;
  assign n17920 = ~n17918 & ~n17919;
  assign n17921 = pi0568 & ~n17920;
  assign n17922 = ~n17917 & ~n17921;
  assign n17923 = pi0663 & n10149;
  assign n17924 = pi0663 & n9951;
  assign n17925 = ~n10017 & n17924;
  assign n17926 = ~n17923 & ~n17925;
  assign n17927 = ~n17922 & n17926;
  assign n17928 = n9829 & ~n17927;
  assign n17929 = ~n17900 & ~n17928;
  assign n17930 = ~n9830 & ~n17929;
  assign n17931 = ~pi0776 & n9850;
  assign n17932 = pi2556 & po3871;
  assign n17933 = pi0874 & n9853;
  assign n17934 = ~n17932 & ~n17933;
  assign n17935 = pi2551 & ~n9903;
  assign n17936 = n17934 & ~n17935;
  assign n17937 = ~n9850 & n17936;
  assign n17938 = ~n17931 & ~n17937;
  assign n17939 = ~n9829 & n17938;
  assign n17940 = pi2260 & n9837;
  assign n17941 = pi2443 & n9834;
  assign n17942 = ~n17940 & ~n17941;
  assign n17943 = pi2265 & n9839;
  assign n17944 = pi1980 & n9832;
  assign n17945 = ~n17943 & ~n17944;
  assign n17946 = n17942 & n17945;
  assign n17947 = n9829 & ~n17946;
  assign n17948 = ~n17939 & ~n17947;
  assign n17949 = n9830 & ~n17948;
  assign n17950 = ~n17930 & ~n17949;
  assign n17951 = ~n9464 & ~n17950;
  assign n17952 = n9464 & ~n14816;
  assign po0205 = n17951 | n17952;
  assign n17954 = pi2264 & n10376;
  assign n17955 = pi2273 & n10381;
  assign n17956 = ~n17954 & ~n17955;
  assign n17957 = pi2259 & n10374;
  assign n17958 = pi1979 & n10379;
  assign n17959 = ~n17957 & ~n17958;
  assign n17960 = n17956 & n17959;
  assign n17961 = ~n9829 & ~n17960;
  assign n17962 = ~n10254 & n10325;
  assign n17963 = n10254 & ~n10325;
  assign n17964 = ~n17962 & ~n17963;
  assign n17965 = n10296 & ~n17964;
  assign n17966 = ~n10257 & n10259;
  assign n17967 = n10257 & ~n10259;
  assign n17968 = ~n17966 & ~n17967;
  assign n17969 = n10203 & ~n17968;
  assign n17970 = ~n10203 & n17968;
  assign n17971 = ~n17969 & ~n17970;
  assign n17972 = ~n10296 & ~n17971;
  assign n17973 = ~n17965 & ~n17972;
  assign n17974 = ~pi0568 & ~n17973;
  assign n17975 = n10362 & ~n17971;
  assign n17976 = ~n10362 & ~n17964;
  assign n17977 = ~n17975 & ~n17976;
  assign n17978 = pi0568 & ~n17977;
  assign n17979 = ~n17974 & ~n17978;
  assign n17980 = pi0662 & n10247;
  assign n17981 = pi0662 & n10249;
  assign n17982 = ~n17980 & ~n17981;
  assign n17983 = n17979 & n17982;
  assign n17984 = n9829 & ~n17983;
  assign n17985 = ~n17961 & ~n17984;
  assign n17986 = ~n9830 & ~n17985;
  assign n17987 = ~pi0775 & n9850;
  assign n17988 = pi2704 & po3871;
  assign n17989 = pi0906 & n9853;
  assign n17990 = ~n17988 & ~n17989;
  assign n17991 = pi2553 & ~n9903;
  assign n17992 = n17990 & ~n17991;
  assign n17993 = ~n9850 & n17992;
  assign n17994 = ~n17987 & ~n17993;
  assign n17995 = ~n9829 & n17994;
  assign n17996 = pi2264 & n9839;
  assign n17997 = pi1979 & n9832;
  assign n17998 = ~n17996 & ~n17997;
  assign n17999 = pi2259 & n9837;
  assign n18000 = pi2273 & n9834;
  assign n18001 = ~n17999 & ~n18000;
  assign n18002 = n17998 & n18001;
  assign n18003 = n9829 & ~n18002;
  assign n18004 = ~n17995 & ~n18003;
  assign n18005 = n9830 & ~n18004;
  assign n18006 = ~n17986 & ~n18005;
  assign n18007 = ~n9464 & ~n18006;
  assign n18008 = n9464 & ~n12415;
  assign po0206 = n18007 | n18008;
  assign n18010 = n9829 & ~n14046;
  assign n18011 = ~n9829 & ~n13735;
  assign n18012 = ~n18010 & ~n18011;
  assign n18013 = ~n9830 & ~n18012;
  assign n18014 = ~pi0774 & n9850;
  assign n18015 = pi0905 & n9853;
  assign n18016 = ~n14051 & ~n18015;
  assign n18017 = pi2645 & ~n9903;
  assign n18018 = n18016 & ~n18017;
  assign n18019 = ~n9850 & n18018;
  assign n18020 = ~n18014 & ~n18019;
  assign n18021 = ~n9829 & n18020;
  assign n18022 = n9829 & ~n13727;
  assign n18023 = ~n18021 & ~n18022;
  assign n18024 = n9830 & ~n18023;
  assign n18025 = ~n18013 & ~n18024;
  assign n18026 = ~n9464 & ~n18025;
  assign n18027 = n9464 & ~n13988;
  assign po0207 = n18026 | n18027;
  assign n18029 = n9829 & ~n13451;
  assign n18030 = ~n9829 & ~n13424;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = ~n9830 & ~n18031;
  assign n18033 = ~pi0773 & n9850;
  assign n18034 = pi0904 & n9853;
  assign n18035 = ~n13456 & ~n18034;
  assign n18036 = pi2797 & ~n9903;
  assign n18037 = n18035 & ~n18036;
  assign n18038 = ~n9850 & n18037;
  assign n18039 = ~n18033 & ~n18038;
  assign n18040 = ~n9829 & n18039;
  assign n18041 = n9829 & ~n13416;
  assign n18042 = ~n18040 & ~n18041;
  assign n18043 = n9830 & ~n18042;
  assign n18044 = ~n18032 & ~n18043;
  assign n18045 = ~n9464 & ~n18044;
  assign n18046 = n9464 & ~n13398;
  assign po0208 = n18045 | n18046;
  assign n18048 = n9829 & ~n12785;
  assign n18049 = ~n9829 & ~n12801;
  assign n18050 = ~n18048 & ~n18049;
  assign n18051 = ~n9830 & ~n18050;
  assign n18052 = ~pi0861 & n9850;
  assign n18053 = pi0876 & n9853;
  assign n18054 = ~n12805 & ~n18053;
  assign n18055 = pi2644 & ~n9903;
  assign n18056 = n18054 & ~n18055;
  assign n18057 = ~n9850 & n18056;
  assign n18058 = ~n18052 & ~n18057;
  assign n18059 = ~n9829 & n18058;
  assign n18060 = n9829 & ~n12793;
  assign n18061 = ~n18059 & ~n18060;
  assign n18062 = n9830 & ~n18061;
  assign n18063 = ~n18051 & ~n18062;
  assign n18064 = ~n9464 & ~n18063;
  assign n18065 = n9464 & ~n13121;
  assign po0209 = n18064 | n18065;
  assign n18067 = n9464 & ~n13701;
  assign n18068 = ~pi0862 & n9850;
  assign n18069 = pi0903 & n9853;
  assign n18070 = ~n14158 & ~n18069;
  assign n18071 = pi2796 & ~n9903;
  assign n18072 = n18070 & ~n18071;
  assign n18073 = ~n9850 & n18072;
  assign n18074 = ~n18068 & ~n18073;
  assign n18075 = ~n9829 & n18074;
  assign n18076 = n9829 & ~n14144;
  assign n18077 = ~n18075 & ~n18076;
  assign n18078 = n9830 & ~n18077;
  assign n18079 = n9829 & ~n14134;
  assign n18080 = ~n9829 & ~n14152;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = ~n9830 & ~n18081;
  assign n18083 = ~n18078 & ~n18082;
  assign n18084 = ~n9464 & ~n18083;
  assign po0210 = n18067 | n18084;
  assign n18086 = n9464 & ~n12726;
  assign n18087 = ~pi0845 & n9850;
  assign n18088 = pi0902 & n9853;
  assign n18089 = ~n12453 & ~n18088;
  assign n18090 = pi2794 & ~n9903;
  assign n18091 = n18089 & ~n18090;
  assign n18092 = ~n9850 & n18091;
  assign n18093 = ~n18087 & ~n18092;
  assign n18094 = ~n9829 & n18093;
  assign n18095 = n9829 & ~n12155;
  assign n18096 = ~n18094 & ~n18095;
  assign n18097 = n9830 & ~n18096;
  assign n18098 = n9829 & ~n12445;
  assign n18099 = ~n9829 & ~n12163;
  assign n18100 = ~n18098 & ~n18099;
  assign n18101 = ~n9830 & ~n18100;
  assign n18102 = ~n18097 & ~n18101;
  assign n18103 = ~n9464 & ~n18102;
  assign po0211 = n18086 | n18103;
  assign n18105 = n9464 & ~n14403;
  assign n18106 = ~pi0781 & n9850;
  assign n18107 = pi0910 & n9853;
  assign n18108 = ~n14463 & ~n18107;
  assign n18109 = pi2788 & ~n9903;
  assign n18110 = n18108 & ~n18109;
  assign n18111 = ~n9850 & n18110;
  assign n18112 = ~n18106 & ~n18111;
  assign n18113 = ~n9829 & n18112;
  assign n18114 = n9829 & ~n14494;
  assign n18115 = ~n18113 & ~n18114;
  assign n18116 = n9830 & ~n18115;
  assign n18117 = n9829 & ~n14458;
  assign n18118 = ~n9829 & ~n14502;
  assign n18119 = ~n18117 & ~n18118;
  assign n18120 = ~n9830 & ~n18119;
  assign n18121 = ~n18116 & ~n18120;
  assign n18122 = ~n9464 & ~n18121;
  assign po0212 = n18105 | n18122;
  assign n18124 = n9464 & ~n15426;
  assign n18125 = ~pi0780 & n9850;
  assign n18126 = pi0820 & n9853;
  assign n18127 = ~n15150 & ~n18126;
  assign n18128 = pi2953 & ~n9903;
  assign n18129 = n18127 & ~n18128;
  assign n18130 = ~n9850 & n18129;
  assign n18131 = ~n18125 & ~n18130;
  assign n18132 = ~n9829 & n18131;
  assign n18133 = n9829 & ~n14849;
  assign n18134 = ~n18132 & ~n18133;
  assign n18135 = n9830 & ~n18134;
  assign n18136 = n9829 & ~n15146;
  assign n18137 = ~n9829 & ~n14857;
  assign n18138 = ~n18136 & ~n18137;
  assign n18139 = ~n9830 & ~n18138;
  assign n18140 = ~n18135 & ~n18139;
  assign n18141 = ~n9464 & ~n18140;
  assign po0213 = n18124 | n18141;
  assign n18143 = n10914 & n11752;
  assign n18144 = ~n10914 & n11214;
  assign n18145 = ~n18143 & ~n18144;
  assign n18146 = n10902 & n18145;
  assign n18147 = ~n11186 & ~n17751;
  assign n18148 = pi0749 & n11700;
  assign n18149 = n10886 & ~n11692;
  assign n18150 = pi0408 & n11714;
  assign n18151 = ~n18149 & ~n18150;
  assign n18152 = pi0873 & n11709;
  assign n18153 = pi1039 & ~n11706;
  assign n18154 = n9424 & ~n17734;
  assign n18155 = ~n9424 & ~n17770;
  assign n18156 = ~n18154 & ~n18155;
  assign n18157 = n11701 & ~n18156;
  assign n18158 = ~n18153 & ~n18157;
  assign n18159 = ~n18152 & n18158;
  assign n18160 = ~n17756 & n18159;
  assign n18161 = n18151 & n18160;
  assign n18162 = ~n11700 & ~n18161;
  assign n18163 = ~n18148 & ~n18162;
  assign n18164 = n11186 & ~n18163;
  assign n18165 = ~n18147 & ~n18164;
  assign n18166 = ~n10902 & ~n18165;
  assign n18167 = ~n18146 & ~n18166;
  assign n18168 = ~n10885 & ~n18167;
  assign n18169 = ~n11181 & ~n11186;
  assign n18170 = n11186 & ~n11674;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = n10902 & n18171;
  assign n18173 = ~n9825 & n11186;
  assign n18174 = n11692 & n18156;
  assign n18175 = ~n11186 & ~n18174;
  assign n18176 = ~n18173 & ~n18175;
  assign n18177 = ~n10902 & n18176;
  assign n18178 = ~n18172 & ~n18177;
  assign n18179 = n10885 & n18178;
  assign po0216 = n18168 | n18179;
  assign n18181 = ~n9424 & ~n17828;
  assign n18182 = n9424 & ~n17784;
  assign n18183 = ~n18181 & ~n18182;
  assign n18184 = n10914 & n18183;
  assign n18185 = n12124 & n18184;
  assign n18186 = n10608 & ~n10914;
  assign n18187 = ~n10902 & ~n18186;
  assign n18188 = ~n18185 & n18187;
  assign n18189 = ~n10914 & ~n12106;
  assign n18190 = n10914 & ~n12061;
  assign n18191 = ~n18189 & ~n18190;
  assign n18192 = n10902 & ~n18191;
  assign n18193 = ~n18188 & ~n18192;
  assign n18194 = n10885 & ~n18193;
  assign n18195 = n10914 & n11781;
  assign n18196 = ~n10914 & n11805;
  assign n18197 = ~n18195 & ~n18196;
  assign n18198 = n10902 & ~n18197;
  assign n18199 = pi0778 & n11700;
  assign n18200 = n11701 & ~n18183;
  assign n18201 = pi1012 & ~n11706;
  assign n18202 = ~n18200 & ~n18201;
  assign n18203 = pi0908 & n11709;
  assign n18204 = ~n17814 & ~n18203;
  assign n18205 = n18202 & n18204;
  assign n18206 = pi0413 & n11714;
  assign n18207 = n18205 & ~n18206;
  assign n18208 = n10886 & ~n12124;
  assign n18209 = n18207 & ~n18208;
  assign n18210 = ~n11700 & ~n18209;
  assign n18211 = ~n18199 & ~n18210;
  assign n18212 = ~n10914 & ~n18211;
  assign n18213 = n10914 & ~n17809;
  assign n18214 = ~n18212 & ~n18213;
  assign n18215 = ~n10902 & n18214;
  assign n18216 = ~n18198 & ~n18215;
  assign n18217 = ~n10885 & n18216;
  assign po0217 = n18194 | n18217;
  assign n18219 = n9424 & ~n17842;
  assign n18220 = ~n9424 & ~n17885;
  assign n18221 = ~n18219 & ~n18220;
  assign n18222 = n10914 & n18221;
  assign n18223 = n15205 & n18222;
  assign n18224 = ~n10914 & n15426;
  assign n18225 = ~n10902 & ~n18224;
  assign n18226 = ~n18223 & n18225;
  assign n18227 = ~n11186 & ~n15115;
  assign n18228 = n11186 & ~n15187;
  assign n18229 = ~n18227 & ~n18228;
  assign n18230 = n10902 & ~n18229;
  assign n18231 = ~n18226 & ~n18230;
  assign n18232 = n10885 & ~n18231;
  assign n18233 = n10914 & n15454;
  assign n18234 = ~n10914 & n14842;
  assign n18235 = ~n18233 & ~n18234;
  assign n18236 = n10902 & ~n18235;
  assign n18237 = pi0777 & n11700;
  assign n18238 = n11701 & ~n18221;
  assign n18239 = pi1034 & ~n11706;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = pi0907 & n11709;
  assign n18242 = ~n17871 & ~n18241;
  assign n18243 = n18240 & n18242;
  assign n18244 = pi0412 & n11714;
  assign n18245 = n18243 & ~n18244;
  assign n18246 = n10886 & ~n15205;
  assign n18247 = n18245 & ~n18246;
  assign n18248 = ~n11700 & ~n18247;
  assign n18249 = ~n18237 & ~n18248;
  assign n18250 = n11186 & ~n18249;
  assign n18251 = n10914 & ~n17866;
  assign n18252 = ~n18250 & ~n18251;
  assign n18253 = ~n10902 & n18252;
  assign n18254 = ~n18236 & ~n18253;
  assign n18255 = ~n10885 & n18254;
  assign po0218 = n18232 | n18255;
  assign n18257 = n10914 & n14430;
  assign n18258 = ~n10914 & n14485;
  assign n18259 = ~n18257 & ~n18258;
  assign n18260 = n10902 & n18259;
  assign n18261 = n10914 & ~n17927;
  assign n18262 = n9424 & ~n17899;
  assign n18263 = ~n9424 & ~n17946;
  assign n18264 = ~n18262 & ~n18263;
  assign n18265 = n11701 & ~n18264;
  assign n18266 = pi1033 & ~n11706;
  assign n18267 = ~n18265 & ~n18266;
  assign n18268 = pi0874 & n11709;
  assign n18269 = ~n17932 & ~n18268;
  assign n18270 = n18267 & n18269;
  assign n18271 = pi0411 & n11714;
  assign n18272 = n18270 & ~n18271;
  assign n18273 = n10886 & ~n14555;
  assign n18274 = n18272 & ~n18273;
  assign n18275 = ~n11700 & ~n18274;
  assign n18276 = pi0776 & n11700;
  assign n18277 = ~n18275 & ~n18276;
  assign n18278 = ~n10914 & ~n18277;
  assign n18279 = ~n18261 & ~n18278;
  assign n18280 = ~n10902 & ~n18279;
  assign n18281 = ~n18260 & ~n18280;
  assign n18282 = ~n10885 & ~n18281;
  assign n18283 = ~n11186 & ~n14816;
  assign n18284 = n11186 & ~n14537;
  assign n18285 = ~n18283 & ~n18284;
  assign n18286 = n10902 & n18285;
  assign n18287 = n14555 & n18264;
  assign n18288 = ~n11186 & ~n18287;
  assign n18289 = n11186 & ~n14403;
  assign n18290 = ~n18288 & ~n18289;
  assign n18291 = ~n10902 & n18290;
  assign n18292 = ~n18286 & ~n18291;
  assign n18293 = n10885 & n18292;
  assign po0219 = n18282 | n18293;
  assign n18295 = n10914 & n12751;
  assign n18296 = ~n10914 & n12148;
  assign n18297 = ~n18295 & ~n18296;
  assign n18298 = n10902 & n18297;
  assign n18299 = ~n11186 & ~n17983;
  assign n18300 = pi0775 & n11700;
  assign n18301 = pi1032 & ~n11706;
  assign n18302 = n9424 & ~n17960;
  assign n18303 = ~n9424 & ~n18002;
  assign n18304 = ~n18302 & ~n18303;
  assign n18305 = n11701 & ~n18304;
  assign n18306 = ~n18301 & ~n18305;
  assign n18307 = pi0906 & n11709;
  assign n18308 = n10886 & ~n12503;
  assign n18309 = pi0410 & n11714;
  assign n18310 = ~n18308 & ~n18309;
  assign n18311 = ~n17988 & n18310;
  assign n18312 = ~n18307 & n18311;
  assign n18313 = n18306 & n18312;
  assign n18314 = ~n11700 & ~n18313;
  assign n18315 = ~n18300 & ~n18314;
  assign n18316 = n11186 & ~n18315;
  assign n18317 = ~n18299 & ~n18316;
  assign n18318 = ~n10902 & ~n18317;
  assign n18319 = ~n18298 & ~n18318;
  assign n18320 = ~n10885 & ~n18319;
  assign n18321 = ~n11186 & ~n12415;
  assign n18322 = n11186 & ~n12485;
  assign n18323 = ~n18321 & ~n18322;
  assign n18324 = n10902 & n18323;
  assign n18325 = n12503 & n18304;
  assign n18326 = ~n11186 & ~n18325;
  assign n18327 = n11186 & ~n12726;
  assign n18328 = ~n18326 & ~n18327;
  assign n18329 = ~n10902 & n18328;
  assign n18330 = ~n18324 & ~n18329;
  assign n18331 = n10885 & n18330;
  assign po0220 = n18320 | n18331;
  assign n18333 = ~pi3460 & n16006;
  assign n18334 = pi1119 & n15846;
  assign n18335 = pi1315 & n15848;
  assign n18336 = ~n18334 & ~n18335;
  assign n18337 = pi1329 & n15841;
  assign n18338 = pi1189 & n15843;
  assign n18339 = ~n18337 & ~n18338;
  assign n18340 = pi1147 & n15831;
  assign n18341 = pi1161 & n15833;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = pi1273 & n15836;
  assign n18344 = pi1245 & n15838;
  assign n18345 = ~n18343 & ~n18344;
  assign n18346 = n18342 & n18345;
  assign n18347 = n18339 & n18346;
  assign n18348 = n18336 & n18347;
  assign n18349 = pi1175 & n15823;
  assign n18350 = pi1217 & n15825;
  assign n18351 = ~n18349 & ~n18350;
  assign n18352 = pi1301 & n15802;
  assign n18353 = pi1259 & n15806;
  assign n18354 = ~n18352 & ~n18353;
  assign n18355 = pi1287 & n15810;
  assign n18356 = pi1133 & n15812;
  assign n18357 = ~n18355 & ~n18356;
  assign n18358 = pi1231 & n15817;
  assign n18359 = pi1203 & n15819;
  assign n18360 = ~n18358 & ~n18359;
  assign n18361 = n18357 & n18360;
  assign n18362 = n18354 & n18361;
  assign n18363 = n18351 & n18362;
  assign n18364 = n18348 & n18363;
  assign n18365 = n15794 & ~n18364;
  assign n18366 = ~n9028 & n15940;
  assign n18367 = ~n18365 & ~n18366;
  assign n18368 = ~pi3400 & n15562;
  assign n18369 = pi0818 & n15579;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = pi2016 & n15945;
  assign n18372 = ~n9028 & ~n15945;
  assign n18373 = ~n18371 & ~n18372;
  assign n18374 = n15944 & ~n18373;
  assign n18375 = pi0014 & n15993;
  assign n18376 = ~n18374 & ~n18375;
  assign n18377 = n18370 & n18376;
  assign n18378 = n18367 & n18377;
  assign n18379 = ~n18333 & n18378;
  assign n18380 = n15552 & ~n18379;
  assign n18381 = pi0873 & n8589;
  assign n18382 = pi0749 & n16113;
  assign n18383 = ~n18381 & ~n18382;
  assign n18384 = po3841 & ~n18383;
  assign n18385 = ~n15552 & n18384;
  assign n18386 = ~n18380 & ~n18385;
  assign n18387 = pi3520 & n8561;
  assign n18388 = pi0408 & ~n8561;
  assign po3846 = n18387 | n18388;
  assign n18390 = ~n16035 & po3846;
  assign n18391 = pi3460 & n16035;
  assign n18392 = ~n18390 & ~n18391;
  assign n18393 = n16034 & ~n18392;
  assign po0230 = ~n18386 | n18393;
  assign n18395 = pi0908 & n8589;
  assign n18396 = pi0778 & n16113;
  assign n18397 = ~n18395 & ~n18396;
  assign n18398 = po3841 & ~n18397;
  assign n18399 = ~n15552 & n18398;
  assign n18400 = pi3400 & ~pi3403;
  assign n18401 = ~pi3400 & pi3403;
  assign n18402 = ~n18400 & ~n18401;
  assign n18403 = n15562 & ~n18402;
  assign n18404 = pi0813 & n15579;
  assign n18405 = ~n18403 & ~n18404;
  assign n18406 = pi1324 & n15841;
  assign n18407 = pi1184 & n15843;
  assign n18408 = ~n18406 & ~n18407;
  assign n18409 = pi1114 & n15846;
  assign n18410 = pi1310 & n15848;
  assign n18411 = ~n18409 & ~n18410;
  assign n18412 = pi1142 & n15831;
  assign n18413 = pi1156 & n15833;
  assign n18414 = ~n18412 & ~n18413;
  assign n18415 = pi1268 & n15836;
  assign n18416 = pi1240 & n15838;
  assign n18417 = ~n18415 & ~n18416;
  assign n18418 = n18414 & n18417;
  assign n18419 = n18411 & n18418;
  assign n18420 = n18408 & n18419;
  assign n18421 = pi1296 & n15802;
  assign n18422 = pi1254 & n15806;
  assign n18423 = ~n18421 & ~n18422;
  assign n18424 = pi1282 & n15810;
  assign n18425 = pi1128 & n15812;
  assign n18426 = ~n18424 & ~n18425;
  assign n18427 = pi1226 & n15817;
  assign n18428 = pi1198 & n15819;
  assign n18429 = ~n18427 & ~n18428;
  assign n18430 = pi1170 & n15823;
  assign n18431 = pi1212 & n15825;
  assign n18432 = ~n18430 & ~n18431;
  assign n18433 = n18429 & n18432;
  assign n18434 = n18426 & n18433;
  assign n18435 = n18423 & n18434;
  assign n18436 = n18420 & n18435;
  assign n18437 = n15794 & ~n18436;
  assign n18438 = ~n8802 & n15940;
  assign n18439 = ~n18437 & ~n18438;
  assign n18440 = pi2015 & n15945;
  assign n18441 = ~n8802 & ~n15945;
  assign n18442 = ~n18440 & ~n18441;
  assign n18443 = n15944 & ~n18442;
  assign n18444 = pi0015 & n15993;
  assign n18445 = ~n18443 & ~n18444;
  assign n18446 = ~pi3437 & pi3460;
  assign n18447 = pi3437 & ~pi3460;
  assign n18448 = ~n18446 & ~n18447;
  assign n18449 = n16006 & ~n18448;
  assign n18450 = n18445 & ~n18449;
  assign n18451 = n18439 & n18450;
  assign n18452 = n18405 & n18451;
  assign n18453 = n15552 & ~n18452;
  assign n18454 = ~n18399 & ~n18453;
  assign n18455 = pi3511 & n8561;
  assign n18456 = pi0413 & ~n8561;
  assign po3837 = n18455 | n18456;
  assign n18458 = ~n16035 & po3837;
  assign n18459 = pi3437 & n16035;
  assign n18460 = ~n18458 & ~n18459;
  assign n18461 = n16034 & ~n18460;
  assign po0231 = ~n18454 | n18461;
  assign n18463 = pi0907 & n8589;
  assign n18464 = pi0777 & n16113;
  assign n18465 = ~n18463 & ~n18464;
  assign n18466 = po3841 & ~n18465;
  assign n18467 = ~n15552 & n18466;
  assign n18468 = ~pi3433 & ~n16009;
  assign n18469 = ~n16045 & ~n18468;
  assign n18470 = n16006 & n18469;
  assign n18471 = ~pi1330 & ~pi3269;
  assign n18472 = ~pi1597 & ~pi2019;
  assign n18473 = ~pi2474 & n18472;
  assign n18474 = ~pi1048 & n18473;
  assign n18475 = n18471 & n18474;
  assign n18476 = n9873 & ~n15553;
  assign n18477 = ~n18475 & n18476;
  assign n18478 = ~n18470 & ~n18477;
  assign n18479 = pi2014 & n15945;
  assign n18480 = ~n9065 & ~n15945;
  assign n18481 = ~n18479 & ~n18480;
  assign n18482 = n15944 & ~n18481;
  assign n18483 = pi0016 & n15993;
  assign n18484 = ~n18482 & ~n18483;
  assign n18485 = pi1113 & n15846;
  assign n18486 = pi1309 & n15848;
  assign n18487 = ~n18485 & ~n18486;
  assign n18488 = pi1141 & n15831;
  assign n18489 = pi1155 & n15833;
  assign n18490 = ~n18488 & ~n18489;
  assign n18491 = pi1323 & n15841;
  assign n18492 = pi1183 & n15843;
  assign n18493 = ~n18491 & ~n18492;
  assign n18494 = pi1267 & n15836;
  assign n18495 = pi1239 & n15838;
  assign n18496 = ~n18494 & ~n18495;
  assign n18497 = n18493 & n18496;
  assign n18498 = n18490 & n18497;
  assign n18499 = n18487 & n18498;
  assign n18500 = pi1295 & n15802;
  assign n18501 = pi1253 & n15806;
  assign n18502 = ~n18500 & ~n18501;
  assign n18503 = pi1169 & n15823;
  assign n18504 = pi1211 & n15825;
  assign n18505 = ~n18503 & ~n18504;
  assign n18506 = pi1225 & n15817;
  assign n18507 = pi1197 & n15819;
  assign n18508 = ~n18506 & ~n18507;
  assign n18509 = pi1281 & n15810;
  assign n18510 = pi1127 & n15812;
  assign n18511 = ~n18509 & ~n18510;
  assign n18512 = n18508 & n18511;
  assign n18513 = n18505 & n18512;
  assign n18514 = n18502 & n18513;
  assign n18515 = n18499 & n18514;
  assign n18516 = n15794 & ~n18515;
  assign n18517 = ~n9065 & n15940;
  assign n18518 = ~n18516 & ~n18517;
  assign n18519 = ~pi3402 & ~n15564;
  assign n18520 = ~n15565 & ~n18519;
  assign n18521 = n15562 & n18520;
  assign n18522 = pi0812 & n15579;
  assign n18523 = ~n18521 & ~n18522;
  assign n18524 = n18518 & n18523;
  assign n18525 = n18484 & n18524;
  assign n18526 = n18478 & n18525;
  assign n18527 = n15552 & ~n18526;
  assign n18528 = ~n18467 & ~n18527;
  assign n18529 = pi3510 & n8561;
  assign n18530 = pi0412 & ~n8561;
  assign po3836 = n18529 | n18530;
  assign n18532 = ~n16035 & po3836;
  assign n18533 = pi3433 & n16035;
  assign n18534 = ~n18532 & ~n18533;
  assign n18535 = n16034 & ~n18534;
  assign po0232 = ~n18528 | n18535;
  assign n18537 = pi0874 & n8589;
  assign n18538 = pi0776 & n16113;
  assign n18539 = ~n18537 & ~n18538;
  assign n18540 = po3841 & ~n18539;
  assign n18541 = ~n15552 & n18540;
  assign n18542 = ~pi3457 & ~n16045;
  assign n18543 = ~n16046 & ~n18542;
  assign n18544 = n16006 & n18543;
  assign n18545 = ~pi1048 & ~pi2018;
  assign n18546 = ~pi1049 & ~pi3269;
  assign n18547 = ~pi1597 & ~pi2777;
  assign n18548 = n18546 & n18547;
  assign n18549 = n18545 & n18548;
  assign n18550 = n18476 & ~n18549;
  assign n18551 = ~n18544 & ~n18550;
  assign n18552 = pi2013 & n15945;
  assign n18553 = ~n8839 & ~n15945;
  assign n18554 = ~n18552 & ~n18553;
  assign n18555 = n15944 & ~n18554;
  assign n18556 = pi0017 & n15993;
  assign n18557 = ~n18555 & ~n18556;
  assign n18558 = pi1280 & n15810;
  assign n18559 = pi1126 & n15812;
  assign n18560 = ~n18558 & ~n18559;
  assign n18561 = pi1168 & n15823;
  assign n18562 = pi1210 & n15825;
  assign n18563 = ~n18561 & ~n18562;
  assign n18564 = pi1224 & n15817;
  assign n18565 = pi1196 & n15819;
  assign n18566 = ~n18564 & ~n18565;
  assign n18567 = pi1294 & n15802;
  assign n18568 = pi1252 & n15806;
  assign n18569 = ~n18567 & ~n18568;
  assign n18570 = n18566 & n18569;
  assign n18571 = n18563 & n18570;
  assign n18572 = n18560 & n18571;
  assign n18573 = pi1140 & n15831;
  assign n18574 = pi1154 & n15833;
  assign n18575 = ~n18573 & ~n18574;
  assign n18576 = pi1322 & n15841;
  assign n18577 = pi1182 & n15843;
  assign n18578 = ~n18576 & ~n18577;
  assign n18579 = pi1266 & n15836;
  assign n18580 = pi1238 & n15838;
  assign n18581 = ~n18579 & ~n18580;
  assign n18582 = pi1112 & n15846;
  assign n18583 = pi1308 & n15848;
  assign n18584 = ~n18582 & ~n18583;
  assign n18585 = n18581 & n18584;
  assign n18586 = n18578 & n18585;
  assign n18587 = n18575 & n18586;
  assign n18588 = n18572 & n18587;
  assign n18589 = n15794 & ~n18588;
  assign n18590 = ~n8839 & n15940;
  assign n18591 = ~n18589 & ~n18590;
  assign n18592 = ~pi3404 & ~n15565;
  assign n18593 = ~n15566 & ~n18592;
  assign n18594 = n15562 & n18593;
  assign n18595 = pi0811 & n15579;
  assign n18596 = ~n18594 & ~n18595;
  assign n18597 = n18591 & n18596;
  assign n18598 = n18557 & n18597;
  assign n18599 = n18551 & n18598;
  assign n18600 = n15552 & ~n18599;
  assign n18601 = ~n18541 & ~n18600;
  assign n18602 = pi3521 & n8561;
  assign n18603 = pi0411 & ~n8561;
  assign po3847 = n18602 | n18603;
  assign n18605 = ~n16035 & po3847;
  assign n18606 = pi3457 & n16035;
  assign n18607 = ~n18605 & ~n18606;
  assign n18608 = n16034 & ~n18607;
  assign po0233 = ~n18601 | n18608;
  assign n18610 = pi2012 & n15945;
  assign n18611 = ~n8950 & ~n15945;
  assign n18612 = ~n18610 & ~n18611;
  assign n18613 = n15944 & ~n18612;
  assign n18614 = pi0018 & n15993;
  assign n18615 = ~n18613 & ~n18614;
  assign n18616 = pi3456 & n16046;
  assign n18617 = ~pi3456 & ~n16046;
  assign n18618 = ~n18616 & ~n18617;
  assign n18619 = n16006 & n18618;
  assign n18620 = n18615 & ~n18619;
  assign n18621 = ~pi2017 & ~pi2019;
  assign n18622 = n18545 & n18621;
  assign n18623 = n18476 & ~n18622;
  assign n18624 = n18620 & ~n18623;
  assign n18625 = ~pi3414 & ~n15566;
  assign n18626 = ~n15567 & ~n18625;
  assign n18627 = n15562 & n18626;
  assign n18628 = pi0810 & n15579;
  assign n18629 = ~n18627 & ~n18628;
  assign n18630 = pi1223 & n15817;
  assign n18631 = pi1195 & n15819;
  assign n18632 = ~n18630 & ~n18631;
  assign n18633 = pi1293 & n15802;
  assign n18634 = pi1251 & n15806;
  assign n18635 = ~n18633 & ~n18634;
  assign n18636 = pi1167 & n15823;
  assign n18637 = pi1209 & n15825;
  assign n18638 = ~n18636 & ~n18637;
  assign n18639 = pi1279 & n15810;
  assign n18640 = pi1125 & n15812;
  assign n18641 = ~n18639 & ~n18640;
  assign n18642 = n18638 & n18641;
  assign n18643 = n18635 & n18642;
  assign n18644 = n18632 & n18643;
  assign n18645 = pi1139 & n15831;
  assign n18646 = pi1153 & n15833;
  assign n18647 = ~n18645 & ~n18646;
  assign n18648 = pi1111 & n15846;
  assign n18649 = pi1307 & n15848;
  assign n18650 = ~n18648 & ~n18649;
  assign n18651 = pi1321 & n15841;
  assign n18652 = pi1181 & n15843;
  assign n18653 = ~n18651 & ~n18652;
  assign n18654 = pi1265 & n15836;
  assign n18655 = pi1237 & n15838;
  assign n18656 = ~n18654 & ~n18655;
  assign n18657 = n18653 & n18656;
  assign n18658 = n18650 & n18657;
  assign n18659 = n18647 & n18658;
  assign n18660 = n18644 & n18659;
  assign n18661 = n15794 & ~n18660;
  assign n18662 = ~n8950 & n15940;
  assign n18663 = ~n18661 & ~n18662;
  assign n18664 = n18629 & n18663;
  assign n18665 = n18624 & n18664;
  assign n18666 = n15552 & ~n18665;
  assign n18667 = pi0906 & n8589;
  assign n18668 = pi0775 & n16113;
  assign n18669 = ~n18667 & ~n18668;
  assign n18670 = po3841 & ~n18669;
  assign n18671 = ~n15552 & n18670;
  assign n18672 = ~n18666 & ~n18671;
  assign n18673 = pi3509 & n8561;
  assign n18674 = pi0410 & ~n8561;
  assign po3835 = n18673 | n18674;
  assign n18676 = ~n16035 & po3835;
  assign n18677 = pi3456 & n16035;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 = n16034 & ~n18678;
  assign po0234 = ~n18672 | n18679;
  assign n18681 = pi2011 & n15945;
  assign n18682 = ~n8876 & ~n15945;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = n15944 & ~n18683;
  assign n18685 = pi0019 & n15993;
  assign n18686 = ~n18684 & ~n18685;
  assign n18687 = ~pi3434 & ~n16012;
  assign n18688 = pi3434 & n16012;
  assign n18689 = ~n18687 & ~n18688;
  assign n18690 = n16006 & n18689;
  assign n18691 = n18686 & ~n18690;
  assign n18692 = ~pi1330 & n18546;
  assign n18693 = ~pi1598 & n18692;
  assign n18694 = n18476 & ~n18693;
  assign n18695 = n18691 & ~n18694;
  assign n18696 = ~pi3405 & ~n15567;
  assign n18697 = pi3405 & n15567;
  assign n18698 = ~n18696 & ~n18697;
  assign n18699 = n15562 & n18698;
  assign n18700 = pi0809 & n15579;
  assign n18701 = ~n18699 & ~n18700;
  assign n18702 = pi1110 & n15846;
  assign n18703 = pi1306 & n15848;
  assign n18704 = ~n18702 & ~n18703;
  assign n18705 = pi1264 & n15836;
  assign n18706 = pi1236 & n15838;
  assign n18707 = ~n18705 & ~n18706;
  assign n18708 = pi1138 & n15831;
  assign n18709 = pi1152 & n15833;
  assign n18710 = ~n18708 & ~n18709;
  assign n18711 = pi1320 & n15841;
  assign n18712 = pi1180 & n15843;
  assign n18713 = ~n18711 & ~n18712;
  assign n18714 = n18710 & n18713;
  assign n18715 = n18707 & n18714;
  assign n18716 = n18704 & n18715;
  assign n18717 = pi1292 & n15802;
  assign n18718 = pi1250 & n15806;
  assign n18719 = ~n18717 & ~n18718;
  assign n18720 = pi1222 & n15817;
  assign n18721 = pi1194 & n15819;
  assign n18722 = ~n18720 & ~n18721;
  assign n18723 = pi1166 & n15823;
  assign n18724 = pi1208 & n15825;
  assign n18725 = ~n18723 & ~n18724;
  assign n18726 = pi1278 & n15810;
  assign n18727 = pi1124 & n15812;
  assign n18728 = ~n18726 & ~n18727;
  assign n18729 = n18725 & n18728;
  assign n18730 = n18722 & n18729;
  assign n18731 = n18719 & n18730;
  assign n18732 = n18716 & n18731;
  assign n18733 = n15794 & ~n18732;
  assign n18734 = ~n8876 & n15940;
  assign n18735 = ~n18733 & ~n18734;
  assign n18736 = n18701 & n18735;
  assign n18737 = n18695 & n18736;
  assign n18738 = n15552 & ~n18737;
  assign n18739 = pi0905 & n8589;
  assign n18740 = pi0774 & n16113;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = po3841 & ~n18741;
  assign n18743 = ~n15552 & n18742;
  assign n18744 = ~n18738 & ~n18743;
  assign n18745 = pi3508 & n8561;
  assign n18746 = pi0409 & ~n8561;
  assign po3834 = n18745 | n18746;
  assign n18748 = ~n16035 & po3834;
  assign n18749 = pi3434 & n16035;
  assign n18750 = ~n18748 & ~n18749;
  assign n18751 = n16034 & ~n18750;
  assign po0235 = ~n18744 | n18751;
  assign n18753 = ~pi3413 & ~n18697;
  assign n18754 = pi3413 & n18697;
  assign n18755 = ~n18753 & ~n18754;
  assign n18756 = n15562 & n18755;
  assign n18757 = pi0808 & n15579;
  assign n18758 = ~n18756 & ~n18757;
  assign n18759 = pi1137 & n15831;
  assign n18760 = pi1151 & n15833;
  assign n18761 = ~n18759 & ~n18760;
  assign n18762 = pi1263 & n15836;
  assign n18763 = pi1235 & n15838;
  assign n18764 = ~n18762 & ~n18763;
  assign n18765 = pi1109 & n15846;
  assign n18766 = pi1305 & n15848;
  assign n18767 = ~n18765 & ~n18766;
  assign n18768 = pi1319 & n15841;
  assign n18769 = pi1179 & n15843;
  assign n18770 = ~n18768 & ~n18769;
  assign n18771 = n18767 & n18770;
  assign n18772 = n18764 & n18771;
  assign n18773 = n18761 & n18772;
  assign n18774 = pi1165 & n15823;
  assign n18775 = pi1207 & n15825;
  assign n18776 = ~n18774 & ~n18775;
  assign n18777 = pi1221 & n15817;
  assign n18778 = pi1193 & n15819;
  assign n18779 = ~n18777 & ~n18778;
  assign n18780 = pi1277 & n15810;
  assign n18781 = pi1123 & n15812;
  assign n18782 = ~n18780 & ~n18781;
  assign n18783 = pi1291 & n15802;
  assign n18784 = pi1249 & n15806;
  assign n18785 = ~n18783 & ~n18784;
  assign n18786 = n18782 & n18785;
  assign n18787 = n18779 & n18786;
  assign n18788 = n18776 & n18787;
  assign n18789 = n18773 & n18788;
  assign n18790 = n15794 & ~n18789;
  assign n18791 = ~n8987 & n15940;
  assign n18792 = ~n18790 & ~n18791;
  assign n18793 = pi2374 & n15945;
  assign n18794 = ~n8987 & ~n15945;
  assign n18795 = ~n18793 & ~n18794;
  assign n18796 = n15944 & ~n18795;
  assign n18797 = pi0020 & n15993;
  assign n18798 = ~n18796 & ~n18797;
  assign n18799 = pi3434 & n16009;
  assign n18800 = n16011 & n18799;
  assign n18801 = ~pi3455 & n18800;
  assign n18802 = pi3455 & ~n18800;
  assign n18803 = ~n18801 & ~n18802;
  assign n18804 = n16006 & ~n18803;
  assign n18805 = n18798 & ~n18804;
  assign n18806 = n18792 & n18805;
  assign n18807 = n18758 & n18806;
  assign n18808 = n15552 & ~n18807;
  assign n18809 = pi0904 & n8589;
  assign n18810 = pi0773 & n16113;
  assign n18811 = ~n18809 & ~n18810;
  assign n18812 = po3841 & ~n18811;
  assign n18813 = ~n15552 & n18812;
  assign n18814 = ~n18808 & ~n18813;
  assign n18815 = pi3517 & n8561;
  assign n18816 = pi0426 & ~n8561;
  assign po3843 = n18815 | n18816;
  assign n18818 = ~n16035 & po3843;
  assign n18819 = pi3455 & n16035;
  assign n18820 = ~n18818 & ~n18819;
  assign n18821 = n16034 & ~n18820;
  assign po0236 = ~n18814 | n18821;
  assign n18823 = pi0876 & n8589;
  assign n18824 = pi0861 & n16113;
  assign n18825 = ~n18823 & ~n18824;
  assign n18826 = po3841 & ~n18825;
  assign n18827 = ~n15552 & n18826;
  assign n18828 = ~pi3406 & ~n15569;
  assign n18829 = ~n16092 & ~n18828;
  assign n18830 = n15562 & n18829;
  assign n18831 = pi0807 & n15579;
  assign n18832 = ~n18830 & ~n18831;
  assign n18833 = pi1164 & n15823;
  assign n18834 = pi1206 & n15825;
  assign n18835 = ~n18833 & ~n18834;
  assign n18836 = pi1220 & n15817;
  assign n18837 = pi1192 & n15819;
  assign n18838 = ~n18836 & ~n18837;
  assign n18839 = pi1276 & n15810;
  assign n18840 = pi1122 & n15812;
  assign n18841 = ~n18839 & ~n18840;
  assign n18842 = pi1290 & n15802;
  assign n18843 = pi1248 & n15806;
  assign n18844 = ~n18842 & ~n18843;
  assign n18845 = n18841 & n18844;
  assign n18846 = n18838 & n18845;
  assign n18847 = n18835 & n18846;
  assign n18848 = pi1318 & n15841;
  assign n18849 = pi1178 & n15843;
  assign n18850 = ~n18848 & ~n18849;
  assign n18851 = pi1136 & n15831;
  assign n18852 = pi1150 & n15833;
  assign n18853 = ~n18851 & ~n18852;
  assign n18854 = pi1262 & n15836;
  assign n18855 = pi1234 & n15838;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = pi1108 & n15846;
  assign n18858 = pi1304 & n15848;
  assign n18859 = ~n18857 & ~n18858;
  assign n18860 = n18856 & n18859;
  assign n18861 = n18853 & n18860;
  assign n18862 = n18850 & n18861;
  assign n18863 = n18847 & n18862;
  assign n18864 = n15794 & ~n18863;
  assign n18865 = ~n8913 & n15940;
  assign n18866 = ~n18864 & ~n18865;
  assign n18867 = pi2010 & n15945;
  assign n18868 = ~n8913 & ~n15945;
  assign n18869 = ~n18867 & ~n18868;
  assign n18870 = n15944 & ~n18869;
  assign n18871 = pi0021 & n15993;
  assign n18872 = ~n18870 & ~n18871;
  assign n18873 = n16008 & n16045;
  assign n18874 = pi3456 & n18873;
  assign n18875 = pi3457 & n18874;
  assign n18876 = pi3454 & n18875;
  assign n18877 = ~pi3454 & ~n18875;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = n16006 & n18878;
  assign n18880 = n18872 & ~n18879;
  assign n18881 = n18866 & n18880;
  assign n18882 = n18832 & n18881;
  assign n18883 = n15552 & ~n18882;
  assign n18884 = ~n18827 & ~n18883;
  assign n18885 = pi3516 & n8561;
  assign n18886 = pi0425 & ~n8561;
  assign po3842 = n18885 | n18886;
  assign n18888 = ~n16035 & po3842;
  assign n18889 = pi3454 & n16035;
  assign n18890 = ~n18888 & ~n18889;
  assign n18891 = n16034 & ~n18890;
  assign po0237 = ~n18884 | n18891;
  assign n18893 = pi0903 & n8589;
  assign n18894 = pi0862 & n16113;
  assign n18895 = ~n18893 & ~n18894;
  assign n18896 = po3841 & ~n18895;
  assign n18897 = ~n15552 & n18896;
  assign n18898 = ~pi3411 & ~n16092;
  assign n18899 = pi3411 & n16092;
  assign n18900 = ~n18898 & ~n18899;
  assign n18901 = n15562 & n18900;
  assign n18902 = pi0806 & n15579;
  assign n18903 = ~n18901 & ~n18902;
  assign n18904 = pi1275 & n15810;
  assign n18905 = pi1121 & n15812;
  assign n18906 = ~n18904 & ~n18905;
  assign n18907 = pi1219 & n15817;
  assign n18908 = pi1191 & n15819;
  assign n18909 = ~n18907 & ~n18908;
  assign n18910 = pi1163 & n15823;
  assign n18911 = pi1205 & n15825;
  assign n18912 = ~n18910 & ~n18911;
  assign n18913 = pi1289 & n15802;
  assign n18914 = pi1247 & n15806;
  assign n18915 = ~n18913 & ~n18914;
  assign n18916 = n18912 & n18915;
  assign n18917 = n18909 & n18916;
  assign n18918 = n18906 & n18917;
  assign n18919 = pi1261 & n15836;
  assign n18920 = pi1233 & n15838;
  assign n18921 = ~n18919 & ~n18920;
  assign n18922 = pi1107 & n15846;
  assign n18923 = pi1303 & n15848;
  assign n18924 = ~n18922 & ~n18923;
  assign n18925 = pi1135 & n15831;
  assign n18926 = pi1149 & n15833;
  assign n18927 = ~n18925 & ~n18926;
  assign n18928 = pi1317 & n15841;
  assign n18929 = pi1177 & n15843;
  assign n18930 = ~n18928 & ~n18929;
  assign n18931 = n18927 & n18930;
  assign n18932 = n18924 & n18931;
  assign n18933 = n18921 & n18932;
  assign n18934 = n18918 & n18933;
  assign n18935 = n15794 & ~n18934;
  assign n18936 = ~n9142 & n15940;
  assign n18937 = ~n18935 & ~n18936;
  assign n18938 = pi2373 & n15945;
  assign n18939 = ~n9142 & ~n15945;
  assign n18940 = ~n18938 & ~n18939;
  assign n18941 = n15944 & ~n18940;
  assign n18942 = pi0022 & n15993;
  assign n18943 = ~n18941 & ~n18942;
  assign n18944 = pi3453 & n16049;
  assign n18945 = ~pi3453 & ~n16049;
  assign n18946 = ~n18944 & ~n18945;
  assign n18947 = n16006 & n18946;
  assign n18948 = n18943 & ~n18947;
  assign n18949 = n18937 & n18948;
  assign n18950 = n18903 & n18949;
  assign n18951 = n15552 & ~n18950;
  assign n18952 = ~n18897 & ~n18951;
  assign n18953 = pi3518 & n8561;
  assign n18954 = pi0406 & ~n8561;
  assign po3844 = n18953 | n18954;
  assign n18956 = ~n16035 & po3844;
  assign n18957 = pi3453 & n16035;
  assign n18958 = ~n18956 & ~n18957;
  assign n18959 = n16034 & ~n18958;
  assign po0238 = ~n18952 | n18959;
  assign n18961 = pi0902 & n8589;
  assign n18962 = pi0845 & n16113;
  assign n18963 = ~n18961 & ~n18962;
  assign n18964 = po3841 & ~n18963;
  assign n18965 = ~n15552 & n18964;
  assign n18966 = ~pi3420 & n15571;
  assign n18967 = pi3420 & ~n15571;
  assign n18968 = ~n18966 & ~n18967;
  assign n18969 = n15562 & ~n18968;
  assign n18970 = pi0788 & n15579;
  assign n18971 = ~n18969 & ~n18970;
  assign n18972 = pi1106 & n15846;
  assign n18973 = pi1302 & n15848;
  assign n18974 = ~n18972 & ~n18973;
  assign n18975 = pi1134 & n15831;
  assign n18976 = pi1148 & n15833;
  assign n18977 = ~n18975 & ~n18976;
  assign n18978 = pi1260 & n15836;
  assign n18979 = pi1232 & n15838;
  assign n18980 = ~n18978 & ~n18979;
  assign n18981 = pi1316 & n15841;
  assign n18982 = pi1176 & n15843;
  assign n18983 = ~n18981 & ~n18982;
  assign n18984 = n18980 & n18983;
  assign n18985 = n18977 & n18984;
  assign n18986 = n18974 & n18985;
  assign n18987 = pi1218 & n15817;
  assign n18988 = pi1190 & n15819;
  assign n18989 = ~n18987 & ~n18988;
  assign n18990 = pi1288 & n15802;
  assign n18991 = pi1246 & n15806;
  assign n18992 = ~n18990 & ~n18991;
  assign n18993 = pi1274 & n15810;
  assign n18994 = pi1120 & n15812;
  assign n18995 = ~n18993 & ~n18994;
  assign n18996 = pi1162 & n15823;
  assign n18997 = pi1204 & n15825;
  assign n18998 = ~n18996 & ~n18997;
  assign n18999 = n18995 & n18998;
  assign n19000 = n18992 & n18999;
  assign n19001 = n18989 & n19000;
  assign n19002 = n18986 & n19001;
  assign n19003 = n15794 & ~n19002;
  assign n19004 = ~n9105 & n15940;
  assign n19005 = ~n19003 & ~n19004;
  assign n19006 = pi2392 & n15945;
  assign n19007 = ~n9105 & ~n15945;
  assign n19008 = ~n19006 & ~n19007;
  assign n19009 = n15944 & ~n19008;
  assign n19010 = pi0023 & n15993;
  assign n19011 = ~n19009 & ~n19010;
  assign n19012 = ~pi3432 & n16015;
  assign n19013 = pi3432 & ~n16015;
  assign n19014 = ~n19012 & ~n19013;
  assign n19015 = n16006 & ~n19014;
  assign n19016 = n19011 & ~n19015;
  assign n19017 = n19005 & n19016;
  assign n19018 = n18971 & n19017;
  assign n19019 = n15552 & ~n19018;
  assign n19020 = ~n18965 & ~n19019;
  assign n19021 = pi3514 & n8561;
  assign n19022 = pi0424 & ~n8561;
  assign po3840 = n19021 | n19022;
  assign n19024 = ~n16035 & po3840;
  assign n19025 = pi3432 & n16035;
  assign n19026 = ~n19024 & ~n19025;
  assign n19027 = n16034 & ~n19026;
  assign po0239 = ~n19020 | n19027;
  assign n19029 = n16013 & n18800;
  assign n19030 = pi3432 & n19029;
  assign n19031 = pi3455 & n19030;
  assign n19032 = pi3459 & n19031;
  assign n19033 = ~pi3459 & ~n19031;
  assign n19034 = ~n19032 & ~n19033;
  assign n19035 = n16006 & n19034;
  assign n19036 = pi1118 & n15846;
  assign n19037 = pi1314 & n15848;
  assign n19038 = ~n19036 & ~n19037;
  assign n19039 = pi1146 & n15831;
  assign n19040 = pi1160 & n15833;
  assign n19041 = ~n19039 & ~n19040;
  assign n19042 = pi1328 & n15841;
  assign n19043 = pi1188 & n15843;
  assign n19044 = ~n19042 & ~n19043;
  assign n19045 = pi1272 & n15836;
  assign n19046 = pi1244 & n15838;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = n19044 & n19047;
  assign n19049 = n19041 & n19048;
  assign n19050 = n19038 & n19049;
  assign n19051 = pi1174 & n15823;
  assign n19052 = pi1216 & n15825;
  assign n19053 = ~n19051 & ~n19052;
  assign n19054 = pi1300 & n15802;
  assign n19055 = pi1258 & n15806;
  assign n19056 = ~n19054 & ~n19055;
  assign n19057 = pi1230 & n15817;
  assign n19058 = pi1202 & n15819;
  assign n19059 = ~n19057 & ~n19058;
  assign n19060 = pi1286 & n15810;
  assign n19061 = pi1132 & n15812;
  assign n19062 = ~n19060 & ~n19061;
  assign n19063 = n19059 & n19062;
  assign n19064 = n19056 & n19063;
  assign n19065 = n19053 & n19064;
  assign n19066 = n19050 & n19065;
  assign n19067 = n15794 & ~n19066;
  assign n19068 = ~n9179 & n15940;
  assign n19069 = ~n19067 & ~n19068;
  assign n19070 = n15570 & n18697;
  assign n19071 = pi3420 & n19070;
  assign n19072 = pi3413 & n19071;
  assign n19073 = ~pi3401 & ~n19072;
  assign n19074 = pi3401 & n19072;
  assign n19075 = ~n19073 & ~n19074;
  assign n19076 = n15562 & n19075;
  assign n19077 = pi0817 & n15579;
  assign n19078 = ~n19076 & ~n19077;
  assign n19079 = pi2378 & n15945;
  assign n19080 = ~n9179 & ~n15945;
  assign n19081 = ~n19079 & ~n19080;
  assign n19082 = n15944 & ~n19081;
  assign n19083 = pi0024 & n15993;
  assign n19084 = ~n19082 & ~n19083;
  assign n19085 = n19078 & n19084;
  assign n19086 = n19069 & n19085;
  assign n19087 = ~n19035 & n19086;
  assign n19088 = n15552 & ~n19087;
  assign n19089 = pi0910 & n8589;
  assign n19090 = pi0781 & n16113;
  assign n19091 = ~n19089 & ~n19090;
  assign n19092 = po3841 & ~n19091;
  assign n19093 = ~n15552 & n19092;
  assign n19094 = ~n19088 & ~n19093;
  assign n19095 = pi3504 & n8561;
  assign n19096 = pi0423 & ~n8561;
  assign po3830 = n19095 | n19096;
  assign n19098 = ~n16035 & po3830;
  assign n19099 = pi3459 & n16035;
  assign n19100 = ~n19098 & ~n19099;
  assign n19101 = n16034 & ~n19100;
  assign po0240 = ~n19094 | n19101;
  assign n19103 = n16013 & n18875;
  assign n19104 = pi3459 & n19103;
  assign n19105 = pi3432 & n19104;
  assign n19106 = pi3478 & n19105;
  assign n19107 = ~pi3478 & ~n19105;
  assign n19108 = ~n19106 & ~n19107;
  assign n19109 = n16006 & n19108;
  assign n19110 = pi1229 & n15817;
  assign n19111 = pi1201 & n15819;
  assign n19112 = ~n19110 & ~n19111;
  assign n19113 = pi1299 & n15802;
  assign n19114 = pi1257 & n15806;
  assign n19115 = ~n19113 & ~n19114;
  assign n19116 = pi1173 & n15823;
  assign n19117 = pi1215 & n15825;
  assign n19118 = ~n19116 & ~n19117;
  assign n19119 = pi1285 & n15810;
  assign n19120 = pi1131 & n15812;
  assign n19121 = ~n19119 & ~n19120;
  assign n19122 = n19118 & n19121;
  assign n19123 = n19115 & n19122;
  assign n19124 = n19112 & n19123;
  assign n19125 = pi1327 & n15841;
  assign n19126 = pi1187 & n15843;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = pi1117 & n15846;
  assign n19129 = pi1313 & n15848;
  assign n19130 = ~n19128 & ~n19129;
  assign n19131 = pi1271 & n15836;
  assign n19132 = pi1243 & n15838;
  assign n19133 = ~n19131 & ~n19132;
  assign n19134 = pi1145 & n15831;
  assign n19135 = pi1159 & n15833;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = n19133 & n19136;
  assign n19138 = n19130 & n19137;
  assign n19139 = n19127 & n19138;
  assign n19140 = n19124 & n19139;
  assign n19141 = n15794 & ~n19140;
  assign n19142 = ~n9216 & n15940;
  assign n19143 = ~n19141 & ~n19142;
  assign n19144 = pi3401 & n15571;
  assign n19145 = pi3420 & n19144;
  assign n19146 = ~pi3422 & ~n19145;
  assign n19147 = pi3422 & n19145;
  assign n19148 = ~n19146 & ~n19147;
  assign n19149 = n15562 & n19148;
  assign n19150 = pi0816 & n15579;
  assign n19151 = ~n19149 & ~n19150;
  assign n19152 = pi2377 & n15945;
  assign n19153 = ~n9216 & ~n15945;
  assign n19154 = ~n19152 & ~n19153;
  assign n19155 = n15944 & ~n19154;
  assign n19156 = pi0025 & n15993;
  assign n19157 = ~n19155 & ~n19156;
  assign n19158 = n19151 & n19157;
  assign n19159 = n19143 & n19158;
  assign n19160 = ~n19109 & n19159;
  assign n19161 = n15552 & ~n19160;
  assign n19162 = pi0820 & n8589;
  assign n19163 = pi0780 & n16113;
  assign n19164 = ~n19162 & ~n19163;
  assign n19165 = po3841 & ~n19164;
  assign n19166 = ~n15552 & n19165;
  assign n19167 = ~n19161 & ~n19166;
  assign n19168 = pi3513 & n8561;
  assign n19169 = pi0422 & ~n8561;
  assign po3839 = n19168 | n19169;
  assign n19171 = ~n16035 & po3839;
  assign n19172 = pi3478 & n16035;
  assign n19173 = ~n19171 & ~n19172;
  assign n19174 = n16034 & ~n19173;
  assign po0241 = ~n19167 | n19174;
  assign n19176 = pi0434 & n8589;
  assign n19177 = pi0393 & ~n16215;
  assign n19178 = pi0844 & n16215;
  assign n19179 = ~n19177 & ~n19178;
  assign n19180 = ~n8589 & ~n19179;
  assign po0244 = n19176 | n19180;
  assign n19182 = pi0433 & n8589;
  assign n19183 = pi0390 & ~n16215;
  assign n19184 = pi0843 & n16215;
  assign n19185 = ~n19183 & ~n19184;
  assign n19186 = ~n8589 & ~n19185;
  assign po0245 = n19182 | n19186;
  assign n19188 = pi0432 & n8589;
  assign n19189 = pi0389 & ~n16215;
  assign n19190 = pi0842 & n16215;
  assign n19191 = ~n19189 & ~n19190;
  assign n19192 = ~n8589 & ~n19191;
  assign po0246 = n19188 | n19192;
  assign n19194 = pi0431 & n8589;
  assign n19195 = pi0388 & ~n16215;
  assign n19196 = pi0864 & n16215;
  assign n19197 = ~n19195 & ~n19196;
  assign n19198 = ~n8589 & ~n19197;
  assign po0247 = n19194 | n19198;
  assign n19200 = pi0430 & n8589;
  assign n19201 = pi0387 & ~n16215;
  assign n19202 = pi0841 & n16215;
  assign n19203 = ~n19201 & ~n19202;
  assign n19204 = ~n8589 & ~n19203;
  assign po0248 = n19200 | n19204;
  assign n19206 = pi0429 & n8589;
  assign n19207 = pi0386 & ~n16215;
  assign n19208 = pi0865 & n16215;
  assign n19209 = ~n19207 & ~n19208;
  assign n19210 = ~n8589 & ~n19209;
  assign po0249 = n19206 | n19210;
  assign n19212 = pi0428 & n8589;
  assign n19213 = pi0385 & ~n16215;
  assign n19214 = pi0840 & n16215;
  assign n19215 = ~n19213 & ~n19214;
  assign n19216 = ~n8589 & ~n19215;
  assign po0250 = n19212 | n19216;
  assign n19218 = pi0435 & n8589;
  assign n19219 = pi0384 & ~n16215;
  assign n19220 = pi0839 & n16215;
  assign n19221 = ~n19219 & ~n19220;
  assign n19222 = ~n8589 & ~n19221;
  assign po0251 = n19218 | n19222;
  assign n19224 = pi0366 & n8589;
  assign n19225 = pi0383 & ~n16215;
  assign n19226 = pi1092 & n16215;
  assign n19227 = ~n19225 & ~n19226;
  assign n19228 = ~n8589 & ~n19227;
  assign po0252 = n19224 | n19228;
  assign n19230 = pi0359 & n8589;
  assign n19231 = pi0382 & ~n16215;
  assign n19232 = pi1060 & n16215;
  assign n19233 = ~n19231 & ~n19232;
  assign n19234 = ~n8589 & ~n19233;
  assign po0253 = n19230 | n19234;
  assign n19236 = pi0358 & n8589;
  assign n19237 = pi0392 & ~n16215;
  assign n19238 = pi1089 & n16215;
  assign n19239 = ~n19237 & ~n19238;
  assign n19240 = ~n8589 & ~n19239;
  assign po0254 = n19236 | n19240;
  assign n19242 = pi0357 & n8589;
  assign n19243 = pi0391 & ~n16215;
  assign n19244 = pi1065 & n16215;
  assign n19245 = ~n19243 & ~n19244;
  assign n19246 = ~n8589 & ~n19245;
  assign po0255 = n19242 | n19246;
  assign n19248 = pi0356 & n8589;
  assign n19249 = pi0381 & ~n16215;
  assign n19250 = pi1064 & n16215;
  assign n19251 = ~n19249 & ~n19250;
  assign n19252 = ~n8589 & ~n19251;
  assign po0256 = n19248 | n19252;
  assign n19254 = pi0355 & n8589;
  assign n19255 = pi0378 & ~n16215;
  assign n19256 = pi1063 & n16215;
  assign n19257 = ~n19255 & ~n19256;
  assign n19258 = ~n8589 & ~n19257;
  assign po0257 = n19254 | n19258;
  assign n19260 = pi0354 & n8589;
  assign n19261 = pi0377 & ~n16215;
  assign n19262 = pi1062 & n16215;
  assign n19263 = ~n19261 & ~n19262;
  assign n19264 = ~n8589 & ~n19263;
  assign po0258 = n19260 | n19264;
  assign n19266 = pi0353 & n8589;
  assign n19267 = pi0376 & ~n16215;
  assign n19268 = pi1061 & n16215;
  assign n19269 = ~n19267 & ~n19268;
  assign n19270 = ~n8589 & ~n19269;
  assign po0259 = n19266 | n19270;
  assign n19272 = pi0352 & n8589;
  assign n19273 = pi0375 & ~n16215;
  assign n19274 = pi3106 & n16215;
  assign n19275 = ~n19273 & ~n19274;
  assign n19276 = ~n8589 & ~n19275;
  assign po0260 = n19272 | n19276;
  assign n19278 = pi0351 & n8589;
  assign n19279 = pi0374 & ~n16215;
  assign n19280 = pi3105 & n16215;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~n8589 & ~n19281;
  assign po0261 = n19278 | n19282;
  assign n19284 = pi0365 & n8589;
  assign n19285 = pi0373 & ~n16215;
  assign n19286 = pi3104 & n16215;
  assign n19287 = ~n19285 & ~n19286;
  assign n19288 = ~n8589 & ~n19287;
  assign po0262 = n19284 | n19288;
  assign n19290 = pi0364 & n8589;
  assign n19291 = pi0372 & ~n16215;
  assign n19292 = pi2985 & n16215;
  assign n19293 = ~n19291 & ~n19292;
  assign n19294 = ~n8589 & ~n19293;
  assign po0263 = n19290 | n19294;
  assign n19296 = pi0363 & n8589;
  assign n19297 = pi0371 & ~n16215;
  assign n19298 = pi3102 & n16215;
  assign n19299 = ~n19297 & ~n19298;
  assign n19300 = ~n8589 & ~n19299;
  assign po0264 = n19296 | n19300;
  assign n19302 = pi0362 & n8589;
  assign n19303 = pi0369 & ~n16215;
  assign n19304 = pi3109 & n16215;
  assign n19305 = ~n19303 & ~n19304;
  assign n19306 = ~n8589 & ~n19305;
  assign po0265 = n19302 | n19306;
  assign n19308 = pi0361 & n8589;
  assign n19309 = pi0380 & ~n16215;
  assign n19310 = pi3111 & n16215;
  assign n19311 = ~n19309 & ~n19310;
  assign n19312 = ~n8589 & ~n19311;
  assign po0266 = n19308 | n19312;
  assign n19314 = pi0360 & n8589;
  assign n19315 = pi0379 & ~n16215;
  assign n19316 = pi3112 & n16215;
  assign n19317 = ~n19315 & ~n19316;
  assign n19318 = ~n8589 & ~n19317;
  assign po0267 = n19314 | n19318;
  assign n19320 = pi3460 & n15546;
  assign n19321 = ~n15546 & ~n18379;
  assign po0268 = n19320 | n19321;
  assign n19323 = pi3437 & n15546;
  assign n19324 = ~n15546 & ~n18452;
  assign po0269 = n19323 | n19324;
  assign n19326 = pi3433 & n15546;
  assign n19327 = ~n15546 & ~n18526;
  assign po0270 = n19326 | n19327;
  assign n19329 = pi3457 & n15546;
  assign n19330 = ~n15546 & ~n18599;
  assign po0271 = n19329 | n19330;
  assign n19332 = pi3456 & n15546;
  assign n19333 = ~n15546 & ~n18665;
  assign po0272 = n19332 | n19333;
  assign n19335 = ~pi3114 & pi3118;
  assign n19336 = ~n8670 & ~n19335;
  assign n19337 = pi3114 & ~pi3118;
  assign po0278 = n19336 | n19337;
  assign n19339 = ~pi3114 & ~pi3118;
  assign n19340 = ~n8670 & ~n19339;
  assign n19341 = pi3114 & pi3118;
  assign po0279 = n19340 | n19341;
  assign n19343 = pi2952 & ~pi3209;
  assign n19344 = ~pi2763 & ~n19343;
  assign n19345 = pi2951 & ~pi3076;
  assign n19346 = n8670 & n19345;
  assign n19347 = ~n8670 & n19345;
  assign n19348 = ~n19346 & ~n19347;
  assign n19349 = pi2951 & pi3076;
  assign n19350 = n8670 & n19349;
  assign n19351 = ~n8670 & n19349;
  assign n19352 = ~n8670 & ~n9265;
  assign n19353 = n8670 & ~n9336;
  assign n19354 = ~n19352 & ~n19353;
  assign n19355 = n19351 & ~n19354;
  assign n19356 = n19351 & n19354;
  assign n19357 = ~n19355 & ~n19356;
  assign n19358 = ~n19350 & n19357;
  assign n19359 = n19348 & n19358;
  assign n19360 = pi3209 & ~n19359;
  assign n19361 = pi2951 & ~n19360;
  assign n19362 = pi2763 & ~n19361;
  assign po0280 = n19344 | n19362;
  assign n19364 = pi3208 & ~n19359;
  assign n19365 = ~pi2951 & pi3405;
  assign n19366 = ~n19364 & ~n19365;
  assign n19367 = pi2763 & ~n19366;
  assign n19368 = pi2952 & pi3208;
  assign n19369 = ~pi2952 & pi3405;
  assign n19370 = ~n19368 & ~n19369;
  assign n19371 = ~pi2763 & ~n19370;
  assign po0281 = n19367 | n19371;
  assign n19373 = pi3235 & ~n19359;
  assign n19374 = ~pi2951 & pi3413;
  assign n19375 = ~n19373 & ~n19374;
  assign n19376 = pi2763 & ~n19375;
  assign n19377 = pi2952 & pi3235;
  assign n19378 = ~pi2952 & pi3413;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = ~pi2763 & ~n19379;
  assign po0282 = n19376 | n19380;
  assign n19382 = pi3234 & ~n19359;
  assign n19383 = ~pi2951 & pi3406;
  assign n19384 = ~n19382 & ~n19383;
  assign n19385 = pi2763 & ~n19384;
  assign n19386 = pi2952 & pi3234;
  assign n19387 = ~pi2952 & pi3406;
  assign n19388 = ~n19386 & ~n19387;
  assign n19389 = ~pi2763 & ~n19388;
  assign po0283 = n19385 | n19389;
  assign n19391 = pi3207 & ~n19359;
  assign n19392 = ~pi2951 & pi3411;
  assign n19393 = ~n19391 & ~n19392;
  assign n19394 = pi2763 & ~n19393;
  assign n19395 = pi2952 & pi3207;
  assign n19396 = ~pi2952 & pi3411;
  assign n19397 = ~n19395 & ~n19396;
  assign n19398 = ~pi2763 & ~n19397;
  assign po0284 = n19394 | n19398;
  assign n19400 = pi3206 & ~n19359;
  assign n19401 = ~pi2951 & pi3420;
  assign n19402 = ~n19400 & ~n19401;
  assign n19403 = pi2763 & ~n19402;
  assign n19404 = pi2952 & pi3206;
  assign n19405 = ~pi2952 & pi3420;
  assign n19406 = ~n19404 & ~n19405;
  assign n19407 = ~pi2763 & ~n19406;
  assign po0285 = n19403 | n19407;
  assign n19409 = pi3231 & ~n19359;
  assign n19410 = ~pi2951 & pi3401;
  assign n19411 = ~n19409 & ~n19410;
  assign n19412 = pi2763 & ~n19411;
  assign n19413 = pi2952 & pi3231;
  assign n19414 = ~pi2952 & pi3401;
  assign n19415 = ~n19413 & ~n19414;
  assign n19416 = ~pi2763 & ~n19415;
  assign po0286 = n19412 | n19416;
  assign n19418 = pi3230 & ~n19359;
  assign n19419 = ~pi2951 & pi3422;
  assign n19420 = ~n19418 & ~n19419;
  assign n19421 = pi2763 & ~n19420;
  assign n19422 = pi2952 & pi3230;
  assign n19423 = ~pi2952 & pi3422;
  assign n19424 = ~n19422 & ~n19423;
  assign n19425 = ~pi2763 & ~n19424;
  assign po0287 = n19421 | n19425;
  assign n19427 = pi3229 & ~n19359;
  assign n19428 = ~pi2951 & pi3421;
  assign n19429 = ~n19427 & ~n19428;
  assign n19430 = pi2763 & ~n19429;
  assign n19431 = pi2952 & pi3229;
  assign n19432 = ~pi2952 & pi3421;
  assign n19433 = ~n19431 & ~n19432;
  assign n19434 = ~pi2763 & ~n19433;
  assign po0288 = n19430 | n19434;
  assign n19436 = pi3228 & ~n19359;
  assign n19437 = ~pi2951 & pi3430;
  assign n19438 = ~n19436 & ~n19437;
  assign n19439 = pi2763 & ~n19438;
  assign n19440 = ~pi2952 & pi3430;
  assign n19441 = pi2952 & pi3228;
  assign n19442 = ~n19440 & ~n19441;
  assign n19443 = ~pi2763 & ~n19442;
  assign po0289 = n19439 | n19443;
  assign n19445 = ~pi2952 & n8670;
  assign n19446 = ~n9352 & ~n19445;
  assign po0290 = ~pi3121 | ~n19446;
  assign n19448 = pi1930 & ~pi2492;
  assign po0291 = ~pi0939 & n19448;
  assign n19450 = ~n19347 & ~n19355;
  assign n19451 = pi2951 & n19450;
  assign n19452 = ~n18373 & ~n19451;
  assign n19453 = ~n19350 & ~n19356;
  assign n19454 = ~n19346 & n19453;
  assign n19455 = pi3195 & ~n19454;
  assign n19456 = ~n19452 & ~n19455;
  assign n19457 = pi2763 & ~n19456;
  assign n19458 = ~pi2763 & pi2952;
  assign n19459 = pi3195 & n19458;
  assign po0293 = n19457 | n19459;
  assign n19461 = pi3124 & ~n19454;
  assign n19462 = ~n18442 & ~n19451;
  assign n19463 = ~n19461 & ~n19462;
  assign n19464 = pi2763 & ~n19463;
  assign n19465 = pi3124 & n19458;
  assign po0294 = n19464 | n19465;
  assign n19467 = ~n18481 & ~n19451;
  assign n19468 = pi3194 & ~n19454;
  assign n19469 = ~n19467 & ~n19468;
  assign n19470 = pi2763 & ~n19469;
  assign n19471 = pi3194 & n19458;
  assign po0295 = n19470 | n19471;
  assign n19473 = pi3139 & ~n19454;
  assign n19474 = ~n18554 & ~n19451;
  assign n19475 = ~n19473 & ~n19474;
  assign n19476 = pi2763 & ~n19475;
  assign n19477 = pi3139 & n19458;
  assign po0296 = n19476 | n19477;
  assign n19479 = ~n18612 & ~n19451;
  assign n19480 = pi3135 & ~n19454;
  assign n19481 = ~n19479 & ~n19480;
  assign n19482 = pi2763 & ~n19481;
  assign n19483 = pi3135 & n19458;
  assign po0297 = n19482 | n19483;
  assign n19485 = ~n18683 & ~n19451;
  assign n19486 = pi3187 & ~n19454;
  assign n19487 = ~n19485 & ~n19486;
  assign n19488 = pi2763 & ~n19487;
  assign n19489 = pi3187 & n19458;
  assign po0298 = n19488 | n19489;
  assign n19491 = pi3193 & ~n19454;
  assign n19492 = ~n18795 & ~n19451;
  assign n19493 = ~n19491 & ~n19492;
  assign n19494 = pi2763 & ~n19493;
  assign n19495 = pi3193 & n19458;
  assign po0299 = n19494 | n19495;
  assign n19497 = pi3192 & ~n19454;
  assign n19498 = ~n18869 & ~n19451;
  assign n19499 = ~n19497 & ~n19498;
  assign n19500 = pi2763 & ~n19499;
  assign n19501 = pi3192 & n19458;
  assign po0300 = n19500 | n19501;
  assign n19503 = ~n18940 & ~n19451;
  assign n19504 = pi3117 & ~n19454;
  assign n19505 = ~n19503 & ~n19504;
  assign n19506 = pi2763 & ~n19505;
  assign n19507 = pi3117 & n19458;
  assign po0301 = n19506 | n19507;
  assign n19509 = ~n19008 & ~n19451;
  assign n19510 = pi3116 & ~n19454;
  assign n19511 = ~n19509 & ~n19510;
  assign n19512 = pi2763 & ~n19511;
  assign n19513 = pi3116 & n19458;
  assign po0302 = n19512 | n19513;
  assign n19515 = pi3198 & ~n19454;
  assign n19516 = ~n19081 & ~n19451;
  assign n19517 = ~n19515 & ~n19516;
  assign n19518 = pi2763 & ~n19517;
  assign n19519 = pi3198 & n19458;
  assign po0303 = n19518 | n19519;
  assign n19521 = pi3115 & ~n19454;
  assign n19522 = ~n19154 & ~n19451;
  assign n19523 = ~n19521 & ~n19522;
  assign n19524 = pi2763 & ~n19523;
  assign n19525 = pi3115 & n19458;
  assign po0304 = n19524 | n19525;
  assign n19527 = ~n16104 & ~n19451;
  assign n19528 = pi3197 & ~n19454;
  assign n19529 = ~n19527 & ~n19528;
  assign n19530 = pi2763 & ~n19529;
  assign n19531 = pi3197 & n19458;
  assign po0305 = n19530 | n19531;
  assign n19533 = pi3196 & ~n19454;
  assign n19534 = ~n15948 & ~n19451;
  assign n19535 = ~n19533 & ~n19534;
  assign n19536 = pi2763 & ~n19535;
  assign n19537 = pi3196 & n19458;
  assign po0306 = n19536 | n19537;
  assign n19539 = pi2763 & pi2951;
  assign n19540 = ~n15945 & ~n19539;
  assign po0307 = n9352 | n19540;
  assign n19542 = pi0038 & n8561;
  assign n19543 = ~pi0835 & n9365;
  assign n19544 = ~pi2487 & ~pi3330;
  assign n19545 = ~pi3394 & n19544;
  assign n19546 = pi3210 & ~n8670;
  assign n19547 = ~n19545 & ~n19546;
  assign n19548 = ~pi1042 & ~pi1093;
  assign n19549 = ~pi1041 & n19548;
  assign n19550 = ~n19547 & ~n19549;
  assign n19551 = ~n9352 & n19550;
  assign n19552 = ~pi1824 & n8670;
  assign n19553 = ~pi3426 & ~n19552;
  assign n19554 = ~pi2142 & n19553;
  assign n19555 = ~n9352 & n19554;
  assign n19556 = ~n19551 & ~n19555;
  assign n19557 = ~n19543 & n19556;
  assign n19558 = ~pi0407 & ~pi0414;
  assign n19559 = pi0415 & pi0427;
  assign n19560 = n19558 & n19559;
  assign n19561 = pi1974 & ~pi1975;
  assign n19562 = pi1972 & ~pi1973;
  assign n19563 = n19561 & n19562;
  assign n19564 = ~pi1974 & pi1975;
  assign n19565 = n19562 & n19564;
  assign n19566 = ~n19563 & ~n19565;
  assign n19567 = ~pi1974 & ~pi1975;
  assign n19568 = n19562 & n19567;
  assign n19569 = pi2758 & pi3065;
  assign n19570 = pi2142 & n19569;
  assign n19571 = pi1974 & pi1975;
  assign n19572 = n19562 & n19571;
  assign n19573 = ~n19570 & ~n19572;
  assign n19574 = ~n19568 & n19573;
  assign n19575 = n19566 & n19574;
  assign n19576 = ~pi1972 & pi1973;
  assign n19577 = n19567 & n19576;
  assign n19578 = ~pi1972 & ~pi1973;
  assign n19579 = n19567 & n19578;
  assign n19580 = ~n19570 & ~n19579;
  assign n19581 = ~n19577 & n19580;
  assign n19582 = ~pi3520 & ~pi3521;
  assign n19583 = ~pi3510 & n19582;
  assign n19584 = ~pi3511 & n19583;
  assign n19585 = ~pi2982 & ~n19584;
  assign n19586 = pi1793 & n19585;
  assign n19587 = ~pi3516 & pi3518;
  assign n19588 = pi3518 & n19587;
  assign n19589 = ~pi0230 & pi0979;
  assign n19590 = ~pi0231 & ~pi0979;
  assign n19591 = ~n19589 & ~n19590;
  assign n19592 = n19588 & ~n19591;
  assign n19593 = pi3516 & ~n17230;
  assign n19594 = ~pi3516 & ~n17234;
  assign n19595 = ~n19593 & ~n19594;
  assign n19596 = ~pi3518 & ~n19595;
  assign n19597 = ~n19592 & ~n19596;
  assign n19598 = ~n19585 & n19597;
  assign n19599 = ~n19586 & ~n19598;
  assign n19600 = n19581 & n19599;
  assign n19601 = n19575 & ~n19600;
  assign n19602 = ~n19575 & n19600;
  assign n19603 = ~n19601 & ~n19602;
  assign n19604 = ~pi3509 & ~n17243;
  assign n19605 = pi3509 & ~n17239;
  assign n19606 = ~n19604 & ~n19605;
  assign n19607 = ~pi3508 & ~pi3517;
  assign n19608 = ~n19606 & n19607;
  assign n19609 = ~pi3508 & pi3517;
  assign n19610 = pi3509 & n19609;
  assign n19611 = ~n9498 & n19610;
  assign n19612 = ~pi3509 & n19609;
  assign n19613 = ~n17327 & n19612;
  assign n19614 = pi3508 & pi3509;
  assign n19615 = ~pi3517 & n19614;
  assign n19616 = ~n17331 & n19615;
  assign n19617 = ~n19613 & ~n19616;
  assign n19618 = pi3508 & ~pi3509;
  assign n19619 = ~pi3517 & n19618;
  assign n19620 = ~n17248 & n19619;
  assign n19621 = ~pi3509 & ~n17221;
  assign n19622 = pi3509 & ~n17217;
  assign n19623 = ~n19621 & ~n19622;
  assign n19624 = pi3508 & pi3517;
  assign n19625 = ~n19623 & n19624;
  assign n19626 = ~n19620 & ~n19625;
  assign n19627 = n19617 & n19626;
  assign n19628 = ~n19611 & n19627;
  assign n19629 = ~n19607 & ~n19628;
  assign n19630 = ~n19608 & ~n19629;
  assign n19631 = n19564 & n19576;
  assign n19632 = pi1974 & n19576;
  assign n19633 = pi3065 & n19632;
  assign n19634 = pi1975 & n19633;
  assign n19635 = n19561 & n19576;
  assign n19636 = ~n19634 & ~n19635;
  assign n19637 = ~n19631 & n19636;
  assign n19638 = ~pi0143 & ~pi3065;
  assign n19639 = ~n19577 & ~n19638;
  assign n19640 = ~n19570 & n19639;
  assign n19641 = n19637 & n19640;
  assign n19642 = n19630 & ~n19641;
  assign n19643 = n19580 & n19639;
  assign n19644 = n19637 & n19643;
  assign n19645 = ~n19630 & ~n19644;
  assign n19646 = ~n19642 & ~n19645;
  assign n19647 = pi1973 & pi1974;
  assign n19648 = pi1972 & n19647;
  assign n19649 = pi1975 & n19648;
  assign n19650 = ~n19634 & ~n19649;
  assign n19651 = ~pi1975 & n19648;
  assign n19652 = n19650 & ~n19651;
  assign n19653 = ~n19572 & n19652;
  assign n19654 = ~n19563 & n19653;
  assign n19655 = ~n19570 & n19654;
  assign n19656 = ~pi3509 & ~n17040;
  assign n19657 = pi3509 & ~n17036;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = n19607 & ~n19658;
  assign n19660 = ~n17045 & n19619;
  assign n19661 = ~pi3509 & ~n17018;
  assign n19662 = pi3509 & ~n17014;
  assign n19663 = ~n19661 & ~n19662;
  assign n19664 = n19624 & ~n19663;
  assign n19665 = ~n19660 & ~n19664;
  assign n19666 = ~n17071 & n19612;
  assign n19667 = ~n17075 & n19615;
  assign n19668 = ~n19666 & ~n19667;
  assign n19669 = n19665 & n19668;
  assign n19670 = ~n19611 & n19669;
  assign n19671 = ~n19607 & ~n19670;
  assign n19672 = ~n19659 & ~n19671;
  assign n19673 = n19655 & ~n19672;
  assign n19674 = ~n19646 & ~n19673;
  assign n19675 = n19646 & n19673;
  assign n19676 = ~n19674 & ~n19675;
  assign n19677 = pi1794 & n19585;
  assign n19678 = ~pi0242 & pi0979;
  assign n19679 = ~pi0244 & ~pi0979;
  assign n19680 = ~n19678 & ~n19679;
  assign n19681 = n19588 & ~n19680;
  assign n19682 = ~pi3516 & ~n17031;
  assign n19683 = pi3516 & ~n17027;
  assign n19684 = ~n19682 & ~n19683;
  assign n19685 = ~pi3518 & ~n19684;
  assign n19686 = ~n19681 & ~n19685;
  assign n19687 = ~n19585 & n19686;
  assign n19688 = ~n19677 & ~n19687;
  assign n19689 = n19581 & n19688;
  assign n19690 = n19575 & ~n19689;
  assign n19691 = ~n19575 & n19689;
  assign n19692 = ~n19690 & ~n19691;
  assign n19693 = ~n19676 & n19692;
  assign n19694 = ~pi3509 & ~n15303;
  assign n19695 = pi3509 & ~n15299;
  assign n19696 = ~n19694 & ~n19695;
  assign n19697 = n19607 & ~n19696;
  assign n19698 = ~n15259 & n19612;
  assign n19699 = ~n15263 & n19615;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = ~n15308 & n19619;
  assign n19702 = ~pi3509 & ~n15281;
  assign n19703 = pi3509 & ~n15277;
  assign n19704 = ~n19702 & ~n19703;
  assign n19705 = n19624 & ~n19704;
  assign n19706 = ~n19701 & ~n19705;
  assign n19707 = n19700 & n19706;
  assign n19708 = ~n19611 & n19707;
  assign n19709 = ~n19607 & ~n19708;
  assign n19710 = ~n19697 & ~n19709;
  assign n19711 = n19655 & ~n19710;
  assign n19712 = n19646 & ~n19711;
  assign n19713 = ~n19646 & n19711;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = pi2081 & n19585;
  assign n19716 = ~pi0274 & pi0979;
  assign n19717 = ~pi0276 & ~pi0979;
  assign n19718 = ~n19716 & ~n19717;
  assign n19719 = n19588 & ~n19718;
  assign n19720 = ~pi3516 & ~n15294;
  assign n19721 = pi3516 & ~n15290;
  assign n19722 = ~n19720 & ~n19721;
  assign n19723 = ~pi3518 & ~n19722;
  assign n19724 = ~n19719 & ~n19723;
  assign n19725 = ~n19585 & n19724;
  assign n19726 = ~n19715 & ~n19725;
  assign n19727 = n19581 & n19726;
  assign n19728 = n19575 & ~n19727;
  assign n19729 = ~n19575 & n19727;
  assign n19730 = ~n19728 & ~n19729;
  assign n19731 = n19714 & n19730;
  assign n19732 = ~n12547 & n19619;
  assign n19733 = pi3509 & ~n12516;
  assign n19734 = ~pi3509 & ~n12520;
  assign n19735 = ~n19733 & ~n19734;
  assign n19736 = n19624 & ~n19735;
  assign n19737 = ~n19732 & ~n19736;
  assign n19738 = ~n19611 & n19737;
  assign n19739 = ~n12609 & n19612;
  assign n19740 = ~n12613 & n19615;
  assign n19741 = ~n19739 & ~n19740;
  assign n19742 = n19738 & n19741;
  assign n19743 = ~n19607 & ~n19742;
  assign n19744 = ~pi3509 & ~n12529;
  assign n19745 = pi3509 & ~n12533;
  assign n19746 = ~n19744 & ~n19745;
  assign n19747 = n19607 & ~n19746;
  assign n19748 = ~n19743 & ~n19747;
  assign n19749 = n19655 & ~n19748;
  assign n19750 = ~n19646 & ~n19749;
  assign n19751 = n19646 & n19749;
  assign n19752 = ~n19750 & ~n19751;
  assign n19753 = pi2194 & n19585;
  assign n19754 = ~pi0301 & pi0979;
  assign n19755 = ~pi0302 & ~pi0979;
  assign n19756 = ~n19754 & ~n19755;
  assign n19757 = n19588 & ~n19756;
  assign n19758 = ~pi3516 & ~n12542;
  assign n19759 = pi3516 & ~n12538;
  assign n19760 = ~n19758 & ~n19759;
  assign n19761 = ~pi3518 & ~n19760;
  assign n19762 = ~n19757 & ~n19761;
  assign n19763 = ~n19585 & n19762;
  assign n19764 = ~n19753 & ~n19763;
  assign n19765 = n19581 & n19764;
  assign n19766 = n19575 & ~n19765;
  assign n19767 = ~n19575 & n19765;
  assign n19768 = ~n19766 & ~n19767;
  assign n19769 = n19752 & ~n19768;
  assign n19770 = ~pi3509 & ~n14272;
  assign n19771 = pi3509 & ~n14268;
  assign n19772 = ~n19770 & ~n19771;
  assign n19773 = n19607 & ~n19772;
  assign n19774 = ~n14219 & n19612;
  assign n19775 = ~n14223 & n19615;
  assign n19776 = ~n19774 & ~n19775;
  assign n19777 = ~n19611 & n19776;
  assign n19778 = ~n14286 & n19619;
  assign n19779 = pi3509 & ~n14255;
  assign n19780 = ~pi3509 & ~n14259;
  assign n19781 = ~n19779 & ~n19780;
  assign n19782 = n19624 & ~n19781;
  assign n19783 = ~n19778 & ~n19782;
  assign n19784 = n19777 & n19783;
  assign n19785 = ~n19607 & ~n19784;
  assign n19786 = ~n19773 & ~n19785;
  assign n19787 = n19655 & ~n19786;
  assign n19788 = ~n19646 & ~n19787;
  assign n19789 = n19646 & n19787;
  assign n19790 = ~n19788 & ~n19789;
  assign n19791 = pi2080 & n19585;
  assign n19792 = ~pi0295 & pi0979;
  assign n19793 = ~pi0296 & ~pi0979;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = n19588 & ~n19794;
  assign n19796 = ~pi3516 & ~n14277;
  assign n19797 = pi3516 & ~n14281;
  assign n19798 = ~n19796 & ~n19797;
  assign n19799 = ~pi3518 & ~n19798;
  assign n19800 = ~n19795 & ~n19799;
  assign n19801 = ~n19585 & n19800;
  assign n19802 = ~n19791 & ~n19801;
  assign n19803 = n19581 & n19802;
  assign n19804 = n19575 & ~n19803;
  assign n19805 = ~n19575 & n19803;
  assign n19806 = ~n19804 & ~n19805;
  assign n19807 = ~n19790 & n19806;
  assign n19808 = ~n19769 & n19807;
  assign n19809 = ~n19731 & ~n19808;
  assign n19810 = ~n19752 & n19768;
  assign n19811 = ~n19714 & ~n19730;
  assign n19812 = ~pi3509 & ~n13569;
  assign n19813 = pi3509 & ~n13565;
  assign n19814 = ~n19812 & ~n19813;
  assign n19815 = n19607 & ~n19814;
  assign n19816 = ~n13534 & n19612;
  assign n19817 = ~n13538 & n19615;
  assign n19818 = ~n19816 & ~n19817;
  assign n19819 = ~n13583 & n19619;
  assign n19820 = pi3509 & ~n13552;
  assign n19821 = ~pi3509 & ~n13556;
  assign n19822 = ~n19820 & ~n19821;
  assign n19823 = n19624 & ~n19822;
  assign n19824 = ~n19611 & ~n19823;
  assign n19825 = ~n19819 & n19824;
  assign n19826 = n19818 & n19825;
  assign n19827 = ~n19607 & ~n19826;
  assign n19828 = ~n19815 & ~n19827;
  assign n19829 = n19655 & ~n19828;
  assign n19830 = ~n19646 & ~n19829;
  assign n19831 = n19646 & n19829;
  assign n19832 = ~n19830 & ~n19831;
  assign n19833 = pi2086 & n19585;
  assign n19834 = ~pi0321 & pi0979;
  assign n19835 = ~pi0322 & ~pi0979;
  assign n19836 = ~n19834 & ~n19835;
  assign n19837 = n19588 & ~n19836;
  assign n19838 = ~pi3516 & ~n13578;
  assign n19839 = pi3516 & ~n13574;
  assign n19840 = ~n19838 & ~n19839;
  assign n19841 = ~pi3518 & ~n19840;
  assign n19842 = ~n19837 & ~n19841;
  assign n19843 = ~n19585 & n19842;
  assign n19844 = ~n19833 & ~n19843;
  assign n19845 = n19581 & n19844;
  assign n19846 = ~n19575 & n19845;
  assign n19847 = n19575 & ~n19845;
  assign n19848 = ~n19846 & ~n19847;
  assign n19849 = ~n19832 & n19848;
  assign n19850 = ~n19811 & n19849;
  assign n19851 = ~n19810 & ~n19850;
  assign n19852 = n19790 & ~n19806;
  assign n19853 = ~n19811 & ~n19852;
  assign n19854 = ~n19851 & n19853;
  assign n19855 = n19809 & ~n19854;
  assign n19856 = ~n9511 & n19612;
  assign n19857 = ~n9515 & n19615;
  assign n19858 = ~n19856 & ~n19857;
  assign n19859 = ~n9570 & n19619;
  assign n19860 = ~pi3509 & ~n9542;
  assign n19861 = pi3509 & ~n9538;
  assign n19862 = ~n19860 & ~n19861;
  assign n19863 = n19624 & ~n19862;
  assign n19864 = ~n19859 & ~n19863;
  assign n19865 = n19858 & n19864;
  assign n19866 = ~n19611 & n19865;
  assign n19867 = ~n19607 & ~n19866;
  assign n19868 = ~pi3509 & ~n9565;
  assign n19869 = pi3509 & ~n9561;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = n19607 & ~n19870;
  assign n19872 = ~n19867 & ~n19871;
  assign n19873 = n19655 & ~n19872;
  assign n19874 = n19646 & n19873;
  assign n19875 = ~n19646 & n19872;
  assign n19876 = ~n19874 & ~n19875;
  assign n19877 = ~n19646 & ~n19655;
  assign n19878 = n19876 & ~n19877;
  assign n19879 = ~pi1795 & n19585;
  assign n19880 = ~pi3516 & ~n9556;
  assign n19881 = pi3516 & ~n9552;
  assign n19882 = ~n19880 & ~n19881;
  assign n19883 = ~pi3518 & ~n19882;
  assign n19884 = ~pi0243 & pi0979;
  assign n19885 = ~pi0245 & ~pi0979;
  assign n19886 = ~n19884 & ~n19885;
  assign n19887 = n19588 & ~n19886;
  assign n19888 = ~n19883 & ~n19887;
  assign n19889 = ~n19585 & ~n19888;
  assign n19890 = ~n19879 & ~n19889;
  assign n19891 = ~n19575 & n19890;
  assign n19892 = n19575 & n19581;
  assign n19893 = ~n19890 & n19892;
  assign n19894 = ~n19891 & ~n19893;
  assign n19895 = ~n19575 & ~n19581;
  assign n19896 = n19894 & ~n19895;
  assign n19897 = n19878 & n19896;
  assign n19898 = ~pi3509 & ~n10473;
  assign n19899 = pi3509 & ~n10469;
  assign n19900 = ~n19898 & ~n19899;
  assign n19901 = n19607 & ~n19900;
  assign n19902 = ~n10420 & n19612;
  assign n19903 = ~n10424 & n19615;
  assign n19904 = ~n19902 & ~n19903;
  assign n19905 = ~n10487 & n19619;
  assign n19906 = ~pi3509 & ~n10460;
  assign n19907 = pi3509 & ~n10456;
  assign n19908 = ~n19906 & ~n19907;
  assign n19909 = n19624 & ~n19908;
  assign n19910 = ~n19905 & ~n19909;
  assign n19911 = n19904 & n19910;
  assign n19912 = ~n19611 & n19911;
  assign n19913 = ~n19607 & ~n19912;
  assign n19914 = ~n19901 & ~n19913;
  assign n19915 = n19655 & ~n19914;
  assign n19916 = ~n19646 & ~n19915;
  assign n19917 = n19646 & n19915;
  assign n19918 = ~n19916 & ~n19917;
  assign n19919 = pi1796 & n19585;
  assign n19920 = ~pi0273 & pi0979;
  assign n19921 = ~pi0275 & ~pi0979;
  assign n19922 = ~n19920 & ~n19921;
  assign n19923 = n19588 & ~n19922;
  assign n19924 = ~pi3516 & ~n10482;
  assign n19925 = pi3516 & ~n10478;
  assign n19926 = ~n19924 & ~n19925;
  assign n19927 = ~pi3518 & ~n19926;
  assign n19928 = ~n19923 & ~n19927;
  assign n19929 = ~n19585 & n19928;
  assign n19930 = ~n19919 & ~n19929;
  assign n19931 = n19581 & n19930;
  assign n19932 = n19575 & ~n19931;
  assign n19933 = ~n19575 & n19931;
  assign n19934 = ~n19932 & ~n19933;
  assign n19935 = n19918 & ~n19934;
  assign n19936 = ~n19897 & ~n19935;
  assign n19937 = ~n19855 & n19936;
  assign n19938 = ~n19630 & n19655;
  assign n19939 = ~n19646 & ~n19938;
  assign n19940 = n19646 & n19938;
  assign n19941 = ~n19939 & ~n19940;
  assign n19942 = ~n19603 & n19941;
  assign n19943 = ~n19918 & n19934;
  assign n19944 = ~n19942 & n19943;
  assign n19945 = ~n19878 & ~n19896;
  assign n19946 = ~n19944 & ~n19945;
  assign n19947 = n19768 & ~n19832;
  assign n19948 = ~n19752 & n19848;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = n19768 & n19848;
  assign n19951 = ~n19752 & ~n19832;
  assign n19952 = ~n19950 & ~n19951;
  assign n19953 = n19949 & n19952;
  assign n19954 = ~pi3509 & ~n12975;
  assign n19955 = pi3509 & ~n12971;
  assign n19956 = ~n19954 & ~n19955;
  assign n19957 = n19607 & ~n19956;
  assign n19958 = ~n12940 & n19612;
  assign n19959 = ~n12944 & n19615;
  assign n19960 = ~n19958 & ~n19959;
  assign n19961 = ~n12989 & n19619;
  assign n19962 = ~pi3509 & ~n12962;
  assign n19963 = pi3509 & ~n12958;
  assign n19964 = ~n19962 & ~n19963;
  assign n19965 = n19624 & ~n19964;
  assign n19966 = ~n19961 & ~n19965;
  assign n19967 = n19960 & n19966;
  assign n19968 = ~n19611 & n19967;
  assign n19969 = ~n19607 & ~n19968;
  assign n19970 = ~n19957 & ~n19969;
  assign n19971 = n19655 & ~n19970;
  assign n19972 = n19646 & ~n19971;
  assign n19973 = ~n19646 & n19971;
  assign n19974 = ~n19972 & ~n19973;
  assign n19975 = pi2195 & n19585;
  assign n19976 = ~pi0325 & pi0979;
  assign n19977 = ~pi0326 & ~pi0979;
  assign n19978 = ~n19976 & ~n19977;
  assign n19979 = n19588 & ~n19978;
  assign n19980 = ~pi3516 & ~n12984;
  assign n19981 = pi3516 & ~n12980;
  assign n19982 = ~n19980 & ~n19981;
  assign n19983 = ~pi3518 & ~n19982;
  assign n19984 = ~n19979 & ~n19983;
  assign n19985 = ~n19585 & n19984;
  assign n19986 = ~n19975 & ~n19985;
  assign n19987 = n19581 & n19986;
  assign n19988 = n19575 & ~n19987;
  assign n19989 = ~n19575 & n19987;
  assign n19990 = ~n19988 & ~n19989;
  assign n19991 = ~n19974 & ~n19990;
  assign n19992 = ~n13173 & n19619;
  assign n19993 = ~n13182 & n19610;
  assign n19994 = ~n19992 & ~n19993;
  assign n19995 = ~n13204 & n19612;
  assign n19996 = ~n13208 & n19615;
  assign n19997 = ~n19995 & ~n19996;
  assign n19998 = n19994 & n19997;
  assign n19999 = ~pi3509 & ~n13297;
  assign n20000 = pi3509 & ~n13293;
  assign n20001 = ~n19999 & ~n20000;
  assign n20002 = n19624 & ~n20001;
  assign n20003 = n19998 & ~n20002;
  assign n20004 = ~n19607 & ~n20003;
  assign n20005 = ~pi3509 & ~n13159;
  assign n20006 = pi3509 & ~n13155;
  assign n20007 = ~n20005 & ~n20006;
  assign n20008 = n19607 & ~n20007;
  assign n20009 = ~n20004 & ~n20008;
  assign n20010 = n19655 & ~n20009;
  assign n20011 = ~n19646 & ~n20010;
  assign n20012 = n19646 & n20010;
  assign n20013 = ~n20011 & ~n20012;
  assign n20014 = pi2196 & n19585;
  assign n20015 = ~pi0337 & pi0979;
  assign n20016 = ~pi0339 & ~pi0979;
  assign n20017 = ~n20015 & ~n20016;
  assign n20018 = n19588 & ~n20017;
  assign n20019 = ~pi3516 & ~n13168;
  assign n20020 = pi3516 & ~n13164;
  assign n20021 = ~n20019 & ~n20020;
  assign n20022 = ~pi3518 & ~n20021;
  assign n20023 = ~n20018 & ~n20022;
  assign n20024 = ~n19585 & n20023;
  assign n20025 = ~n20014 & ~n20024;
  assign n20026 = n19581 & n20025;
  assign n20027 = n19575 & ~n20026;
  assign n20028 = ~n19575 & n20026;
  assign n20029 = ~n20027 & ~n20028;
  assign n20030 = n20013 & ~n20029;
  assign n20031 = ~n19991 & ~n20030;
  assign n20032 = ~pi2199 & n19585;
  assign n20033 = ~pi3516 & ~n14644;
  assign n20034 = pi3516 & ~n14640;
  assign n20035 = ~n20033 & ~n20034;
  assign n20036 = ~pi3518 & ~n20035;
  assign n20037 = ~pi0347 & pi0979;
  assign n20038 = ~pi0349 & ~pi0979;
  assign n20039 = ~n20037 & ~n20038;
  assign n20040 = n19588 & ~n20039;
  assign n20041 = ~n20036 & ~n20040;
  assign n20042 = ~n19585 & ~n20041;
  assign n20043 = ~n20032 & ~n20042;
  assign n20044 = ~n19575 & n20043;
  assign n20045 = n19892 & ~n20043;
  assign n20046 = ~n20044 & ~n20045;
  assign n20047 = ~n19895 & n20046;
  assign n20048 = pi3509 & ~n14605;
  assign n20049 = ~pi3509 & ~n14609;
  assign n20050 = ~n20048 & ~n20049;
  assign n20051 = n19624 & ~n20050;
  assign n20052 = ~n14649 & n19619;
  assign n20053 = ~n14685 & n19610;
  assign n20054 = ~n14676 & n19612;
  assign n20055 = ~n14680 & n19615;
  assign n20056 = ~n20054 & ~n20055;
  assign n20057 = ~n20053 & n20056;
  assign n20058 = ~n20052 & n20057;
  assign n20059 = ~n20051 & n20058;
  assign n20060 = ~n19607 & ~n20059;
  assign n20061 = ~pi3509 & ~n14635;
  assign n20062 = pi3509 & ~n14631;
  assign n20063 = ~n20061 & ~n20062;
  assign n20064 = n19607 & ~n20063;
  assign n20065 = ~n20060 & ~n20064;
  assign n20066 = n19655 & ~n20065;
  assign n20067 = n19646 & n20066;
  assign n20068 = ~n19646 & n20065;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = ~n19877 & n20069;
  assign n20071 = ~n20047 & ~n20070;
  assign n20072 = ~pi2197 & n19585;
  assign n20073 = ~pi3516 & ~n13816;
  assign n20074 = pi3516 & ~n13812;
  assign n20075 = ~n20073 & ~n20074;
  assign n20076 = ~pi3518 & ~n20075;
  assign n20077 = ~pi0338 & pi0979;
  assign n20078 = ~pi0340 & ~pi0979;
  assign n20079 = ~n20077 & ~n20078;
  assign n20080 = n19588 & ~n20079;
  assign n20081 = ~n20076 & ~n20080;
  assign n20082 = ~n19585 & ~n20081;
  assign n20083 = ~n20072 & ~n20082;
  assign n20084 = ~n19575 & n20083;
  assign n20085 = n19892 & ~n20083;
  assign n20086 = ~n20084 & ~n20085;
  assign n20087 = ~n19895 & n20086;
  assign n20088 = ~n13839 & n19612;
  assign n20089 = ~n13843 & n19615;
  assign n20090 = ~n20088 & ~n20089;
  assign n20091 = ~n13821 & n19619;
  assign n20092 = ~n13848 & n19610;
  assign n20093 = ~n20091 & ~n20092;
  assign n20094 = n20090 & n20093;
  assign n20095 = ~pi3509 & ~n13794;
  assign n20096 = pi3509 & ~n13790;
  assign n20097 = ~n20095 & ~n20096;
  assign n20098 = n19624 & ~n20097;
  assign n20099 = n20094 & ~n20098;
  assign n20100 = ~n19607 & ~n20099;
  assign n20101 = ~pi3509 & ~n13807;
  assign n20102 = pi3509 & ~n13803;
  assign n20103 = ~n20101 & ~n20102;
  assign n20104 = n19607 & ~n20103;
  assign n20105 = ~n20100 & ~n20104;
  assign n20106 = n19655 & ~n20105;
  assign n20107 = n19646 & n20106;
  assign n20108 = ~n19646 & n20105;
  assign n20109 = ~n20107 & ~n20108;
  assign n20110 = ~n19877 & n20109;
  assign n20111 = n20087 & n20110;
  assign n20112 = ~pi3509 & ~n14868;
  assign n20113 = pi3509 & ~n14864;
  assign n20114 = ~n20112 & ~n20113;
  assign n20115 = n19607 & ~n20114;
  assign n20116 = ~n14913 & n19612;
  assign n20117 = ~n14917 & n19615;
  assign n20118 = ~n20116 & ~n20117;
  assign n20119 = pi3509 & ~n14993;
  assign n20120 = ~pi3509 & ~n14997;
  assign n20121 = ~n20119 & ~n20120;
  assign n20122 = n19624 & ~n20121;
  assign n20123 = ~n14882 & n19619;
  assign n20124 = ~n14891 & n19610;
  assign n20125 = ~n20123 & ~n20124;
  assign n20126 = ~n20122 & n20125;
  assign n20127 = n20118 & n20126;
  assign n20128 = ~n19607 & ~n20127;
  assign n20129 = ~n20115 & ~n20128;
  assign n20130 = n19655 & ~n20129;
  assign n20131 = ~n19646 & ~n20130;
  assign n20132 = n19646 & n20130;
  assign n20133 = ~n20131 & ~n20132;
  assign n20134 = pi2198 & n19585;
  assign n20135 = ~pi0401 & pi0979;
  assign n20136 = ~pi0402 & ~pi0979;
  assign n20137 = ~n20135 & ~n20136;
  assign n20138 = n19588 & ~n20137;
  assign n20139 = ~pi3516 & ~n14877;
  assign n20140 = pi3516 & ~n14873;
  assign n20141 = ~n20139 & ~n20140;
  assign n20142 = ~pi3518 & ~n20141;
  assign n20143 = ~n20138 & ~n20142;
  assign n20144 = ~n19585 & n20143;
  assign n20145 = ~n20134 & ~n20144;
  assign n20146 = n19581 & n20145;
  assign n20147 = n19575 & ~n20146;
  assign n20148 = ~n19575 & n20146;
  assign n20149 = ~n20147 & ~n20148;
  assign n20150 = ~n20133 & n20149;
  assign n20151 = ~n20111 & n20150;
  assign n20152 = ~n20071 & ~n20151;
  assign n20153 = n20133 & ~n20149;
  assign n20154 = n20047 & n20070;
  assign n20155 = ~n20153 & ~n20154;
  assign n20156 = ~pi3509 & ~n11810;
  assign n20157 = pi3509 & ~n11814;
  assign n20158 = ~n20156 & ~n20157;
  assign n20159 = n19607 & ~n20158;
  assign n20160 = ~n11929 & n19612;
  assign n20161 = ~n11933 & n19615;
  assign n20162 = ~n20160 & ~n20161;
  assign n20163 = pi3509 & ~n11855;
  assign n20164 = ~pi3509 & ~n11837;
  assign n20165 = ~n20163 & ~n20164;
  assign n20166 = n19624 & ~n20165;
  assign n20167 = ~n11819 & n19619;
  assign n20168 = ~n11947 & n19610;
  assign n20169 = ~n20167 & ~n20168;
  assign n20170 = ~n20166 & n20169;
  assign n20171 = n20162 & n20170;
  assign n20172 = ~n19607 & ~n20171;
  assign n20173 = ~n20159 & ~n20172;
  assign n20174 = n19655 & ~n20173;
  assign n20175 = ~n19646 & n20174;
  assign n20176 = n19646 & ~n20174;
  assign n20177 = ~n20175 & ~n20176;
  assign n20178 = pi2083 & n19585;
  assign n20179 = ~pi0436 & pi0979;
  assign n20180 = ~pi0437 & ~pi0979;
  assign n20181 = ~n20179 & ~n20180;
  assign n20182 = n19588 & ~n20181;
  assign n20183 = ~pi3516 & ~n11829;
  assign n20184 = pi3516 & ~n11825;
  assign n20185 = ~n20183 & ~n20184;
  assign n20186 = ~pi3518 & ~n20185;
  assign n20187 = ~n20182 & ~n20186;
  assign n20188 = ~n19585 & n20187;
  assign n20189 = ~n20178 & ~n20188;
  assign n20190 = n19581 & n20189;
  assign n20191 = n19575 & ~n20190;
  assign n20192 = ~n19575 & n20190;
  assign n20193 = ~n20191 & ~n20192;
  assign n20194 = n20177 & n20193;
  assign n20195 = ~pi3509 & ~n10997;
  assign n20196 = pi3509 & ~n10993;
  assign n20197 = ~n20195 & ~n20196;
  assign n20198 = n19607 & ~n20197;
  assign n20199 = ~n10966 & n19612;
  assign n20200 = ~n10970 & n19615;
  assign n20201 = ~n20199 & ~n20200;
  assign n20202 = pi3509 & ~n11020;
  assign n20203 = ~pi3509 & ~n11038;
  assign n20204 = ~n20202 & ~n20203;
  assign n20205 = n19624 & ~n20204;
  assign n20206 = ~n11011 & n19619;
  assign n20207 = ~n20205 & ~n20206;
  assign n20208 = n20201 & n20207;
  assign n20209 = ~n10975 & n19610;
  assign n20210 = n20208 & ~n20209;
  assign n20211 = ~n19607 & ~n20210;
  assign n20212 = ~n20198 & ~n20211;
  assign n20213 = n19655 & ~n20212;
  assign n20214 = ~n19646 & n20213;
  assign n20215 = n19646 & ~n20213;
  assign n20216 = ~n20214 & ~n20215;
  assign n20217 = ~pi2200 & n19585;
  assign n20218 = pi3516 & ~n11002;
  assign n20219 = ~pi3516 & ~n11006;
  assign n20220 = ~n20218 & ~n20219;
  assign n20221 = ~pi3518 & ~n20220;
  assign n20222 = ~pi0463 & pi0979;
  assign n20223 = ~pi0464 & ~pi0979;
  assign n20224 = ~n20222 & ~n20223;
  assign n20225 = n19588 & ~n20224;
  assign n20226 = ~n20221 & ~n20225;
  assign n20227 = ~n19585 & ~n20226;
  assign n20228 = ~n20217 & ~n20227;
  assign n20229 = n19581 & ~n20228;
  assign n20230 = n19575 & ~n20229;
  assign n20231 = ~n19575 & n20229;
  assign n20232 = ~n20230 & ~n20231;
  assign n20233 = n20216 & n20232;
  assign n20234 = ~n20177 & ~n20193;
  assign n20235 = pi0196 & n19631;
  assign n20236 = pi0196 & n19565;
  assign n20237 = ~n19563 & ~n20236;
  assign n20238 = n19580 & n20237;
  assign n20239 = pi1972 & pi1973;
  assign n20240 = ~pi1974 & n20239;
  assign n20241 = pi0196 & n20240;
  assign n20242 = pi1975 & n20241;
  assign n20243 = ~n19651 & ~n20242;
  assign n20244 = ~n19638 & n20243;
  assign n20245 = n20238 & n20244;
  assign n20246 = ~n19568 & n20245;
  assign n20247 = ~n20235 & n20246;
  assign n20248 = ~n19635 & n20247;
  assign n20249 = ~n19630 & ~n20248;
  assign n20250 = ~n19568 & ~n19635;
  assign n20251 = pi2142 & pi3065;
  assign n20252 = pi2758 & n20251;
  assign n20253 = ~n20235 & ~n20252;
  assign n20254 = n20237 & n20244;
  assign n20255 = n20253 & n20254;
  assign n20256 = n20250 & n20255;
  assign n20257 = n19630 & ~n20256;
  assign n20258 = ~n20249 & ~n20257;
  assign n20259 = ~n20234 & ~n20258;
  assign n20260 = ~n20233 & ~n20259;
  assign n20261 = ~n20216 & ~n20232;
  assign n20262 = ~n20260 & ~n20261;
  assign n20263 = ~n20194 & ~n20262;
  assign n20264 = n20155 & ~n20263;
  assign n20265 = n20152 & ~n20264;
  assign n20266 = ~pi3509 & ~n12234;
  assign n20267 = pi3509 & ~n12230;
  assign n20268 = ~n20266 & ~n20267;
  assign n20269 = n19607 & ~n20268;
  assign n20270 = pi3509 & ~n12217;
  assign n20271 = ~pi3509 & ~n12221;
  assign n20272 = ~n20270 & ~n20271;
  assign n20273 = n19624 & ~n20272;
  assign n20274 = ~n12248 & n19619;
  assign n20275 = ~n12257 & n19610;
  assign n20276 = ~n12270 & n19612;
  assign n20277 = ~n12274 & n19615;
  assign n20278 = ~n20276 & ~n20277;
  assign n20279 = ~n20275 & n20278;
  assign n20280 = ~n20274 & n20279;
  assign n20281 = ~n20273 & n20280;
  assign n20282 = ~n19607 & ~n20281;
  assign n20283 = ~n20269 & ~n20282;
  assign n20284 = n19655 & ~n20283;
  assign n20285 = ~n19646 & ~n20284;
  assign n20286 = n19646 & n20284;
  assign n20287 = ~n20285 & ~n20286;
  assign n20288 = ~n20087 & ~n20287;
  assign n20289 = pi2079 & n19585;
  assign n20290 = ~pi0346 & pi0979;
  assign n20291 = ~pi0348 & ~pi0979;
  assign n20292 = ~n20290 & ~n20291;
  assign n20293 = n19588 & ~n20292;
  assign n20294 = ~pi3516 & ~n12243;
  assign n20295 = pi3516 & ~n12239;
  assign n20296 = ~n20294 & ~n20295;
  assign n20297 = ~pi3518 & ~n20296;
  assign n20298 = ~n20293 & ~n20297;
  assign n20299 = ~n19585 & n20298;
  assign n20300 = ~n20289 & ~n20299;
  assign n20301 = n19581 & n20300;
  assign n20302 = n19575 & ~n20301;
  assign n20303 = ~n19575 & n20301;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = ~n20110 & n20304;
  assign n20306 = ~n20288 & ~n20305;
  assign n20307 = ~n20087 & n20304;
  assign n20308 = ~n20110 & ~n20287;
  assign n20309 = ~n20307 & ~n20308;
  assign n20310 = n20306 & n20309;
  assign n20311 = ~n20265 & ~n20310;
  assign n20312 = ~n20087 & ~n20110;
  assign n20313 = ~n20287 & n20304;
  assign n20314 = ~n20154 & n20313;
  assign n20315 = ~n20312 & ~n20314;
  assign n20316 = ~n20311 & n20315;
  assign n20317 = n20031 & ~n20316;
  assign n20318 = ~n20013 & n20029;
  assign n20319 = ~n19991 & n20318;
  assign n20320 = ~n20317 & ~n20319;
  assign n20321 = n19974 & n19990;
  assign n20322 = n20320 & ~n20321;
  assign n20323 = ~n19953 & ~n20322;
  assign n20324 = n19853 & n20323;
  assign n20325 = n19936 & n20324;
  assign n20326 = n19946 & ~n20325;
  assign n20327 = ~n19937 & n20326;
  assign n20328 = n19676 & ~n19692;
  assign n20329 = ~n20327 & ~n20328;
  assign n20330 = ~n19693 & ~n20329;
  assign n20331 = n19603 & n20330;
  assign n20332 = ~n19603 & ~n20330;
  assign n20333 = ~n20331 & ~n20332;
  assign n20334 = ~n19567 & n19578;
  assign n20335 = n19603 & ~n19941;
  assign n20336 = ~n19942 & ~n20335;
  assign n20337 = ~n20334 & ~n20336;
  assign n20338 = ~n20333 & n20337;
  assign n20339 = pi0152 & pi0829;
  assign n20340 = ~n20338 & ~n20339;
  assign n20341 = n19554 & ~n20340;
  assign n20342 = ~pi0835 & ~n15115;
  assign n20343 = ~n20341 & ~n20342;
  assign n20344 = pi1042 & pi1093;
  assign n20345 = ~pi1041 & n20344;
  assign n20346 = ~pi1517 & n20345;
  assign n20347 = pi1041 & n19548;
  assign n20348 = ~pi1417 & n20347;
  assign n20349 = ~n20346 & ~n20348;
  assign n20350 = pi1041 & n20344;
  assign n20351 = ~pi1585 & n20350;
  assign n20352 = ~pi1042 & pi1093;
  assign n20353 = pi1041 & n20352;
  assign n20354 = ~pi1570 & n20353;
  assign n20355 = pi1041 & pi1042;
  assign n20356 = ~pi1093 & n20355;
  assign n20357 = ~pi1553 & n20356;
  assign n20358 = ~n20354 & ~n20357;
  assign n20359 = ~pi1041 & ~pi1042;
  assign n20360 = pi1093 & n20359;
  assign n20361 = ~pi1499 & n20360;
  assign n20362 = pi1042 & ~pi1093;
  assign n20363 = ~pi1041 & n20362;
  assign n20364 = ~pi1481 & n20363;
  assign n20365 = ~n20361 & ~n20364;
  assign n20366 = n20358 & n20365;
  assign n20367 = ~n20351 & n20366;
  assign n20368 = n20349 & n20367;
  assign n20369 = n19550 & ~n20368;
  assign n20370 = n20343 & ~n20369;
  assign n20371 = n19560 & ~n20370;
  assign n20372 = pi0415 & ~pi0427;
  assign n20373 = n19558 & n20372;
  assign n20374 = n20370 & n20373;
  assign n20375 = pi0407 & ~pi0414;
  assign n20376 = n19559 & n20375;
  assign n20377 = ~pi0835 & ~n12061;
  assign n20378 = ~n20330 & ~n20334;
  assign n20379 = pi1974 & n19578;
  assign n20380 = pi1975 & n20379;
  assign n20381 = n20336 & ~n20380;
  assign n20382 = n19603 & n20379;
  assign n20383 = ~n19941 & n20382;
  assign n20384 = ~n20381 & ~n20383;
  assign n20385 = n20378 & ~n20384;
  assign n20386 = ~n20378 & n20384;
  assign n20387 = ~n20385 & ~n20386;
  assign n20388 = pi0828 & n20338;
  assign n20389 = n20387 & ~n20388;
  assign n20390 = ~n20387 & n20388;
  assign n20391 = ~n20389 & ~n20390;
  assign n20392 = n19554 & ~n20391;
  assign n20393 = ~n20377 & ~n20392;
  assign n20394 = ~pi1521 & n20345;
  assign n20395 = ~pi1540 & n20347;
  assign n20396 = ~n20394 & ~n20395;
  assign n20397 = ~pi1588 & n20350;
  assign n20398 = ~pi1625 & n20353;
  assign n20399 = ~pi1557 & n20356;
  assign n20400 = ~n20398 & ~n20399;
  assign n20401 = ~pi1620 & n20360;
  assign n20402 = ~pi1485 & n20363;
  assign n20403 = ~n20401 & ~n20402;
  assign n20404 = n20400 & n20403;
  assign n20405 = ~n20397 & n20404;
  assign n20406 = n20396 & n20405;
  assign n20407 = n19550 & ~n20406;
  assign n20408 = n20393 & ~n20407;
  assign n20409 = n20370 & n20408;
  assign n20410 = ~n20370 & ~n20408;
  assign n20411 = ~n20409 & ~n20410;
  assign n20412 = n20376 & n20411;
  assign n20413 = n20372 & n20375;
  assign n20414 = ~n20411 & n20413;
  assign n20415 = ~n20412 & ~n20414;
  assign n20416 = pi0414 & ~pi0427;
  assign n20417 = pi0407 & ~pi0415;
  assign n20418 = n20416 & n20417;
  assign n20419 = ~n19942 & ~n20328;
  assign n20420 = ~n19855 & n20419;
  assign n20421 = n19936 & n20420;
  assign n20422 = ~n20326 & n20419;
  assign n20423 = n19693 & ~n19897;
  assign n20424 = ~n20422 & ~n20423;
  assign n20425 = ~n20421 & n20424;
  assign n20426 = ~n20335 & n20425;
  assign n20427 = ~n20334 & ~n20426;
  assign n20428 = n19554 & n20427;
  assign n20429 = ~pi1516 & n20345;
  assign n20430 = ~pi1535 & n20347;
  assign n20431 = ~n20429 & ~n20430;
  assign n20432 = ~pi1584 & n20350;
  assign n20433 = ~pi1569 & n20353;
  assign n20434 = ~pi1409 & n20356;
  assign n20435 = ~n20433 & ~n20434;
  assign n20436 = ~pi1498 & n20360;
  assign n20437 = ~pi1406 & n20363;
  assign n20438 = ~n20436 & ~n20437;
  assign n20439 = n20435 & n20438;
  assign n20440 = ~n20432 & n20439;
  assign n20441 = n20431 & n20440;
  assign n20442 = n19550 & ~n20441;
  assign n20443 = ~n20428 & ~n20442;
  assign n20444 = ~pi0835 & ~n14816;
  assign n20445 = n20443 & ~n20444;
  assign n20446 = n20418 & n20445;
  assign n20447 = pi0414 & pi0427;
  assign n20448 = n20417 & n20447;
  assign n20449 = ~n20445 & n20448;
  assign n20450 = ~n20446 & ~n20449;
  assign n20451 = n20415 & n20450;
  assign n20452 = ~n20374 & n20451;
  assign n20453 = ~n20371 & n20452;
  assign n20454 = ~n19557 & ~n20453;
  assign n20455 = n19554 & n19579;
  assign n20456 = ~pi1971 & n20455;
  assign n20457 = ~n9352 & n20456;
  assign n20458 = ~n19551 & ~n20457;
  assign n20459 = ~n19543 & n20458;
  assign n20460 = ~pi0407 & ~pi0415;
  assign n20461 = n20447 & n20460;
  assign n20462 = ~pi1515 & n20345;
  assign n20463 = ~pi1534 & n20347;
  assign n20464 = ~n20462 & ~n20463;
  assign n20465 = ~pi1583 & n20350;
  assign n20466 = ~pi1394 & n20353;
  assign n20467 = ~pi1552 & n20356;
  assign n20468 = ~n20466 & ~n20467;
  assign n20469 = ~pi1626 & n20360;
  assign n20470 = ~pi1480 & n20363;
  assign n20471 = ~n20469 & ~n20470;
  assign n20472 = n20468 & n20471;
  assign n20473 = ~n20465 & n20472;
  assign n20474 = n20464 & n20473;
  assign n20475 = n19550 & ~n20474;
  assign n20476 = ~n19630 & n20456;
  assign n20477 = ~n20475 & ~n20476;
  assign n20478 = ~pi0835 & ~n12415;
  assign n20479 = n20477 & ~n20478;
  assign n20480 = n20461 & ~n20479;
  assign n20481 = n20416 & n20460;
  assign n20482 = n20479 & n20481;
  assign n20483 = ~n20480 & ~n20482;
  assign n20484 = ~n20459 & ~n20483;
  assign n20485 = ~n20454 & ~n20484;
  assign n20486 = pi0152 & n19560;
  assign n20487 = ~pi0152 & n20373;
  assign n20488 = ~n20486 & ~n20487;
  assign n20489 = n8640 & n20376;
  assign n20490 = ~n8640 & n20413;
  assign n20491 = ~n20489 & ~n20490;
  assign n20492 = n20488 & n20491;
  assign n20493 = ~pi0196 & n20418;
  assign n20494 = pi0196 & n20448;
  assign n20495 = ~n20493 & ~n20494;
  assign n20496 = n20492 & n20495;
  assign n20497 = n19557 & ~n20496;
  assign n20498 = ~pi0407 & ~pi0427;
  assign n20499 = pi0415 & n20498;
  assign n20500 = pi0414 & n20499;
  assign n20501 = pi0659 & n20461;
  assign n20502 = ~pi0659 & n20481;
  assign n20503 = ~n20501 & ~n20502;
  assign n20504 = n20459 & ~n20503;
  assign n20505 = ~n20500 & ~n20504;
  assign n20506 = ~n20497 & n20505;
  assign n20507 = n20485 & n20506;
  assign n20508 = ~n8561 & ~n20507;
  assign n20509 = ~n19542 & ~n20508;
  assign po0493 = ~pi3377 & pi3642;
  assign po0308 = ~n20509 & po0493;
  assign n20512 = pi0979 & ~pi1666;
  assign n20513 = ~pi0714 & ~pi3426;
  assign n20514 = ~pi2757 & ~pi3633;
  assign n20515 = ~pi3426 & n20514;
  assign n20516 = ~n20513 & ~n20515;
  assign n20517 = pi0979 & ~n20516;
  assign n20518 = ~n20512 & ~n20517;
  assign n20519 = ~pi0713 & ~pi3426;
  assign n20520 = pi0979 & n20519;
  assign n20521 = n20518 & ~n20520;
  assign n20522 = ~n9352 & n19553;
  assign n20523 = n20512 & n20522;
  assign n20524 = ~n20521 & n20523;
  assign n20525 = pi0039 & ~n20524;
  assign n20526 = n20521 & n20525;
  assign n20527 = pi0066 & pi0104;
  assign n20528 = ~pi1473 & n20527;
  assign n20529 = pi0081 & pi1640;
  assign n20530 = n20528 & n20529;
  assign n20531 = pi0104 & pi1473;
  assign n20532 = pi0066 & n20531;
  assign n20533 = ~n20529 & n20532;
  assign n20534 = ~n20530 & ~n20533;
  assign n20535 = ~pi0066 & ~pi0104;
  assign n20536 = pi1473 & n20535;
  assign n20537 = pi0066 & ~pi0104;
  assign n20538 = ~pi1473 & n20537;
  assign n20539 = ~n20536 & ~n20538;
  assign n20540 = n20529 & n20539;
  assign n20541 = pi1473 & n20537;
  assign n20542 = ~pi1473 & n20535;
  assign n20543 = ~n20541 & ~n20542;
  assign n20544 = ~n20529 & n20543;
  assign n20545 = ~n20540 & ~n20544;
  assign n20546 = n20534 & ~n20545;
  assign n20547 = pi0055 & ~pi0097;
  assign n20548 = ~pi0066 & n20547;
  assign n20549 = ~pi1424 & n20548;
  assign n20550 = ~pi0055 & pi0097;
  assign n20551 = pi0066 & n20550;
  assign n20552 = pi1424 & n20551;
  assign n20553 = ~n20549 & ~n20552;
  assign n20554 = n20529 & n20553;
  assign n20555 = pi1424 & ~n20548;
  assign n20556 = ~pi1424 & ~n20551;
  assign n20557 = ~n20555 & ~n20556;
  assign n20558 = ~n20529 & ~n20557;
  assign n20559 = ~n20554 & ~n20558;
  assign n20560 = pi0055 & pi0066;
  assign n20561 = ~pi0055 & ~pi0066;
  assign n20562 = ~n20560 & ~n20561;
  assign n20563 = pi0097 & ~n20562;
  assign n20564 = pi1424 & n20563;
  assign n20565 = ~pi0097 & ~n20562;
  assign n20566 = ~pi1424 & n20565;
  assign n20567 = ~n20564 & ~n20566;
  assign n20568 = n20529 & n20567;
  assign n20569 = pi1424 & n20565;
  assign n20570 = ~pi1424 & n20563;
  assign n20571 = ~n20569 & ~n20570;
  assign n20572 = ~n20529 & n20571;
  assign n20573 = ~n20568 & ~n20572;
  assign n20574 = ~n20559 & ~n20573;
  assign n20575 = ~pi0075 & pi0076;
  assign n20576 = pi0097 & n20575;
  assign n20577 = ~pi1468 & n20576;
  assign n20578 = pi0075 & ~pi0076;
  assign n20579 = ~pi0097 & n20578;
  assign n20580 = pi1468 & n20579;
  assign n20581 = ~n20577 & ~n20580;
  assign n20582 = n20529 & n20581;
  assign n20583 = pi1468 & ~n20576;
  assign n20584 = ~pi1468 & ~n20579;
  assign n20585 = ~n20583 & ~n20584;
  assign n20586 = ~n20529 & ~n20585;
  assign n20587 = ~n20582 & ~n20586;
  assign n20588 = pi0076 & ~pi0097;
  assign n20589 = ~pi0076 & pi0097;
  assign n20590 = ~n20588 & ~n20589;
  assign n20591 = pi0075 & ~n20590;
  assign n20592 = pi1468 & n20591;
  assign n20593 = ~pi0075 & ~n20590;
  assign n20594 = ~pi1468 & n20593;
  assign n20595 = ~n20592 & ~n20594;
  assign n20596 = n20529 & ~n20595;
  assign n20597 = pi1468 & n20593;
  assign n20598 = ~pi1468 & n20591;
  assign n20599 = ~n20597 & ~n20598;
  assign n20600 = ~n20529 & ~n20599;
  assign n20601 = ~n20596 & ~n20600;
  assign n20602 = ~n20587 & n20601;
  assign n20603 = ~n20574 & n20602;
  assign n20604 = n20574 & ~n20602;
  assign n20605 = ~n20603 & ~n20604;
  assign n20606 = pi0074 & ~pi0075;
  assign n20607 = ~pi0074 & pi0075;
  assign n20608 = ~n20606 & ~n20607;
  assign n20609 = pi0096 & ~n20608;
  assign n20610 = pi1469 & n20609;
  assign n20611 = ~pi0096 & ~n20608;
  assign n20612 = ~pi1469 & n20611;
  assign n20613 = ~n20610 & ~n20612;
  assign n20614 = n20529 & n20613;
  assign n20615 = pi1469 & n20611;
  assign n20616 = ~pi1469 & n20609;
  assign n20617 = ~n20615 & ~n20616;
  assign n20618 = ~n20529 & n20617;
  assign n20619 = ~n20614 & ~n20618;
  assign n20620 = ~pi0074 & ~pi0075;
  assign n20621 = pi0096 & n20620;
  assign n20622 = pi1469 & n20621;
  assign n20623 = pi0074 & pi0075;
  assign n20624 = ~pi0096 & n20623;
  assign n20625 = ~pi1469 & n20624;
  assign n20626 = ~n20622 & ~n20625;
  assign n20627 = n20529 & n20626;
  assign n20628 = pi1469 & ~n20624;
  assign n20629 = ~pi1469 & ~n20621;
  assign n20630 = ~n20628 & ~n20629;
  assign n20631 = ~n20529 & ~n20630;
  assign n20632 = ~n20627 & ~n20631;
  assign n20633 = ~n20619 & ~n20632;
  assign n20634 = n20605 & ~n20633;
  assign n20635 = ~n20605 & n20633;
  assign n20636 = ~n20634 & ~n20635;
  assign n20637 = ~n20574 & ~n20602;
  assign n20638 = n20574 & n20602;
  assign n20639 = ~n20633 & ~n20638;
  assign n20640 = ~n20637 & ~n20639;
  assign n20641 = n20636 & n20640;
  assign n20642 = ~n20636 & ~n20640;
  assign n20643 = ~n20641 & ~n20642;
  assign n20644 = n20546 & ~n20643;
  assign n20645 = ~n20546 & n20643;
  assign n20646 = ~n20644 & ~n20645;
  assign n20647 = ~n20546 & ~n20636;
  assign n20648 = ~n20546 & ~n20640;
  assign n20649 = ~n20647 & ~n20648;
  assign n20650 = n20646 & ~n20649;
  assign n20651 = ~n20646 & n20649;
  assign n20652 = ~n20650 & ~n20651;
  assign n20653 = ~n20642 & ~n20646;
  assign n20654 = n20646 & n20649;
  assign n20655 = ~n20653 & ~n20654;
  assign n20656 = ~n20652 & ~n20655;
  assign n20657 = ~pi0077 & pi0099;
  assign n20658 = pi0100 & n20657;
  assign n20659 = pi1471 & ~n20658;
  assign n20660 = pi0077 & ~pi0099;
  assign n20661 = ~pi0100 & n20660;
  assign n20662 = ~pi1471 & ~n20661;
  assign n20663 = ~n20659 & ~n20662;
  assign n20664 = ~pi0109 & n20663;
  assign n20665 = pi0099 & ~pi0100;
  assign n20666 = ~pi0099 & pi0100;
  assign n20667 = ~n20665 & ~n20666;
  assign n20668 = pi0077 & ~n20667;
  assign n20669 = pi1471 & n20668;
  assign n20670 = ~pi0077 & ~n20667;
  assign n20671 = ~pi1471 & n20670;
  assign n20672 = ~n20669 & ~n20671;
  assign n20673 = pi0081 & ~n20672;
  assign n20674 = ~n20664 & ~n20673;
  assign n20675 = pi1471 & n20670;
  assign n20676 = ~pi1471 & n20668;
  assign n20677 = ~n20675 & ~n20676;
  assign n20678 = ~pi0081 & ~n20677;
  assign n20679 = ~pi1471 & n20658;
  assign n20680 = pi1471 & n20661;
  assign n20681 = ~n20679 & ~n20680;
  assign n20682 = pi0109 & ~n20681;
  assign n20683 = ~n20678 & ~n20682;
  assign n20684 = n20674 & n20683;
  assign n20685 = ~pi0077 & ~pi1647;
  assign n20686 = ~pi1424 & n20685;
  assign n20687 = ~pi0110 & ~n20686;
  assign n20688 = pi1473 & n20685;
  assign n20689 = pi0110 & ~n20688;
  assign n20690 = ~n20687 & ~n20689;
  assign n20691 = pi2384 & ~n17071;
  assign n20692 = ~pi0868 & n20691;
  assign n20693 = pi2384 & ~n9511;
  assign n20694 = pi0868 & n20693;
  assign n20695 = ~n20692 & ~n20694;
  assign n20696 = pi1472 & ~n20695;
  assign n20697 = ~n20690 & ~n20696;
  assign n20698 = ~n20684 & ~n20697;
  assign n20699 = n20690 & n20696;
  assign n20700 = ~n20698 & ~n20699;
  assign n20701 = ~pi0109 & ~n20686;
  assign n20702 = pi0109 & ~n20688;
  assign n20703 = ~n20701 & ~n20702;
  assign n20704 = ~pi0081 & n20663;
  assign n20705 = pi0081 & ~n20681;
  assign n20706 = ~n20704 & ~n20705;
  assign n20707 = n20529 & ~n20672;
  assign n20708 = ~n20529 & ~n20677;
  assign n20709 = ~n20707 & ~n20708;
  assign n20710 = n20706 & n20709;
  assign n20711 = n20703 & n20710;
  assign n20712 = ~n20703 & ~n20710;
  assign n20713 = ~n20711 & ~n20712;
  assign n20714 = pi2384 & ~n17327;
  assign n20715 = ~pi0868 & n20714;
  assign n20716 = pi0868 & n20691;
  assign n20717 = ~n20715 & ~n20716;
  assign n20718 = pi1472 & ~n20717;
  assign n20719 = ~n20713 & ~n20718;
  assign n20720 = n20713 & n20718;
  assign n20721 = ~n20719 & ~n20720;
  assign n20722 = n20700 & n20721;
  assign n20723 = pi0095 & ~pi0096;
  assign n20724 = ~pi0095 & pi0096;
  assign n20725 = ~n20723 & ~n20724;
  assign n20726 = pi0098 & ~n20725;
  assign n20727 = pi1425 & n20726;
  assign n20728 = ~pi0098 & ~n20725;
  assign n20729 = ~pi1425 & n20728;
  assign n20730 = ~n20727 & ~n20729;
  assign n20731 = n20529 & n20730;
  assign n20732 = pi1425 & n20728;
  assign n20733 = ~pi1425 & n20726;
  assign n20734 = ~n20732 & ~n20733;
  assign n20735 = ~n20529 & n20734;
  assign n20736 = ~n20731 & ~n20735;
  assign n20737 = pi0095 & pi0096;
  assign n20738 = ~pi0098 & n20737;
  assign n20739 = ~pi1425 & n20738;
  assign n20740 = ~pi0095 & ~pi0096;
  assign n20741 = pi0098 & n20740;
  assign n20742 = pi1425 & n20741;
  assign n20743 = ~n20739 & ~n20742;
  assign n20744 = n20529 & n20743;
  assign n20745 = pi1425 & ~n20738;
  assign n20746 = ~pi1425 & ~n20741;
  assign n20747 = ~n20745 & ~n20746;
  assign n20748 = ~n20529 & ~n20747;
  assign n20749 = ~n20744 & ~n20748;
  assign n20750 = ~n20736 & ~n20749;
  assign n20751 = ~pi0098 & pi0103;
  assign n20752 = pi0098 & ~pi0103;
  assign n20753 = ~n20751 & ~n20752;
  assign n20754 = pi0102 & ~n20753;
  assign n20755 = pi1470 & n20754;
  assign n20756 = ~pi0102 & ~n20753;
  assign n20757 = ~pi1470 & n20756;
  assign n20758 = ~n20755 & ~n20757;
  assign n20759 = n20529 & n20758;
  assign n20760 = pi1470 & n20756;
  assign n20761 = ~pi1470 & n20754;
  assign n20762 = ~n20760 & ~n20761;
  assign n20763 = ~n20529 & n20762;
  assign n20764 = ~n20759 & ~n20763;
  assign n20765 = pi0098 & pi0103;
  assign n20766 = ~pi0102 & n20765;
  assign n20767 = ~pi1470 & n20766;
  assign n20768 = ~pi0098 & ~pi0103;
  assign n20769 = pi0102 & n20768;
  assign n20770 = pi1470 & n20769;
  assign n20771 = ~n20767 & ~n20770;
  assign n20772 = n20529 & n20771;
  assign n20773 = pi1470 & ~n20766;
  assign n20774 = ~pi1470 & ~n20769;
  assign n20775 = ~n20773 & ~n20774;
  assign n20776 = ~n20529 & ~n20775;
  assign n20777 = ~n20772 & ~n20776;
  assign n20778 = ~n20764 & ~n20777;
  assign n20779 = n20750 & ~n20778;
  assign n20780 = ~n20750 & n20778;
  assign n20781 = ~n20779 & ~n20780;
  assign n20782 = pi0101 & ~pi0102;
  assign n20783 = ~pi0101 & pi0102;
  assign n20784 = ~n20782 & ~n20783;
  assign n20785 = pi0100 & ~n20784;
  assign n20786 = pi1418 & n20785;
  assign n20787 = ~pi0100 & ~n20784;
  assign n20788 = ~pi1418 & n20787;
  assign n20789 = ~n20786 & ~n20788;
  assign n20790 = n20529 & n20789;
  assign n20791 = pi1418 & n20787;
  assign n20792 = ~pi1418 & n20785;
  assign n20793 = ~n20791 & ~n20792;
  assign n20794 = ~n20529 & n20793;
  assign n20795 = ~n20790 & ~n20794;
  assign n20796 = pi0100 & ~pi0101;
  assign n20797 = ~pi0102 & n20796;
  assign n20798 = pi1418 & n20797;
  assign n20799 = ~pi0100 & pi0101;
  assign n20800 = pi0102 & n20799;
  assign n20801 = ~pi1418 & n20800;
  assign n20802 = ~n20798 & ~n20801;
  assign n20803 = n20529 & n20802;
  assign n20804 = pi1418 & ~n20800;
  assign n20805 = ~pi1418 & ~n20797;
  assign n20806 = ~n20804 & ~n20805;
  assign n20807 = ~n20529 & ~n20806;
  assign n20808 = ~n20803 & ~n20807;
  assign n20809 = ~n20795 & ~n20808;
  assign n20810 = n20781 & ~n20809;
  assign n20811 = ~n20781 & n20809;
  assign n20812 = ~n20810 & ~n20811;
  assign n20813 = ~n20750 & ~n20778;
  assign n20814 = n20750 & n20778;
  assign n20815 = ~n20809 & ~n20814;
  assign n20816 = ~n20813 & ~n20815;
  assign n20817 = n20812 & n20816;
  assign n20818 = ~n20722 & ~n20817;
  assign n20819 = ~n20812 & ~n20816;
  assign n20820 = ~n20817 & ~n20819;
  assign n20821 = ~n20703 & ~n20718;
  assign n20822 = ~n20710 & ~n20821;
  assign n20823 = n20703 & n20718;
  assign n20824 = ~n20822 & ~n20823;
  assign n20825 = ~pi0081 & ~n20686;
  assign n20826 = pi0081 & ~n20688;
  assign n20827 = ~n20825 & ~n20826;
  assign n20828 = n20529 & ~n20681;
  assign n20829 = ~n20529 & n20663;
  assign n20830 = ~n20828 & ~n20829;
  assign n20831 = n20709 & n20830;
  assign n20832 = n20827 & n20831;
  assign n20833 = ~n20827 & ~n20831;
  assign n20834 = ~n20832 & ~n20833;
  assign n20835 = pi2384 & ~n10975;
  assign n20836 = ~pi0868 & n20835;
  assign n20837 = pi0868 & n20714;
  assign n20838 = ~n20836 & ~n20837;
  assign n20839 = pi1472 & ~n20838;
  assign n20840 = ~n20834 & ~n20839;
  assign n20841 = n20834 & n20839;
  assign n20842 = ~n20840 & ~n20841;
  assign n20843 = n20824 & n20842;
  assign n20844 = ~n20824 & ~n20842;
  assign n20845 = ~n20843 & ~n20844;
  assign n20846 = n20820 & ~n20845;
  assign n20847 = ~n20820 & n20845;
  assign n20848 = ~n20846 & ~n20847;
  assign n20849 = n20818 & n20848;
  assign n20850 = ~n20818 & ~n20848;
  assign n20851 = ~n20849 & ~n20850;
  assign n20852 = pi0111 & n20688;
  assign n20853 = ~pi0111 & n20686;
  assign n20854 = ~n20852 & ~n20853;
  assign n20855 = ~pi0868 & n20693;
  assign n20856 = pi2384 & ~n10420;
  assign n20857 = pi0868 & n20856;
  assign n20858 = ~n20855 & ~n20857;
  assign n20859 = pi1472 & ~n20858;
  assign n20860 = ~n20854 & n20859;
  assign n20861 = ~pi0109 & ~n20677;
  assign n20862 = pi0109 & ~n20672;
  assign n20863 = pi0110 & ~n20681;
  assign n20864 = ~n20862 & ~n20863;
  assign n20865 = ~pi0110 & n20663;
  assign n20866 = n20864 & ~n20865;
  assign n20867 = ~n20861 & n20866;
  assign n20868 = n20854 & ~n20859;
  assign n20869 = ~n20867 & ~n20868;
  assign n20870 = ~n20860 & ~n20869;
  assign n20871 = ~pi0081 & ~n20806;
  assign n20872 = pi0081 & n20802;
  assign n20873 = ~n20871 & ~n20872;
  assign n20874 = ~n20795 & ~n20873;
  assign n20875 = ~n20814 & ~n20874;
  assign n20876 = ~n20813 & ~n20875;
  assign n20877 = ~n20870 & ~n20876;
  assign n20878 = n20684 & n20690;
  assign n20879 = ~n20684 & ~n20690;
  assign n20880 = ~n20878 & ~n20879;
  assign n20881 = ~n20696 & ~n20880;
  assign n20882 = n20696 & n20880;
  assign n20883 = ~n20881 & ~n20882;
  assign n20884 = ~n20812 & ~n20883;
  assign n20885 = ~n20877 & ~n20884;
  assign n20886 = ~n20812 & ~n20870;
  assign n20887 = ~n20876 & ~n20883;
  assign n20888 = ~n20886 & ~n20887;
  assign n20889 = n20885 & n20888;
  assign n20890 = ~n20700 & ~n20721;
  assign n20891 = ~n20722 & ~n20890;
  assign n20892 = n20820 & ~n20891;
  assign n20893 = ~n20820 & n20891;
  assign n20894 = ~n20892 & ~n20893;
  assign n20895 = n20889 & ~n20894;
  assign n20896 = ~n20819 & n20894;
  assign n20897 = ~n20890 & n20896;
  assign n20898 = ~n20895 & ~n20897;
  assign n20899 = n20851 & ~n20898;
  assign n20900 = ~n20656 & ~n20899;
  assign n20901 = n20652 & ~n20655;
  assign n20902 = ~n20652 & n20655;
  assign n20903 = ~n20901 & ~n20902;
  assign n20904 = ~n20844 & n20848;
  assign n20905 = ~n20819 & n20904;
  assign n20906 = ~n20850 & ~n20905;
  assign n20907 = pi2384 & ~n11947;
  assign n20908 = ~pi0868 & n20907;
  assign n20909 = pi0868 & n20835;
  assign n20910 = ~n20908 & ~n20909;
  assign n20911 = pi1472 & ~n20910;
  assign n20912 = n20529 & ~n20688;
  assign n20913 = ~n20529 & ~n20686;
  assign n20914 = ~n20912 & ~n20913;
  assign n20915 = ~n20831 & n20914;
  assign n20916 = n20831 & ~n20914;
  assign n20917 = ~n20915 & ~n20916;
  assign n20918 = n20911 & n20917;
  assign n20919 = ~n20911 & ~n20917;
  assign n20920 = ~n20918 & ~n20919;
  assign n20921 = ~n20827 & ~n20839;
  assign n20922 = ~n20831 & ~n20921;
  assign n20923 = n20827 & n20839;
  assign n20924 = ~n20922 & ~n20923;
  assign n20925 = ~n20920 & ~n20924;
  assign n20926 = n20920 & n20924;
  assign n20927 = ~n20925 & ~n20926;
  assign n20928 = n20820 & ~n20927;
  assign n20929 = ~n20820 & n20927;
  assign n20930 = ~n20928 & ~n20929;
  assign n20931 = ~n20817 & ~n20843;
  assign n20932 = n20930 & ~n20931;
  assign n20933 = ~n20930 & n20931;
  assign n20934 = ~n20932 & ~n20933;
  assign n20935 = n20906 & n20934;
  assign n20936 = ~n20906 & ~n20934;
  assign n20937 = ~n20935 & ~n20936;
  assign n20938 = n20903 & ~n20937;
  assign n20939 = ~n20903 & n20937;
  assign n20940 = ~n20938 & ~n20939;
  assign n20941 = ~n20900 & ~n20940;
  assign n20942 = n20652 & n20655;
  assign n20943 = n20940 & ~n20942;
  assign n20944 = n20906 & ~n20934;
  assign n20945 = n20943 & ~n20944;
  assign n20946 = ~n20941 & ~n20945;
  assign n20947 = ~n20906 & n20934;
  assign n20948 = n20655 & ~n20947;
  assign n20949 = n20652 & ~n20934;
  assign n20950 = ~n20948 & ~n20949;
  assign n20951 = n20652 & n20906;
  assign n20952 = n20950 & ~n20951;
  assign n20953 = n20920 & ~n20924;
  assign n20954 = ~n20930 & ~n20953;
  assign n20955 = ~n20819 & n20954;
  assign n20956 = ~n20932 & ~n20955;
  assign n20957 = ~n20920 & n20924;
  assign n20958 = ~n20817 & ~n20957;
  assign n20959 = pi2384 & ~n14891;
  assign n20960 = ~pi0868 & n20959;
  assign n20961 = pi0868 & n20907;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = pi1472 & ~n20962;
  assign n20964 = n20917 & n20963;
  assign n20965 = ~n20917 & ~n20963;
  assign n20966 = ~n20964 & ~n20965;
  assign n20967 = n20911 & ~n20916;
  assign n20968 = ~n20915 & ~n20967;
  assign n20969 = ~n20966 & ~n20968;
  assign n20970 = n20966 & n20968;
  assign n20971 = ~n20969 & ~n20970;
  assign n20972 = n20820 & ~n20971;
  assign n20973 = ~n20820 & n20971;
  assign n20974 = ~n20972 & ~n20973;
  assign n20975 = n20958 & n20974;
  assign n20976 = ~n20958 & ~n20974;
  assign n20977 = ~n20975 & ~n20976;
  assign n20978 = ~n20956 & n20977;
  assign n20979 = n20956 & ~n20977;
  assign n20980 = ~n20978 & ~n20979;
  assign n20981 = n20903 & ~n20980;
  assign n20982 = ~n20903 & n20980;
  assign n20983 = ~n20981 & ~n20982;
  assign n20984 = ~n20952 & n20983;
  assign n20985 = n20952 & ~n20983;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = n20946 & ~n20986;
  assign n20988 = ~n20889 & n20894;
  assign n20989 = ~n20895 & ~n20988;
  assign n20990 = ~pi0110 & ~n20677;
  assign n20991 = pi0110 & ~n20672;
  assign n20992 = pi0111 & ~n20681;
  assign n20993 = ~n20991 & ~n20992;
  assign n20994 = ~pi0111 & n20663;
  assign n20995 = n20993 & ~n20994;
  assign n20996 = ~n20990 & n20995;
  assign n20997 = ~pi0112 & ~n20686;
  assign n20998 = pi0112 & ~n20688;
  assign n20999 = ~n20997 & ~n20998;
  assign n21000 = ~pi0868 & n20856;
  assign n21001 = pi2384 & ~n15259;
  assign n21002 = pi0868 & n21001;
  assign n21003 = ~n21000 & ~n21002;
  assign n21004 = pi1472 & ~n21003;
  assign n21005 = ~n20999 & ~n21004;
  assign n21006 = ~n20996 & ~n21005;
  assign n21007 = n20999 & n21004;
  assign n21008 = ~n21006 & ~n21007;
  assign n21009 = ~pi0109 & ~n20806;
  assign n21010 = pi0109 & n20802;
  assign n21011 = ~n21009 & ~n21010;
  assign n21012 = ~pi0081 & n20793;
  assign n21013 = pi0081 & n20789;
  assign n21014 = ~n21012 & ~n21013;
  assign n21015 = ~n21011 & ~n21014;
  assign n21016 = ~n20814 & ~n21015;
  assign n21017 = ~n20813 & ~n21016;
  assign n21018 = ~n21008 & ~n21017;
  assign n21019 = ~n20860 & ~n20868;
  assign n21020 = ~n20867 & ~n21019;
  assign n21021 = n20854 & n20859;
  assign n21022 = ~n20854 & ~n20859;
  assign n21023 = ~n21021 & ~n21022;
  assign n21024 = n20867 & ~n21023;
  assign n21025 = ~n21020 & ~n21024;
  assign n21026 = n20781 & ~n20874;
  assign n21027 = ~n20781 & n20874;
  assign n21028 = ~n21026 & ~n21027;
  assign n21029 = ~n21025 & ~n21028;
  assign n21030 = ~n21018 & ~n21029;
  assign n21031 = ~n21008 & ~n21028;
  assign n21032 = ~n21017 & ~n21025;
  assign n21033 = ~n21031 & ~n21032;
  assign n21034 = n21030 & n21033;
  assign n21035 = ~n20870 & n20883;
  assign n21036 = n20870 & ~n20883;
  assign n21037 = ~n21035 & ~n21036;
  assign n21038 = n20812 & n20876;
  assign n21039 = ~n20812 & ~n20876;
  assign n21040 = ~n21038 & ~n21039;
  assign n21041 = ~n21037 & n21040;
  assign n21042 = n21037 & ~n21040;
  assign n21043 = ~n21041 & ~n21042;
  assign n21044 = n21034 & n21043;
  assign n21045 = ~n20870 & ~n20883;
  assign n21046 = ~n21039 & ~n21045;
  assign n21047 = ~n21043 & n21046;
  assign n21048 = ~n21044 & ~n21047;
  assign n21049 = n20989 & ~n21048;
  assign n21050 = ~n20656 & ~n21049;
  assign n21051 = ~n20851 & ~n20898;
  assign n21052 = n20851 & n20898;
  assign n21053 = ~n21051 & ~n21052;
  assign n21054 = n20903 & ~n21053;
  assign n21055 = ~n20903 & n21053;
  assign n21056 = ~n21054 & ~n21055;
  assign n21057 = n21050 & n21056;
  assign n21058 = ~n21050 & ~n21056;
  assign n21059 = ~n21057 & ~n21058;
  assign n21060 = ~n20989 & ~n21048;
  assign n21061 = n20989 & n21048;
  assign n21062 = ~n21060 & ~n21061;
  assign n21063 = n20903 & ~n21062;
  assign n21064 = ~n20903 & n21062;
  assign n21065 = ~n21063 & ~n21064;
  assign n21066 = ~n20942 & n21065;
  assign n21067 = ~n20989 & n21048;
  assign n21068 = n21066 & ~n21067;
  assign n21069 = ~n21034 & ~n21043;
  assign n21070 = ~n21044 & ~n21069;
  assign n21071 = n20655 & ~n21070;
  assign n21072 = n20996 & ~n20999;
  assign n21073 = ~n20996 & n20999;
  assign n21074 = ~n21072 & ~n21073;
  assign n21075 = ~n21004 & ~n21074;
  assign n21076 = n21004 & n21074;
  assign n21077 = ~n21075 & ~n21076;
  assign n21078 = ~pi0081 & n20775;
  assign n21079 = pi0081 & ~n20771;
  assign n21080 = ~n21078 & ~n21079;
  assign n21081 = ~n20764 & n21080;
  assign n21082 = ~pi0110 & ~n20806;
  assign n21083 = pi0110 & n20802;
  assign n21084 = ~n21082 & ~n21083;
  assign n21085 = ~pi0109 & n20793;
  assign n21086 = pi0109 & n20789;
  assign n21087 = ~n21085 & ~n21086;
  assign n21088 = ~n21084 & ~n21087;
  assign n21089 = ~n21081 & ~n21088;
  assign n21090 = n21081 & n21088;
  assign n21091 = ~n20750 & ~n21090;
  assign n21092 = ~n21089 & ~n21091;
  assign n21093 = n20781 & ~n21015;
  assign n21094 = ~n20781 & n21015;
  assign n21095 = ~n21093 & ~n21094;
  assign n21096 = n21092 & n21095;
  assign n21097 = n21077 & ~n21096;
  assign n21098 = pi0113 & n20688;
  assign n21099 = ~pi0113 & n20686;
  assign n21100 = ~n21098 & ~n21099;
  assign n21101 = ~pi0868 & n21001;
  assign n21102 = pi2384 & ~n14219;
  assign n21103 = pi0868 & n21102;
  assign n21104 = ~n21101 & ~n21103;
  assign n21105 = pi1472 & ~n21104;
  assign n21106 = ~n21100 & n21105;
  assign n21107 = ~pi0111 & ~n20677;
  assign n21108 = pi0111 & ~n20672;
  assign n21109 = pi0112 & ~n20681;
  assign n21110 = ~n21108 & ~n21109;
  assign n21111 = ~pi0112 & n20663;
  assign n21112 = n21110 & ~n21111;
  assign n21113 = ~n21107 & n21112;
  assign n21114 = n21100 & ~n21105;
  assign n21115 = ~n21113 & ~n21114;
  assign n21116 = ~n21106 & ~n21115;
  assign n21117 = ~n21095 & ~n21116;
  assign n21118 = ~n21097 & ~n21117;
  assign n21119 = ~n21092 & ~n21116;
  assign n21120 = n21118 & ~n21119;
  assign n21121 = n21008 & ~n21025;
  assign n21122 = ~n21008 & n21025;
  assign n21123 = ~n21121 & ~n21122;
  assign n21124 = n21017 & n21028;
  assign n21125 = ~n21017 & ~n21028;
  assign n21126 = ~n21124 & ~n21125;
  assign n21127 = ~n21123 & n21126;
  assign n21128 = n21123 & ~n21126;
  assign n21129 = ~n21127 & ~n21128;
  assign n21130 = n21120 & n21129;
  assign n21131 = ~n21008 & ~n21025;
  assign n21132 = ~n21125 & ~n21131;
  assign n21133 = ~n21129 & n21132;
  assign n21134 = ~n21130 & ~n21133;
  assign n21135 = n21070 & ~n21134;
  assign n21136 = n20652 & ~n21135;
  assign n21137 = ~n21071 & ~n21136;
  assign n21138 = n20655 & n21134;
  assign n21139 = n21137 & ~n21138;
  assign n21140 = ~n21065 & n21139;
  assign n21141 = ~n21068 & ~n21140;
  assign n21142 = ~n21059 & n21141;
  assign n21143 = n21070 & n21134;
  assign n21144 = ~n21070 & ~n21134;
  assign n21145 = ~n21143 & ~n21144;
  assign n21146 = n20903 & ~n21145;
  assign n21147 = ~n20903 & n21145;
  assign n21148 = ~n21146 & ~n21147;
  assign n21149 = ~n20942 & n21148;
  assign n21150 = ~n21070 & n21134;
  assign n21151 = n21149 & ~n21150;
  assign n21152 = ~pi0081 & ~n20762;
  assign n21153 = pi0109 & ~n20771;
  assign n21154 = ~n21152 & ~n21153;
  assign n21155 = ~pi0109 & n20775;
  assign n21156 = pi0081 & ~n20758;
  assign n21157 = ~n21155 & ~n21156;
  assign n21158 = n21154 & n21157;
  assign n21159 = ~pi0111 & ~n20806;
  assign n21160 = pi0111 & n20802;
  assign n21161 = ~n21159 & ~n21160;
  assign n21162 = ~pi0110 & n20793;
  assign n21163 = pi0110 & n20789;
  assign n21164 = ~n21162 & ~n21163;
  assign n21165 = ~n21161 & ~n21164;
  assign n21166 = ~n21158 & ~n21165;
  assign n21167 = n21158 & n21165;
  assign n21168 = ~n20750 & ~n21167;
  assign n21169 = ~n21166 & ~n21168;
  assign n21170 = ~n21089 & ~n21090;
  assign n21171 = ~n20750 & ~n21170;
  assign n21172 = n21081 & ~n21088;
  assign n21173 = ~n21081 & n21088;
  assign n21174 = ~n21172 & ~n21173;
  assign n21175 = n20750 & ~n21174;
  assign n21176 = ~n21171 & ~n21175;
  assign n21177 = n21169 & n21176;
  assign n21178 = ~n21106 & ~n21114;
  assign n21179 = ~n21113 & ~n21178;
  assign n21180 = n21100 & n21105;
  assign n21181 = ~n21100 & ~n21105;
  assign n21182 = ~n21180 & ~n21181;
  assign n21183 = n21113 & ~n21182;
  assign n21184 = ~n21179 & ~n21183;
  assign n21185 = ~n21177 & ~n21184;
  assign n21186 = ~pi0113 & n20663;
  assign n21187 = pi0113 & ~n20681;
  assign n21188 = ~n21186 & ~n21187;
  assign n21189 = ~pi0112 & ~n20677;
  assign n21190 = pi0112 & ~n20672;
  assign n21191 = ~n21189 & ~n21190;
  assign n21192 = n21188 & n21191;
  assign n21193 = ~pi0105 & ~n20686;
  assign n21194 = pi0105 & ~n20688;
  assign n21195 = ~n21193 & ~n21194;
  assign n21196 = ~pi0868 & n21102;
  assign n21197 = pi2384 & ~n12609;
  assign n21198 = pi0868 & n21197;
  assign n21199 = ~n21196 & ~n21198;
  assign n21200 = pi1472 & ~n21199;
  assign n21201 = ~n21195 & ~n21200;
  assign n21202 = ~n21192 & ~n21201;
  assign n21203 = n21195 & n21200;
  assign n21204 = ~n21202 & ~n21203;
  assign n21205 = ~n21169 & ~n21204;
  assign n21206 = ~n21185 & ~n21205;
  assign n21207 = ~n21176 & ~n21204;
  assign n21208 = n21206 & ~n21207;
  assign n21209 = n21077 & ~n21116;
  assign n21210 = ~n21077 & n21116;
  assign n21211 = ~n21209 & ~n21210;
  assign n21212 = n21092 & ~n21095;
  assign n21213 = ~n21092 & n21095;
  assign n21214 = ~n21212 & ~n21213;
  assign n21215 = ~n21211 & ~n21214;
  assign n21216 = n21211 & n21214;
  assign n21217 = ~n21215 & ~n21216;
  assign n21218 = n21208 & ~n21217;
  assign n21219 = ~n21092 & ~n21095;
  assign n21220 = ~n21209 & ~n21219;
  assign n21221 = n21217 & n21220;
  assign n21222 = ~n21218 & ~n21221;
  assign n21223 = ~n21120 & ~n21129;
  assign n21224 = ~n21130 & ~n21223;
  assign n21225 = ~n21222 & n21224;
  assign n21226 = ~n20656 & ~n21225;
  assign n21227 = ~n21148 & ~n21226;
  assign n21228 = ~n21151 & ~n21227;
  assign n21229 = n21148 & n21226;
  assign n21230 = ~n21227 & ~n21229;
  assign n21231 = n21228 & ~n21230;
  assign n21232 = ~n21208 & n21217;
  assign n21233 = ~n21218 & ~n21232;
  assign n21234 = n20652 & ~n21233;
  assign n21235 = ~pi0112 & ~n20806;
  assign n21236 = pi0112 & n20802;
  assign n21237 = ~n21235 & ~n21236;
  assign n21238 = ~pi0111 & n20793;
  assign n21239 = pi0111 & n20789;
  assign n21240 = ~n21238 & ~n21239;
  assign n21241 = ~n21237 & ~n21240;
  assign n21242 = ~pi0081 & n20747;
  assign n21243 = pi0081 & ~n20743;
  assign n21244 = ~n21242 & ~n21243;
  assign n21245 = ~n20736 & n21244;
  assign n21246 = ~n21241 & ~n21245;
  assign n21247 = ~pi0109 & ~n20762;
  assign n21248 = pi0109 & ~n20758;
  assign n21249 = pi0110 & ~n20771;
  assign n21250 = ~n21248 & ~n21249;
  assign n21251 = ~pi0110 & n20775;
  assign n21252 = n21250 & ~n21251;
  assign n21253 = ~n21247 & n21252;
  assign n21254 = n21241 & n21245;
  assign n21255 = ~n21253 & ~n21254;
  assign n21256 = ~n21246 & ~n21255;
  assign n21257 = pi0113 & ~n20672;
  assign n21258 = pi0105 & ~n20681;
  assign n21259 = ~n21257 & ~n21258;
  assign n21260 = ~pi0113 & ~n20677;
  assign n21261 = ~pi0105 & n20663;
  assign n21262 = ~n21260 & ~n21261;
  assign n21263 = n21259 & n21262;
  assign n21264 = ~pi0107 & ~n20686;
  assign n21265 = pi0107 & ~n20688;
  assign n21266 = ~n21264 & ~n21265;
  assign n21267 = ~pi0868 & n21197;
  assign n21268 = pi2384 & ~n13534;
  assign n21269 = pi0868 & n21268;
  assign n21270 = ~n21267 & ~n21269;
  assign n21271 = pi1472 & ~n21270;
  assign n21272 = ~n21266 & ~n21271;
  assign n21273 = ~n21263 & ~n21272;
  assign n21274 = n21266 & n21271;
  assign n21275 = ~n21273 & ~n21274;
  assign n21276 = ~n21256 & ~n21275;
  assign n21277 = ~n21166 & ~n21167;
  assign n21278 = ~n20750 & ~n21277;
  assign n21279 = n21158 & ~n21165;
  assign n21280 = ~n21158 & n21165;
  assign n21281 = ~n21279 & ~n21280;
  assign n21282 = n20750 & ~n21281;
  assign n21283 = ~n21278 & ~n21282;
  assign n21284 = n21192 & ~n21195;
  assign n21285 = ~n21192 & n21195;
  assign n21286 = ~n21284 & ~n21285;
  assign n21287 = ~n21200 & ~n21286;
  assign n21288 = n21200 & n21286;
  assign n21289 = ~n21287 & ~n21288;
  assign n21290 = n21275 & ~n21289;
  assign n21291 = ~n21283 & ~n21290;
  assign n21292 = ~n21276 & ~n21291;
  assign n21293 = ~n21256 & n21289;
  assign n21294 = n21292 & ~n21293;
  assign n21295 = ~n21169 & ~n21176;
  assign n21296 = ~n21177 & ~n21295;
  assign n21297 = ~n21184 & n21204;
  assign n21298 = n21184 & ~n21204;
  assign n21299 = ~n21297 & ~n21298;
  assign n21300 = ~n21296 & n21299;
  assign n21301 = n21296 & ~n21299;
  assign n21302 = ~n21300 & ~n21301;
  assign n21303 = n21294 & n21302;
  assign n21304 = ~n21184 & ~n21204;
  assign n21305 = ~n21295 & ~n21304;
  assign n21306 = ~n21302 & n21305;
  assign n21307 = ~n21303 & ~n21306;
  assign n21308 = n21233 & ~n21307;
  assign n21309 = n20655 & ~n21308;
  assign n21310 = ~n21234 & ~n21309;
  assign n21311 = n20652 & n21307;
  assign n21312 = n21310 & ~n21311;
  assign n21313 = n21222 & n21224;
  assign n21314 = ~n21222 & ~n21224;
  assign n21315 = ~n21313 & ~n21314;
  assign n21316 = n20903 & n21315;
  assign n21317 = ~n20903 & ~n21315;
  assign n21318 = ~n21316 & ~n21317;
  assign n21319 = n21312 & n21318;
  assign n21320 = ~n20942 & ~n21318;
  assign n21321 = n21222 & ~n21224;
  assign n21322 = n21320 & ~n21321;
  assign n21323 = ~n21319 & ~n21322;
  assign n21324 = n21065 & n21139;
  assign n21325 = ~n21065 & ~n21139;
  assign n21326 = ~n21324 & ~n21325;
  assign n21327 = n21323 & n21326;
  assign n21328 = ~n21231 & ~n21327;
  assign n21329 = n21228 & n21323;
  assign n21330 = ~n21230 & n21326;
  assign n21331 = ~n21329 & ~n21330;
  assign n21332 = n21328 & n21331;
  assign n21333 = ~pi0113 & ~n20806;
  assign n21334 = pi0113 & n20802;
  assign n21335 = ~n21333 & ~n21334;
  assign n21336 = ~pi0112 & n20793;
  assign n21337 = pi0112 & n20789;
  assign n21338 = ~n21336 & ~n21337;
  assign n21339 = ~n21335 & ~n21338;
  assign n21340 = ~pi0081 & ~n20734;
  assign n21341 = pi0081 & ~n20730;
  assign n21342 = pi0109 & ~n20743;
  assign n21343 = ~n21341 & ~n21342;
  assign n21344 = ~pi0109 & n20747;
  assign n21345 = n21343 & ~n21344;
  assign n21346 = ~n21340 & n21345;
  assign n21347 = ~n21339 & ~n21346;
  assign n21348 = ~pi0110 & ~n20762;
  assign n21349 = pi0110 & ~n20758;
  assign n21350 = pi0111 & ~n20771;
  assign n21351 = ~n21349 & ~n21350;
  assign n21352 = ~pi0111 & n20775;
  assign n21353 = n21351 & ~n21352;
  assign n21354 = ~n21348 & n21353;
  assign n21355 = n21339 & n21346;
  assign n21356 = ~n21354 & ~n21355;
  assign n21357 = ~n21347 & ~n21356;
  assign n21358 = ~n21246 & ~n21254;
  assign n21359 = ~n21253 & ~n21358;
  assign n21360 = n21241 & ~n21245;
  assign n21361 = ~n21241 & n21245;
  assign n21362 = ~n21360 & ~n21361;
  assign n21363 = n21253 & ~n21362;
  assign n21364 = ~n21359 & ~n21363;
  assign n21365 = n21357 & n21364;
  assign n21366 = ~n21357 & ~n21364;
  assign n21367 = ~n21365 & ~n21366;
  assign n21368 = pi0108 & n20688;
  assign n21369 = ~pi0108 & n20686;
  assign n21370 = ~n21368 & ~n21369;
  assign n21371 = ~pi0868 & n21268;
  assign n21372 = pi2384 & ~n12940;
  assign n21373 = pi0868 & n21372;
  assign n21374 = ~n21371 & ~n21373;
  assign n21375 = pi1472 & ~n21374;
  assign n21376 = ~n21370 & n21375;
  assign n21377 = ~pi0107 & n20663;
  assign n21378 = pi0107 & ~n20681;
  assign n21379 = ~n21377 & ~n21378;
  assign n21380 = ~pi0105 & ~n20677;
  assign n21381 = pi0105 & ~n20672;
  assign n21382 = ~n21380 & ~n21381;
  assign n21383 = n21379 & n21382;
  assign n21384 = n21370 & ~n21375;
  assign n21385 = ~n21383 & ~n21384;
  assign n21386 = ~n21376 & ~n21385;
  assign n21387 = n21263 & n21266;
  assign n21388 = ~n21263 & ~n21266;
  assign n21389 = ~n21387 & ~n21388;
  assign n21390 = ~n21271 & ~n21389;
  assign n21391 = n21271 & n21389;
  assign n21392 = ~n21390 & ~n21391;
  assign n21393 = ~n21386 & n21392;
  assign n21394 = n21386 & ~n21392;
  assign n21395 = ~n21393 & ~n21394;
  assign n21396 = ~n21367 & n21395;
  assign n21397 = n21367 & ~n21395;
  assign n21398 = ~n21396 & ~n21397;
  assign n21399 = ~pi0107 & ~n20677;
  assign n21400 = pi0107 & ~n20672;
  assign n21401 = pi0108 & ~n20681;
  assign n21402 = ~n21400 & ~n21401;
  assign n21403 = ~pi0108 & n20663;
  assign n21404 = n21402 & ~n21403;
  assign n21405 = ~n21399 & n21404;
  assign n21406 = ~pi0868 & n21372;
  assign n21407 = pi2384 & ~n13204;
  assign n21408 = pi0868 & n21407;
  assign n21409 = ~n21406 & ~n21408;
  assign n21410 = pi1472 & ~n21409;
  assign n21411 = ~pi0078 & ~n20686;
  assign n21412 = pi0078 & ~n20688;
  assign n21413 = ~n21411 & ~n21412;
  assign n21414 = ~n21410 & ~n21413;
  assign n21415 = ~n21405 & ~n21414;
  assign n21416 = n21410 & n21413;
  assign n21417 = ~n21415 & ~n21416;
  assign n21418 = ~pi0105 & ~n20806;
  assign n21419 = pi0105 & n20802;
  assign n21420 = ~n21418 & ~n21419;
  assign n21421 = ~pi0113 & n20793;
  assign n21422 = pi0113 & n20789;
  assign n21423 = ~n21421 & ~n21422;
  assign n21424 = ~n21420 & ~n21423;
  assign n21425 = ~pi0110 & n20747;
  assign n21426 = pi0109 & ~n20730;
  assign n21427 = ~n21425 & ~n21426;
  assign n21428 = ~pi0109 & ~n20734;
  assign n21429 = pi0110 & ~n20743;
  assign n21430 = ~n21428 & ~n21429;
  assign n21431 = n21427 & n21430;
  assign n21432 = ~n21424 & ~n21431;
  assign n21433 = ~pi0111 & ~n20762;
  assign n21434 = pi0111 & ~n20758;
  assign n21435 = pi0112 & ~n20771;
  assign n21436 = ~n21434 & ~n21435;
  assign n21437 = ~pi0112 & n20775;
  assign n21438 = n21436 & ~n21437;
  assign n21439 = ~n21433 & n21438;
  assign n21440 = n21424 & n21431;
  assign n21441 = ~n21439 & ~n21440;
  assign n21442 = ~n21432 & ~n21441;
  assign n21443 = ~n21417 & ~n21442;
  assign n21444 = ~n21376 & ~n21384;
  assign n21445 = ~n21383 & ~n21444;
  assign n21446 = n21370 & n21375;
  assign n21447 = ~n21370 & ~n21375;
  assign n21448 = ~n21446 & ~n21447;
  assign n21449 = n21383 & ~n21448;
  assign n21450 = ~n21445 & ~n21449;
  assign n21451 = ~n21347 & ~n21355;
  assign n21452 = ~n21354 & ~n21451;
  assign n21453 = n21339 & ~n21346;
  assign n21454 = ~n21339 & n21346;
  assign n21455 = ~n21453 & ~n21454;
  assign n21456 = n21354 & ~n21455;
  assign n21457 = ~n21452 & ~n21456;
  assign n21458 = n21442 & n21457;
  assign n21459 = ~n21450 & ~n21458;
  assign n21460 = ~n21443 & ~n21459;
  assign n21461 = ~n21417 & ~n21457;
  assign n21462 = n21460 & ~n21461;
  assign n21463 = n21398 & n21462;
  assign n21464 = ~n21386 & ~n21392;
  assign n21465 = ~n21366 & ~n21464;
  assign n21466 = ~n21398 & n21465;
  assign n21467 = ~n21463 & ~n21466;
  assign n21468 = n20652 & n21467;
  assign n21469 = ~n21357 & ~n21386;
  assign n21470 = ~n21364 & ~n21392;
  assign n21471 = ~n21469 & ~n21470;
  assign n21472 = ~n21364 & ~n21386;
  assign n21473 = ~n21357 & ~n21392;
  assign n21474 = ~n21472 & ~n21473;
  assign n21475 = n21471 & n21474;
  assign n21476 = n21256 & n21283;
  assign n21477 = ~n21256 & ~n21283;
  assign n21478 = ~n21476 & ~n21477;
  assign n21479 = ~n21275 & ~n21289;
  assign n21480 = n21275 & n21289;
  assign n21481 = ~n21479 & ~n21480;
  assign n21482 = ~n21478 & n21481;
  assign n21483 = n21478 & ~n21481;
  assign n21484 = ~n21482 & ~n21483;
  assign n21485 = n21475 & n21484;
  assign n21486 = ~n21475 & ~n21484;
  assign n21487 = ~n21485 & ~n21486;
  assign n21488 = ~n21467 & n21487;
  assign n21489 = ~pi0081 & ~n20630;
  assign n21490 = pi0081 & n20626;
  assign n21491 = ~n21489 & ~n21490;
  assign n21492 = ~n20619 & ~n21491;
  assign n21493 = ~n20638 & ~n21492;
  assign n21494 = ~n20637 & ~n21493;
  assign n21495 = ~n20546 & ~n21494;
  assign n21496 = ~n20647 & ~n21495;
  assign n21497 = n20646 & n21496;
  assign n21498 = ~n20653 & ~n21497;
  assign n21499 = ~n21488 & n21498;
  assign n21500 = n20652 & ~n21487;
  assign n21501 = ~n21499 & ~n21500;
  assign n21502 = ~n21468 & n21501;
  assign n21503 = ~n21294 & ~n21302;
  assign n21504 = ~n21303 & ~n21503;
  assign n21505 = ~n21275 & n21289;
  assign n21506 = ~n21477 & ~n21505;
  assign n21507 = ~n21484 & n21506;
  assign n21508 = ~n21485 & ~n21507;
  assign n21509 = ~n21504 & ~n21508;
  assign n21510 = n21504 & n21508;
  assign n21511 = ~n21509 & ~n21510;
  assign n21512 = n20903 & ~n21511;
  assign n21513 = ~n20903 & n21511;
  assign n21514 = ~n21512 & ~n21513;
  assign n21515 = n21502 & ~n21514;
  assign n21516 = ~n20942 & n21514;
  assign n21517 = ~n21504 & n21508;
  assign n21518 = n21516 & ~n21517;
  assign n21519 = ~n21515 & ~n21518;
  assign n21520 = n20655 & ~n21504;
  assign n21521 = n21504 & ~n21508;
  assign n21522 = n20652 & ~n21521;
  assign n21523 = ~n21520 & ~n21522;
  assign n21524 = n20655 & n21508;
  assign n21525 = n21523 & ~n21524;
  assign n21526 = ~n21233 & ~n21307;
  assign n21527 = n21233 & n21307;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = n20903 & ~n21528;
  assign n21530 = ~n20903 & n21528;
  assign n21531 = ~n21529 & ~n21530;
  assign n21532 = n21525 & n21531;
  assign n21533 = ~n21525 & ~n21531;
  assign n21534 = ~n21532 & ~n21533;
  assign n21535 = ~n21312 & ~n21318;
  assign n21536 = ~n21319 & ~n21535;
  assign n21537 = n21534 & ~n21536;
  assign n21538 = ~n20942 & n21531;
  assign n21539 = ~n21233 & n21307;
  assign n21540 = n21538 & ~n21539;
  assign n21541 = n21525 & ~n21531;
  assign n21542 = ~n21540 & ~n21541;
  assign n21543 = n21534 & n21542;
  assign n21544 = ~n21537 & ~n21543;
  assign n21545 = n21519 & ~n21544;
  assign n21546 = ~n21536 & n21542;
  assign n21547 = ~n21545 & ~n21546;
  assign n21548 = ~n21332 & ~n21547;
  assign n21549 = n21228 & n21326;
  assign n21550 = ~n21548 & ~n21549;
  assign n21551 = ~n21228 & ~n21326;
  assign n21552 = ~n21230 & n21323;
  assign n21553 = ~n21551 & n21552;
  assign n21554 = n21550 & ~n21553;
  assign n21555 = ~n21398 & ~n21462;
  assign n21556 = ~n21463 & ~n21555;
  assign n21557 = ~pi0109 & ~n20630;
  assign n21558 = pi0109 & n20626;
  assign n21559 = ~n21557 & ~n21558;
  assign n21560 = ~pi0081 & n20617;
  assign n21561 = pi0081 & n20613;
  assign n21562 = ~n21560 & ~n21561;
  assign n21563 = ~n21559 & ~n21562;
  assign n21564 = ~n20638 & ~n21563;
  assign n21565 = ~n20637 & ~n21564;
  assign n21566 = n20605 & ~n21492;
  assign n21567 = ~n20605 & n21492;
  assign n21568 = ~n21566 & ~n21567;
  assign n21569 = n21565 & n21568;
  assign n21570 = ~n20546 & ~n21569;
  assign n21571 = n20636 & ~n21494;
  assign n21572 = ~n20636 & n21494;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = n20546 & ~n21573;
  assign n21575 = ~n20546 & n21573;
  assign n21576 = ~n21574 & ~n21575;
  assign n21577 = ~n21570 & ~n21576;
  assign n21578 = ~n20636 & ~n21494;
  assign n21579 = n21576 & ~n21578;
  assign n21580 = ~n21577 & ~n21579;
  assign n21581 = ~n21556 & n21580;
  assign n21582 = n21417 & n21450;
  assign n21583 = ~n21417 & ~n21450;
  assign n21584 = ~n21582 & ~n21583;
  assign n21585 = ~n21442 & ~n21457;
  assign n21586 = ~n21458 & ~n21585;
  assign n21587 = ~n21584 & n21586;
  assign n21588 = n21584 & ~n21586;
  assign n21589 = ~n21587 & ~n21588;
  assign n21590 = ~pi0107 & ~n20806;
  assign n21591 = pi0107 & n20802;
  assign n21592 = ~n21590 & ~n21591;
  assign n21593 = ~pi0105 & n20793;
  assign n21594 = pi0105 & n20789;
  assign n21595 = ~n21593 & ~n21594;
  assign n21596 = ~n21592 & ~n21595;
  assign n21597 = ~pi0110 & ~n20734;
  assign n21598 = pi0111 & ~n20743;
  assign n21599 = ~n21597 & ~n21598;
  assign n21600 = ~pi0111 & n20747;
  assign n21601 = pi0110 & ~n20730;
  assign n21602 = ~n21600 & ~n21601;
  assign n21603 = n21599 & n21602;
  assign n21604 = ~n21596 & ~n21603;
  assign n21605 = ~pi0113 & n20775;
  assign n21606 = pi0112 & ~n20758;
  assign n21607 = ~n21605 & ~n21606;
  assign n21608 = ~pi0112 & ~n20762;
  assign n21609 = pi0113 & ~n20771;
  assign n21610 = ~n21608 & ~n21609;
  assign n21611 = n21607 & n21610;
  assign n21612 = n21596 & n21603;
  assign n21613 = ~n21611 & ~n21612;
  assign n21614 = ~n21604 & ~n21613;
  assign n21615 = n21405 & ~n21413;
  assign n21616 = ~n21405 & n21413;
  assign n21617 = ~n21615 & ~n21616;
  assign n21618 = ~n21410 & ~n21617;
  assign n21619 = n21410 & n21617;
  assign n21620 = ~n21618 & ~n21619;
  assign n21621 = ~n21614 & n21620;
  assign n21622 = ~pi0078 & n20663;
  assign n21623 = pi0108 & ~n20672;
  assign n21624 = ~n21622 & ~n21623;
  assign n21625 = ~pi0108 & ~n20677;
  assign n21626 = pi0078 & ~n20681;
  assign n21627 = ~n21625 & ~n21626;
  assign n21628 = n21624 & n21627;
  assign n21629 = pi2384 & ~n13839;
  assign n21630 = pi0868 & n21629;
  assign n21631 = ~pi0868 & n21407;
  assign n21632 = ~n21630 & ~n21631;
  assign n21633 = pi1472 & ~n21632;
  assign n21634 = ~pi0079 & ~n20686;
  assign n21635 = pi0079 & ~n20688;
  assign n21636 = ~n21634 & ~n21635;
  assign n21637 = ~n21633 & ~n21636;
  assign n21638 = ~n21628 & ~n21637;
  assign n21639 = n21633 & n21636;
  assign n21640 = ~n21638 & ~n21639;
  assign n21641 = ~n21620 & n21640;
  assign n21642 = ~n21432 & ~n21440;
  assign n21643 = ~n21439 & ~n21642;
  assign n21644 = n21424 & ~n21431;
  assign n21645 = ~n21424 & n21431;
  assign n21646 = ~n21644 & ~n21645;
  assign n21647 = n21439 & ~n21646;
  assign n21648 = ~n21643 & ~n21647;
  assign n21649 = ~n21641 & ~n21648;
  assign n21650 = ~n21621 & ~n21649;
  assign n21651 = ~n21614 & ~n21640;
  assign n21652 = n21650 & ~n21651;
  assign n21653 = ~n21589 & n21652;
  assign n21654 = ~n21583 & ~n21585;
  assign n21655 = n21589 & n21654;
  assign n21656 = ~n21653 & ~n21655;
  assign n21657 = ~n20646 & ~n21496;
  assign n21658 = ~n21497 & ~n21657;
  assign n21659 = n21656 & ~n21658;
  assign n21660 = ~n21581 & ~n21659;
  assign n21661 = n21580 & n21656;
  assign n21662 = ~n21556 & ~n21658;
  assign n21663 = ~n21661 & ~n21662;
  assign n21664 = n21660 & n21663;
  assign n21665 = n21467 & ~n21487;
  assign n21666 = ~n21488 & ~n21665;
  assign n21667 = n20652 & ~n21498;
  assign n21668 = ~n20652 & n21498;
  assign n21669 = ~n21667 & ~n21668;
  assign n21670 = ~n21666 & n21669;
  assign n21671 = n21666 & ~n21669;
  assign n21672 = ~n21670 & ~n21671;
  assign n21673 = ~n21664 & n21672;
  assign n21674 = n21664 & ~n21672;
  assign n21675 = ~n21673 & ~n21674;
  assign n21676 = n21664 & n21672;
  assign n21677 = n20652 & n21498;
  assign n21678 = ~n21665 & ~n21677;
  assign n21679 = ~n21672 & n21678;
  assign n21680 = ~n21676 & ~n21679;
  assign n21681 = n21675 & n21680;
  assign n21682 = ~n21502 & n21514;
  assign n21683 = ~n21515 & ~n21682;
  assign n21684 = n21675 & ~n21683;
  assign n21685 = ~n21565 & ~n21568;
  assign n21686 = ~n21569 & ~n21685;
  assign n21687 = n20546 & ~n21686;
  assign n21688 = ~n20546 & n21686;
  assign n21689 = ~n21687 & ~n21688;
  assign n21690 = ~n21685 & ~n21689;
  assign n21691 = ~pi0110 & ~n20630;
  assign n21692 = pi0110 & n20626;
  assign n21693 = ~n21691 & ~n21692;
  assign n21694 = ~pi0109 & n20617;
  assign n21695 = pi0109 & n20613;
  assign n21696 = ~n21694 & ~n21695;
  assign n21697 = ~n21693 & ~n21696;
  assign n21698 = ~pi0081 & n20585;
  assign n21699 = pi0081 & ~n20581;
  assign n21700 = ~n21698 & ~n21699;
  assign n21701 = n20601 & n21700;
  assign n21702 = ~n21697 & ~n21701;
  assign n21703 = n21697 & n21701;
  assign n21704 = ~n20574 & ~n21703;
  assign n21705 = ~n21702 & ~n21704;
  assign n21706 = n20605 & ~n21563;
  assign n21707 = ~n20605 & n21563;
  assign n21708 = ~n21706 & ~n21707;
  assign n21709 = n21705 & n21708;
  assign n21710 = ~n20546 & ~n21709;
  assign n21711 = n21689 & ~n21710;
  assign n21712 = ~n21690 & ~n21711;
  assign n21713 = n21589 & ~n21652;
  assign n21714 = ~n21653 & ~n21713;
  assign n21715 = n21712 & ~n21714;
  assign n21716 = n21570 & n21576;
  assign n21717 = ~n21577 & ~n21716;
  assign n21718 = ~n21614 & ~n21648;
  assign n21719 = n21614 & n21648;
  assign n21720 = ~n21718 & ~n21719;
  assign n21721 = ~n21620 & ~n21640;
  assign n21722 = n21620 & n21640;
  assign n21723 = ~n21721 & ~n21722;
  assign n21724 = ~n21720 & n21723;
  assign n21725 = n21720 & ~n21723;
  assign n21726 = ~n21724 & ~n21725;
  assign n21727 = pi0080 & n20688;
  assign n21728 = ~pi0080 & n20686;
  assign n21729 = ~n21727 & ~n21728;
  assign n21730 = pi2384 & ~n12270;
  assign n21731 = pi0868 & n21730;
  assign n21732 = ~pi0868 & n21629;
  assign n21733 = ~n21731 & ~n21732;
  assign n21734 = pi1472 & ~n21733;
  assign n21735 = ~n21729 & n21734;
  assign n21736 = ~pi0079 & n20663;
  assign n21737 = pi0079 & ~n20681;
  assign n21738 = ~n21736 & ~n21737;
  assign n21739 = ~pi0078 & ~n20677;
  assign n21740 = pi0078 & ~n20672;
  assign n21741 = ~n21739 & ~n21740;
  assign n21742 = n21738 & n21741;
  assign n21743 = n21729 & ~n21734;
  assign n21744 = ~n21742 & ~n21743;
  assign n21745 = ~n21735 & ~n21744;
  assign n21746 = ~pi0108 & ~n20806;
  assign n21747 = pi0108 & n20802;
  assign n21748 = ~n21746 & ~n21747;
  assign n21749 = ~pi0107 & n20793;
  assign n21750 = pi0107 & n20789;
  assign n21751 = ~n21749 & ~n21750;
  assign n21752 = ~n21748 & ~n21751;
  assign n21753 = ~pi0113 & ~n20762;
  assign n21754 = pi0113 & ~n20758;
  assign n21755 = pi0105 & ~n20771;
  assign n21756 = ~n21754 & ~n21755;
  assign n21757 = ~pi0105 & n20775;
  assign n21758 = n21756 & ~n21757;
  assign n21759 = ~n21753 & n21758;
  assign n21760 = ~n21752 & ~n21759;
  assign n21761 = ~pi0111 & ~n20734;
  assign n21762 = pi0111 & ~n20730;
  assign n21763 = pi0112 & ~n20743;
  assign n21764 = ~n21762 & ~n21763;
  assign n21765 = ~pi0112 & n20747;
  assign n21766 = n21764 & ~n21765;
  assign n21767 = ~n21761 & n21766;
  assign n21768 = n21752 & n21759;
  assign n21769 = ~n21767 & ~n21768;
  assign n21770 = ~n21760 & ~n21769;
  assign n21771 = ~n21745 & ~n21770;
  assign n21772 = ~n21604 & ~n21612;
  assign n21773 = ~n21611 & ~n21772;
  assign n21774 = n21596 & ~n21603;
  assign n21775 = ~n21596 & n21603;
  assign n21776 = ~n21774 & ~n21775;
  assign n21777 = n21611 & ~n21776;
  assign n21778 = ~n21773 & ~n21777;
  assign n21779 = n21628 & n21636;
  assign n21780 = ~n21628 & ~n21636;
  assign n21781 = ~n21779 & ~n21780;
  assign n21782 = ~n21633 & ~n21781;
  assign n21783 = n21633 & n21781;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = ~n21778 & ~n21784;
  assign n21786 = ~n21771 & ~n21785;
  assign n21787 = ~n21745 & ~n21778;
  assign n21788 = ~n21770 & ~n21784;
  assign n21789 = ~n21787 & ~n21788;
  assign n21790 = n21786 & n21789;
  assign n21791 = n21726 & n21790;
  assign n21792 = n21620 & ~n21640;
  assign n21793 = ~n21718 & ~n21792;
  assign n21794 = ~n21726 & n21793;
  assign n21795 = ~n21791 & ~n21794;
  assign n21796 = ~n21717 & n21795;
  assign n21797 = ~n21715 & ~n21796;
  assign n21798 = n21712 & n21795;
  assign n21799 = ~n21714 & ~n21717;
  assign n21800 = ~n21798 & ~n21799;
  assign n21801 = n21797 & n21800;
  assign n21802 = n21556 & ~n21656;
  assign n21803 = ~n21556 & n21656;
  assign n21804 = ~n21802 & ~n21803;
  assign n21805 = ~n21580 & ~n21658;
  assign n21806 = n21580 & n21658;
  assign n21807 = ~n21805 & ~n21806;
  assign n21808 = ~n21804 & n21807;
  assign n21809 = n21804 & ~n21807;
  assign n21810 = ~n21808 & ~n21809;
  assign n21811 = n21801 & n21810;
  assign n21812 = n21580 & ~n21658;
  assign n21813 = ~n21803 & ~n21812;
  assign n21814 = ~n21810 & n21813;
  assign n21815 = ~n21811 & ~n21814;
  assign n21816 = ~n21680 & n21683;
  assign n21817 = n21815 & ~n21816;
  assign n21818 = ~n21684 & ~n21817;
  assign n21819 = ~n21681 & n21818;
  assign n21820 = ~n21714 & ~n21795;
  assign n21821 = n21714 & n21795;
  assign n21822 = ~n21820 & ~n21821;
  assign n21823 = n21712 & ~n21717;
  assign n21824 = ~n21712 & n21717;
  assign n21825 = ~n21823 & ~n21824;
  assign n21826 = ~n21822 & n21825;
  assign n21827 = n21822 & ~n21825;
  assign n21828 = ~n21826 & ~n21827;
  assign n21829 = ~n21705 & ~n21708;
  assign n21830 = ~n21709 & ~n21829;
  assign n21831 = n20546 & ~n21830;
  assign n21832 = ~n20546 & n21830;
  assign n21833 = ~n21831 & ~n21832;
  assign n21834 = ~n21829 & ~n21833;
  assign n21835 = ~pi0111 & ~n20630;
  assign n21836 = pi0111 & n20626;
  assign n21837 = ~n21835 & ~n21836;
  assign n21838 = ~pi0110 & n20617;
  assign n21839 = pi0110 & n20613;
  assign n21840 = ~n21838 & ~n21839;
  assign n21841 = ~n21837 & ~n21840;
  assign n21842 = ~pi0081 & ~n20599;
  assign n21843 = pi0081 & ~n20595;
  assign n21844 = pi0109 & ~n20581;
  assign n21845 = ~n21843 & ~n21844;
  assign n21846 = ~pi0109 & n20585;
  assign n21847 = n21845 & ~n21846;
  assign n21848 = ~n21842 & n21847;
  assign n21849 = ~n21841 & ~n21848;
  assign n21850 = n21841 & n21848;
  assign n21851 = ~n20574 & ~n21850;
  assign n21852 = ~n21849 & ~n21851;
  assign n21853 = ~n21702 & ~n21703;
  assign n21854 = ~n20574 & ~n21853;
  assign n21855 = n21697 & ~n21701;
  assign n21856 = ~n21697 & n21701;
  assign n21857 = ~n21855 & ~n21856;
  assign n21858 = n20574 & ~n21857;
  assign n21859 = ~n21854 & ~n21858;
  assign n21860 = n21852 & n21859;
  assign n21861 = ~n20546 & ~n21860;
  assign n21862 = n21833 & ~n21861;
  assign n21863 = ~n21834 & ~n21862;
  assign n21864 = ~n21770 & ~n21778;
  assign n21865 = n21770 & n21778;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = ~n21745 & ~n21784;
  assign n21868 = n21745 & n21784;
  assign n21869 = ~n21867 & ~n21868;
  assign n21870 = ~n21866 & n21869;
  assign n21871 = n21866 & ~n21869;
  assign n21872 = ~n21870 & ~n21871;
  assign n21873 = ~pi0078 & ~n20806;
  assign n21874 = pi0078 & n20802;
  assign n21875 = ~n21873 & ~n21874;
  assign n21876 = ~pi0108 & n20793;
  assign n21877 = pi0108 & n20789;
  assign n21878 = ~n21876 & ~n21877;
  assign n21879 = ~n21875 & ~n21878;
  assign n21880 = ~pi0112 & ~n20734;
  assign n21881 = pi0112 & ~n20730;
  assign n21882 = pi0113 & ~n20743;
  assign n21883 = ~n21881 & ~n21882;
  assign n21884 = ~pi0113 & n20747;
  assign n21885 = n21883 & ~n21884;
  assign n21886 = ~n21880 & n21885;
  assign n21887 = ~n21879 & ~n21886;
  assign n21888 = ~pi0105 & ~n20762;
  assign n21889 = pi0105 & ~n20758;
  assign n21890 = pi0107 & ~n20771;
  assign n21891 = ~n21889 & ~n21890;
  assign n21892 = ~pi0107 & n20775;
  assign n21893 = n21891 & ~n21892;
  assign n21894 = ~n21888 & n21893;
  assign n21895 = n21879 & n21886;
  assign n21896 = ~n21894 & ~n21895;
  assign n21897 = ~n21887 & ~n21896;
  assign n21898 = ~n21735 & ~n21743;
  assign n21899 = ~n21742 & ~n21898;
  assign n21900 = n21729 & n21734;
  assign n21901 = ~n21729 & ~n21734;
  assign n21902 = ~n21900 & ~n21901;
  assign n21903 = n21742 & ~n21902;
  assign n21904 = ~n21899 & ~n21903;
  assign n21905 = ~n21897 & ~n21904;
  assign n21906 = ~pi0080 & n20663;
  assign n21907 = pi0080 & ~n20681;
  assign n21908 = ~n21906 & ~n21907;
  assign n21909 = ~pi0079 & ~n20677;
  assign n21910 = pi0079 & ~n20672;
  assign n21911 = ~n21909 & ~n21910;
  assign n21912 = n21908 & n21911;
  assign n21913 = pi2384 & ~n14676;
  assign n21914 = pi0868 & n21913;
  assign n21915 = ~pi0868 & n21730;
  assign n21916 = ~n21914 & ~n21915;
  assign n21917 = pi1472 & ~n21916;
  assign n21918 = ~pi0106 & ~n20686;
  assign n21919 = pi0106 & ~n20688;
  assign n21920 = ~n21918 & ~n21919;
  assign n21921 = ~n21917 & ~n21920;
  assign n21922 = ~n21912 & ~n21921;
  assign n21923 = n21917 & n21920;
  assign n21924 = ~n21922 & ~n21923;
  assign n21925 = n21904 & n21924;
  assign n21926 = ~n21760 & ~n21768;
  assign n21927 = ~n21767 & ~n21926;
  assign n21928 = n21752 & ~n21759;
  assign n21929 = ~n21752 & n21759;
  assign n21930 = ~n21928 & ~n21929;
  assign n21931 = n21767 & ~n21930;
  assign n21932 = ~n21927 & ~n21931;
  assign n21933 = ~n21925 & ~n21932;
  assign n21934 = ~n21905 & ~n21933;
  assign n21935 = ~n21897 & ~n21924;
  assign n21936 = n21934 & ~n21935;
  assign n21937 = ~n21872 & n21936;
  assign n21938 = ~n21864 & ~n21867;
  assign n21939 = n21872 & n21938;
  assign n21940 = ~n21937 & ~n21939;
  assign n21941 = n21863 & n21940;
  assign n21942 = ~n21726 & ~n21790;
  assign n21943 = ~n21791 & ~n21942;
  assign n21944 = ~n21689 & n21710;
  assign n21945 = ~n21711 & ~n21944;
  assign n21946 = ~n21943 & ~n21945;
  assign n21947 = ~n21941 & ~n21946;
  assign n21948 = n21863 & ~n21943;
  assign n21949 = n21940 & ~n21945;
  assign n21950 = ~n21948 & ~n21949;
  assign n21951 = n21947 & n21950;
  assign n21952 = n21828 & n21951;
  assign n21953 = ~n21714 & n21795;
  assign n21954 = ~n21823 & ~n21953;
  assign n21955 = ~n21828 & n21954;
  assign n21956 = ~n21952 & ~n21955;
  assign n21957 = ~n21801 & n21810;
  assign n21958 = n21801 & ~n21810;
  assign n21959 = ~n21957 & ~n21958;
  assign n21960 = ~n21956 & ~n21959;
  assign n21961 = n21828 & ~n21951;
  assign n21962 = ~n21828 & n21951;
  assign n21963 = ~n21961 & ~n21962;
  assign n21964 = n21940 & n21943;
  assign n21965 = ~n21940 & ~n21943;
  assign n21966 = ~n21964 & ~n21965;
  assign n21967 = n21863 & ~n21945;
  assign n21968 = ~n21863 & n21945;
  assign n21969 = ~n21967 & ~n21968;
  assign n21970 = ~n21966 & n21969;
  assign n21971 = n21966 & ~n21969;
  assign n21972 = ~n21970 & ~n21971;
  assign n21973 = ~n21852 & ~n21859;
  assign n21974 = ~n21860 & ~n21973;
  assign n21975 = n20546 & ~n21974;
  assign n21976 = ~n20546 & n21974;
  assign n21977 = ~n21975 & ~n21976;
  assign n21978 = ~n21973 & ~n21977;
  assign n21979 = ~pi0081 & n20557;
  assign n21980 = pi0081 & ~n20553;
  assign n21981 = ~n21979 & ~n21980;
  assign n21982 = ~n20573 & n21981;
  assign n21983 = ~pi0112 & ~n20630;
  assign n21984 = pi0112 & n20626;
  assign n21985 = ~n21983 & ~n21984;
  assign n21986 = ~pi0111 & n20617;
  assign n21987 = pi0111 & n20613;
  assign n21988 = ~n21986 & ~n21987;
  assign n21989 = ~n21985 & ~n21988;
  assign n21990 = ~n21982 & ~n21989;
  assign n21991 = ~pi0109 & ~n20599;
  assign n21992 = pi0109 & ~n20595;
  assign n21993 = pi0110 & ~n20581;
  assign n21994 = ~n21992 & ~n21993;
  assign n21995 = ~pi0110 & n20585;
  assign n21996 = n21994 & ~n21995;
  assign n21997 = ~n21991 & n21996;
  assign n21998 = n21982 & n21989;
  assign n21999 = ~n21997 & ~n21998;
  assign n22000 = ~n21990 & ~n21999;
  assign n22001 = ~n21849 & ~n21850;
  assign n22002 = ~n20574 & ~n22001;
  assign n22003 = n21841 & ~n21848;
  assign n22004 = ~n21841 & n21848;
  assign n22005 = ~n22003 & ~n22004;
  assign n22006 = n20574 & ~n22005;
  assign n22007 = ~n22002 & ~n22006;
  assign n22008 = n22000 & n22007;
  assign n22009 = ~n20546 & ~n22008;
  assign n22010 = n21977 & ~n22009;
  assign n22011 = ~n21978 & ~n22010;
  assign n22012 = n21872 & ~n21936;
  assign n22013 = ~n21937 & ~n22012;
  assign n22014 = n22011 & ~n22013;
  assign n22015 = ~n21904 & ~n21924;
  assign n22016 = ~n21897 & ~n21932;
  assign n22017 = ~n22015 & ~n22016;
  assign n22018 = n21897 & n21932;
  assign n22019 = ~n22016 & ~n22018;
  assign n22020 = ~n21925 & ~n22015;
  assign n22021 = ~n22019 & n22020;
  assign n22022 = n22019 & ~n22020;
  assign n22023 = ~n22021 & ~n22022;
  assign n22024 = n22017 & n22023;
  assign n22025 = n21912 & n21920;
  assign n22026 = ~n21912 & ~n21920;
  assign n22027 = ~n22025 & ~n22026;
  assign n22028 = ~n21917 & ~n22027;
  assign n22029 = n21917 & n22027;
  assign n22030 = ~n22028 & ~n22029;
  assign n22031 = ~pi0079 & ~n20806;
  assign n22032 = pi0079 & n20802;
  assign n22033 = ~n22031 & ~n22032;
  assign n22034 = ~pi0078 & n20793;
  assign n22035 = pi0078 & n20789;
  assign n22036 = ~n22034 & ~n22035;
  assign n22037 = ~n22033 & ~n22036;
  assign n22038 = ~pi0105 & n20747;
  assign n22039 = pi0105 & ~n20743;
  assign n22040 = ~n22038 & ~n22039;
  assign n22041 = ~pi0113 & ~n20734;
  assign n22042 = pi0113 & ~n20730;
  assign n22043 = ~n22041 & ~n22042;
  assign n22044 = n22040 & n22043;
  assign n22045 = ~n22037 & ~n22044;
  assign n22046 = ~pi0107 & ~n20762;
  assign n22047 = pi0107 & ~n20758;
  assign n22048 = pi0108 & ~n20771;
  assign n22049 = ~n22047 & ~n22048;
  assign n22050 = ~pi0108 & n20775;
  assign n22051 = n22049 & ~n22050;
  assign n22052 = ~n22046 & n22051;
  assign n22053 = n22037 & n22044;
  assign n22054 = ~n22052 & ~n22053;
  assign n22055 = ~n22045 & ~n22054;
  assign n22056 = ~n22030 & ~n22055;
  assign n22057 = ~n21887 & ~n21895;
  assign n22058 = ~n21894 & ~n22057;
  assign n22059 = n21879 & ~n21886;
  assign n22060 = ~n21879 & n21886;
  assign n22061 = ~n22059 & ~n22060;
  assign n22062 = n21894 & ~n22061;
  assign n22063 = ~n22058 & ~n22062;
  assign n22064 = n22055 & n22063;
  assign n22065 = pi0056 & n20688;
  assign n22066 = ~pi0056 & n20686;
  assign n22067 = ~n22065 & ~n22066;
  assign n22068 = pi2384 & ~n14913;
  assign n22069 = pi0868 & n22068;
  assign n22070 = ~pi0868 & n21913;
  assign n22071 = ~n22069 & ~n22070;
  assign n22072 = pi1472 & ~n22071;
  assign n22073 = ~n22067 & n22072;
  assign n22074 = ~pi0080 & ~n20677;
  assign n22075 = pi0080 & ~n20672;
  assign n22076 = pi0106 & ~n20681;
  assign n22077 = ~n22075 & ~n22076;
  assign n22078 = ~pi0106 & n20663;
  assign n22079 = n22077 & ~n22078;
  assign n22080 = ~n22074 & n22079;
  assign n22081 = n22067 & ~n22072;
  assign n22082 = ~n22080 & ~n22081;
  assign n22083 = ~n22073 & ~n22082;
  assign n22084 = ~n22064 & ~n22083;
  assign n22085 = ~n22056 & ~n22084;
  assign n22086 = ~n22030 & ~n22063;
  assign n22087 = n22085 & ~n22086;
  assign n22088 = ~n22023 & n22087;
  assign n22089 = ~n22024 & ~n22088;
  assign n22090 = ~n21833 & n21861;
  assign n22091 = ~n21862 & ~n22090;
  assign n22092 = n22089 & ~n22091;
  assign n22093 = ~n22014 & ~n22092;
  assign n22094 = n22011 & n22089;
  assign n22095 = ~n22013 & ~n22091;
  assign n22096 = ~n22094 & ~n22095;
  assign n22097 = n22093 & n22096;
  assign n22098 = n21972 & n22097;
  assign n22099 = n21940 & ~n21943;
  assign n22100 = ~n21967 & ~n22099;
  assign n22101 = ~n21972 & n22100;
  assign n22102 = ~n22098 & ~n22101;
  assign n22103 = n21963 & n22102;
  assign n22104 = ~n21960 & n22103;
  assign n22105 = n21956 & n21959;
  assign n22106 = ~n22104 & ~n22105;
  assign n22107 = ~n21819 & ~n22106;
  assign n22108 = ~n21963 & ~n22102;
  assign n22109 = ~n21960 & ~n22108;
  assign n22110 = ~n21819 & n22109;
  assign n22111 = n22011 & ~n22091;
  assign n22112 = ~n22013 & n22089;
  assign n22113 = ~n22111 & ~n22112;
  assign n22114 = n22013 & ~n22089;
  assign n22115 = ~n22112 & ~n22114;
  assign n22116 = n22011 & n22091;
  assign n22117 = ~n22011 & ~n22091;
  assign n22118 = ~n22116 & ~n22117;
  assign n22119 = ~n22115 & n22118;
  assign n22120 = n22115 & ~n22118;
  assign n22121 = ~n22119 & ~n22120;
  assign n22122 = n22113 & ~n22121;
  assign n22123 = ~n21977 & n22009;
  assign n22124 = ~n22010 & ~n22123;
  assign n22125 = n22023 & n22087;
  assign n22126 = ~n22023 & ~n22087;
  assign n22127 = ~n22125 & ~n22126;
  assign n22128 = ~n22124 & n22127;
  assign n22129 = ~n22000 & ~n22007;
  assign n22130 = ~n22008 & ~n22129;
  assign n22131 = n20546 & ~n22130;
  assign n22132 = ~n20546 & n22130;
  assign n22133 = ~n22131 & ~n22132;
  assign n22134 = ~n22129 & ~n22133;
  assign n22135 = ~pi0113 & ~n20630;
  assign n22136 = pi0113 & n20626;
  assign n22137 = ~n22135 & ~n22136;
  assign n22138 = ~pi0112 & n20617;
  assign n22139 = pi0112 & n20613;
  assign n22140 = ~n22138 & ~n22139;
  assign n22141 = ~n22137 & ~n22140;
  assign n22142 = ~pi0110 & ~n20599;
  assign n22143 = pi0110 & ~n20595;
  assign n22144 = pi0111 & ~n20581;
  assign n22145 = ~n22143 & ~n22144;
  assign n22146 = ~pi0111 & n20585;
  assign n22147 = n22145 & ~n22146;
  assign n22148 = ~n22142 & n22147;
  assign n22149 = ~n22141 & ~n22148;
  assign n22150 = ~pi0109 & n20557;
  assign n22151 = pi0081 & ~n20567;
  assign n22152 = ~n22150 & ~n22151;
  assign n22153 = ~pi0081 & ~n20571;
  assign n22154 = pi0109 & ~n20553;
  assign n22155 = ~n22153 & ~n22154;
  assign n22156 = n22152 & n22155;
  assign n22157 = n22141 & n22148;
  assign n22158 = ~n22156 & ~n22157;
  assign n22159 = ~n22149 & ~n22158;
  assign n22160 = ~n21990 & ~n21998;
  assign n22161 = ~n21997 & ~n22160;
  assign n22162 = n21982 & ~n21989;
  assign n22163 = ~n21982 & n21989;
  assign n22164 = ~n22162 & ~n22163;
  assign n22165 = n21997 & ~n22164;
  assign n22166 = ~n22161 & ~n22165;
  assign n22167 = n22159 & n22166;
  assign n22168 = ~n20546 & ~n22167;
  assign n22169 = n22133 & ~n22168;
  assign n22170 = ~n22134 & ~n22169;
  assign n22171 = ~n22055 & ~n22063;
  assign n22172 = ~n22064 & ~n22171;
  assign n22173 = n22030 & ~n22083;
  assign n22174 = ~n22030 & n22083;
  assign n22175 = ~n22173 & ~n22174;
  assign n22176 = ~n22172 & n22175;
  assign n22177 = n22172 & ~n22175;
  assign n22178 = ~n22176 & ~n22177;
  assign n22179 = pi0067 & n20688;
  assign n22180 = ~pi0067 & n20686;
  assign n22181 = ~n22179 & ~n22180;
  assign n22182 = ~pi0868 & n22068;
  assign n22183 = pi2384 & ~n11929;
  assign n22184 = pi0868 & n22183;
  assign n22185 = ~n22182 & ~n22184;
  assign n22186 = pi1472 & ~n22185;
  assign n22187 = ~n22181 & n22186;
  assign n22188 = ~pi0106 & ~n20677;
  assign n22189 = pi0106 & ~n20672;
  assign n22190 = pi0056 & ~n20681;
  assign n22191 = ~n22189 & ~n22190;
  assign n22192 = ~pi0056 & n20663;
  assign n22193 = n22191 & ~n22192;
  assign n22194 = ~n22188 & n22193;
  assign n22195 = n22181 & ~n22186;
  assign n22196 = ~n22194 & ~n22195;
  assign n22197 = ~n22187 & ~n22196;
  assign n22198 = ~pi0078 & n20775;
  assign n22199 = pi0078 & ~n20771;
  assign n22200 = ~n22198 & ~n22199;
  assign n22201 = ~pi0108 & ~n20762;
  assign n22202 = pi0108 & ~n20758;
  assign n22203 = ~n22201 & ~n22202;
  assign n22204 = n22200 & n22203;
  assign n22205 = ~pi0107 & n20747;
  assign n22206 = pi0107 & ~n20743;
  assign n22207 = ~n22205 & ~n22206;
  assign n22208 = ~pi0105 & ~n20734;
  assign n22209 = pi0105 & ~n20730;
  assign n22210 = ~n22208 & ~n22209;
  assign n22211 = n22207 & n22210;
  assign n22212 = ~n22204 & ~n22211;
  assign n22213 = ~pi0080 & ~n20806;
  assign n22214 = pi0080 & n20802;
  assign n22215 = ~n22213 & ~n22214;
  assign n22216 = ~pi0079 & n20793;
  assign n22217 = pi0079 & n20789;
  assign n22218 = ~n22216 & ~n22217;
  assign n22219 = ~n22215 & ~n22218;
  assign n22220 = n22204 & n22211;
  assign n22221 = ~n22219 & ~n22220;
  assign n22222 = ~n22212 & ~n22221;
  assign n22223 = ~n22197 & ~n22222;
  assign n22224 = ~n22073 & ~n22081;
  assign n22225 = ~n22080 & ~n22224;
  assign n22226 = n22067 & n22072;
  assign n22227 = ~n22067 & ~n22072;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = n22080 & ~n22228;
  assign n22230 = ~n22225 & ~n22229;
  assign n22231 = ~n22045 & ~n22053;
  assign n22232 = ~n22052 & ~n22231;
  assign n22233 = n22037 & ~n22044;
  assign n22234 = ~n22037 & n22044;
  assign n22235 = ~n22233 & ~n22234;
  assign n22236 = n22052 & ~n22235;
  assign n22237 = ~n22232 & ~n22236;
  assign n22238 = ~n22230 & ~n22237;
  assign n22239 = ~n22223 & ~n22238;
  assign n22240 = ~n22197 & ~n22237;
  assign n22241 = ~n22222 & ~n22230;
  assign n22242 = ~n22240 & ~n22241;
  assign n22243 = n22239 & n22242;
  assign n22244 = n22178 & n22243;
  assign n22245 = ~n22030 & ~n22083;
  assign n22246 = ~n22171 & ~n22245;
  assign n22247 = ~n22178 & n22246;
  assign n22248 = ~n22244 & ~n22247;
  assign n22249 = ~n22127 & ~n22248;
  assign n22250 = n22170 & ~n22249;
  assign n22251 = ~n22128 & ~n22250;
  assign n22252 = ~n22124 & n22248;
  assign n22253 = n22251 & ~n22252;
  assign n22254 = n22121 & n22253;
  assign n22255 = ~n22122 & ~n22254;
  assign n22256 = n22121 & ~n22253;
  assign n22257 = ~n22121 & n22253;
  assign n22258 = ~n22256 & ~n22257;
  assign n22259 = n22255 & n22258;
  assign n22260 = ~n21972 & ~n22097;
  assign n22261 = ~n22098 & ~n22260;
  assign n22262 = n22258 & ~n22261;
  assign n22263 = n22127 & n22248;
  assign n22264 = ~n22249 & ~n22263;
  assign n22265 = ~n22124 & ~n22170;
  assign n22266 = n22124 & n22170;
  assign n22267 = ~n22265 & ~n22266;
  assign n22268 = ~n22264 & n22267;
  assign n22269 = n22264 & ~n22267;
  assign n22270 = ~n22268 & ~n22269;
  assign n22271 = ~n22159 & n22166;
  assign n22272 = n22159 & ~n22166;
  assign n22273 = ~n22271 & ~n22272;
  assign n22274 = n20546 & ~n22273;
  assign n22275 = ~n20546 & n22273;
  assign n22276 = ~n22274 & ~n22275;
  assign n22277 = ~n22159 & ~n22166;
  assign n22278 = n22276 & ~n22277;
  assign n22279 = ~n22149 & ~n22157;
  assign n22280 = ~n22156 & ~n22279;
  assign n22281 = n22141 & ~n22148;
  assign n22282 = ~n22141 & n22148;
  assign n22283 = ~n22281 & ~n22282;
  assign n22284 = n22156 & ~n22283;
  assign n22285 = ~n22280 & ~n22284;
  assign n22286 = ~n20546 & ~n22285;
  assign n22287 = ~pi0105 & ~n20630;
  assign n22288 = pi0105 & n20626;
  assign n22289 = ~n22287 & ~n22288;
  assign n22290 = ~pi0113 & n20617;
  assign n22291 = pi0113 & n20613;
  assign n22292 = ~n22290 & ~n22291;
  assign n22293 = ~n22289 & ~n22292;
  assign n22294 = ~pi0111 & ~n20599;
  assign n22295 = pi0111 & ~n20595;
  assign n22296 = pi0112 & ~n20581;
  assign n22297 = ~n22295 & ~n22296;
  assign n22298 = ~pi0112 & n20585;
  assign n22299 = n22297 & ~n22298;
  assign n22300 = ~n22294 & n22299;
  assign n22301 = ~n22293 & ~n22300;
  assign n22302 = ~pi0109 & ~n20571;
  assign n22303 = pi0109 & ~n20567;
  assign n22304 = pi0110 & ~n20553;
  assign n22305 = ~n22303 & ~n22304;
  assign n22306 = ~pi0110 & n20557;
  assign n22307 = n22305 & ~n22306;
  assign n22308 = ~n22302 & n22307;
  assign n22309 = n22293 & n22300;
  assign n22310 = ~n22308 & ~n22309;
  assign n22311 = ~n22301 & ~n22310;
  assign n22312 = ~pi0081 & ~n20532;
  assign n22313 = pi0081 & ~n20528;
  assign n22314 = ~n22312 & ~n22313;
  assign n22315 = ~n20545 & ~n22314;
  assign n22316 = n20686 & ~n22315;
  assign n22317 = ~n22311 & n22316;
  assign n22318 = ~n22286 & ~n22317;
  assign n22319 = ~n20546 & ~n22311;
  assign n22320 = ~n22285 & n22316;
  assign n22321 = ~n22319 & ~n22320;
  assign n22322 = n22318 & n22321;
  assign n22323 = ~n22276 & n22322;
  assign n22324 = ~n22278 & ~n22323;
  assign n22325 = ~n22178 & ~n22243;
  assign n22326 = ~n22244 & ~n22325;
  assign n22327 = n22324 & ~n22326;
  assign n22328 = ~n22133 & n22168;
  assign n22329 = ~n22169 & ~n22328;
  assign n22330 = ~n22222 & ~n22237;
  assign n22331 = n22222 & n22237;
  assign n22332 = ~n22330 & ~n22331;
  assign n22333 = ~n22197 & n22230;
  assign n22334 = n22197 & ~n22230;
  assign n22335 = ~n22333 & ~n22334;
  assign n22336 = ~n22332 & n22335;
  assign n22337 = n22332 & ~n22335;
  assign n22338 = ~n22336 & ~n22337;
  assign n22339 = pi0114 & n20688;
  assign n22340 = ~pi0114 & n20686;
  assign n22341 = ~n22339 & ~n22340;
  assign n22342 = ~pi0868 & n22183;
  assign n22343 = pi2384 & ~n10966;
  assign n22344 = pi0868 & n22343;
  assign n22345 = ~n22342 & ~n22344;
  assign n22346 = pi1472 & ~n22345;
  assign n22347 = ~n22341 & n22346;
  assign n22348 = ~pi0056 & ~n20677;
  assign n22349 = pi0056 & ~n20672;
  assign n22350 = pi0067 & ~n20681;
  assign n22351 = ~n22349 & ~n22350;
  assign n22352 = ~pi0067 & n20663;
  assign n22353 = n22351 & ~n22352;
  assign n22354 = ~n22348 & n22353;
  assign n22355 = n22341 & ~n22346;
  assign n22356 = ~n22354 & ~n22355;
  assign n22357 = ~n22347 & ~n22356;
  assign n22358 = ~pi0106 & ~n20806;
  assign n22359 = pi0106 & n20802;
  assign n22360 = ~n22358 & ~n22359;
  assign n22361 = ~pi0080 & n20793;
  assign n22362 = pi0080 & n20789;
  assign n22363 = ~n22361 & ~n22362;
  assign n22364 = ~n22360 & ~n22363;
  assign n22365 = ~pi0078 & ~n20762;
  assign n22366 = pi0078 & ~n20758;
  assign n22367 = pi0079 & ~n20771;
  assign n22368 = ~n22366 & ~n22367;
  assign n22369 = ~pi0079 & n20775;
  assign n22370 = n22368 & ~n22369;
  assign n22371 = ~n22365 & n22370;
  assign n22372 = ~n22364 & ~n22371;
  assign n22373 = ~pi0107 & ~n20734;
  assign n22374 = pi0107 & ~n20730;
  assign n22375 = pi0108 & ~n20743;
  assign n22376 = ~n22374 & ~n22375;
  assign n22377 = ~pi0108 & n20747;
  assign n22378 = n22376 & ~n22377;
  assign n22379 = ~n22373 & n22378;
  assign n22380 = n22364 & n22371;
  assign n22381 = ~n22379 & ~n22380;
  assign n22382 = ~n22372 & ~n22381;
  assign n22383 = ~n22357 & ~n22382;
  assign n22384 = ~n22212 & ~n22220;
  assign n22385 = ~n22219 & ~n22384;
  assign n22386 = n22204 & ~n22211;
  assign n22387 = ~n22204 & n22211;
  assign n22388 = ~n22386 & ~n22387;
  assign n22389 = n22219 & ~n22388;
  assign n22390 = ~n22385 & ~n22389;
  assign n22391 = ~n22187 & ~n22195;
  assign n22392 = ~n22194 & ~n22391;
  assign n22393 = n22181 & n22186;
  assign n22394 = ~n22181 & ~n22186;
  assign n22395 = ~n22393 & ~n22394;
  assign n22396 = n22194 & ~n22395;
  assign n22397 = ~n22392 & ~n22396;
  assign n22398 = ~n22390 & ~n22397;
  assign n22399 = ~n22383 & ~n22398;
  assign n22400 = ~n22357 & ~n22390;
  assign n22401 = ~n22382 & ~n22397;
  assign n22402 = ~n22400 & ~n22401;
  assign n22403 = n22399 & n22402;
  assign n22404 = n22338 & n22403;
  assign n22405 = ~n22197 & ~n22230;
  assign n22406 = ~n22330 & ~n22405;
  assign n22407 = ~n22338 & n22406;
  assign n22408 = ~n22404 & ~n22407;
  assign n22409 = ~n22329 & n22408;
  assign n22410 = ~n22327 & ~n22409;
  assign n22411 = n22324 & n22408;
  assign n22412 = ~n22326 & ~n22329;
  assign n22413 = ~n22411 & ~n22412;
  assign n22414 = n22410 & n22413;
  assign n22415 = n22270 & n22414;
  assign n22416 = ~n22124 & n22170;
  assign n22417 = ~n22263 & ~n22416;
  assign n22418 = ~n22270 & n22417;
  assign n22419 = ~n22415 & ~n22418;
  assign n22420 = n22255 & n22419;
  assign n22421 = ~n22262 & ~n22420;
  assign n22422 = ~n22261 & n22419;
  assign n22423 = n22421 & ~n22422;
  assign n22424 = ~n22259 & n22423;
  assign n22425 = n22276 & n22322;
  assign n22426 = ~n22276 & ~n22322;
  assign n22427 = ~n22425 & ~n22426;
  assign n22428 = ~n22285 & ~n22311;
  assign n22429 = n22285 & n22311;
  assign n22430 = ~n22428 & ~n22429;
  assign n22431 = n20546 & n22316;
  assign n22432 = ~n20546 & ~n22316;
  assign n22433 = ~n22431 & ~n22432;
  assign n22434 = ~n22430 & n22433;
  assign n22435 = n22430 & ~n22433;
  assign n22436 = ~n22434 & ~n22435;
  assign n22437 = pi2384 & ~n17331;
  assign n22438 = pi1472 & n22437;
  assign n22439 = pi0868 & n22438;
  assign n22440 = n20663 & n22439;
  assign n22441 = ~pi0109 & ~n20532;
  assign n22442 = pi0109 & ~n20528;
  assign n22443 = ~n22441 & ~n22442;
  assign n22444 = ~pi0081 & n20543;
  assign n22445 = pi0081 & n20539;
  assign n22446 = ~n22444 & ~n22445;
  assign n22447 = ~n22443 & ~n22446;
  assign n22448 = ~n20663 & ~n22439;
  assign n22449 = ~n22447 & ~n22448;
  assign n22450 = ~n22440 & ~n22449;
  assign n22451 = ~pi0107 & ~n20630;
  assign n22452 = pi0107 & n20626;
  assign n22453 = ~n22451 & ~n22452;
  assign n22454 = ~pi0105 & n20617;
  assign n22455 = pi0105 & n20613;
  assign n22456 = ~n22454 & ~n22455;
  assign n22457 = ~n22453 & ~n22456;
  assign n22458 = ~pi0112 & ~n20599;
  assign n22459 = pi0112 & ~n20595;
  assign n22460 = pi0113 & ~n20581;
  assign n22461 = ~n22459 & ~n22460;
  assign n22462 = ~pi0113 & n20585;
  assign n22463 = n22461 & ~n22462;
  assign n22464 = ~n22458 & n22463;
  assign n22465 = ~n22457 & ~n22464;
  assign n22466 = ~pi0110 & ~n20571;
  assign n22467 = pi0110 & ~n20567;
  assign n22468 = pi0111 & ~n20553;
  assign n22469 = ~n22467 & ~n22468;
  assign n22470 = ~pi0111 & n20557;
  assign n22471 = n22469 & ~n22470;
  assign n22472 = ~n22466 & n22471;
  assign n22473 = n22457 & n22464;
  assign n22474 = ~n22472 & ~n22473;
  assign n22475 = ~n22465 & ~n22474;
  assign n22476 = ~n22450 & ~n22475;
  assign n22477 = ~n22301 & ~n22309;
  assign n22478 = ~n22308 & ~n22477;
  assign n22479 = n22293 & ~n22300;
  assign n22480 = ~n22293 & n22300;
  assign n22481 = ~n22479 & ~n22480;
  assign n22482 = n22308 & ~n22481;
  assign n22483 = ~n22478 & ~n22482;
  assign n22484 = n20686 & n22315;
  assign n22485 = ~n20686 & ~n22315;
  assign n22486 = ~n22484 & ~n22485;
  assign n22487 = ~n22483 & ~n22486;
  assign n22488 = ~n22476 & ~n22487;
  assign n22489 = ~n22450 & ~n22483;
  assign n22490 = ~n22475 & ~n22486;
  assign n22491 = ~n22489 & ~n22490;
  assign n22492 = n22488 & n22491;
  assign n22493 = n22436 & n22492;
  assign n22494 = ~n20546 & n22316;
  assign n22495 = ~n22428 & ~n22494;
  assign n22496 = ~n22436 & n22495;
  assign n22497 = ~n22493 & ~n22496;
  assign n22498 = n22427 & n22497;
  assign n22499 = ~n22427 & ~n22497;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = ~n22382 & ~n22390;
  assign n22502 = n22382 & n22390;
  assign n22503 = ~n22501 & ~n22502;
  assign n22504 = ~n22357 & ~n22397;
  assign n22505 = n22357 & n22397;
  assign n22506 = ~n22504 & ~n22505;
  assign n22507 = ~n22503 & n22506;
  assign n22508 = n22503 & ~n22506;
  assign n22509 = ~n22507 & ~n22508;
  assign n22510 = ~n22347 & ~n22355;
  assign n22511 = ~n22354 & ~n22510;
  assign n22512 = n22341 & n22346;
  assign n22513 = ~n22341 & ~n22346;
  assign n22514 = ~n22512 & ~n22513;
  assign n22515 = n22354 & ~n22514;
  assign n22516 = ~n22511 & ~n22515;
  assign n22517 = ~pi0868 & pi1472;
  assign n22518 = n22343 & n22517;
  assign n22519 = pi0868 & ~pi1789;
  assign n22520 = ~n22518 & ~n22519;
  assign n22521 = ~pi0067 & ~n20677;
  assign n22522 = ~pi0114 & n20663;
  assign n22523 = ~n22521 & ~n22522;
  assign n22524 = pi0067 & ~n20672;
  assign n22525 = pi0114 & ~n20681;
  assign n22526 = ~n22524 & ~n22525;
  assign n22527 = n22523 & n22526;
  assign n22528 = ~n22520 & ~n22527;
  assign n22529 = n22516 & ~n22528;
  assign n22530 = ~pi0056 & ~n20806;
  assign n22531 = pi0056 & n20802;
  assign n22532 = ~n22530 & ~n22531;
  assign n22533 = ~pi0106 & n20793;
  assign n22534 = pi0106 & n20789;
  assign n22535 = ~n22533 & ~n22534;
  assign n22536 = ~n22532 & ~n22535;
  assign n22537 = ~pi0079 & ~n20762;
  assign n22538 = pi0079 & ~n20758;
  assign n22539 = pi0080 & ~n20771;
  assign n22540 = ~n22538 & ~n22539;
  assign n22541 = ~pi0080 & n20775;
  assign n22542 = n22540 & ~n22541;
  assign n22543 = ~n22537 & n22542;
  assign n22544 = ~n22536 & ~n22543;
  assign n22545 = ~pi0108 & ~n20734;
  assign n22546 = pi0108 & ~n20730;
  assign n22547 = pi0078 & ~n20743;
  assign n22548 = ~n22546 & ~n22547;
  assign n22549 = ~pi0078 & n20747;
  assign n22550 = n22548 & ~n22549;
  assign n22551 = ~n22545 & n22550;
  assign n22552 = n22536 & n22543;
  assign n22553 = ~n22551 & ~n22552;
  assign n22554 = ~n22544 & ~n22553;
  assign n22555 = ~n22529 & ~n22554;
  assign n22556 = ~n22372 & ~n22380;
  assign n22557 = ~n22379 & ~n22556;
  assign n22558 = n22364 & ~n22371;
  assign n22559 = ~n22364 & n22371;
  assign n22560 = ~n22558 & ~n22559;
  assign n22561 = n22379 & ~n22560;
  assign n22562 = ~n22557 & ~n22561;
  assign n22563 = n22528 & ~n22562;
  assign n22564 = ~n22555 & ~n22563;
  assign n22565 = ~n22516 & ~n22562;
  assign n22566 = n22564 & ~n22565;
  assign n22567 = ~n22509 & n22566;
  assign n22568 = ~n22501 & ~n22504;
  assign n22569 = n22509 & n22568;
  assign n22570 = ~n22567 & ~n22569;
  assign n22571 = ~n22338 & ~n22403;
  assign n22572 = ~n22404 & ~n22571;
  assign n22573 = ~n22570 & ~n22572;
  assign n22574 = n22570 & n22572;
  assign n22575 = ~n22573 & ~n22574;
  assign n22576 = ~n22500 & n22575;
  assign n22577 = n22500 & ~n22575;
  assign n22578 = ~n22576 & ~n22577;
  assign n22579 = n22436 & ~n22492;
  assign n22580 = ~n22436 & n22492;
  assign n22581 = ~n22579 & ~n22580;
  assign n22582 = ~n22475 & ~n22483;
  assign n22583 = n22475 & n22483;
  assign n22584 = ~n22582 & ~n22583;
  assign n22585 = ~n22450 & n22486;
  assign n22586 = n22450 & ~n22486;
  assign n22587 = ~n22585 & ~n22586;
  assign n22588 = ~n22584 & n22587;
  assign n22589 = n22584 & ~n22587;
  assign n22590 = ~n22588 & ~n22589;
  assign n22591 = pi2384 & ~n17075;
  assign n22592 = pi0868 & n22591;
  assign n22593 = ~pi0868 & n22437;
  assign n22594 = ~n22592 & ~n22593;
  assign n22595 = pi1472 & ~n22594;
  assign n22596 = ~n20677 & n22595;
  assign n22597 = ~pi0110 & ~n20532;
  assign n22598 = pi0110 & ~n20528;
  assign n22599 = ~n22597 & ~n22598;
  assign n22600 = ~pi0109 & n20543;
  assign n22601 = pi0109 & n20539;
  assign n22602 = ~n22600 & ~n22601;
  assign n22603 = ~n22599 & ~n22602;
  assign n22604 = n20677 & ~n22595;
  assign n22605 = ~n22603 & ~n22604;
  assign n22606 = ~n22596 & ~n22605;
  assign n22607 = ~pi0108 & ~n20630;
  assign n22608 = pi0108 & n20626;
  assign n22609 = ~n22607 & ~n22608;
  assign n22610 = ~pi0107 & n20617;
  assign n22611 = pi0107 & n20613;
  assign n22612 = ~n22610 & ~n22611;
  assign n22613 = ~n22609 & ~n22612;
  assign n22614 = ~pi0113 & ~n20599;
  assign n22615 = pi0113 & ~n20595;
  assign n22616 = pi0105 & ~n20581;
  assign n22617 = ~n22615 & ~n22616;
  assign n22618 = ~pi0105 & n20585;
  assign n22619 = n22617 & ~n22618;
  assign n22620 = ~n22614 & n22619;
  assign n22621 = ~n22613 & ~n22620;
  assign n22622 = ~pi0111 & ~n20571;
  assign n22623 = pi0111 & ~n20567;
  assign n22624 = pi0112 & ~n20553;
  assign n22625 = ~n22623 & ~n22624;
  assign n22626 = ~pi0112 & n20557;
  assign n22627 = n22625 & ~n22626;
  assign n22628 = ~n22622 & n22627;
  assign n22629 = n22613 & n22620;
  assign n22630 = ~n22628 & ~n22629;
  assign n22631 = ~n22621 & ~n22630;
  assign n22632 = ~n22606 & ~n22631;
  assign n22633 = ~n22465 & ~n22473;
  assign n22634 = ~n22472 & ~n22633;
  assign n22635 = n22457 & ~n22464;
  assign n22636 = ~n22457 & n22464;
  assign n22637 = ~n22635 & ~n22636;
  assign n22638 = n22472 & ~n22637;
  assign n22639 = ~n22634 & ~n22638;
  assign n22640 = ~n22440 & ~n22448;
  assign n22641 = ~n22447 & ~n22640;
  assign n22642 = n20663 & ~n22439;
  assign n22643 = ~n20663 & n22439;
  assign n22644 = ~n22642 & ~n22643;
  assign n22645 = n22447 & ~n22644;
  assign n22646 = ~n22641 & ~n22645;
  assign n22647 = ~n22639 & ~n22646;
  assign n22648 = ~n22632 & ~n22647;
  assign n22649 = ~n22606 & ~n22639;
  assign n22650 = ~n22631 & ~n22646;
  assign n22651 = ~n22649 & ~n22650;
  assign n22652 = n22648 & n22651;
  assign n22653 = n22590 & n22652;
  assign n22654 = ~n22450 & ~n22486;
  assign n22655 = ~n22582 & ~n22654;
  assign n22656 = ~n22590 & n22655;
  assign n22657 = ~n22653 & ~n22656;
  assign n22658 = ~n22581 & ~n22657;
  assign n22659 = ~n22554 & ~n22562;
  assign n22660 = n22554 & n22562;
  assign n22661 = ~n22659 & ~n22660;
  assign n22662 = ~n22516 & ~n22528;
  assign n22663 = n22516 & n22528;
  assign n22664 = ~n22662 & ~n22663;
  assign n22665 = ~n22661 & n22664;
  assign n22666 = n22661 & ~n22664;
  assign n22667 = ~n22665 & ~n22666;
  assign n22668 = ~pi0067 & ~n20806;
  assign n22669 = pi0067 & n20802;
  assign n22670 = ~n22668 & ~n22669;
  assign n22671 = ~pi0056 & n20793;
  assign n22672 = pi0056 & n20789;
  assign n22673 = ~n22671 & ~n22672;
  assign n22674 = ~n22670 & ~n22673;
  assign n22675 = ~pi0080 & ~n20762;
  assign n22676 = pi0080 & ~n20758;
  assign n22677 = pi0106 & ~n20771;
  assign n22678 = ~n22676 & ~n22677;
  assign n22679 = ~pi0106 & n20775;
  assign n22680 = n22678 & ~n22679;
  assign n22681 = ~n22675 & n22680;
  assign n22682 = ~n22674 & ~n22681;
  assign n22683 = ~pi0078 & ~n20734;
  assign n22684 = pi0078 & ~n20730;
  assign n22685 = pi0079 & ~n20743;
  assign n22686 = ~n22684 & ~n22685;
  assign n22687 = ~pi0079 & n20747;
  assign n22688 = n22686 & ~n22687;
  assign n22689 = ~n22683 & n22688;
  assign n22690 = n22674 & n22681;
  assign n22691 = ~n22689 & ~n22690;
  assign n22692 = ~n22682 & ~n22691;
  assign n22693 = ~n22520 & n22527;
  assign n22694 = n22520 & ~n22527;
  assign n22695 = ~n22693 & ~n22694;
  assign n22696 = ~n22692 & ~n22695;
  assign n22697 = ~pi0868 & ~pi1789;
  assign n22698 = ~pi0114 & ~n20677;
  assign n22699 = pi0114 & ~n20672;
  assign n22700 = ~n22698 & ~n22699;
  assign n22701 = n22697 & ~n22700;
  assign n22702 = ~n22544 & ~n22552;
  assign n22703 = ~n22551 & ~n22702;
  assign n22704 = n22536 & ~n22543;
  assign n22705 = ~n22536 & n22543;
  assign n22706 = ~n22704 & ~n22705;
  assign n22707 = n22551 & ~n22706;
  assign n22708 = ~n22703 & ~n22707;
  assign n22709 = n22701 & ~n22708;
  assign n22710 = ~n22696 & ~n22709;
  assign n22711 = ~n22692 & n22701;
  assign n22712 = ~n22695 & ~n22708;
  assign n22713 = ~n22711 & ~n22712;
  assign n22714 = n22710 & n22713;
  assign n22715 = n22667 & n22714;
  assign n22716 = ~n22516 & n22528;
  assign n22717 = ~n22659 & ~n22716;
  assign n22718 = ~n22667 & n22717;
  assign n22719 = ~n22715 & ~n22718;
  assign n22720 = ~n22658 & n22719;
  assign n22721 = ~n22509 & ~n22566;
  assign n22722 = n22509 & n22566;
  assign n22723 = ~n22721 & ~n22722;
  assign n22724 = n22657 & n22723;
  assign n22725 = ~n22720 & ~n22724;
  assign n22726 = n22581 & n22723;
  assign n22727 = n22725 & ~n22726;
  assign n22728 = n22578 & n22727;
  assign n22729 = n22570 & ~n22572;
  assign n22730 = ~n22498 & ~n22729;
  assign n22731 = ~n22578 & n22730;
  assign n22732 = ~n22728 & ~n22731;
  assign n22733 = n22427 & ~n22572;
  assign n22734 = ~n22570 & n22572;
  assign n22735 = n22497 & ~n22734;
  assign n22736 = ~n22733 & ~n22735;
  assign n22737 = n22427 & n22570;
  assign n22738 = n22736 & ~n22737;
  assign n22739 = n22326 & n22408;
  assign n22740 = ~n22326 & ~n22408;
  assign n22741 = ~n22739 & ~n22740;
  assign n22742 = ~n22324 & ~n22329;
  assign n22743 = n22324 & n22329;
  assign n22744 = ~n22742 & ~n22743;
  assign n22745 = ~n22741 & n22744;
  assign n22746 = n22741 & ~n22744;
  assign n22747 = ~n22745 & ~n22746;
  assign n22748 = n22738 & ~n22747;
  assign n22749 = ~n22738 & n22747;
  assign n22750 = ~n22748 & ~n22749;
  assign n22751 = ~n22732 & n22750;
  assign n22752 = n22270 & ~n22414;
  assign n22753 = ~n22270 & n22414;
  assign n22754 = ~n22752 & ~n22753;
  assign n22755 = n22324 & ~n22329;
  assign n22756 = ~n22326 & n22408;
  assign n22757 = ~n22755 & ~n22756;
  assign n22758 = n22747 & n22757;
  assign n22759 = ~n22748 & ~n22758;
  assign n22760 = ~n22754 & ~n22759;
  assign n22761 = ~n22751 & ~n22760;
  assign n22762 = ~n22424 & n22761;
  assign n22763 = n22110 & n22762;
  assign n22764 = ~n22719 & n22723;
  assign n22765 = n22719 & ~n22723;
  assign n22766 = ~n22764 & ~n22765;
  assign n22767 = n22581 & n22657;
  assign n22768 = ~n22658 & ~n22767;
  assign n22769 = ~n22766 & n22768;
  assign n22770 = n22766 & ~n22768;
  assign n22771 = ~n22769 & ~n22770;
  assign n22772 = n22667 & ~n22714;
  assign n22773 = ~n22667 & n22714;
  assign n22774 = ~n22772 & ~n22773;
  assign n22775 = n22590 & ~n22652;
  assign n22776 = ~n22590 & n22652;
  assign n22777 = ~n22775 & ~n22776;
  assign n22778 = n22774 & n22777;
  assign n22779 = n22631 & n22639;
  assign n22780 = ~n22631 & ~n22639;
  assign n22781 = ~n22779 & ~n22780;
  assign n22782 = n22606 & n22646;
  assign n22783 = ~n22606 & ~n22646;
  assign n22784 = ~n22782 & ~n22783;
  assign n22785 = ~n22781 & n22784;
  assign n22786 = n22781 & ~n22784;
  assign n22787 = ~n22785 & ~n22786;
  assign n22788 = ~pi0078 & ~n20630;
  assign n22789 = pi0078 & n20626;
  assign n22790 = ~n22788 & ~n22789;
  assign n22791 = ~pi0108 & n20617;
  assign n22792 = pi0108 & n20613;
  assign n22793 = ~n22791 & ~n22792;
  assign n22794 = ~n22790 & ~n22793;
  assign n22795 = ~pi0105 & ~n20599;
  assign n22796 = pi0105 & ~n20595;
  assign n22797 = pi0107 & ~n20581;
  assign n22798 = ~n22796 & ~n22797;
  assign n22799 = ~pi0107 & n20585;
  assign n22800 = n22798 & ~n22799;
  assign n22801 = ~n22795 & n22800;
  assign n22802 = ~n22794 & ~n22801;
  assign n22803 = ~pi0112 & ~n20571;
  assign n22804 = pi0112 & ~n20567;
  assign n22805 = pi0113 & ~n20553;
  assign n22806 = ~n22804 & ~n22805;
  assign n22807 = ~pi0113 & n20557;
  assign n22808 = n22806 & ~n22807;
  assign n22809 = ~n22803 & n22808;
  assign n22810 = n22794 & n22801;
  assign n22811 = ~n22809 & ~n22810;
  assign n22812 = ~n22802 & ~n22811;
  assign n22813 = pi2384 & ~n9515;
  assign n22814 = pi0868 & n22813;
  assign n22815 = ~pi0868 & n22591;
  assign n22816 = ~n22814 & ~n22815;
  assign n22817 = pi1472 & ~n22816;
  assign n22818 = n20806 & n22817;
  assign n22819 = ~pi0111 & ~n20532;
  assign n22820 = pi0111 & ~n20528;
  assign n22821 = ~n22819 & ~n22820;
  assign n22822 = ~pi0110 & n20543;
  assign n22823 = pi0110 & n20539;
  assign n22824 = ~n22822 & ~n22823;
  assign n22825 = ~n22821 & ~n22824;
  assign n22826 = ~n20806 & ~n22817;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~n22818 & ~n22827;
  assign n22829 = ~n22596 & ~n22604;
  assign n22830 = ~n22603 & ~n22829;
  assign n22831 = n20677 & n22595;
  assign n22832 = ~n20677 & ~n22595;
  assign n22833 = ~n22831 & ~n22832;
  assign n22834 = n22603 & ~n22833;
  assign n22835 = ~n22830 & ~n22834;
  assign n22836 = n22828 & n22835;
  assign n22837 = ~n22812 & ~n22836;
  assign n22838 = ~n22621 & ~n22629;
  assign n22839 = ~n22628 & ~n22838;
  assign n22840 = n22613 & ~n22620;
  assign n22841 = ~n22613 & n22620;
  assign n22842 = ~n22840 & ~n22841;
  assign n22843 = n22628 & ~n22842;
  assign n22844 = ~n22839 & ~n22843;
  assign n22845 = ~n22828 & ~n22844;
  assign n22846 = ~n22837 & ~n22845;
  assign n22847 = ~n22835 & ~n22844;
  assign n22848 = n22846 & ~n22847;
  assign n22849 = ~n22787 & n22848;
  assign n22850 = ~n22780 & ~n22783;
  assign n22851 = n22787 & n22850;
  assign n22852 = ~n22849 & ~n22851;
  assign n22853 = ~pi0114 & ~n20806;
  assign n22854 = pi0114 & n20802;
  assign n22855 = ~n22853 & ~n22854;
  assign n22856 = ~pi0067 & n20793;
  assign n22857 = pi0067 & n20789;
  assign n22858 = ~n22856 & ~n22857;
  assign n22859 = ~n22855 & ~n22858;
  assign n22860 = ~pi0106 & ~n20762;
  assign n22861 = pi0106 & ~n20758;
  assign n22862 = pi0056 & ~n20771;
  assign n22863 = ~n22861 & ~n22862;
  assign n22864 = ~pi0056 & n20775;
  assign n22865 = n22863 & ~n22864;
  assign n22866 = ~n22860 & n22865;
  assign n22867 = ~n22859 & ~n22866;
  assign n22868 = ~pi0079 & ~n20734;
  assign n22869 = pi0079 & ~n20730;
  assign n22870 = pi0080 & ~n20743;
  assign n22871 = ~n22869 & ~n22870;
  assign n22872 = ~pi0080 & n20747;
  assign n22873 = n22871 & ~n22872;
  assign n22874 = ~n22868 & n22873;
  assign n22875 = n22859 & n22866;
  assign n22876 = ~n22874 & ~n22875;
  assign n22877 = ~n22867 & ~n22876;
  assign n22878 = ~n22682 & ~n22690;
  assign n22879 = ~n22689 & ~n22878;
  assign n22880 = n22674 & ~n22681;
  assign n22881 = ~n22674 & n22681;
  assign n22882 = ~n22880 & ~n22881;
  assign n22883 = n22689 & ~n22882;
  assign n22884 = ~n22879 & ~n22883;
  assign n22885 = n22877 & n22884;
  assign n22886 = ~n22697 & n22700;
  assign n22887 = ~n22701 & ~n22886;
  assign n22888 = ~n22885 & n22887;
  assign n22889 = n22692 & n22708;
  assign n22890 = ~n22692 & ~n22708;
  assign n22891 = ~n22889 & ~n22890;
  assign n22892 = n22695 & ~n22701;
  assign n22893 = ~n22695 & n22701;
  assign n22894 = ~n22892 & ~n22893;
  assign n22895 = ~n22891 & n22894;
  assign n22896 = n22891 & ~n22894;
  assign n22897 = ~n22895 & ~n22896;
  assign n22898 = ~n22888 & ~n22897;
  assign n22899 = ~n22890 & ~n22893;
  assign n22900 = n22897 & n22899;
  assign n22901 = ~n22898 & ~n22900;
  assign n22902 = ~n22774 & ~n22901;
  assign n22903 = n22852 & ~n22902;
  assign n22904 = ~n22778 & ~n22903;
  assign n22905 = n22777 & n22901;
  assign n22906 = n22904 & ~n22905;
  assign n22907 = n22771 & n22906;
  assign n22908 = n22719 & n22723;
  assign n22909 = ~n22767 & ~n22908;
  assign n22910 = ~n22771 & n22909;
  assign n22911 = ~n22907 & ~n22910;
  assign n22912 = ~n22578 & n22727;
  assign n22913 = n22578 & ~n22727;
  assign n22914 = ~n22912 & ~n22913;
  assign n22915 = ~n22911 & ~n22914;
  assign n22916 = ~pi0079 & ~n20630;
  assign n22917 = pi0079 & n20626;
  assign n22918 = ~n22916 & ~n22917;
  assign n22919 = ~pi0078 & n20617;
  assign n22920 = pi0078 & n20613;
  assign n22921 = ~n22919 & ~n22920;
  assign n22922 = ~n22918 & ~n22921;
  assign n22923 = ~pi0113 & ~n20571;
  assign n22924 = pi0113 & ~n20567;
  assign n22925 = pi0105 & ~n20553;
  assign n22926 = ~n22924 & ~n22925;
  assign n22927 = ~pi0105 & n20557;
  assign n22928 = n22926 & ~n22927;
  assign n22929 = ~n22923 & n22928;
  assign n22930 = ~n22922 & ~n22929;
  assign n22931 = ~pi0107 & ~n20599;
  assign n22932 = pi0107 & ~n20595;
  assign n22933 = pi0108 & ~n20581;
  assign n22934 = ~n22932 & ~n22933;
  assign n22935 = ~pi0108 & n20585;
  assign n22936 = n22934 & ~n22935;
  assign n22937 = ~n22931 & n22936;
  assign n22938 = n22922 & n22929;
  assign n22939 = ~n22937 & ~n22938;
  assign n22940 = ~n22930 & ~n22939;
  assign n22941 = ~n22802 & ~n22810;
  assign n22942 = ~n22809 & ~n22941;
  assign n22943 = n22794 & ~n22801;
  assign n22944 = ~n22794 & n22801;
  assign n22945 = ~n22943 & ~n22944;
  assign n22946 = n22809 & ~n22945;
  assign n22947 = ~n22942 & ~n22946;
  assign n22948 = n22940 & n22947;
  assign n22949 = pi2384 & ~n10424;
  assign n22950 = pi0868 & n22949;
  assign n22951 = ~pi0868 & n22813;
  assign n22952 = ~n22950 & ~n22951;
  assign n22953 = pi1472 & ~n22952;
  assign n22954 = n20793 & ~n22953;
  assign n22955 = ~pi0112 & ~n20532;
  assign n22956 = pi0112 & ~n20528;
  assign n22957 = ~n22955 & ~n22956;
  assign n22958 = ~pi0111 & n20543;
  assign n22959 = pi0111 & n20539;
  assign n22960 = ~n22958 & ~n22959;
  assign n22961 = ~n22957 & ~n22960;
  assign n22962 = ~n20793 & n22953;
  assign n22963 = n22961 & ~n22962;
  assign n22964 = ~n22954 & ~n22963;
  assign n22965 = ~n22818 & ~n22826;
  assign n22966 = ~n22825 & n22965;
  assign n22967 = n22825 & ~n22965;
  assign n22968 = ~n22966 & ~n22967;
  assign n22969 = ~n22964 & ~n22968;
  assign n22970 = ~n22948 & ~n22969;
  assign n22971 = n22812 & n22844;
  assign n22972 = ~n22812 & ~n22844;
  assign n22973 = ~n22971 & ~n22972;
  assign n22974 = ~n22828 & n22835;
  assign n22975 = n22828 & ~n22835;
  assign n22976 = ~n22974 & ~n22975;
  assign n22977 = ~n22973 & n22976;
  assign n22978 = n22973 & ~n22976;
  assign n22979 = ~n22977 & ~n22978;
  assign n22980 = ~n22970 & n22979;
  assign n22981 = ~n22828 & ~n22835;
  assign n22982 = ~n22972 & ~n22981;
  assign n22983 = ~n22979 & n22982;
  assign n22984 = ~n22980 & ~n22983;
  assign n22985 = ~n22877 & ~n22884;
  assign n22986 = ~n22885 & ~n22985;
  assign n22987 = n22887 & ~n22986;
  assign n22988 = ~n22887 & n22986;
  assign n22989 = ~n22987 & ~n22988;
  assign n22990 = ~n22884 & n22989;
  assign n22991 = ~n22877 & n22990;
  assign n22992 = n22984 & n22991;
  assign n22993 = n22888 & n22897;
  assign n22994 = ~n22898 & ~n22993;
  assign n22995 = n22787 & ~n22848;
  assign n22996 = ~n22849 & ~n22995;
  assign n22997 = ~n22994 & ~n22996;
  assign n22998 = ~n22992 & ~n22997;
  assign n22999 = n22984 & ~n22994;
  assign n23000 = n22991 & ~n22996;
  assign n23001 = ~n22999 & ~n23000;
  assign n23002 = n22998 & n23001;
  assign n23003 = n22774 & ~n22901;
  assign n23004 = ~n22774 & n22901;
  assign n23005 = ~n23003 & ~n23004;
  assign n23006 = n22777 & n22852;
  assign n23007 = ~n22777 & ~n22852;
  assign n23008 = ~n23006 & ~n23007;
  assign n23009 = ~n23005 & n23008;
  assign n23010 = n23005 & ~n23008;
  assign n23011 = ~n23009 & ~n23010;
  assign n23012 = n23002 & n23011;
  assign n23013 = n22774 & n22901;
  assign n23014 = ~n23006 & ~n23013;
  assign n23015 = ~n23011 & n23014;
  assign n23016 = ~n23012 & ~n23015;
  assign n23017 = n22771 & ~n22906;
  assign n23018 = ~n22771 & n22906;
  assign n23019 = ~n23017 & ~n23018;
  assign n23020 = ~n23016 & ~n23019;
  assign n23021 = ~n22915 & ~n23020;
  assign n23022 = ~pi0080 & ~n20630;
  assign n23023 = pi0080 & n20626;
  assign n23024 = ~n23022 & ~n23023;
  assign n23025 = ~pi0079 & n20617;
  assign n23026 = pi0079 & n20613;
  assign n23027 = ~n23025 & ~n23026;
  assign n23028 = ~n23024 & ~n23027;
  assign n23029 = ~pi0108 & ~n20599;
  assign n23030 = pi0108 & ~n20595;
  assign n23031 = pi0078 & ~n20581;
  assign n23032 = ~n23030 & ~n23031;
  assign n23033 = ~pi0078 & n20585;
  assign n23034 = n23032 & ~n23033;
  assign n23035 = ~n23029 & n23034;
  assign n23036 = ~n23028 & ~n23035;
  assign n23037 = ~pi0105 & ~n20571;
  assign n23038 = pi0105 & ~n20567;
  assign n23039 = pi0107 & ~n20553;
  assign n23040 = ~n23038 & ~n23039;
  assign n23041 = ~pi0107 & n20557;
  assign n23042 = n23040 & ~n23041;
  assign n23043 = ~n23037 & n23042;
  assign n23044 = n23028 & n23035;
  assign n23045 = ~n23043 & ~n23044;
  assign n23046 = ~n23036 & ~n23045;
  assign n23047 = ~n22930 & ~n22938;
  assign n23048 = ~n22937 & ~n23047;
  assign n23049 = n22922 & ~n22929;
  assign n23050 = ~n22922 & n22929;
  assign n23051 = ~n23049 & ~n23050;
  assign n23052 = n22937 & ~n23051;
  assign n23053 = ~n23048 & ~n23052;
  assign n23054 = n23046 & n23053;
  assign n23055 = ~pi0868 & n22949;
  assign n23056 = pi2384 & ~n15263;
  assign n23057 = pi0868 & n23056;
  assign n23058 = ~n23055 & ~n23057;
  assign n23059 = pi1472 & ~n23058;
  assign n23060 = ~n20775 & ~n23059;
  assign n23061 = pi0113 & ~n20528;
  assign n23062 = ~pi0113 & ~n20532;
  assign n23063 = ~n23061 & ~n23062;
  assign n23064 = ~pi0112 & n20543;
  assign n23065 = pi0112 & n20539;
  assign n23066 = ~n23064 & ~n23065;
  assign n23067 = ~n23063 & ~n23066;
  assign n23068 = n20775 & n23059;
  assign n23069 = n23067 & ~n23068;
  assign n23070 = ~n23060 & ~n23069;
  assign n23071 = ~n22954 & ~n22962;
  assign n23072 = n22961 & ~n23071;
  assign n23073 = ~n20793 & ~n22953;
  assign n23074 = n20793 & n22953;
  assign n23075 = ~n23073 & ~n23074;
  assign n23076 = ~n22961 & ~n23075;
  assign n23077 = ~n23072 & ~n23076;
  assign n23078 = ~n23070 & ~n23077;
  assign n23079 = ~n23054 & ~n23078;
  assign n23080 = ~n22940 & ~n22947;
  assign n23081 = ~n22948 & ~n23080;
  assign n23082 = ~n22964 & n22968;
  assign n23083 = n22964 & ~n22968;
  assign n23084 = ~n23082 & ~n23083;
  assign n23085 = ~n23081 & n23084;
  assign n23086 = n23081 & ~n23084;
  assign n23087 = ~n23085 & ~n23086;
  assign n23088 = n23079 & n23087;
  assign n23089 = ~n23079 & ~n23087;
  assign n23090 = ~n23088 & ~n23089;
  assign n23091 = ~pi0067 & ~n20762;
  assign n23092 = pi0067 & ~n20758;
  assign n23093 = pi0114 & ~n20771;
  assign n23094 = ~n23092 & ~n23093;
  assign n23095 = ~pi0114 & n20775;
  assign n23096 = n23094 & ~n23095;
  assign n23097 = ~n23091 & n23096;
  assign n23098 = ~pi0106 & ~n20734;
  assign n23099 = pi0106 & ~n20730;
  assign n23100 = pi0056 & ~n20743;
  assign n23101 = ~n23099 & ~n23100;
  assign n23102 = ~pi0056 & n20747;
  assign n23103 = n23101 & ~n23102;
  assign n23104 = ~n23098 & n23103;
  assign n23105 = ~n23097 & ~n23104;
  assign n23106 = ~pi0080 & ~n20734;
  assign n23107 = pi0080 & ~n20730;
  assign n23108 = pi0106 & ~n20743;
  assign n23109 = ~n23107 & ~n23108;
  assign n23110 = ~pi0106 & n20747;
  assign n23111 = n23109 & ~n23110;
  assign n23112 = ~n23106 & n23111;
  assign n23113 = pi0114 & ~n20789;
  assign n23114 = ~pi0114 & ~n20793;
  assign n23115 = ~n23113 & ~n23114;
  assign n23116 = ~pi0056 & ~n20762;
  assign n23117 = pi0056 & ~n20758;
  assign n23118 = pi0067 & ~n20771;
  assign n23119 = ~n23117 & ~n23118;
  assign n23120 = ~pi0067 & n20775;
  assign n23121 = n23119 & ~n23120;
  assign n23122 = ~n23116 & n23121;
  assign n23123 = ~n23115 & ~n23122;
  assign n23124 = n23115 & n23122;
  assign n23125 = ~n23123 & ~n23124;
  assign n23126 = ~n23112 & ~n23125;
  assign n23127 = n23115 & ~n23122;
  assign n23128 = ~n23115 & n23122;
  assign n23129 = ~n23127 & ~n23128;
  assign n23130 = n23112 & ~n23129;
  assign n23131 = ~n23126 & ~n23130;
  assign n23132 = ~n23105 & n23131;
  assign n23133 = n23105 & ~n23131;
  assign n23134 = ~n23132 & ~n23133;
  assign n23135 = ~n23131 & ~n23134;
  assign n23136 = n23105 & n23135;
  assign n23137 = n23090 & n23136;
  assign n23138 = ~n23046 & ~n23053;
  assign n23139 = ~n23054 & ~n23138;
  assign n23140 = n23070 & ~n23077;
  assign n23141 = ~n23070 & n23077;
  assign n23142 = ~n23140 & ~n23141;
  assign n23143 = ~n23139 & n23142;
  assign n23144 = n23139 & ~n23142;
  assign n23145 = ~n23143 & ~n23144;
  assign n23146 = ~pi0106 & ~n20630;
  assign n23147 = pi0106 & n20626;
  assign n23148 = ~n23146 & ~n23147;
  assign n23149 = ~pi0080 & n20617;
  assign n23150 = pi0080 & n20613;
  assign n23151 = ~n23149 & ~n23150;
  assign n23152 = ~n23148 & ~n23151;
  assign n23153 = ~pi0078 & ~n20599;
  assign n23154 = pi0078 & ~n20595;
  assign n23155 = pi0079 & ~n20581;
  assign n23156 = ~n23154 & ~n23155;
  assign n23157 = ~pi0079 & n20585;
  assign n23158 = n23156 & ~n23157;
  assign n23159 = ~n23153 & n23158;
  assign n23160 = ~n23152 & ~n23159;
  assign n23161 = ~pi0107 & ~n20571;
  assign n23162 = pi0107 & ~n20567;
  assign n23163 = pi0108 & ~n20553;
  assign n23164 = ~n23162 & ~n23163;
  assign n23165 = ~pi0108 & n20557;
  assign n23166 = n23164 & ~n23165;
  assign n23167 = ~n23161 & n23166;
  assign n23168 = n23152 & n23159;
  assign n23169 = ~n23167 & ~n23168;
  assign n23170 = ~n23160 & ~n23169;
  assign n23171 = ~n23036 & ~n23044;
  assign n23172 = ~n23043 & ~n23171;
  assign n23173 = n23028 & ~n23035;
  assign n23174 = ~n23028 & n23035;
  assign n23175 = ~n23173 & ~n23174;
  assign n23176 = n23043 & ~n23175;
  assign n23177 = ~n23172 & ~n23176;
  assign n23178 = n23170 & n23177;
  assign n23179 = ~pi0868 & n23056;
  assign n23180 = pi2384 & ~n14223;
  assign n23181 = pi0868 & n23180;
  assign n23182 = ~n23179 & ~n23181;
  assign n23183 = pi1472 & ~n23182;
  assign n23184 = n20762 & ~n23183;
  assign n23185 = ~pi0105 & ~n20532;
  assign n23186 = pi0105 & ~n20528;
  assign n23187 = ~n23185 & ~n23186;
  assign n23188 = ~pi0113 & n20543;
  assign n23189 = pi0113 & n20539;
  assign n23190 = ~n23188 & ~n23189;
  assign n23191 = ~n23187 & ~n23190;
  assign n23192 = ~n20762 & n23183;
  assign n23193 = n23191 & ~n23192;
  assign n23194 = ~n23184 & ~n23193;
  assign n23195 = ~n23060 & ~n23068;
  assign n23196 = n23067 & ~n23195;
  assign n23197 = n20775 & ~n23059;
  assign n23198 = ~n20775 & n23059;
  assign n23199 = ~n23197 & ~n23198;
  assign n23200 = ~n23067 & ~n23199;
  assign n23201 = ~n23196 & ~n23200;
  assign n23202 = ~n23194 & ~n23201;
  assign n23203 = ~n23178 & ~n23202;
  assign n23204 = n23145 & ~n23203;
  assign n23205 = n23070 & n23077;
  assign n23206 = ~n23138 & ~n23205;
  assign n23207 = ~n23145 & n23206;
  assign n23208 = ~n23204 & ~n23207;
  assign n23209 = ~n22867 & ~n22875;
  assign n23210 = ~n22874 & ~n23209;
  assign n23211 = n22859 & ~n22866;
  assign n23212 = ~n22859 & n22866;
  assign n23213 = ~n23211 & ~n23212;
  assign n23214 = n22874 & ~n23213;
  assign n23215 = ~n23210 & ~n23214;
  assign n23216 = ~n23112 & ~n23124;
  assign n23217 = ~n23123 & ~n23216;
  assign n23218 = ~n23215 & n23217;
  assign n23219 = n23215 & ~n23217;
  assign n23220 = ~n23218 & ~n23219;
  assign n23221 = n23208 & ~n23220;
  assign n23222 = ~n23137 & ~n23221;
  assign n23223 = n23090 & ~n23220;
  assign n23224 = n23136 & n23208;
  assign n23225 = ~n23223 & ~n23224;
  assign n23226 = n23222 & n23225;
  assign n23227 = n22970 & ~n22979;
  assign n23228 = ~n22980 & ~n23227;
  assign n23229 = ~n23079 & n23087;
  assign n23230 = n22964 & n22968;
  assign n23231 = ~n23080 & ~n23230;
  assign n23232 = ~n23087 & n23231;
  assign n23233 = ~n23229 & ~n23232;
  assign n23234 = ~n23228 & ~n23233;
  assign n23235 = n23228 & n23233;
  assign n23236 = ~n23234 & ~n23235;
  assign n23237 = ~n23217 & n23220;
  assign n23238 = ~n23215 & n23237;
  assign n23239 = n22989 & ~n23238;
  assign n23240 = ~n22989 & n23238;
  assign n23241 = ~n23239 & ~n23240;
  assign n23242 = ~n23236 & n23241;
  assign n23243 = n23236 & ~n23241;
  assign n23244 = ~n23242 & ~n23243;
  assign n23245 = n23226 & n23244;
  assign n23246 = ~n23228 & n23233;
  assign n23247 = ~n23240 & ~n23246;
  assign n23248 = ~n23244 & n23247;
  assign n23249 = ~n23245 & ~n23248;
  assign n23250 = ~n23002 & ~n23011;
  assign n23251 = ~n23012 & ~n23250;
  assign n23252 = ~n22989 & ~n23228;
  assign n23253 = n23233 & n23238;
  assign n23254 = ~n23252 & ~n23253;
  assign n23255 = ~n23228 & n23238;
  assign n23256 = ~n22989 & n23233;
  assign n23257 = ~n23255 & ~n23256;
  assign n23258 = n23254 & n23257;
  assign n23259 = ~n22984 & n22996;
  assign n23260 = n22984 & ~n22996;
  assign n23261 = ~n23259 & ~n23260;
  assign n23262 = n22991 & n22994;
  assign n23263 = ~n22991 & ~n22994;
  assign n23264 = ~n23262 & ~n23263;
  assign n23265 = ~n23261 & n23264;
  assign n23266 = n23261 & ~n23264;
  assign n23267 = ~n23265 & ~n23266;
  assign n23268 = n23258 & n23267;
  assign n23269 = ~n23258 & ~n23267;
  assign n23270 = ~n23268 & ~n23269;
  assign n23271 = ~n23251 & ~n23270;
  assign n23272 = n22991 & ~n22994;
  assign n23273 = ~n23260 & ~n23272;
  assign n23274 = ~n23267 & n23273;
  assign n23275 = ~n23268 & ~n23274;
  assign n23276 = ~n23270 & n23275;
  assign n23277 = ~n23271 & ~n23276;
  assign n23278 = n23249 & ~n23277;
  assign n23279 = ~n23251 & n23275;
  assign n23280 = ~n23278 & ~n23279;
  assign n23281 = n23021 & ~n23280;
  assign n23282 = n22911 & n22914;
  assign n23283 = ~n23281 & ~n23282;
  assign n23284 = n23016 & n23019;
  assign n23285 = ~n22915 & n23284;
  assign n23286 = n23283 & ~n23285;
  assign n23287 = n22763 & ~n23286;
  assign n23288 = n22259 & n22419;
  assign n23289 = n22258 & n22422;
  assign n23290 = ~n23288 & ~n23289;
  assign n23291 = n22732 & ~n22750;
  assign n23292 = ~n22754 & ~n23291;
  assign n23293 = n22759 & ~n23292;
  assign n23294 = ~n22750 & n22754;
  assign n23295 = n22732 & n23294;
  assign n23296 = ~n23293 & ~n23295;
  assign n23297 = ~n22424 & ~n23296;
  assign n23298 = n22255 & ~n22261;
  assign n23299 = ~n23297 & ~n23298;
  assign n23300 = n23290 & n23299;
  assign n23301 = n22110 & ~n23300;
  assign n23302 = ~n23287 & ~n23301;
  assign n23303 = ~n21681 & ~n21684;
  assign n23304 = n21815 & ~n23303;
  assign n23305 = n21680 & ~n21683;
  assign n23306 = ~n23304 & ~n23305;
  assign n23307 = n23302 & n23306;
  assign n23308 = ~n22107 & n23307;
  assign n23309 = ~n23226 & ~n23244;
  assign n23310 = ~n23245 & ~n23309;
  assign n23311 = ~pi0056 & ~n20734;
  assign n23312 = pi0056 & ~n20730;
  assign n23313 = pi0067 & ~n20743;
  assign n23314 = ~n23312 & ~n23313;
  assign n23315 = ~pi0067 & n20747;
  assign n23316 = n23314 & ~n23315;
  assign n23317 = ~n23311 & n23316;
  assign n23318 = ~pi0114 & ~n20762;
  assign n23319 = pi0114 & ~n20758;
  assign n23320 = ~n23318 & ~n23319;
  assign n23321 = ~n23317 & ~n23320;
  assign n23322 = n23097 & ~n23104;
  assign n23323 = ~n23097 & n23104;
  assign n23324 = ~n23322 & ~n23323;
  assign n23325 = ~n23321 & n23324;
  assign n23326 = n23321 & ~n23324;
  assign n23327 = ~n23325 & ~n23326;
  assign n23328 = ~n23324 & ~n23327;
  assign n23329 = n23321 & n23328;
  assign n23330 = ~n23134 & ~n23329;
  assign n23331 = ~n23145 & n23203;
  assign n23332 = ~n23204 & ~n23331;
  assign n23333 = ~n23330 & ~n23332;
  assign n23334 = ~n23170 & ~n23177;
  assign n23335 = ~n23178 & ~n23334;
  assign n23336 = n23194 & ~n23201;
  assign n23337 = ~n23194 & n23201;
  assign n23338 = ~n23336 & ~n23337;
  assign n23339 = ~n23335 & n23338;
  assign n23340 = n23335 & ~n23338;
  assign n23341 = ~n23339 & ~n23340;
  assign n23342 = ~pi0056 & ~n20630;
  assign n23343 = pi0056 & n20626;
  assign n23344 = ~n23342 & ~n23343;
  assign n23345 = ~pi0106 & n20617;
  assign n23346 = pi0106 & n20613;
  assign n23347 = ~n23345 & ~n23346;
  assign n23348 = ~n23344 & ~n23347;
  assign n23349 = ~pi0108 & ~n20571;
  assign n23350 = pi0108 & ~n20567;
  assign n23351 = pi0078 & ~n20553;
  assign n23352 = ~n23350 & ~n23351;
  assign n23353 = ~pi0078 & n20557;
  assign n23354 = n23352 & ~n23353;
  assign n23355 = ~n23349 & n23354;
  assign n23356 = ~n23348 & ~n23355;
  assign n23357 = ~pi0079 & ~n20599;
  assign n23358 = pi0079 & ~n20595;
  assign n23359 = pi0080 & ~n20581;
  assign n23360 = ~n23358 & ~n23359;
  assign n23361 = ~pi0080 & n20585;
  assign n23362 = n23360 & ~n23361;
  assign n23363 = ~n23357 & n23362;
  assign n23364 = n23348 & n23355;
  assign n23365 = ~n23363 & ~n23364;
  assign n23366 = ~n23356 & ~n23365;
  assign n23367 = ~n23160 & ~n23168;
  assign n23368 = ~n23167 & ~n23367;
  assign n23369 = n23152 & ~n23159;
  assign n23370 = ~n23152 & n23159;
  assign n23371 = ~n23369 & ~n23370;
  assign n23372 = n23167 & ~n23371;
  assign n23373 = ~n23368 & ~n23372;
  assign n23374 = n23366 & n23373;
  assign n23375 = ~pi0868 & n23180;
  assign n23376 = pi2384 & ~n12613;
  assign n23377 = pi0868 & n23376;
  assign n23378 = ~n23375 & ~n23377;
  assign n23379 = pi1472 & ~n23378;
  assign n23380 = ~n20747 & ~n23379;
  assign n23381 = ~pi0107 & ~n20532;
  assign n23382 = pi0107 & ~n20528;
  assign n23383 = ~n23381 & ~n23382;
  assign n23384 = ~pi0105 & n20543;
  assign n23385 = pi0105 & n20539;
  assign n23386 = ~n23384 & ~n23385;
  assign n23387 = ~n23383 & ~n23386;
  assign n23388 = n20747 & n23379;
  assign n23389 = n23387 & ~n23388;
  assign n23390 = ~n23380 & ~n23389;
  assign n23391 = ~n23184 & ~n23192;
  assign n23392 = n23191 & ~n23391;
  assign n23393 = ~n20762 & ~n23183;
  assign n23394 = n20762 & n23183;
  assign n23395 = ~n23393 & ~n23394;
  assign n23396 = ~n23191 & ~n23395;
  assign n23397 = ~n23392 & ~n23396;
  assign n23398 = ~n23390 & ~n23397;
  assign n23399 = ~n23374 & ~n23398;
  assign n23400 = n23341 & ~n23399;
  assign n23401 = n23194 & n23201;
  assign n23402 = ~n23334 & ~n23401;
  assign n23403 = ~n23341 & n23402;
  assign n23404 = ~n23400 & ~n23403;
  assign n23405 = n23134 & n23404;
  assign n23406 = ~n23333 & ~n23405;
  assign n23407 = n23329 & n23404;
  assign n23408 = n23406 & ~n23407;
  assign n23409 = ~n23090 & ~n23208;
  assign n23410 = n23090 & n23208;
  assign n23411 = ~n23409 & ~n23410;
  assign n23412 = n23136 & n23220;
  assign n23413 = ~n23136 & ~n23220;
  assign n23414 = ~n23412 & ~n23413;
  assign n23415 = ~n23411 & n23414;
  assign n23416 = n23411 & ~n23414;
  assign n23417 = ~n23415 & ~n23416;
  assign n23418 = n23408 & n23417;
  assign n23419 = n23136 & ~n23220;
  assign n23420 = ~n23410 & ~n23419;
  assign n23421 = ~n23417 & n23420;
  assign n23422 = ~n23418 & ~n23421;
  assign n23423 = ~n23408 & ~n23417;
  assign n23424 = ~n23418 & ~n23423;
  assign n23425 = ~n23332 & n23404;
  assign n23426 = n23332 & ~n23404;
  assign n23427 = ~n23425 & ~n23426;
  assign n23428 = n23134 & ~n23329;
  assign n23429 = ~n23134 & n23329;
  assign n23430 = ~n23428 & ~n23429;
  assign n23431 = ~n23427 & n23430;
  assign n23432 = n23427 & ~n23430;
  assign n23433 = ~n23431 & ~n23432;
  assign n23434 = n23341 & n23399;
  assign n23435 = ~n23341 & ~n23399;
  assign n23436 = ~n23434 & ~n23435;
  assign n23437 = ~n23366 & ~n23373;
  assign n23438 = ~n23374 & ~n23437;
  assign n23439 = n23390 & ~n23397;
  assign n23440 = ~n23390 & n23397;
  assign n23441 = ~n23439 & ~n23440;
  assign n23442 = ~n23438 & n23441;
  assign n23443 = n23438 & ~n23441;
  assign n23444 = ~n23442 & ~n23443;
  assign n23445 = ~pi0067 & ~n20630;
  assign n23446 = pi0067 & n20626;
  assign n23447 = ~n23445 & ~n23446;
  assign n23448 = ~pi0056 & n20617;
  assign n23449 = pi0056 & n20613;
  assign n23450 = ~n23448 & ~n23449;
  assign n23451 = ~n23447 & ~n23450;
  assign n23452 = ~pi0078 & ~n20571;
  assign n23453 = pi0078 & ~n20567;
  assign n23454 = pi0079 & ~n20553;
  assign n23455 = ~n23453 & ~n23454;
  assign n23456 = ~pi0079 & n20557;
  assign n23457 = n23455 & ~n23456;
  assign n23458 = ~n23452 & n23457;
  assign n23459 = ~n23451 & ~n23458;
  assign n23460 = ~pi0080 & ~n20599;
  assign n23461 = pi0080 & ~n20595;
  assign n23462 = pi0106 & ~n20581;
  assign n23463 = ~n23461 & ~n23462;
  assign n23464 = ~pi0106 & n20585;
  assign n23465 = n23463 & ~n23464;
  assign n23466 = ~n23460 & n23465;
  assign n23467 = n23451 & n23458;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = ~n23459 & ~n23468;
  assign n23470 = ~n23356 & ~n23364;
  assign n23471 = ~n23363 & ~n23470;
  assign n23472 = n23348 & ~n23355;
  assign n23473 = ~n23348 & n23355;
  assign n23474 = ~n23472 & ~n23473;
  assign n23475 = n23363 & ~n23474;
  assign n23476 = ~n23471 & ~n23475;
  assign n23477 = n23469 & n23476;
  assign n23478 = ~pi0868 & n23376;
  assign n23479 = pi2384 & ~n13538;
  assign n23480 = pi0868 & n23479;
  assign n23481 = ~n23478 & ~n23480;
  assign n23482 = pi1472 & ~n23481;
  assign n23483 = n20734 & ~n23482;
  assign n23484 = pi0108 & ~n20528;
  assign n23485 = ~pi0108 & ~n20532;
  assign n23486 = ~n23484 & ~n23485;
  assign n23487 = ~pi0107 & n20543;
  assign n23488 = pi0107 & n20539;
  assign n23489 = ~n23487 & ~n23488;
  assign n23490 = ~n23486 & ~n23489;
  assign n23491 = ~n20734 & n23482;
  assign n23492 = n23490 & ~n23491;
  assign n23493 = ~n23483 & ~n23492;
  assign n23494 = ~n23380 & ~n23388;
  assign n23495 = n23387 & ~n23494;
  assign n23496 = n20747 & ~n23379;
  assign n23497 = ~n20747 & n23379;
  assign n23498 = ~n23496 & ~n23497;
  assign n23499 = ~n23387 & ~n23498;
  assign n23500 = ~n23495 & ~n23499;
  assign n23501 = ~n23493 & ~n23500;
  assign n23502 = ~n23477 & ~n23501;
  assign n23503 = n23444 & ~n23502;
  assign n23504 = n23390 & n23397;
  assign n23505 = ~n23437 & ~n23504;
  assign n23506 = ~n23444 & n23505;
  assign n23507 = ~n23503 & ~n23506;
  assign n23508 = ~n23436 & ~n23507;
  assign n23509 = n23327 & ~n23508;
  assign n23510 = n23433 & ~n23509;
  assign n23511 = n23134 & n23329;
  assign n23512 = ~n23425 & ~n23511;
  assign n23513 = ~n23433 & n23512;
  assign n23514 = ~n23510 & ~n23513;
  assign n23515 = ~n23424 & n23514;
  assign n23516 = ~n23422 & ~n23515;
  assign n23517 = ~n23310 & ~n23516;
  assign n23518 = n23422 & n23514;
  assign n23519 = ~n23424 & n23518;
  assign n23520 = ~n23517 & ~n23519;
  assign n23521 = ~n23444 & n23502;
  assign n23522 = ~n23503 & ~n23521;
  assign n23523 = ~n23469 & ~n23476;
  assign n23524 = ~n23477 & ~n23523;
  assign n23525 = n23493 & ~n23500;
  assign n23526 = ~n23493 & n23500;
  assign n23527 = ~n23525 & ~n23526;
  assign n23528 = ~n23524 & n23527;
  assign n23529 = n23524 & ~n23527;
  assign n23530 = ~n23528 & ~n23529;
  assign n23531 = ~pi0114 & ~n20630;
  assign n23532 = pi0114 & n20626;
  assign n23533 = ~n23531 & ~n23532;
  assign n23534 = ~pi0067 & n20617;
  assign n23535 = pi0067 & n20613;
  assign n23536 = ~n23534 & ~n23535;
  assign n23537 = ~n23533 & ~n23536;
  assign n23538 = ~pi0079 & ~n20571;
  assign n23539 = pi0079 & ~n20567;
  assign n23540 = pi0080 & ~n20553;
  assign n23541 = ~n23539 & ~n23540;
  assign n23542 = ~pi0080 & n20557;
  assign n23543 = n23541 & ~n23542;
  assign n23544 = ~n23538 & n23543;
  assign n23545 = ~n23537 & ~n23544;
  assign n23546 = ~pi0106 & ~n20599;
  assign n23547 = pi0106 & ~n20595;
  assign n23548 = pi0056 & ~n20581;
  assign n23549 = ~n23547 & ~n23548;
  assign n23550 = ~pi0056 & n20585;
  assign n23551 = n23549 & ~n23550;
  assign n23552 = ~n23546 & n23551;
  assign n23553 = n23537 & n23544;
  assign n23554 = ~n23552 & ~n23553;
  assign n23555 = ~n23545 & ~n23554;
  assign n23556 = ~n23459 & ~n23467;
  assign n23557 = ~n23466 & ~n23556;
  assign n23558 = n23451 & ~n23458;
  assign n23559 = ~n23451 & n23458;
  assign n23560 = ~n23558 & ~n23559;
  assign n23561 = n23466 & ~n23560;
  assign n23562 = ~n23557 & ~n23561;
  assign n23563 = n23555 & n23562;
  assign n23564 = ~n23483 & ~n23491;
  assign n23565 = n23490 & ~n23564;
  assign n23566 = ~n20734 & ~n23482;
  assign n23567 = n20734 & n23482;
  assign n23568 = ~n23566 & ~n23567;
  assign n23569 = ~n23490 & ~n23568;
  assign n23570 = ~n23565 & ~n23569;
  assign n23571 = ~pi0868 & n23479;
  assign n23572 = pi2384 & ~n12944;
  assign n23573 = pi0868 & n23572;
  assign n23574 = ~n23571 & ~n23573;
  assign n23575 = pi1472 & ~n23574;
  assign n23576 = ~n20630 & ~n23575;
  assign n23577 = ~pi0078 & ~n20532;
  assign n23578 = pi0078 & ~n20528;
  assign n23579 = ~n23577 & ~n23578;
  assign n23580 = ~pi0108 & n20543;
  assign n23581 = pi0108 & n20539;
  assign n23582 = ~n23580 & ~n23581;
  assign n23583 = ~n23579 & ~n23582;
  assign n23584 = n20630 & n23575;
  assign n23585 = n23583 & ~n23584;
  assign n23586 = ~n23576 & ~n23585;
  assign n23587 = ~n23570 & ~n23586;
  assign n23588 = ~n23563 & ~n23587;
  assign n23589 = n23530 & ~n23588;
  assign n23590 = n23493 & n23500;
  assign n23591 = ~n23523 & ~n23590;
  assign n23592 = ~n23530 & n23591;
  assign n23593 = ~n23589 & ~n23592;
  assign n23594 = ~n23522 & ~n23593;
  assign n23595 = n23522 & n23593;
  assign n23596 = ~n23594 & ~n23595;
  assign n23597 = n23317 & n23320;
  assign n23598 = ~n23321 & ~n23597;
  assign n23599 = ~n23596 & n23598;
  assign n23600 = n23596 & ~n23598;
  assign n23601 = ~n23599 & ~n23600;
  assign n23602 = ~n23522 & n23593;
  assign n23603 = ~n23601 & ~n23602;
  assign n23604 = ~pi0067 & ~n20734;
  assign n23605 = pi0067 & ~n20730;
  assign n23606 = pi0114 & ~n20743;
  assign n23607 = ~n23605 & ~n23606;
  assign n23608 = ~pi0114 & n20747;
  assign n23609 = n23607 & ~n23608;
  assign n23610 = ~n23604 & n23609;
  assign n23611 = ~n23530 & n23588;
  assign n23612 = ~n23589 & ~n23611;
  assign n23613 = pi0114 & ~n20613;
  assign n23614 = ~pi0114 & ~n20617;
  assign n23615 = ~n23613 & ~n23614;
  assign n23616 = ~pi0080 & ~n20571;
  assign n23617 = pi0080 & ~n20567;
  assign n23618 = pi0106 & ~n20553;
  assign n23619 = ~n23617 & ~n23618;
  assign n23620 = ~pi0106 & n20557;
  assign n23621 = n23619 & ~n23620;
  assign n23622 = ~n23616 & n23621;
  assign n23623 = ~n23615 & ~n23622;
  assign n23624 = ~pi0056 & ~n20599;
  assign n23625 = pi0056 & ~n20595;
  assign n23626 = pi0067 & ~n20581;
  assign n23627 = ~n23625 & ~n23626;
  assign n23628 = ~pi0067 & n20585;
  assign n23629 = n23627 & ~n23628;
  assign n23630 = ~n23624 & n23629;
  assign n23631 = n23615 & n23622;
  assign n23632 = ~n23630 & ~n23631;
  assign n23633 = ~n23623 & ~n23632;
  assign n23634 = ~n23545 & ~n23553;
  assign n23635 = ~n23552 & ~n23634;
  assign n23636 = n23537 & ~n23544;
  assign n23637 = ~n23537 & n23544;
  assign n23638 = ~n23636 & ~n23637;
  assign n23639 = n23552 & ~n23638;
  assign n23640 = ~n23635 & ~n23639;
  assign n23641 = n23633 & n23640;
  assign n23642 = ~n23576 & ~n23584;
  assign n23643 = n23583 & ~n23642;
  assign n23644 = n20630 & ~n23575;
  assign n23645 = ~n20630 & n23575;
  assign n23646 = ~n23644 & ~n23645;
  assign n23647 = ~n23583 & ~n23646;
  assign n23648 = ~n23643 & ~n23647;
  assign n23649 = ~pi0868 & n23572;
  assign n23650 = pi2384 & ~n13208;
  assign n23651 = pi0868 & n23650;
  assign n23652 = ~n23649 & ~n23651;
  assign n23653 = pi1472 & ~n23652;
  assign n23654 = n20617 & ~n23653;
  assign n23655 = ~pi0079 & ~n20532;
  assign n23656 = pi0079 & ~n20528;
  assign n23657 = ~n23655 & ~n23656;
  assign n23658 = ~pi0078 & n20543;
  assign n23659 = pi0078 & n20539;
  assign n23660 = ~n23658 & ~n23659;
  assign n23661 = ~n23657 & ~n23660;
  assign n23662 = ~n20617 & n23653;
  assign n23663 = n23661 & ~n23662;
  assign n23664 = ~n23654 & ~n23663;
  assign n23665 = ~n23648 & ~n23664;
  assign n23666 = ~n23641 & ~n23665;
  assign n23667 = ~n23555 & ~n23562;
  assign n23668 = ~n23563 & ~n23667;
  assign n23669 = ~n23570 & n23586;
  assign n23670 = n23570 & ~n23586;
  assign n23671 = ~n23669 & ~n23670;
  assign n23672 = ~n23668 & n23671;
  assign n23673 = n23668 & ~n23671;
  assign n23674 = ~n23672 & ~n23673;
  assign n23675 = ~n23666 & n23674;
  assign n23676 = n23570 & n23586;
  assign n23677 = ~n23667 & ~n23676;
  assign n23678 = ~n23674 & n23677;
  assign n23679 = ~n23675 & ~n23678;
  assign n23680 = n23612 & ~n23679;
  assign n23681 = ~n23610 & ~n23680;
  assign n23682 = n23601 & ~n23681;
  assign n23683 = ~n23603 & ~n23682;
  assign n23684 = n23522 & ~n23593;
  assign n23685 = n23598 & ~n23684;
  assign n23686 = n23436 & n23507;
  assign n23687 = ~n23508 & ~n23686;
  assign n23688 = n23327 & ~n23687;
  assign n23689 = ~n23327 & n23687;
  assign n23690 = ~n23688 & ~n23689;
  assign n23691 = ~n23685 & n23690;
  assign n23692 = n23685 & ~n23690;
  assign n23693 = ~n23691 & ~n23692;
  assign n23694 = ~n23683 & ~n23693;
  assign n23695 = ~n23686 & n23690;
  assign n23696 = ~n23685 & ~n23690;
  assign n23697 = ~n23695 & ~n23696;
  assign n23698 = ~n23433 & n23509;
  assign n23699 = ~n23510 & ~n23698;
  assign n23700 = ~n23697 & n23699;
  assign n23701 = ~n23694 & ~n23700;
  assign n23702 = ~n23310 & ~n23424;
  assign n23703 = ~n23310 & n23514;
  assign n23704 = n23422 & ~n23424;
  assign n23705 = ~n23703 & ~n23704;
  assign n23706 = ~n23702 & n23705;
  assign n23707 = ~n23518 & n23706;
  assign n23708 = ~n23612 & ~n23679;
  assign n23709 = n23612 & n23679;
  assign n23710 = ~n23708 & ~n23709;
  assign n23711 = n23610 & ~n23710;
  assign n23712 = ~n23610 & n23710;
  assign n23713 = ~n23711 & ~n23712;
  assign n23714 = ~n23612 & n23679;
  assign n23715 = n23713 & ~n23714;
  assign n23716 = ~pi0114 & ~n20734;
  assign n23717 = pi0114 & ~n20730;
  assign n23718 = ~n23716 & ~n23717;
  assign n23719 = n23666 & ~n23674;
  assign n23720 = ~n23675 & ~n23719;
  assign n23721 = ~n23633 & n23640;
  assign n23722 = n23633 & ~n23640;
  assign n23723 = ~n23721 & ~n23722;
  assign n23724 = ~n23648 & n23664;
  assign n23725 = n23648 & ~n23664;
  assign n23726 = ~n23724 & ~n23725;
  assign n23727 = ~n23723 & n23726;
  assign n23728 = n23723 & ~n23726;
  assign n23729 = ~n23727 & ~n23728;
  assign n23730 = ~pi0868 & n23650;
  assign n23731 = pi2384 & ~n13843;
  assign n23732 = pi0868 & n23731;
  assign n23733 = ~n23730 & ~n23732;
  assign n23734 = pi1472 & ~n23733;
  assign n23735 = ~n20585 & ~n23734;
  assign n23736 = pi0080 & ~n20528;
  assign n23737 = ~pi0080 & ~n20532;
  assign n23738 = ~n23736 & ~n23737;
  assign n23739 = ~pi0079 & n20543;
  assign n23740 = pi0079 & n20539;
  assign n23741 = ~n23739 & ~n23740;
  assign n23742 = ~n23738 & ~n23741;
  assign n23743 = n20585 & n23734;
  assign n23744 = n23742 & ~n23743;
  assign n23745 = ~n23735 & ~n23744;
  assign n23746 = ~n23654 & ~n23662;
  assign n23747 = n23661 & ~n23746;
  assign n23748 = n20617 & n23653;
  assign n23749 = ~n20617 & ~n23653;
  assign n23750 = ~n23748 & ~n23749;
  assign n23751 = ~n23661 & ~n23750;
  assign n23752 = ~n23747 & ~n23751;
  assign n23753 = ~n23745 & ~n23752;
  assign n23754 = ~n23623 & ~n23631;
  assign n23755 = ~n23630 & ~n23754;
  assign n23756 = n23615 & ~n23622;
  assign n23757 = ~n23615 & n23622;
  assign n23758 = ~n23756 & ~n23757;
  assign n23759 = n23630 & ~n23758;
  assign n23760 = ~n23755 & ~n23759;
  assign n23761 = ~pi0067 & ~n20599;
  assign n23762 = pi0067 & ~n20595;
  assign n23763 = pi0114 & ~n20581;
  assign n23764 = ~n23762 & ~n23763;
  assign n23765 = ~pi0114 & n20585;
  assign n23766 = n23764 & ~n23765;
  assign n23767 = ~n23761 & n23766;
  assign n23768 = ~pi0106 & ~n20571;
  assign n23769 = pi0106 & ~n20567;
  assign n23770 = pi0056 & ~n20553;
  assign n23771 = ~n23769 & ~n23770;
  assign n23772 = ~pi0056 & n20557;
  assign n23773 = n23771 & ~n23772;
  assign n23774 = ~n23768 & n23773;
  assign n23775 = ~n23767 & ~n23774;
  assign n23776 = n23760 & ~n23775;
  assign n23777 = ~n23753 & ~n23776;
  assign n23778 = ~n23729 & ~n23777;
  assign n23779 = n23648 & n23664;
  assign n23780 = ~n23633 & ~n23640;
  assign n23781 = ~n23779 & ~n23780;
  assign n23782 = n23729 & n23781;
  assign n23783 = ~n23778 & ~n23782;
  assign n23784 = n23720 & ~n23783;
  assign n23785 = ~n23718 & ~n23784;
  assign n23786 = ~n23713 & ~n23785;
  assign n23787 = ~n23715 & ~n23786;
  assign n23788 = ~n23601 & n23681;
  assign n23789 = ~n23682 & ~n23788;
  assign n23790 = n23787 & ~n23789;
  assign n23791 = n23713 & ~n23785;
  assign n23792 = ~n23713 & n23785;
  assign n23793 = ~n23791 & ~n23792;
  assign n23794 = ~n23720 & ~n23783;
  assign n23795 = n23720 & n23783;
  assign n23796 = ~n23794 & ~n23795;
  assign n23797 = ~n23718 & ~n23796;
  assign n23798 = n23718 & n23796;
  assign n23799 = ~n23797 & ~n23798;
  assign n23800 = ~n23720 & ~n23799;
  assign n23801 = n23783 & n23800;
  assign n23802 = ~n23793 & ~n23801;
  assign n23803 = ~n23787 & n23789;
  assign n23804 = ~n23802 & ~n23803;
  assign n23805 = ~n23760 & n23775;
  assign n23806 = ~n23776 & ~n23805;
  assign n23807 = n23745 & ~n23752;
  assign n23808 = ~n23745 & n23752;
  assign n23809 = ~n23807 & ~n23808;
  assign n23810 = ~n23806 & n23809;
  assign n23811 = n23806 & ~n23809;
  assign n23812 = ~n23810 & ~n23811;
  assign n23813 = ~pi0868 & n23731;
  assign n23814 = pi2384 & ~n12274;
  assign n23815 = pi0868 & n23814;
  assign n23816 = ~n23813 & ~n23815;
  assign n23817 = pi1472 & ~n23816;
  assign n23818 = n20599 & ~n23817;
  assign n23819 = ~pi0106 & ~n20532;
  assign n23820 = pi0106 & ~n20528;
  assign n23821 = ~n23819 & ~n23820;
  assign n23822 = ~pi0080 & n20543;
  assign n23823 = pi0080 & n20539;
  assign n23824 = ~n23822 & ~n23823;
  assign n23825 = ~n23821 & ~n23824;
  assign n23826 = ~n23818 & ~n23825;
  assign n23827 = ~n20599 & n23817;
  assign n23828 = ~n23826 & ~n23827;
  assign n23829 = ~n23735 & ~n23743;
  assign n23830 = n23742 & ~n23829;
  assign n23831 = n20585 & ~n23734;
  assign n23832 = ~n20585 & n23734;
  assign n23833 = ~n23831 & ~n23832;
  assign n23834 = ~n23742 & ~n23833;
  assign n23835 = ~n23830 & ~n23834;
  assign n23836 = n23828 & ~n23835;
  assign n23837 = n23767 & ~n23774;
  assign n23838 = ~n23767 & n23774;
  assign n23839 = ~n23837 & ~n23838;
  assign n23840 = ~pi0056 & ~n20571;
  assign n23841 = pi0056 & ~n20567;
  assign n23842 = pi0067 & ~n20553;
  assign n23843 = ~n23841 & ~n23842;
  assign n23844 = ~pi0067 & n20557;
  assign n23845 = n23843 & ~n23844;
  assign n23846 = ~n23840 & n23845;
  assign n23847 = ~pi0114 & ~n20599;
  assign n23848 = pi0114 & ~n20595;
  assign n23849 = ~n23847 & ~n23848;
  assign n23850 = ~n23846 & ~n23849;
  assign n23851 = n23839 & ~n23850;
  assign n23852 = ~n23836 & ~n23851;
  assign n23853 = n23812 & ~n23852;
  assign n23854 = n23745 & n23752;
  assign n23855 = ~n23805 & ~n23854;
  assign n23856 = ~n23812 & n23855;
  assign n23857 = ~n23853 & ~n23856;
  assign n23858 = n23729 & n23777;
  assign n23859 = ~n23778 & ~n23858;
  assign n23860 = ~n23857 & ~n23859;
  assign n23861 = n23857 & n23859;
  assign n23862 = ~n23860 & ~n23861;
  assign n23863 = ~n23859 & n23862;
  assign n23864 = n23857 & n23863;
  assign n23865 = ~n23799 & ~n23864;
  assign n23866 = ~n23828 & ~n23835;
  assign n23867 = n23828 & n23835;
  assign n23868 = ~n23866 & ~n23867;
  assign n23869 = ~n23839 & ~n23850;
  assign n23870 = n23839 & n23850;
  assign n23871 = ~n23869 & ~n23870;
  assign n23872 = ~n23868 & n23871;
  assign n23873 = n23868 & ~n23871;
  assign n23874 = ~n23872 & ~n23873;
  assign n23875 = n23846 & n23849;
  assign n23876 = ~n23850 & ~n23875;
  assign n23877 = ~pi0868 & n23814;
  assign n23878 = pi2384 & ~n14680;
  assign n23879 = pi0868 & n23878;
  assign n23880 = ~n23877 & ~n23879;
  assign n23881 = pi1472 & ~n23880;
  assign n23882 = ~n20557 & ~n23881;
  assign n23883 = pi0056 & ~n20528;
  assign n23884 = ~pi0056 & ~n20532;
  assign n23885 = ~n23883 & ~n23884;
  assign n23886 = ~pi0106 & n20543;
  assign n23887 = pi0106 & n20539;
  assign n23888 = ~n23886 & ~n23887;
  assign n23889 = ~n23885 & ~n23888;
  assign n23890 = n20557 & n23881;
  assign n23891 = n23889 & ~n23890;
  assign n23892 = ~n23882 & ~n23891;
  assign n23893 = ~n23818 & ~n23827;
  assign n23894 = n23825 & n23893;
  assign n23895 = ~n23825 & ~n23893;
  assign n23896 = ~n23894 & ~n23895;
  assign n23897 = ~n23892 & n23896;
  assign n23898 = n23876 & ~n23897;
  assign n23899 = ~n23874 & ~n23898;
  assign n23900 = ~n23839 & n23850;
  assign n23901 = ~n23828 & n23835;
  assign n23902 = ~n23900 & ~n23901;
  assign n23903 = n23874 & n23902;
  assign n23904 = ~n23899 & ~n23903;
  assign n23905 = ~n23812 & n23852;
  assign n23906 = ~n23853 & ~n23905;
  assign n23907 = ~n23904 & ~n23906;
  assign n23908 = n23904 & n23906;
  assign n23909 = ~n23907 & ~n23908;
  assign n23910 = ~n23906 & n23909;
  assign n23911 = n23904 & n23910;
  assign n23912 = ~n23862 & n23911;
  assign n23913 = ~n23865 & n23912;
  assign n23914 = n23799 & n23864;
  assign n23915 = ~n23913 & ~n23914;
  assign n23916 = n23804 & ~n23915;
  assign n23917 = ~n23790 & ~n23916;
  assign n23918 = n23793 & n23801;
  assign n23919 = ~n23803 & n23918;
  assign n23920 = n23917 & ~n23919;
  assign n23921 = ~n23707 & ~n23920;
  assign n23922 = n23701 & n23921;
  assign n23923 = n23862 & ~n23911;
  assign n23924 = ~n23865 & ~n23923;
  assign n23925 = ~pi0868 & n23878;
  assign n23926 = pi2384 & ~n14917;
  assign n23927 = pi0868 & n23926;
  assign n23928 = ~n23925 & ~n23927;
  assign n23929 = pi1472 & ~n23928;
  assign n23930 = n20571 & ~n23929;
  assign n23931 = ~pi0067 & ~n20532;
  assign n23932 = pi0067 & ~n20528;
  assign n23933 = ~n23931 & ~n23932;
  assign n23934 = ~pi0056 & n20543;
  assign n23935 = pi0056 & n20539;
  assign n23936 = ~n23934 & ~n23935;
  assign n23937 = ~n23933 & ~n23936;
  assign n23938 = ~n20571 & n23929;
  assign n23939 = n23937 & ~n23938;
  assign n23940 = ~n23930 & ~n23939;
  assign n23941 = ~n23882 & ~n23890;
  assign n23942 = n23889 & ~n23941;
  assign n23943 = n20557 & ~n23881;
  assign n23944 = ~n20557 & n23881;
  assign n23945 = ~n23943 & ~n23944;
  assign n23946 = ~n23889 & ~n23945;
  assign n23947 = ~n23942 & ~n23946;
  assign n23948 = n23940 & n23947;
  assign n23949 = n23940 & ~n23947;
  assign n23950 = ~n23940 & n23947;
  assign n23951 = ~n23949 & ~n23950;
  assign n23952 = ~pi0067 & ~n20571;
  assign n23953 = pi0067 & ~n20567;
  assign n23954 = pi0114 & ~n20553;
  assign n23955 = ~n23953 & ~n23954;
  assign n23956 = ~pi0114 & n20557;
  assign n23957 = n23955 & ~n23956;
  assign n23958 = ~n23952 & n23957;
  assign n23959 = ~n23951 & n23958;
  assign n23960 = n23951 & ~n23958;
  assign n23961 = ~n23959 & ~n23960;
  assign n23962 = n23948 & n23961;
  assign n23963 = ~pi0114 & ~n20571;
  assign n23964 = pi0114 & ~n20567;
  assign n23965 = ~n23963 & ~n23964;
  assign n23966 = pi2384 & ~n11933;
  assign n23967 = pi0868 & n23966;
  assign n23968 = ~pi0868 & n23926;
  assign n23969 = ~n23967 & ~n23968;
  assign n23970 = pi1472 & ~n23969;
  assign n23971 = n20532 & n23970;
  assign n23972 = ~pi0114 & ~n20532;
  assign n23973 = pi0114 & ~n20528;
  assign n23974 = ~n23972 & ~n23973;
  assign n23975 = ~pi0067 & n20543;
  assign n23976 = pi0067 & n20539;
  assign n23977 = ~n23975 & ~n23976;
  assign n23978 = ~n23974 & ~n23977;
  assign n23979 = ~n20532 & ~n23970;
  assign n23980 = ~n23978 & ~n23979;
  assign n23981 = ~n23971 & ~n23980;
  assign n23982 = ~n23930 & ~n23938;
  assign n23983 = n23937 & ~n23982;
  assign n23984 = ~n20571 & ~n23929;
  assign n23985 = n20571 & n23929;
  assign n23986 = ~n23984 & ~n23985;
  assign n23987 = ~n23937 & ~n23986;
  assign n23988 = ~n23983 & ~n23987;
  assign n23989 = n23981 & ~n23988;
  assign n23990 = ~n23965 & ~n23989;
  assign n23991 = ~n23961 & n23990;
  assign n23992 = ~n23962 & ~n23991;
  assign n23993 = ~n23940 & ~n23947;
  assign n23994 = ~n23958 & ~n23993;
  assign n23995 = n23892 & ~n23896;
  assign n23996 = ~n23897 & ~n23995;
  assign n23997 = n23876 & ~n23996;
  assign n23998 = ~n23876 & n23996;
  assign n23999 = ~n23997 & ~n23998;
  assign n24000 = n23994 & n23999;
  assign n24001 = ~n23994 & ~n23999;
  assign n24002 = ~n24000 & ~n24001;
  assign n24003 = n23992 & n24002;
  assign n24004 = ~n23992 & ~n24002;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = n23981 & n23988;
  assign n24007 = ~n23981 & ~n23988;
  assign n24008 = ~n24006 & ~n24007;
  assign n24009 = ~n23965 & ~n24008;
  assign n24010 = n23965 & n24008;
  assign n24011 = ~n24009 & ~n24010;
  assign n24012 = n23988 & ~n24011;
  assign n24013 = ~n23981 & n24012;
  assign n24014 = n23961 & n23990;
  assign n24015 = ~n23961 & ~n23990;
  assign n24016 = ~n24014 & ~n24015;
  assign n24017 = ~n24013 & n24016;
  assign n24018 = n24013 & ~n24016;
  assign n24019 = ~n24017 & ~n24018;
  assign n24020 = pi0868 & pi2384;
  assign n24021 = ~n10970 & n24020;
  assign n24022 = ~pi0868 & n23966;
  assign n24023 = ~n24021 & ~n24022;
  assign n24024 = pi1472 & ~n24023;
  assign n24025 = n20543 & ~n24024;
  assign n24026 = ~pi0114 & n20543;
  assign n24027 = pi0114 & n20539;
  assign n24028 = ~n24026 & ~n24027;
  assign n24029 = ~n20543 & n24024;
  assign n24030 = ~n24028 & ~n24029;
  assign n24031 = ~n24025 & ~n24030;
  assign n24032 = ~n23971 & ~n23979;
  assign n24033 = ~n23978 & ~n24032;
  assign n24034 = ~n20532 & n23970;
  assign n24035 = n20532 & ~n23970;
  assign n24036 = ~n24034 & ~n24035;
  assign n24037 = n23978 & ~n24036;
  assign n24038 = ~n24033 & ~n24037;
  assign n24039 = n24031 & ~n24038;
  assign n24040 = ~n24031 & n24038;
  assign n24041 = ~n24039 & ~n24040;
  assign n24042 = ~n24038 & ~n24041;
  assign n24043 = n24031 & n24042;
  assign n24044 = n24011 & n24043;
  assign n24045 = ~n24011 & ~n24043;
  assign n24046 = ~n24044 & ~n24045;
  assign n24047 = n24011 & ~n24046;
  assign n24048 = n24043 & n24047;
  assign n24049 = n24019 & n24048;
  assign n24050 = ~n24005 & ~n24049;
  assign n24051 = n24013 & ~n24019;
  assign n24052 = ~n24016 & n24051;
  assign n24053 = n24005 & n24049;
  assign n24054 = ~n24052 & ~n24053;
  assign n24055 = ~n24050 & ~n24054;
  assign n24056 = ~n23992 & ~n24005;
  assign n24057 = ~n24002 & n24056;
  assign n24058 = n23874 & n23898;
  assign n24059 = ~n23899 & ~n24058;
  assign n24060 = ~n23995 & n23999;
  assign n24061 = ~n24001 & ~n24060;
  assign n24062 = n24059 & ~n24061;
  assign n24063 = ~n24059 & n24061;
  assign n24064 = ~n24062 & ~n24063;
  assign n24065 = n24061 & ~n24064;
  assign n24066 = ~n24059 & n24065;
  assign n24067 = n24057 & n24066;
  assign n24068 = n24064 & n24066;
  assign n24069 = ~n24067 & ~n24068;
  assign n24070 = ~n24057 & ~n24064;
  assign n24071 = ~n23909 & ~n24070;
  assign n24072 = n24069 & ~n24071;
  assign n24073 = n24055 & ~n24072;
  assign n24074 = ~n23909 & n24066;
  assign n24075 = ~n24073 & ~n24074;
  assign n24076 = ~n23909 & n24057;
  assign n24077 = ~n24067 & ~n24076;
  assign n24078 = n24064 & ~n24077;
  assign n24079 = n24075 & ~n24078;
  assign n24080 = n23924 & ~n24079;
  assign n24081 = ~n23707 & n24080;
  assign n24082 = n23701 & n24081;
  assign n24083 = n23804 & n24082;
  assign n24084 = n23683 & n23693;
  assign n24085 = ~n23700 & n24084;
  assign n24086 = n23697 & ~n23699;
  assign n24087 = ~n24085 & ~n24086;
  assign n24088 = ~n23707 & ~n24087;
  assign n24089 = ~n24083 & ~n24088;
  assign n24090 = ~n23922 & n24089;
  assign n24091 = n23520 & n24090;
  assign n24092 = n23251 & ~n23275;
  assign n24093 = n23249 & ~n24092;
  assign n24094 = ~n23271 & ~n24093;
  assign n24095 = ~n23276 & n24094;
  assign n24096 = n23021 & ~n24095;
  assign n24097 = n22763 & n24096;
  assign n24098 = ~n24091 & n24097;
  assign n24099 = n23308 & ~n24098;
  assign n24100 = n21536 & ~n21542;
  assign n24101 = n21519 & ~n24100;
  assign n24102 = ~n21537 & ~n24101;
  assign n24103 = ~n21543 & n24102;
  assign n24104 = ~n21332 & ~n24103;
  assign n24105 = ~n24099 & n24104;
  assign n24106 = n21554 & ~n24105;
  assign n24107 = n21059 & ~n21141;
  assign n24108 = ~n24106 & ~n24107;
  assign n24109 = ~n21142 & ~n24108;
  assign n24110 = ~n20942 & n21056;
  assign n24111 = ~n20851 & n20898;
  assign n24112 = n24110 & ~n24111;
  assign n24113 = ~n21058 & ~n24112;
  assign n24114 = ~n21059 & n24113;
  assign n24115 = n20900 & n20940;
  assign n24116 = ~n20941 & ~n24115;
  assign n24117 = ~n21059 & ~n24116;
  assign n24118 = ~n24113 & n24116;
  assign n24119 = n21141 & ~n24118;
  assign n24120 = ~n24117 & ~n24119;
  assign n24121 = ~n24114 & n24120;
  assign n24122 = ~n24109 & ~n24121;
  assign n24123 = ~n24114 & ~n24117;
  assign n24124 = n21141 & ~n24123;
  assign n24125 = n24113 & ~n24116;
  assign n24126 = ~n24124 & ~n24125;
  assign n24127 = ~n24122 & n24126;
  assign n24128 = ~n20946 & n20986;
  assign n24129 = ~n24127 & ~n24128;
  assign n24130 = ~n20987 & ~n24129;
  assign n24131 = ~n20956 & ~n20977;
  assign n24132 = n20655 & ~n24131;
  assign n24133 = n20652 & n20977;
  assign n24134 = ~n24132 & ~n24133;
  assign n24135 = n20652 & n20956;
  assign n24136 = n24134 & ~n24135;
  assign n24137 = ~n20966 & n20968;
  assign n24138 = ~n20817 & ~n24137;
  assign n24139 = pi2384 & ~n14685;
  assign n24140 = ~pi0868 & n24139;
  assign n24141 = pi0868 & n20959;
  assign n24142 = ~n24140 & ~n24141;
  assign n24143 = pi1472 & ~n24142;
  assign n24144 = n20917 & n24143;
  assign n24145 = ~n20917 & ~n24143;
  assign n24146 = ~n24144 & ~n24145;
  assign n24147 = ~n20916 & n20963;
  assign n24148 = ~n20915 & ~n24147;
  assign n24149 = ~n24146 & ~n24148;
  assign n24150 = n24146 & n24148;
  assign n24151 = ~n24149 & ~n24150;
  assign n24152 = n20820 & ~n24151;
  assign n24153 = ~n20820 & n24151;
  assign n24154 = ~n24152 & ~n24153;
  assign n24155 = n24138 & n24154;
  assign n24156 = ~n24138 & ~n24154;
  assign n24157 = ~n24155 & ~n24156;
  assign n24158 = n20966 & ~n20968;
  assign n24159 = ~n20974 & ~n24158;
  assign n24160 = ~n20819 & n24159;
  assign n24161 = ~n20958 & n20974;
  assign n24162 = ~n24160 & ~n24161;
  assign n24163 = ~n24157 & n24162;
  assign n24164 = n24157 & ~n24162;
  assign n24165 = ~n24163 & ~n24164;
  assign n24166 = n20903 & ~n24165;
  assign n24167 = ~n20903 & n24165;
  assign n24168 = ~n24166 & ~n24167;
  assign n24169 = ~n24136 & n24168;
  assign n24170 = n24136 & ~n24168;
  assign n24171 = ~n24169 & ~n24170;
  assign n24172 = ~n20942 & n20983;
  assign n24173 = n20956 & n20977;
  assign n24174 = n24172 & ~n24173;
  assign n24175 = ~n20985 & ~n24174;
  assign n24176 = ~n24171 & ~n24175;
  assign n24177 = n24171 & n24175;
  assign n24178 = ~n24176 & ~n24177;
  assign n24179 = n24130 & n24178;
  assign n24180 = ~n24130 & ~n24178;
  assign n24181 = ~n24179 & ~n24180;
  assign n24182 = ~pi0868 & n24181;
  assign n24183 = ~n20942 & n24168;
  assign n24184 = n24157 & n24162;
  assign n24185 = n24183 & ~n24184;
  assign n24186 = ~n24170 & ~n24185;
  assign n24187 = n24146 & ~n24148;
  assign n24188 = ~n24154 & ~n24187;
  assign n24189 = ~n20819 & n24188;
  assign n24190 = ~n24138 & n24154;
  assign n24191 = ~n24189 & ~n24190;
  assign n24192 = ~n24146 & n24148;
  assign n24193 = ~n20817 & ~n24192;
  assign n24194 = pi2384 & ~n12257;
  assign n24195 = ~pi0868 & n24194;
  assign n24196 = pi0868 & n24139;
  assign n24197 = ~n24195 & ~n24196;
  assign n24198 = pi1472 & ~n24197;
  assign n24199 = n20917 & n24198;
  assign n24200 = ~n20917 & ~n24198;
  assign n24201 = ~n24199 & ~n24200;
  assign n24202 = ~n20916 & n24143;
  assign n24203 = ~n20915 & ~n24202;
  assign n24204 = ~n24201 & ~n24203;
  assign n24205 = n24201 & n24203;
  assign n24206 = ~n24204 & ~n24205;
  assign n24207 = n20820 & ~n24206;
  assign n24208 = ~n20820 & n24206;
  assign n24209 = ~n24207 & ~n24208;
  assign n24210 = n24193 & n24209;
  assign n24211 = ~n24193 & ~n24209;
  assign n24212 = ~n24210 & ~n24211;
  assign n24213 = ~n24191 & n24212;
  assign n24214 = n24191 & ~n24212;
  assign n24215 = ~n24213 & ~n24214;
  assign n24216 = n20903 & ~n24215;
  assign n24217 = ~n20903 & n24215;
  assign n24218 = ~n24216 & ~n24217;
  assign n24219 = ~n24157 & ~n24162;
  assign n24220 = ~n20656 & ~n24219;
  assign n24221 = n24218 & ~n24220;
  assign n24222 = ~n24218 & n24220;
  assign n24223 = ~n24221 & ~n24222;
  assign n24224 = ~n24186 & n24223;
  assign n24225 = n24186 & ~n24223;
  assign n24226 = ~n24224 & ~n24225;
  assign n24227 = n24171 & ~n24175;
  assign n24228 = ~n24128 & ~n24227;
  assign n24229 = ~n24121 & n24228;
  assign n24230 = ~n21554 & n24229;
  assign n24231 = ~n24126 & n24228;
  assign n24232 = ~n24171 & n24175;
  assign n24233 = ~n24231 & ~n24232;
  assign n24234 = n20987 & ~n24227;
  assign n24235 = n24233 & ~n24234;
  assign n24236 = n24104 & n24229;
  assign n24237 = ~n23308 & n24236;
  assign n24238 = n24235 & ~n24237;
  assign n24239 = ~n24091 & n24229;
  assign n24240 = n24097 & n24239;
  assign n24241 = n24104 & n24240;
  assign n24242 = n24238 & ~n24241;
  assign n24243 = ~n24230 & n24242;
  assign n24244 = ~n24226 & n24243;
  assign n24245 = n24226 & ~n24243;
  assign n24246 = ~n24244 & ~n24245;
  assign n24247 = pi0868 & ~n24246;
  assign n24248 = ~n24182 & ~n24247;
  assign n24249 = n20524 & ~n24248;
  assign n24250 = ~n20526 & ~n24249;
  assign n24251 = pi0979 & ~n9352;
  assign n24252 = n20519 & n24251;
  assign n24253 = pi0039 & ~n24252;
  assign n24254 = ~pi3245 & ~n14816;
  assign n24255 = pi3245 & ~n16640;
  assign n24256 = ~n24254 & ~n24255;
  assign n24257 = n24252 & ~n24256;
  assign n24258 = ~n24253 & ~n24257;
  assign n24259 = n20513 & n24251;
  assign n24260 = n20515 & n24251;
  assign n24261 = ~n24259 & ~n24260;
  assign n24262 = ~n24258 & n24261;
  assign n24263 = ~pi3245 & ~n17368;
  assign n24264 = pi3245 & ~n17397;
  assign n24265 = ~n24263 & ~n24264;
  assign n24266 = n24259 & ~n24265;
  assign n24267 = ~n24260 & n24266;
  assign n24268 = ~n24262 & ~n24267;
  assign n24269 = ~n20521 & ~n24268;
  assign n24270 = pi0051 & n24260;
  assign n24271 = ~n20521 & n24270;
  assign n24272 = ~n24269 & ~n24271;
  assign n24273 = ~n20524 & ~n24272;
  assign po0309 = ~n24250 | n24273;
  assign n24275 = pi0040 & ~n20524;
  assign n24276 = n20521 & n24275;
  assign n24277 = ~n20987 & ~n24128;
  assign n24278 = n24127 & ~n24277;
  assign n24279 = ~n24127 & n24277;
  assign n24280 = ~n24278 & ~n24279;
  assign n24281 = ~pi0868 & n24280;
  assign n24282 = pi0868 & n24181;
  assign n24283 = ~n24281 & ~n24282;
  assign n24284 = n20524 & ~n24283;
  assign n24285 = ~n24276 & ~n24284;
  assign n24286 = pi0040 & ~n24252;
  assign n24287 = ~pi3245 & ~n15115;
  assign n24288 = pi3245 & ~n16604;
  assign n24289 = ~n24287 & ~n24288;
  assign n24290 = n24252 & ~n24289;
  assign n24291 = ~n24286 & ~n24290;
  assign n24292 = n24261 & ~n24291;
  assign n24293 = ~n24267 & ~n24292;
  assign n24294 = ~n20521 & ~n24293;
  assign n24295 = ~n24271 & ~n24294;
  assign n24296 = ~n20524 & ~n24295;
  assign po0310 = ~n24285 | n24296;
  assign n24298 = ~pi0979 & ~pi1666;
  assign n24299 = ~pi0979 & ~n20516;
  assign n24300 = ~n24298 & ~n24299;
  assign n24301 = ~pi0979 & n20519;
  assign n24302 = n24300 & ~n24301;
  assign n24303 = n20522 & n24298;
  assign n24304 = ~n24302 & n24303;
  assign n24305 = pi0041 & ~n24304;
  assign n24306 = n24302 & n24305;
  assign n24307 = ~n24248 & n24304;
  assign n24308 = ~n24306 & ~n24307;
  assign n24309 = ~pi0979 & ~n9352;
  assign n24310 = n20519 & n24309;
  assign n24311 = pi0041 & ~n24310;
  assign n24312 = ~n24256 & n24310;
  assign n24313 = ~n24311 & ~n24312;
  assign n24314 = n20513 & n24309;
  assign n24315 = n20515 & n24309;
  assign n24316 = ~n24314 & ~n24315;
  assign n24317 = ~n24313 & n24316;
  assign n24318 = ~n24265 & n24314;
  assign n24319 = ~n24315 & n24318;
  assign n24320 = ~n24317 & ~n24319;
  assign n24321 = ~n24302 & ~n24320;
  assign n24322 = pi0053 & n24315;
  assign n24323 = ~n24302 & n24322;
  assign n24324 = ~n24321 & ~n24323;
  assign n24325 = ~n24304 & ~n24324;
  assign po0311 = ~n24308 | n24325;
  assign n24327 = pi0042 & ~n24304;
  assign n24328 = n24302 & n24327;
  assign n24329 = ~n24283 & n24304;
  assign n24330 = ~n24328 & ~n24329;
  assign n24331 = pi0042 & ~n24310;
  assign n24332 = ~n24289 & n24310;
  assign n24333 = ~n24331 & ~n24332;
  assign n24334 = n24316 & ~n24333;
  assign n24335 = ~n24319 & ~n24334;
  assign n24336 = ~n24302 & ~n24335;
  assign n24337 = ~n24323 & ~n24336;
  assign n24338 = ~n24304 & ~n24337;
  assign po0312 = ~n24330 | n24338;
  assign n24340 = pi2384 & n20522;
  assign n24341 = ~n24248 & n24340;
  assign n24342 = pi0043 & ~n24340;
  assign po0313 = n24341 | n24342;
  assign n24344 = ~n24283 & n24340;
  assign n24345 = pi0044 & ~n24340;
  assign po0314 = n24344 | n24345;
  assign n24347 = ~pi0045 & n8561;
  assign n24348 = ~pi2335 & n15594;
  assign n24349 = ~pi2358 & n15592;
  assign n24350 = ~n24348 & ~n24349;
  assign n24351 = ~pi2471 & n15599;
  assign n24352 = ~pi2519 & n15597;
  assign n24353 = ~n24351 & ~n24352;
  assign n24354 = n24350 & n24353;
  assign n24355 = ~pi2328 & n15594;
  assign n24356 = ~pi2353 & n15592;
  assign n24357 = ~n24355 & ~n24356;
  assign n24358 = ~pi2407 & n15599;
  assign n24359 = ~pi2406 & n15597;
  assign n24360 = ~n24358 & ~n24359;
  assign n24361 = n24357 & n24360;
  assign n24362 = ~n24354 & ~n24361;
  assign n24363 = ~pi2364 & n15599;
  assign n24364 = ~pi2340 & n15597;
  assign n24365 = ~n24363 & ~n24364;
  assign n24366 = ~pi2329 & n15594;
  assign n24367 = ~pi2354 & n15592;
  assign n24368 = ~n24366 & ~n24367;
  assign n24369 = n24365 & n24368;
  assign n24370 = ~pi1990 & n15594;
  assign n24371 = ~pi2001 & n15592;
  assign n24372 = ~n24370 & ~n24371;
  assign n24373 = ~pi2362 & n15599;
  assign n24374 = ~pi2338 & n15597;
  assign n24375 = ~n24373 & ~n24374;
  assign n24376 = n24372 & n24375;
  assign n24377 = ~n24369 & n24376;
  assign n24378 = n24362 & n24377;
  assign n24379 = ~n20479 & n24378;
  assign n24380 = n24354 & ~n24361;
  assign n24381 = n24377 & n24380;
  assign n24382 = n20479 & n24381;
  assign n24383 = ~n24379 & ~n24382;
  assign n24384 = ~n20459 & ~n24383;
  assign n24385 = pi0659 & n24378;
  assign n24386 = ~pi0659 & n24381;
  assign n24387 = ~n24385 & ~n24386;
  assign n24388 = n20459 & ~n24387;
  assign n24389 = ~n24384 & ~n24388;
  assign n24390 = ~n24354 & n24361;
  assign n24391 = ~n24369 & ~n24376;
  assign n24392 = n24390 & n24391;
  assign n24393 = pi0152 & n24392;
  assign n24394 = n24354 & n24361;
  assign n24395 = n24391 & n24394;
  assign n24396 = ~pi0152 & n24395;
  assign n24397 = ~n24393 & ~n24396;
  assign n24398 = n24369 & ~n24376;
  assign n24399 = n24390 & n24398;
  assign n24400 = n8640 & n24399;
  assign n24401 = n24394 & n24398;
  assign n24402 = ~n8640 & n24401;
  assign n24403 = ~n24400 & ~n24402;
  assign n24404 = n24397 & n24403;
  assign n24405 = n24369 & n24376;
  assign n24406 = n24362 & n24405;
  assign n24407 = pi0196 & n24406;
  assign n24408 = n24380 & n24405;
  assign n24409 = ~pi0196 & n24408;
  assign n24410 = ~n24407 & ~n24409;
  assign n24411 = n24404 & n24410;
  assign n24412 = n19557 & ~n24411;
  assign n24413 = n24389 & ~n24412;
  assign n24414 = n20445 & n24408;
  assign n24415 = ~n20445 & n24406;
  assign n24416 = ~n24414 & ~n24415;
  assign n24417 = ~n20411 & n24401;
  assign n24418 = n20411 & n24399;
  assign n24419 = ~n24417 & ~n24418;
  assign n24420 = n20370 & n24395;
  assign n24421 = ~n20370 & n24392;
  assign n24422 = ~n24420 & ~n24421;
  assign n24423 = n24419 & n24422;
  assign n24424 = n24416 & n24423;
  assign n24425 = ~n19557 & ~n24424;
  assign n24426 = n24413 & ~n24425;
  assign n24427 = ~n8561 & n24426;
  assign n24428 = ~n24347 & ~n24427;
  assign po0315 = po0493 & n24428;
  assign n24430 = pi0046 & ~n20524;
  assign n24431 = n20521 & n24430;
  assign n24432 = pi0868 & n24280;
  assign n24433 = n24113 & n24116;
  assign n24434 = ~n24113 & ~n24116;
  assign n24435 = ~n24433 & ~n24434;
  assign n24436 = n24109 & n24435;
  assign n24437 = ~n24109 & ~n24435;
  assign n24438 = ~n24436 & ~n24437;
  assign n24439 = ~pi0868 & n24438;
  assign n24440 = ~n24432 & ~n24439;
  assign n24441 = n20524 & ~n24440;
  assign n24442 = ~n24431 & ~n24441;
  assign n24443 = pi0046 & ~n24252;
  assign n24444 = ~pi3245 & ~n12061;
  assign n24445 = pi3245 & ~n16568;
  assign n24446 = ~n24444 & ~n24445;
  assign n24447 = n24252 & ~n24446;
  assign n24448 = ~n24443 & ~n24447;
  assign n24449 = n24261 & ~n24448;
  assign n24450 = ~n24267 & ~n24449;
  assign n24451 = ~n20521 & ~n24450;
  assign n24452 = ~n24271 & ~n24451;
  assign n24453 = ~n20524 & ~n24452;
  assign po0316 = ~n24442 | n24453;
  assign n24455 = pi0047 & ~n24304;
  assign n24456 = n24302 & n24455;
  assign n24457 = n24304 & ~n24440;
  assign n24458 = ~n24456 & ~n24457;
  assign n24459 = pi0047 & ~n24310;
  assign n24460 = n24310 & ~n24446;
  assign n24461 = ~n24459 & ~n24460;
  assign n24462 = n24316 & ~n24461;
  assign n24463 = ~n24319 & ~n24462;
  assign n24464 = ~n24302 & ~n24463;
  assign n24465 = ~n24323 & ~n24464;
  assign n24466 = ~n24304 & ~n24465;
  assign po0317 = ~n24458 | n24466;
  assign n24468 = n24340 & ~n24440;
  assign n24469 = pi0048 & ~n24340;
  assign po0318 = n24468 | n24469;
  assign n24471 = pi0049 & ~n20524;
  assign n24472 = n20521 & n24471;
  assign n24473 = pi0868 & n24438;
  assign n24474 = ~n21142 & ~n24107;
  assign n24475 = ~n24106 & ~n24474;
  assign n24476 = n21059 & n21141;
  assign n24477 = ~n21059 & ~n21141;
  assign n24478 = ~n24476 & ~n24477;
  assign n24479 = n24106 & ~n24478;
  assign n24480 = ~n24475 & ~n24479;
  assign n24481 = ~pi0868 & ~n24480;
  assign n24482 = ~n24473 & ~n24481;
  assign n24483 = n20524 & ~n24482;
  assign n24484 = ~n24472 & ~n24483;
  assign n24485 = pi0049 & ~n24252;
  assign n24486 = ~pi3245 & ~n11181;
  assign n24487 = pi3245 & ~n16529;
  assign n24488 = ~n24486 & ~n24487;
  assign n24489 = n24252 & ~n24488;
  assign n24490 = ~n24485 & ~n24489;
  assign n24491 = n24261 & ~n24490;
  assign n24492 = ~n24267 & ~n24491;
  assign n24493 = ~n20521 & ~n24492;
  assign n24494 = ~n24271 & ~n24493;
  assign n24495 = ~n20524 & ~n24494;
  assign po0319 = ~n24484 | n24495;
  assign n24497 = pi0050 & ~n24304;
  assign n24498 = n24302 & n24497;
  assign n24499 = n24304 & ~n24482;
  assign n24500 = ~n24498 & ~n24499;
  assign n24501 = pi0050 & ~n24310;
  assign n24502 = n24310 & ~n24488;
  assign n24503 = ~n24501 & ~n24502;
  assign n24504 = n24316 & ~n24503;
  assign n24505 = ~n24319 & ~n24504;
  assign n24506 = ~n24302 & ~n24505;
  assign n24507 = ~n24323 & ~n24506;
  assign n24508 = ~n24304 & ~n24507;
  assign po0320 = ~n24500 | n24508;
  assign n24510 = pi0051 & ~n20524;
  assign n24511 = n20521 & n24510;
  assign n24512 = pi2384 & ~n13848;
  assign n24513 = ~pi0868 & n24512;
  assign n24514 = pi0868 & n24194;
  assign n24515 = ~n24513 & ~n24514;
  assign n24516 = pi1472 & ~n24515;
  assign n24517 = n20917 & n24516;
  assign n24518 = ~n20917 & ~n24516;
  assign n24519 = ~n24517 & ~n24518;
  assign n24520 = ~n20916 & n24198;
  assign n24521 = ~n20915 & ~n24520;
  assign n24522 = ~n24519 & n24521;
  assign n24523 = ~n20817 & ~n24522;
  assign n24524 = pi2384 & ~n13182;
  assign n24525 = ~pi0868 & n24524;
  assign n24526 = pi0868 & n24512;
  assign n24527 = ~n24525 & ~n24526;
  assign n24528 = pi1472 & ~n24527;
  assign n24529 = n20917 & n24528;
  assign n24530 = ~n20917 & ~n24528;
  assign n24531 = ~n24529 & ~n24530;
  assign n24532 = ~n20916 & n24516;
  assign n24533 = ~n20915 & ~n24532;
  assign n24534 = ~n24531 & ~n24533;
  assign n24535 = n24531 & n24533;
  assign n24536 = ~n24534 & ~n24535;
  assign n24537 = n20820 & ~n24536;
  assign n24538 = ~n20820 & n24536;
  assign n24539 = ~n24537 & ~n24538;
  assign n24540 = n24523 & n24539;
  assign n24541 = ~n24523 & ~n24539;
  assign n24542 = ~n24540 & ~n24541;
  assign n24543 = ~n24519 & ~n24521;
  assign n24544 = n24519 & n24521;
  assign n24545 = ~n24543 & ~n24544;
  assign n24546 = n20820 & ~n24545;
  assign n24547 = ~n20820 & n24545;
  assign n24548 = ~n24546 & ~n24547;
  assign n24549 = n24519 & ~n24521;
  assign n24550 = ~n24548 & ~n24549;
  assign n24551 = ~n20819 & n24550;
  assign n24552 = ~n24201 & n24203;
  assign n24553 = ~n20817 & ~n24552;
  assign n24554 = n24548 & ~n24553;
  assign n24555 = ~n24551 & ~n24554;
  assign n24556 = ~n24542 & n24555;
  assign n24557 = n24542 & ~n24555;
  assign n24558 = ~n24556 & ~n24557;
  assign n24559 = n20903 & ~n24558;
  assign n24560 = ~n20903 & n24558;
  assign n24561 = ~n24559 & ~n24560;
  assign n24562 = ~n20942 & n24561;
  assign n24563 = n24542 & n24555;
  assign n24564 = n24562 & ~n24563;
  assign n24565 = n24201 & ~n24203;
  assign n24566 = ~n24209 & ~n24565;
  assign n24567 = ~n20819 & n24566;
  assign n24568 = ~n24193 & n24209;
  assign n24569 = ~n24567 & ~n24568;
  assign n24570 = n24548 & n24553;
  assign n24571 = ~n24548 & ~n24553;
  assign n24572 = ~n24570 & ~n24571;
  assign n24573 = ~n24569 & ~n24572;
  assign n24574 = n20655 & ~n24573;
  assign n24575 = n20652 & n24572;
  assign n24576 = ~n24574 & ~n24575;
  assign n24577 = n20652 & n24569;
  assign n24578 = n24576 & ~n24577;
  assign n24579 = ~n24561 & n24578;
  assign n24580 = ~n24564 & ~n24579;
  assign n24581 = ~n24542 & ~n24555;
  assign n24582 = n20655 & ~n24581;
  assign n24583 = n20652 & n24542;
  assign n24584 = ~n24582 & ~n24583;
  assign n24585 = n20652 & n24555;
  assign n24586 = n24584 & ~n24585;
  assign n24587 = ~n24531 & n24533;
  assign n24588 = ~n20817 & ~n24587;
  assign n24589 = pi2384 & ~n9498;
  assign n24590 = ~pi0868 & n24589;
  assign n24591 = pi0868 & n24524;
  assign n24592 = ~n24590 & ~n24591;
  assign n24593 = pi1472 & ~n24592;
  assign n24594 = n20917 & n24593;
  assign n24595 = ~n20917 & ~n24593;
  assign n24596 = ~n24594 & ~n24595;
  assign n24597 = ~n20916 & n24528;
  assign n24598 = ~n20915 & ~n24597;
  assign n24599 = ~n24596 & ~n24598;
  assign n24600 = n24596 & n24598;
  assign n24601 = ~n24599 & ~n24600;
  assign n24602 = n20820 & ~n24601;
  assign n24603 = ~n20820 & n24601;
  assign n24604 = ~n24602 & ~n24603;
  assign n24605 = n24588 & n24604;
  assign n24606 = ~n24588 & ~n24604;
  assign n24607 = ~n24605 & ~n24606;
  assign n24608 = n24531 & ~n24533;
  assign n24609 = ~n24539 & ~n24608;
  assign n24610 = ~n20819 & n24609;
  assign n24611 = ~n24523 & n24539;
  assign n24612 = ~n24610 & ~n24611;
  assign n24613 = ~n24607 & n24612;
  assign n24614 = n24607 & ~n24612;
  assign n24615 = ~n24613 & ~n24614;
  assign n24616 = n20903 & ~n24615;
  assign n24617 = ~n20903 & n24615;
  assign n24618 = ~n24616 & ~n24617;
  assign n24619 = ~n24586 & n24618;
  assign n24620 = n24586 & ~n24618;
  assign n24621 = ~n24619 & ~n24620;
  assign n24622 = ~n24580 & n24621;
  assign n24623 = n24580 & ~n24621;
  assign n24624 = ~n24622 & ~n24623;
  assign n24625 = ~n24191 & ~n24212;
  assign n24626 = n20652 & ~n24625;
  assign n24627 = n20655 & n24212;
  assign n24628 = ~n24626 & ~n24627;
  assign n24629 = n20655 & n24191;
  assign n24630 = n24628 & ~n24629;
  assign n24631 = n24569 & ~n24572;
  assign n24632 = ~n24569 & n24572;
  assign n24633 = ~n24631 & ~n24632;
  assign n24634 = n20903 & ~n24633;
  assign n24635 = ~n20903 & n24633;
  assign n24636 = ~n24634 & ~n24635;
  assign n24637 = n24630 & ~n24636;
  assign n24638 = ~n20942 & n24636;
  assign n24639 = n24569 & n24572;
  assign n24640 = n24638 & ~n24639;
  assign n24641 = ~n24637 & ~n24640;
  assign n24642 = n24561 & ~n24578;
  assign n24643 = ~n24579 & ~n24642;
  assign n24644 = n24641 & ~n24643;
  assign n24645 = ~n24630 & n24636;
  assign n24646 = ~n24637 & ~n24645;
  assign n24647 = n24223 & ~n24646;
  assign n24648 = ~n20942 & n24218;
  assign n24649 = n24191 & n24212;
  assign n24650 = n24648 & ~n24649;
  assign n24651 = ~n24218 & ~n24220;
  assign n24652 = ~n24650 & ~n24651;
  assign n24653 = n24223 & n24652;
  assign n24654 = ~n24647 & ~n24653;
  assign n24655 = n24186 & ~n24654;
  assign n24656 = ~n24646 & n24652;
  assign n24657 = ~n24655 & ~n24656;
  assign n24658 = n24646 & ~n24652;
  assign n24659 = n24186 & ~n24658;
  assign n24660 = ~n24647 & ~n24659;
  assign n24661 = ~n24653 & n24660;
  assign n24662 = ~n24243 & ~n24661;
  assign n24663 = n24657 & ~n24662;
  assign n24664 = ~n24641 & n24643;
  assign n24665 = ~n24663 & ~n24664;
  assign n24666 = ~n24644 & ~n24665;
  assign n24667 = ~n24624 & n24666;
  assign n24668 = n24624 & ~n24666;
  assign n24669 = ~n24667 & ~n24668;
  assign n24670 = ~pi0868 & n24669;
  assign n24671 = ~n24596 & n24598;
  assign n24672 = ~n20817 & ~n24671;
  assign n24673 = ~n20916 & n24593;
  assign n24674 = ~n20915 & ~n24673;
  assign n24675 = pi1472 & n24589;
  assign n24676 = n20917 & n24675;
  assign n24677 = ~n20917 & ~n24675;
  assign n24678 = ~n24676 & ~n24677;
  assign n24679 = n24674 & n24678;
  assign n24680 = ~n24674 & ~n24678;
  assign n24681 = ~n24679 & ~n24680;
  assign n24682 = n20820 & ~n24681;
  assign n24683 = ~n20820 & n24681;
  assign n24684 = ~n24682 & ~n24683;
  assign n24685 = n24672 & n24684;
  assign n24686 = ~n24672 & ~n24684;
  assign n24687 = ~n24685 & ~n24686;
  assign n24688 = n24596 & ~n24598;
  assign n24689 = ~n24604 & ~n24688;
  assign n24690 = ~n20819 & n24689;
  assign n24691 = ~n24588 & n24604;
  assign n24692 = ~n24690 & ~n24691;
  assign n24693 = ~n24687 & n24692;
  assign n24694 = n24687 & ~n24692;
  assign n24695 = ~n24693 & ~n24694;
  assign n24696 = n20903 & ~n24695;
  assign n24697 = ~n20903 & n24695;
  assign n24698 = ~n24696 & ~n24697;
  assign n24699 = ~n24607 & ~n24612;
  assign n24700 = n20655 & ~n24699;
  assign n24701 = n20652 & n24607;
  assign n24702 = ~n24700 & ~n24701;
  assign n24703 = n20652 & n24612;
  assign n24704 = n24702 & ~n24703;
  assign n24705 = ~n24698 & n24704;
  assign n24706 = n24698 & ~n24704;
  assign n24707 = ~n24705 & ~n24706;
  assign n24708 = ~n20942 & n24618;
  assign n24709 = n24607 & n24612;
  assign n24710 = n24708 & ~n24709;
  assign n24711 = ~n24620 & ~n24710;
  assign n24712 = ~n24707 & n24711;
  assign n24713 = n24707 & ~n24711;
  assign n24714 = ~n24712 & ~n24713;
  assign n24715 = ~n24622 & ~n24664;
  assign n24716 = ~n24661 & n24715;
  assign n24717 = n24236 & n24716;
  assign n24718 = ~n24091 & n24717;
  assign n24719 = n24097 & n24718;
  assign n24720 = ~n23308 & n24717;
  assign n24721 = n24230 & n24716;
  assign n24722 = ~n24720 & ~n24721;
  assign n24723 = ~n24235 & n24716;
  assign n24724 = ~n24657 & n24715;
  assign n24725 = ~n24723 & ~n24724;
  assign n24726 = n24621 & ~n24644;
  assign n24727 = n24580 & ~n24726;
  assign n24728 = ~n24621 & ~n24643;
  assign n24729 = n24641 & n24728;
  assign n24730 = ~n24727 & ~n24729;
  assign n24731 = n24725 & n24730;
  assign n24732 = n24722 & n24731;
  assign n24733 = ~n24719 & n24732;
  assign n24734 = ~n24714 & n24733;
  assign n24735 = n24714 & ~n24733;
  assign n24736 = ~n24734 & ~n24735;
  assign n24737 = pi0868 & n24736;
  assign n24738 = ~n24670 & ~n24737;
  assign n24739 = n20524 & ~n24738;
  assign n24740 = ~n24511 & ~n24739;
  assign n24741 = pi0051 & ~n24252;
  assign n24742 = pi3245 & ~n16784;
  assign n24743 = ~pi3245 & ~n13121;
  assign n24744 = ~n24742 & ~n24743;
  assign n24745 = n24252 & ~n24744;
  assign n24746 = ~n24741 & ~n24745;
  assign n24747 = n24261 & ~n24746;
  assign n24748 = ~n24267 & ~n24747;
  assign n24749 = ~n20521 & ~n24748;
  assign n24750 = ~n24271 & ~n24749;
  assign n24751 = ~n20524 & ~n24750;
  assign po0321 = ~n24740 | n24751;
  assign n24753 = pi0052 & ~n20524;
  assign n24754 = n20521 & n24753;
  assign n24755 = ~n24641 & ~n24643;
  assign n24756 = n24641 & n24643;
  assign n24757 = ~n24755 & ~n24756;
  assign n24758 = ~n24663 & ~n24757;
  assign n24759 = n24663 & n24757;
  assign n24760 = ~n24758 & ~n24759;
  assign n24761 = ~pi0868 & n24760;
  assign n24762 = pi0868 & n24669;
  assign n24763 = ~n24761 & ~n24762;
  assign n24764 = n20524 & ~n24763;
  assign n24765 = ~n24754 & ~n24764;
  assign n24766 = pi0052 & ~n24252;
  assign n24767 = pi3245 & ~n16748;
  assign n24768 = ~pi3245 & ~n13398;
  assign n24769 = ~n24767 & ~n24768;
  assign n24770 = n24252 & ~n24769;
  assign n24771 = ~n24766 & ~n24770;
  assign n24772 = n24261 & ~n24771;
  assign n24773 = ~n24267 & ~n24772;
  assign n24774 = ~n20521 & ~n24773;
  assign n24775 = ~n24271 & ~n24774;
  assign n24776 = ~n20524 & ~n24775;
  assign po0322 = ~n24765 | n24776;
  assign n24778 = pi0053 & ~n24304;
  assign n24779 = n24302 & n24778;
  assign n24780 = n24304 & ~n24738;
  assign n24781 = ~n24779 & ~n24780;
  assign n24782 = pi0053 & ~n24310;
  assign n24783 = n24310 & ~n24744;
  assign n24784 = ~n24782 & ~n24783;
  assign n24785 = n24316 & ~n24784;
  assign n24786 = ~n24319 & ~n24785;
  assign n24787 = ~n24302 & ~n24786;
  assign n24788 = ~n24323 & ~n24787;
  assign n24789 = ~n24304 & ~n24788;
  assign po0323 = ~n24781 | n24789;
  assign n24791 = pi0054 & ~n24304;
  assign n24792 = n24302 & n24791;
  assign n24793 = n24304 & ~n24763;
  assign n24794 = ~n24792 & ~n24793;
  assign n24795 = pi0054 & ~n24310;
  assign n24796 = n24310 & ~n24769;
  assign n24797 = ~n24795 & ~n24796;
  assign n24798 = n24316 & ~n24797;
  assign n24799 = ~n24319 & ~n24798;
  assign n24800 = ~n24302 & ~n24799;
  assign n24801 = ~n24323 & ~n24800;
  assign n24802 = ~n24304 & ~n24801;
  assign po0324 = ~n24794 | n24802;
  assign n24804 = ~pi0410 & ~pi0426;
  assign n24805 = pi0409 & n24804;
  assign n24806 = ~pi0423 & ~pi0424;
  assign n24807 = ~pi0405 & ~pi0422;
  assign n24808 = n24806 & n24807;
  assign n24809 = ~pi0421 & ~n24808;
  assign n24810 = ~n8615 & ~n10749;
  assign n24811 = ~pi0418 & n8608;
  assign n24812 = ~pi0419 & n24811;
  assign n24813 = pi0403 & n24812;
  assign n24814 = pi0418 & n8608;
  assign n24815 = pi0403 & n24814;
  assign n24816 = ~n24813 & ~n24815;
  assign n24817 = ~n8619 & n24816;
  assign n24818 = n24810 & n24817;
  assign n24819 = n24809 & ~n24818;
  assign n24820 = pi0409 & pi0410;
  assign n24821 = pi0426 & n24820;
  assign n24822 = ~pi2140 & n19553;
  assign n24823 = pi0709 & ~pi3426;
  assign n24824 = ~n24822 & ~n24823;
  assign n24825 = n24821 & ~n24824;
  assign n24826 = pi0408 & n24813;
  assign n24827 = n24809 & n24826;
  assign n24828 = pi0426 & n24827;
  assign n24829 = n24827 & n24828;
  assign n24830 = ~pi0409 & n24827;
  assign n24831 = ~pi0406 & ~n24827;
  assign n24832 = ~n24830 & ~n24831;
  assign n24833 = ~pi0425 & ~n24827;
  assign n24834 = ~pi0410 & n24827;
  assign n24835 = ~n24833 & ~n24834;
  assign n24836 = n24832 & n24835;
  assign n24837 = n24829 & n24836;
  assign n24838 = n24823 & n24837;
  assign n24839 = ~n24825 & ~n24838;
  assign n24840 = n24832 & ~n24835;
  assign n24841 = n24829 & n24840;
  assign n24842 = ~pi0410 & pi0426;
  assign n24843 = pi0409 & n24842;
  assign n24844 = ~n24841 & ~n24843;
  assign n24845 = n24822 & ~n24844;
  assign n24846 = pi0710 & ~pi3426;
  assign n24847 = n24843 & n24846;
  assign n24848 = ~n24845 & ~n24847;
  assign n24849 = n24827 & ~n24828;
  assign n24850 = n24840 & n24849;
  assign n24851 = ~n24805 & ~n24850;
  assign n24852 = ~pi2020 & n19553;
  assign n24853 = pi0715 & ~pi3426;
  assign n24854 = ~n24852 & ~n24853;
  assign n24855 = ~n24851 & ~n24854;
  assign n24856 = n24822 & n24837;
  assign n24857 = n24841 & n24846;
  assign n24858 = ~n24856 & ~n24857;
  assign n24859 = ~n24855 & n24858;
  assign n24860 = n24848 & n24859;
  assign n24861 = n24839 & n24860;
  assign n24862 = pi0410 & ~pi0426;
  assign n24863 = pi0409 & n24862;
  assign n24864 = n20515 & n24863;
  assign n24865 = ~pi0695 & ~pi3426;
  assign n24866 = ~n20515 & ~n24865;
  assign n24867 = n24836 & n24849;
  assign n24868 = ~n24866 & n24867;
  assign n24869 = ~pi0409 & ~pi0410;
  assign n24870 = pi0426 & n24869;
  assign n24871 = ~n24832 & n24835;
  assign n24872 = n24829 & n24871;
  assign n24873 = ~pi0409 & pi0426;
  assign n24874 = pi0410 & n24873;
  assign n24875 = ~n24872 & ~n24874;
  assign n24876 = ~n24832 & ~n24835;
  assign n24877 = n24829 & n24876;
  assign n24878 = n24875 & ~n24877;
  assign n24879 = ~n24870 & n24878;
  assign n24880 = ~n20516 & ~n24879;
  assign n24881 = n20519 & ~n24875;
  assign n24882 = ~n24880 & ~n24881;
  assign n24883 = n24863 & n24865;
  assign n24884 = n24882 & ~n24883;
  assign n24885 = ~n24868 & n24884;
  assign n24886 = ~n24864 & n24885;
  assign n24887 = n24861 & n24886;
  assign n24888 = n24819 & ~n24887;
  assign n24889 = n24805 & n24888;
  assign n24890 = ~pi0715 & ~po3872;
  assign n24891 = n24889 & n24890;
  assign n24892 = ~n20388 & n24891;
  assign n24893 = ~n20263 & ~n20334;
  assign n24894 = n20150 & n20379;
  assign n24895 = ~n20150 & ~n20153;
  assign n24896 = ~n20380 & n24895;
  assign n24897 = ~n24894 & ~n24896;
  assign n24898 = n24893 & n24897;
  assign n24899 = ~n24893 & ~n24897;
  assign n24900 = ~n24898 & ~n24899;
  assign n24901 = n24892 & ~n24900;
  assign n24902 = ~po3872 & n24805;
  assign n24903 = ~n24888 & n24902;
  assign n24904 = po3872 & n19619;
  assign n24905 = ~n24903 & ~n24904;
  assign n24906 = ~n14882 & ~n24905;
  assign n24907 = ~n24901 & ~n24906;
  assign n24908 = n20388 & n24891;
  assign n24909 = ~n20427 & n24908;
  assign n24910 = n24907 & ~n24909;
  assign n24911 = ~po3872 & n24889;
  assign n24912 = pi0715 & pi3245;
  assign n24913 = n24911 & n24912;
  assign n24914 = ~n16604 & n24913;
  assign n24915 = ~pi3245 & n24911;
  assign n24916 = pi0715 & n24915;
  assign n24917 = ~n15115 & n24916;
  assign n24918 = ~n24914 & ~n24917;
  assign n24919 = pi0409 & pi0426;
  assign n24920 = ~po3872 & n24919;
  assign n24921 = ~pi0410 & n24920;
  assign n24922 = ~n24888 & n24921;
  assign n24923 = ~n14997 & n24922;
  assign n24924 = pi0410 & n24920;
  assign n24925 = ~n24888 & n24924;
  assign n24926 = ~n14993 & n24925;
  assign n24927 = ~n24923 & ~n24926;
  assign n24928 = pi3504 & pi3514;
  assign n24929 = ~pi2021 & ~n24928;
  assign n24930 = ~n13288 & n19607;
  assign n24931 = ~n20004 & ~n24930;
  assign n24932 = n24929 & ~n24931;
  assign n24933 = pi3504 & ~pi3514;
  assign n24934 = n11024 & n24933;
  assign n24935 = pi2486 & ~n11024;
  assign n24936 = ~pi2486 & ~pi3394;
  assign n24937 = ~n24935 & ~n24936;
  assign n24938 = ~n24933 & n24937;
  assign n24939 = ~n24934 & ~n24938;
  assign n24940 = n24929 & n24939;
  assign n24941 = pi3518 & n24929;
  assign n24942 = n12208 & n15011;
  assign n24943 = n11024 & n11841;
  assign n24944 = n14623 & n24943;
  assign n24945 = n24942 & n24944;
  assign n24946 = n13781 & n24945;
  assign n24947 = ~n13781 & ~n24945;
  assign n24948 = ~n24946 & ~n24947;
  assign n24949 = n24933 & ~n24948;
  assign n24950 = pi2486 & ~n13781;
  assign n24951 = ~pi2486 & pi3511;
  assign n24952 = ~n24950 & ~n24951;
  assign n24953 = ~n24933 & n24952;
  assign n24954 = ~n24949 & ~n24953;
  assign n24955 = n24929 & n24954;
  assign n24956 = n15011 & n24943;
  assign n24957 = n14623 & n24956;
  assign n24958 = n12208 & n13781;
  assign n24959 = n13284 & n24958;
  assign n24960 = n24957 & n24959;
  assign n24961 = n9530 & ~n24960;
  assign n24962 = ~n9530 & n24960;
  assign n24963 = ~n24961 & ~n24962;
  assign n24964 = n24933 & n24963;
  assign n24965 = pi2486 & ~n9530;
  assign n24966 = ~pi2486 & pi3521;
  assign n24967 = ~n24965 & ~n24966;
  assign n24968 = ~n24933 & n24967;
  assign n24969 = ~n24964 & ~n24968;
  assign n24970 = n24929 & n24969;
  assign n24971 = n24944 & n24958;
  assign n24972 = n15011 & n24971;
  assign n24973 = n13284 & n24972;
  assign n24974 = ~n13284 & ~n24972;
  assign n24975 = ~n24973 & ~n24974;
  assign n24976 = n24933 & ~n24975;
  assign n24977 = pi2486 & n13284;
  assign n24978 = ~pi2486 & ~pi3510;
  assign n24979 = ~n24977 & ~n24978;
  assign n24980 = ~n24933 & ~n24979;
  assign n24981 = ~n24976 & ~n24980;
  assign n24982 = n24929 & n24981;
  assign n24983 = n24970 & n24982;
  assign n24984 = n24955 & n24983;
  assign n24985 = ~n24941 & n24984;
  assign n24986 = ~n14623 & ~n24956;
  assign n24987 = ~n24957 & ~n24986;
  assign n24988 = n24933 & ~n24987;
  assign n24989 = pi2486 & ~n14623;
  assign n24990 = ~pi2486 & pi3398;
  assign n24991 = ~n24989 & ~n24990;
  assign n24992 = ~n24933 & n24991;
  assign n24993 = ~n24988 & ~n24992;
  assign n24994 = n24929 & n24993;
  assign n24995 = ~n11024 & n11841;
  assign n24996 = n11024 & ~n11841;
  assign n24997 = ~n24995 & ~n24996;
  assign n24998 = n24933 & ~n24997;
  assign n24999 = pi2486 & ~n11841;
  assign n25000 = ~pi2486 & ~pi3330;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = ~n24933 & ~n25001;
  assign n25003 = ~n24998 & ~n25002;
  assign n25004 = n24929 & ~n25003;
  assign n25005 = n24994 & ~n25004;
  assign n25006 = n12208 & n24957;
  assign n25007 = ~n12208 & ~n24957;
  assign n25008 = ~n25006 & ~n25007;
  assign n25009 = n24933 & ~n25008;
  assign n25010 = pi2486 & ~n12208;
  assign n25011 = ~pi2486 & pi3520;
  assign n25012 = ~n25010 & ~n25011;
  assign n25013 = ~n24933 & n25012;
  assign n25014 = ~n25009 & ~n25013;
  assign n25015 = n24929 & n25014;
  assign n25016 = ~n15011 & ~n24943;
  assign n25017 = ~n24956 & ~n25016;
  assign n25018 = n24933 & ~n25017;
  assign n25019 = pi2486 & n15011;
  assign n25020 = ~pi2486 & ~pi3392;
  assign n25021 = ~n25019 & ~n25020;
  assign n25022 = ~n24933 & ~n25021;
  assign n25023 = ~n25018 & ~n25022;
  assign n25024 = n24929 & n25023;
  assign n25025 = n25015 & n25024;
  assign n25026 = n25005 & n25025;
  assign n25027 = n24985 & n25026;
  assign n25028 = ~n24940 & n25027;
  assign n25029 = n24932 & n25028;
  assign n25030 = ~n10452 & n19607;
  assign n25031 = ~n19913 & ~n25030;
  assign n25032 = n24929 & ~n25031;
  assign n25033 = ~n24994 & n25004;
  assign n25034 = n25025 & n25033;
  assign n25035 = n24985 & n25034;
  assign n25036 = ~n24940 & n25035;
  assign n25037 = n25032 & n25036;
  assign n25038 = ~n25029 & ~n25037;
  assign n25039 = ~n11846 & n19607;
  assign n25040 = ~n20172 & ~n25039;
  assign n25041 = n24929 & ~n25040;
  assign n25042 = ~n24970 & ~n24982;
  assign n25043 = ~n24941 & ~n24955;
  assign n25044 = n25042 & n25043;
  assign n25045 = ~n25015 & ~n25024;
  assign n25046 = ~n24994 & ~n25004;
  assign n25047 = n25045 & n25046;
  assign n25048 = n25044 & n25047;
  assign n25049 = n24940 & n25048;
  assign n25050 = n25041 & n25049;
  assign n25051 = n25038 & ~n25050;
  assign n25052 = ~n17213 & n19607;
  assign n25053 = ~n19629 & ~n25052;
  assign n25054 = ~pi3504 & pi3514;
  assign n25055 = ~n25053 & n25054;
  assign n25056 = pi0196 & n24933;
  assign n25057 = pi0152 & ~pi3518;
  assign n25058 = n25056 & n25057;
  assign n25059 = ~n25055 & ~n25058;
  assign n25060 = n24929 & ~n25059;
  assign n25061 = n25015 & ~n25024;
  assign n25062 = n25046 & n25061;
  assign n25063 = n24985 & n25062;
  assign n25064 = n24940 & n25063;
  assign n25065 = n25060 & n25064;
  assign n25066 = n24994 & n25004;
  assign n25067 = ~n25015 & n25024;
  assign n25068 = n25066 & n25067;
  assign n25069 = n24985 & n25068;
  assign n25070 = n24940 & n25069;
  assign n25071 = n25060 & n25070;
  assign n25072 = ~n25065 & ~n25071;
  assign n25073 = n24941 & ~n24955;
  assign n25074 = n25042 & n25073;
  assign n25075 = n25047 & n25074;
  assign n25076 = n24940 & n25075;
  assign n25077 = n25060 & n25076;
  assign n25078 = ~n24940 & n25075;
  assign n25079 = n25060 & n25078;
  assign n25080 = ~n25077 & ~n25079;
  assign n25081 = n25072 & n25080;
  assign n25082 = n25005 & n25045;
  assign n25083 = n24985 & n25082;
  assign n25084 = ~n24940 & n25083;
  assign n25085 = n25060 & n25084;
  assign n25086 = n24940 & n25083;
  assign n25087 = n25060 & n25086;
  assign n25088 = ~n25085 & ~n25087;
  assign n25089 = n25045 & n25066;
  assign n25090 = n24985 & n25089;
  assign n25091 = ~n24940 & n25090;
  assign n25092 = n25060 & n25091;
  assign n25093 = n25088 & ~n25092;
  assign n25094 = n25081 & n25093;
  assign n25095 = n25033 & n25067;
  assign n25096 = n25074 & n25095;
  assign n25097 = ~n24940 & n25096;
  assign n25098 = n25032 & n25097;
  assign n25099 = n25074 & n25082;
  assign n25100 = ~n24940 & n25099;
  assign n25101 = ~n14251 & n19607;
  assign n25102 = ~n19785 & ~n25101;
  assign n25103 = n24929 & ~n25102;
  assign n25104 = n25100 & n25103;
  assign n25105 = ~n25098 & ~n25104;
  assign n25106 = pi3516 & ~n14993;
  assign n25107 = n24941 & n24984;
  assign n25108 = n25005 & n25061;
  assign n25109 = n25107 & n25108;
  assign n25110 = n24940 & n25109;
  assign n25111 = n25060 & n25110;
  assign n25112 = n25061 & n25066;
  assign n25113 = n25107 & n25112;
  assign n25114 = ~n24940 & n25113;
  assign n25115 = n25060 & n25114;
  assign n25116 = ~n25111 & ~n25115;
  assign n25117 = ~n24982 & n25060;
  assign n25118 = n24970 & n25117;
  assign n25119 = n24941 & n25118;
  assign n25120 = n25033 & n25061;
  assign n25121 = n25107 & n25120;
  assign n25122 = n24940 & n25121;
  assign n25123 = n25060 & n25122;
  assign n25124 = ~n25119 & ~n25123;
  assign n25125 = n25033 & n25045;
  assign n25126 = n24985 & n25125;
  assign n25127 = ~n24940 & n25126;
  assign n25128 = n25060 & n25127;
  assign n25129 = n24985 & n25095;
  assign n25130 = n24940 & n25129;
  assign n25131 = n25060 & n25130;
  assign n25132 = ~n25128 & ~n25131;
  assign n25133 = n25124 & n25132;
  assign n25134 = n25116 & n25133;
  assign n25135 = ~n25106 & n25134;
  assign n25136 = n25105 & n25135;
  assign n25137 = n25062 & n25107;
  assign n25138 = ~n24940 & n25060;
  assign n25139 = n25137 & n25138;
  assign n25140 = n25025 & n25066;
  assign n25141 = n25107 & n25140;
  assign n25142 = n24940 & n25141;
  assign n25143 = n25060 & n25142;
  assign n25144 = ~n25139 & ~n25143;
  assign n25145 = n24985 & n25112;
  assign n25146 = n24940 & n25145;
  assign n25147 = ~n12954 & n19607;
  assign n25148 = ~n19969 & ~n25147;
  assign n25149 = n24929 & ~n25148;
  assign n25150 = n25146 & n25149;
  assign n25151 = n24929 & ~n25053;
  assign n25152 = n25074 & n25125;
  assign n25153 = n24940 & n25152;
  assign n25154 = n25151 & n25153;
  assign n25155 = ~n25150 & ~n25154;
  assign n25156 = ~n12512 & n19607;
  assign n25157 = ~n19743 & ~n25156;
  assign n25158 = n24929 & ~n25157;
  assign n25159 = n24985 & n25108;
  assign n25160 = n24940 & n25159;
  assign n25161 = n25158 & n25160;
  assign n25162 = ~n24940 & n25145;
  assign n25163 = ~n13548 & n19607;
  assign n25164 = ~n19827 & ~n25163;
  assign n25165 = n24929 & ~n25164;
  assign n25166 = n25162 & n25165;
  assign n25167 = ~n25161 & ~n25166;
  assign n25168 = n24985 & n25120;
  assign n25169 = n24940 & n25168;
  assign n25170 = n25151 & n25169;
  assign n25171 = n25167 & ~n25170;
  assign n25172 = ~n24940 & n25168;
  assign n25173 = n25060 & n25172;
  assign n25174 = n25171 & ~n25173;
  assign n25175 = n25005 & n25067;
  assign n25176 = n24985 & n25175;
  assign n25177 = ~n24940 & n25176;
  assign n25178 = n25060 & n25177;
  assign n25179 = ~n24940 & n25109;
  assign n25180 = n25060 & n25179;
  assign n25181 = ~n25178 & ~n25180;
  assign n25182 = ~n24940 & n25121;
  assign n25183 = n25060 & n25182;
  assign n25184 = ~n24940 & n25159;
  assign n25185 = n25103 & n25184;
  assign n25186 = ~n25183 & ~n25185;
  assign n25187 = n25181 & n25186;
  assign n25188 = n25062 & n25074;
  assign n25189 = n24940 & n25188;
  assign n25190 = n25041 & n25189;
  assign n25191 = n25187 & ~n25190;
  assign n25192 = n25174 & n25191;
  assign n25193 = n25155 & n25192;
  assign n25194 = n25144 & n25193;
  assign n25195 = n24940 & n25027;
  assign n25196 = ~n13785 & n19607;
  assign n25197 = ~n20100 & ~n25196;
  assign n25198 = n24929 & ~n25197;
  assign n25199 = n25195 & n25198;
  assign n25200 = ~n14614 & n19607;
  assign n25201 = ~n20060 & ~n25200;
  assign n25202 = n24929 & ~n25201;
  assign n25203 = n24985 & n25140;
  assign n25204 = n24940 & n25203;
  assign n25205 = n25202 & n25204;
  assign n25206 = ~n25199 & ~n25205;
  assign n25207 = ~n24940 & n25141;
  assign n25208 = n25060 & n25207;
  assign n25209 = ~n24940 & n25063;
  assign n25210 = n25060 & n25209;
  assign n25211 = ~n25208 & ~n25210;
  assign n25212 = n25206 & n25211;
  assign n25213 = n24940 & n25113;
  assign n25214 = n25060 & n25213;
  assign n25215 = n24940 & n25090;
  assign n25216 = n25060 & n25215;
  assign n25217 = ~n25214 & ~n25216;
  assign n25218 = n25046 & n25067;
  assign n25219 = n24985 & n25218;
  assign n25220 = n24940 & n25219;
  assign n25221 = n25060 & n25220;
  assign n25222 = n25025 & n25046;
  assign n25223 = n25107 & n25222;
  assign n25224 = n24940 & n25223;
  assign n25225 = n25060 & n25224;
  assign n25226 = ~n25221 & ~n25225;
  assign n25227 = n25217 & n25226;
  assign n25228 = ~n15002 & n19607;
  assign n25229 = ~n20128 & ~n25228;
  assign n25230 = n24929 & ~n25229;
  assign n25231 = ~n24940 & n25048;
  assign n25232 = n25230 & n25231;
  assign n25233 = n25227 & ~n25232;
  assign n25234 = n24940 & n25096;
  assign n25235 = ~n15273 & n19607;
  assign n25236 = ~n19709 & ~n25235;
  assign n25237 = n24929 & ~n25236;
  assign n25238 = n25234 & n25237;
  assign n25239 = n24940 & n25099;
  assign n25240 = n25158 & n25239;
  assign n25241 = ~n25238 & ~n25240;
  assign n25242 = n24985 & n25222;
  assign n25243 = ~n24940 & n25242;
  assign n25244 = ~n17010 & n19607;
  assign n25245 = ~n19671 & ~n25244;
  assign n25246 = n24929 & ~n25245;
  assign n25247 = n25243 & n25246;
  assign n25248 = n24940 & n25242;
  assign n25249 = ~n9526 & n19607;
  assign n25250 = ~n19867 & ~n25249;
  assign n25251 = n24929 & ~n25250;
  assign n25252 = n25248 & n25251;
  assign n25253 = ~n25247 & ~n25252;
  assign n25254 = ~n24940 & n25152;
  assign n25255 = n25060 & n25254;
  assign n25256 = n25034 & n25107;
  assign n25257 = n24940 & n25256;
  assign n25258 = n25060 & n25257;
  assign n25259 = ~n25255 & ~n25258;
  assign n25260 = n25253 & n25259;
  assign n25261 = ~n24940 & n25188;
  assign n25262 = n25230 & n25261;
  assign n25263 = n25260 & ~n25262;
  assign n25264 = ~n24940 & n25203;
  assign n25265 = ~n12212 & n19607;
  assign n25266 = ~n20282 & ~n25265;
  assign n25267 = n24929 & ~n25266;
  assign n25268 = n25264 & n25267;
  assign n25269 = n25068 & n25074;
  assign n25270 = n24940 & n25269;
  assign n25271 = n25202 & n25270;
  assign n25272 = ~n25268 & ~n25271;
  assign n25273 = n25263 & n25272;
  assign n25274 = n25241 & n25273;
  assign n25275 = n25233 & n25274;
  assign n25276 = ~n24940 & n25069;
  assign n25277 = n25060 & n25276;
  assign n25278 = ~n24940 & n25256;
  assign n25279 = n25060 & n25278;
  assign n25280 = ~n25277 & ~n25279;
  assign n25281 = n24940 & n25035;
  assign n25282 = n25237 & n25281;
  assign n25283 = n25280 & ~n25282;
  assign n25284 = n24940 & n25137;
  assign n25285 = n25060 & n25284;
  assign n25286 = n25074 & n25120;
  assign n25287 = ~n24940 & n25286;
  assign n25288 = ~n11029 & n19607;
  assign n25289 = ~n20211 & ~n25288;
  assign n25290 = n24929 & ~n25289;
  assign n25291 = n25287 & n25290;
  assign n25292 = ~n24940 & n25269;
  assign n25293 = n25267 & n25292;
  assign n25294 = ~n25291 & ~n25293;
  assign n25295 = n25044 & n25125;
  assign n25296 = ~n24940 & n25295;
  assign n25297 = n25290 & n25296;
  assign n25298 = n25294 & ~n25297;
  assign n25299 = ~n25285 & n25298;
  assign n25300 = n25283 & n25299;
  assign n25301 = n25275 & n25300;
  assign n25302 = n25212 & n25301;
  assign n25303 = n25194 & n25302;
  assign n25304 = n25136 & n25303;
  assign n25305 = n25074 & n25175;
  assign n25306 = n24940 & n25305;
  assign n25307 = n25198 & n25306;
  assign n25308 = n25074 & n25218;
  assign n25309 = ~n24940 & n25308;
  assign n25310 = n25246 & n25309;
  assign n25311 = ~n25307 & ~n25310;
  assign n25312 = ~n24940 & n25129;
  assign n25313 = n25060 & n25312;
  assign n25314 = n24940 & n25176;
  assign n25315 = n25060 & n25314;
  assign n25316 = ~n25313 & ~n25315;
  assign n25317 = ~n24940 & n25223;
  assign n25318 = n25060 & n25317;
  assign n25319 = n25026 & n25107;
  assign n25320 = ~n24940 & n25319;
  assign n25321 = n25060 & n25320;
  assign n25322 = ~n25318 & ~n25321;
  assign n25323 = n24940 & n25319;
  assign n25324 = n25060 & n25323;
  assign n25325 = n25322 & ~n25324;
  assign n25326 = n25316 & n25325;
  assign n25327 = ~n24940 & n25219;
  assign n25328 = n25060 & n25327;
  assign n25329 = n24940 & n25126;
  assign n25330 = n25060 & n25329;
  assign n25331 = ~n25328 & ~n25330;
  assign n25332 = ~n24941 & n25118;
  assign n25333 = n24982 & n25060;
  assign n25334 = n25043 & n25333;
  assign n25335 = n24970 & n25334;
  assign n25336 = ~n25332 & ~n25335;
  assign n25337 = ~n25015 & n25060;
  assign n25338 = n25107 & n25337;
  assign n25339 = n25073 & n25333;
  assign n25340 = n24970 & n25339;
  assign n25341 = ~n25338 & ~n25340;
  assign n25342 = n25336 & n25341;
  assign n25343 = n25331 & n25342;
  assign n25344 = n24985 & n25047;
  assign n25345 = n24940 & n25344;
  assign n25346 = n25060 & n25345;
  assign n25347 = n25138 & n25344;
  assign n25348 = ~n25346 & ~n25347;
  assign n25349 = n25343 & n25348;
  assign n25350 = n25326 & n25349;
  assign n25351 = n25311 & n25350;
  assign n25352 = n24940 & n25308;
  assign n25353 = n25251 & n25352;
  assign n25354 = n25074 & n25089;
  assign n25355 = ~n24940 & n25354;
  assign n25356 = n25165 & n25355;
  assign n25357 = ~n25353 & ~n25356;
  assign n25358 = n24940 & n25354;
  assign n25359 = n25149 & n25358;
  assign n25360 = ~n24940 & n25305;
  assign n25361 = n24932 & n25360;
  assign n25362 = ~n25359 & ~n25361;
  assign n25363 = n25357 & n25362;
  assign n25364 = n25351 & n25363;
  assign n25365 = n25304 & n25364;
  assign n25366 = n25094 & n25365;
  assign n25367 = n25051 & n25366;
  assign n25368 = n24888 & n24919;
  assign n25369 = ~po3872 & n25368;
  assign n25370 = pi0410 & ~pi0709;
  assign n25371 = n25369 & n25370;
  assign n25372 = ~n25367 & n25371;
  assign n25373 = n25198 & n25323;
  assign n25374 = n24932 & n25320;
  assign n25375 = ~n25373 & ~n25374;
  assign n25376 = n25254 & n25290;
  assign n25377 = n25032 & n25312;
  assign n25378 = ~n25376 & ~n25377;
  assign n25379 = n25086 & n25158;
  assign n25380 = n25084 & n25103;
  assign n25381 = ~n25379 & ~n25380;
  assign n25382 = n25091 & n25165;
  assign n25383 = n25070 & n25202;
  assign n25384 = ~n25382 & ~n25383;
  assign n25385 = ~n25064 & ~n25076;
  assign n25386 = n25041 & ~n25385;
  assign n25387 = n25078 & n25230;
  assign n25388 = ~n25386 & ~n25387;
  assign n25389 = n25342 & n25348;
  assign n25390 = n25246 & n25327;
  assign n25391 = n25151 & n25329;
  assign n25392 = ~n25390 & ~n25391;
  assign n25393 = n25389 & n25392;
  assign n25394 = n25388 & n25393;
  assign n25395 = n25384 & n25394;
  assign n25396 = n25381 & n25395;
  assign n25397 = n24932 & n25177;
  assign n25398 = n25396 & ~n25397;
  assign n25399 = n25122 & n25151;
  assign n25400 = ~n25128 & ~n25399;
  assign n25401 = ~n25119 & n25400;
  assign n25402 = n25130 & n25237;
  assign n25403 = n25401 & ~n25402;
  assign n25404 = n25110 & n25158;
  assign n25405 = n25114 & n25165;
  assign n25406 = ~n25404 & ~n25405;
  assign n25407 = n25403 & n25406;
  assign n25408 = n25103 & n25179;
  assign n25409 = n25142 & n25202;
  assign n25410 = ~n25408 & ~n25409;
  assign n25411 = ~n25139 & ~n25183;
  assign n25412 = n25410 & n25411;
  assign n25413 = n25407 & n25412;
  assign n25414 = n25398 & n25413;
  assign n25415 = pi3516 & ~n14997;
  assign n25416 = n25414 & ~n25415;
  assign n25417 = n25198 & n25314;
  assign n25418 = n25267 & n25276;
  assign n25419 = ~n25417 & ~n25418;
  assign n25420 = ~n25220 & ~n25224;
  assign n25421 = n25251 & ~n25420;
  assign n25422 = n25207 & n25267;
  assign n25423 = n25149 & n25213;
  assign n25424 = ~n25422 & ~n25423;
  assign n25425 = ~n25421 & n25424;
  assign n25426 = n25172 & n25290;
  assign n25427 = n25425 & ~n25426;
  assign n25428 = n25149 & n25215;
  assign n25429 = n25209 & n25230;
  assign n25430 = ~n25428 & ~n25429;
  assign n25431 = n25246 & n25317;
  assign n25432 = ~n25285 & ~n25431;
  assign n25433 = n25430 & n25432;
  assign n25434 = n25427 & n25433;
  assign n25435 = n25237 & n25257;
  assign n25436 = n25434 & ~n25435;
  assign n25437 = n25419 & n25436;
  assign n25438 = ~n25279 & n25437;
  assign n25439 = n25416 & n25438;
  assign n25440 = n25378 & n25439;
  assign n25441 = n25375 & n25440;
  assign n25442 = ~pi0410 & ~pi0710;
  assign n25443 = n25369 & n25442;
  assign n25444 = ~n25441 & n25443;
  assign n25445 = ~n25372 & ~n25444;
  assign n25446 = n24927 & n25445;
  assign n25447 = n24918 & n25446;
  assign n25448 = n24910 & n25447;
  assign n25449 = pi0341 & ~pi0343;
  assign n25450 = ~n16604 & n25449;
  assign n25451 = pi0341 & ~n24265;
  assign n25452 = pi0343 & n25451;
  assign n25453 = ~n25450 & ~n25452;
  assign n25454 = ~pi0342 & ~n25453;
  assign n25455 = pi0343 & ~n16604;
  assign n25456 = ~pi0343 & ~n15115;
  assign n25457 = ~n25455 & ~n25456;
  assign n25458 = ~pi0341 & ~pi0342;
  assign n25459 = ~n25457 & n25458;
  assign n25460 = ~n25454 & ~n25459;
  assign n25461 = po3872 & n19624;
  assign n25462 = ~pi3509 & n25461;
  assign n25463 = ~n14997 & n25462;
  assign n25464 = pi3509 & po3872;
  assign n25465 = n19624 & n25464;
  assign n25466 = ~n14993 & n25465;
  assign n25467 = ~n25463 & ~n25466;
  assign n25468 = n20515 & n24888;
  assign n25469 = ~po3872 & n24874;
  assign n25470 = ~n9498 & n25469;
  assign n25471 = n25468 & n25470;
  assign n25472 = ~po3872 & n24870;
  assign n25473 = ~n24888 & n25472;
  assign n25474 = po3872 & n19612;
  assign n25475 = ~n25473 & ~n25474;
  assign n25476 = ~n14913 & ~n25475;
  assign n25477 = ~n25471 & ~n25476;
  assign n25478 = n25468 & n25472;
  assign n25479 = n9498 & n25478;
  assign n25480 = ~po3872 & n24863;
  assign n25481 = ~n24888 & n25480;
  assign n25482 = po3872 & n19615;
  assign n25483 = ~n25481 & ~n25482;
  assign n25484 = ~n14917 & ~n25483;
  assign n25485 = ~n24888 & n25469;
  assign n25486 = po3872 & n19610;
  assign n25487 = ~n25485 & ~n25486;
  assign n25488 = ~n14891 & ~n25487;
  assign n25489 = ~n25484 & ~n25488;
  assign n25490 = n9498 & n25468;
  assign n25491 = n25480 & n25490;
  assign n25492 = n25489 & ~n25491;
  assign n25493 = ~n25479 & n25492;
  assign n25494 = n25477 & n25493;
  assign n25495 = ~pi0343 & ~n25494;
  assign n25496 = pi0343 & ~n15115;
  assign n25497 = ~n25495 & ~n25496;
  assign n25498 = ~pi0341 & pi0342;
  assign n25499 = ~n25497 & n25498;
  assign n25500 = n25467 & ~n25499;
  assign n25501 = n25460 & n25500;
  assign n25502 = n25448 & n25501;
  assign n25503 = ~pi0410 & pi0710;
  assign n25504 = pi0410 & pi0709;
  assign n25505 = ~n25503 & ~n25504;
  assign n25506 = n24888 & ~n25505;
  assign n25507 = n24920 & n25506;
  assign n25508 = pi3245 & n25507;
  assign n25509 = ~n16604 & n25508;
  assign n25510 = ~pi3245 & ~po3872;
  assign n25511 = n25506 & n25510;
  assign n25512 = n24919 & n25511;
  assign n25513 = ~n15115 & n25512;
  assign n25514 = ~n25509 & ~n25513;
  assign n25515 = n25502 & n25514;
  assign n25516 = ~n24827 & ~n24828;
  assign n25517 = ~po3872 & n24819;
  assign n25518 = ~n24832 & n25517;
  assign n25519 = n25516 & n25518;
  assign n25520 = ~pi0580 & ~pi3426;
  assign n25521 = ~n24835 & n25520;
  assign n25522 = ~pi0596 & ~pi3426;
  assign n25523 = n24835 & n25522;
  assign n25524 = ~n25521 & ~n25523;
  assign n25525 = n25519 & ~n25524;
  assign n25526 = pi0406 & pi0425;
  assign n25527 = ~po3872 & n25526;
  assign n25528 = pi3516 & pi3518;
  assign n25529 = po3872 & n25528;
  assign n25530 = ~n25527 & ~n25529;
  assign n25531 = ~n25525 & n25530;
  assign n25532 = n8561 & ~po3872;
  assign n25533 = ~pi2384 & ~n24819;
  assign n25534 = ~n25532 & ~n25533;
  assign n25535 = ~po3872 & n24826;
  assign n25536 = ~pi3130 & po3872;
  assign n25537 = ~n25535 & ~n25536;
  assign n25538 = ~pi0409 & ~pi0426;
  assign n25539 = ~po3872 & n25538;
  assign n25540 = po3872 & n19607;
  assign n25541 = ~n25539 & ~n25540;
  assign n25542 = ~n25537 & n25541;
  assign n25543 = n25534 & n25542;
  assign n25544 = n25531 & n25543;
  assign n25545 = ~n25515 & n25544;
  assign n25546 = ~pi0055 & n25533;
  assign n25547 = ~pi3245 & ~pi3344;
  assign n25548 = ~n8561 & ~n25547;
  assign n25549 = n25525 & n25548;
  assign n25550 = n25517 & n25538;
  assign n25551 = ~pi0597 & ~pi3426;
  assign n25552 = pi0410 & n25551;
  assign n25553 = n25550 & n25552;
  assign n25554 = ~pi0579 & ~pi3426;
  assign n25555 = n25517 & n25554;
  assign n25556 = ~pi0426 & n24869;
  assign n25557 = n25555 & n25556;
  assign n25558 = ~n25553 & ~n25557;
  assign n25559 = ~n25537 & ~n25558;
  assign n25560 = n25531 & n25559;
  assign n25561 = ~n25541 & n25560;
  assign n25562 = pi3245 & ~n25532;
  assign n25563 = n25561 & n25562;
  assign n25564 = ~n25549 & ~n25563;
  assign n25565 = ~pi0406 & ~po3872;
  assign n25566 = ~pi3518 & po3872;
  assign n25567 = ~n25565 & ~n25566;
  assign n25568 = ~n25525 & n25537;
  assign n25569 = n25530 & n25568;
  assign n25570 = ~n25532 & n25569;
  assign n25571 = n25567 & n25570;
  assign n25572 = ~pi0220 & pi0979;
  assign n25573 = ~pi0222 & ~pi0979;
  assign n25574 = ~n25572 & ~n25573;
  assign n25575 = n25571 & ~n25574;
  assign n25576 = ~n25532 & ~n25541;
  assign n25577 = ~n25537 & n25558;
  assign n25578 = ~n25525 & n25577;
  assign n25579 = n25530 & n25578;
  assign n25580 = n25576 & n25579;
  assign n25581 = pi0410 & ~po3872;
  assign n25582 = ~n25464 & ~n25581;
  assign n25583 = ~n14895 & ~n25582;
  assign n25584 = ~n14899 & n25582;
  assign n25585 = ~n25583 & ~n25584;
  assign n25586 = n25580 & ~n25585;
  assign n25587 = ~pi0055 & n25532;
  assign n25588 = ~n25586 & ~n25587;
  assign n25589 = n25537 & ~n25567;
  assign n25590 = n25531 & n25589;
  assign n25591 = ~n25532 & n25590;
  assign n25592 = pi0425 & ~po3872;
  assign n25593 = pi3516 & po3872;
  assign n25594 = ~n25592 & ~n25593;
  assign n25595 = n14904 & ~n25594;
  assign n25596 = n14908 & n25594;
  assign n25597 = ~n25595 & ~n25596;
  assign n25598 = n25591 & n25597;
  assign n25599 = n25588 & ~n25598;
  assign n25600 = ~n25575 & n25599;
  assign n25601 = ~pi3245 & n25525;
  assign n25602 = ~pi3344 & ~n8561;
  assign n25603 = n25601 & n25602;
  assign n25604 = ~pi3245 & ~n25532;
  assign n25605 = n25561 & n25604;
  assign n25606 = ~n25603 & ~n25605;
  assign n25607 = ~n25600 & n25606;
  assign n25608 = ~n15115 & ~n25606;
  assign n25609 = ~n25607 & ~n25608;
  assign n25610 = n25564 & ~n25609;
  assign n25611 = ~n16604 & n25606;
  assign n25612 = ~n25600 & ~n25606;
  assign n25613 = ~n25611 & ~n25612;
  assign n25614 = ~n25564 & ~n25613;
  assign n25615 = ~n25610 & ~n25614;
  assign n25616 = ~n25533 & ~n25615;
  assign n25617 = ~n25546 & ~n25616;
  assign n25618 = ~n25544 & ~n25617;
  assign po0325 = n25545 | n25618;
  assign n25620 = n25534 & n25541;
  assign n25621 = ~n25515 & n25620;
  assign n25622 = pi2384 & po3872;
  assign n25623 = ~n8561 & n24819;
  assign n25624 = ~n25622 & ~n25623;
  assign n25625 = ~n25533 & ~n25624;
  assign n25626 = pi0056 & ~n25625;
  assign n25627 = n25558 & ~n25585;
  assign n25628 = ~n24289 & ~n25558;
  assign n25629 = ~n25627 & ~n25628;
  assign n25630 = n25625 & ~n25629;
  assign n25631 = ~n25626 & ~n25630;
  assign n25632 = ~n25620 & ~n25631;
  assign po0326 = n25621 | n25632;
  assign n25634 = n24340 & ~n24482;
  assign n25635 = pi0057 & ~n24340;
  assign po0327 = n25634 | n25635;
  assign n25637 = ~n20518 & n20523;
  assign n25638 = ~n21228 & n21326;
  assign n25639 = n21228 & ~n21326;
  assign n25640 = ~n25638 & ~n25639;
  assign n25641 = n21230 & ~n21323;
  assign n25642 = ~n24099 & ~n24103;
  assign n25643 = n21547 & ~n25642;
  assign n25644 = ~n25641 & ~n25643;
  assign n25645 = ~n21552 & ~n25644;
  assign n25646 = ~n25640 & ~n25645;
  assign n25647 = n25640 & n25645;
  assign n25648 = ~n25646 & ~n25647;
  assign n25649 = ~pi0868 & n25648;
  assign n25650 = pi0868 & ~n24480;
  assign n25651 = ~n25649 & ~n25650;
  assign n25652 = n25637 & ~n25651;
  assign n25653 = pi0058 & ~n25637;
  assign n25654 = n20518 & n25653;
  assign n25655 = ~n25652 & ~n25654;
  assign n25656 = pi0058 & n24261;
  assign n25657 = ~n24267 & ~n25656;
  assign n25658 = ~n20518 & ~n25657;
  assign n25659 = ~n20518 & n24270;
  assign n25660 = ~n25658 & ~n25659;
  assign n25661 = ~n25637 & ~n25660;
  assign po0328 = ~n25655 | n25661;
  assign n25663 = ~n24300 & n24303;
  assign n25664 = ~n25651 & n25663;
  assign n25665 = pi0059 & ~n25663;
  assign n25666 = n24300 & n25665;
  assign n25667 = ~n25664 & ~n25666;
  assign n25668 = pi0059 & n24316;
  assign n25669 = ~n24319 & ~n25668;
  assign n25670 = ~n24300 & ~n25669;
  assign n25671 = ~n24300 & n24322;
  assign n25672 = ~n25670 & ~n25671;
  assign n25673 = ~n25663 & ~n25672;
  assign po0329 = ~n25667 | n25673;
  assign n25675 = n24340 & ~n24738;
  assign n25676 = pi0060 & ~n24340;
  assign po0330 = n25675 | n25676;
  assign n25678 = n24340 & ~n24763;
  assign n25679 = pi0061 & ~n24340;
  assign po0331 = n25678 | n25679;
  assign n25681 = pi0062 & ~n20524;
  assign n25682 = n20521 & n25681;
  assign n25683 = pi0868 & n24760;
  assign n25684 = ~n24656 & ~n24658;
  assign n25685 = ~n24186 & ~n24223;
  assign n25686 = ~n24243 & ~n25685;
  assign n25687 = n24186 & n24223;
  assign n25688 = ~n25686 & ~n25687;
  assign n25689 = ~n25684 & n25688;
  assign n25690 = n25684 & ~n25688;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = ~pi0868 & n25691;
  assign n25693 = ~n25683 & ~n25692;
  assign n25694 = n20524 & ~n25693;
  assign n25695 = ~n25682 & ~n25694;
  assign n25696 = pi0062 & ~n24252;
  assign n25697 = pi3245 & ~n16712;
  assign n25698 = ~pi3245 & ~n13988;
  assign n25699 = ~n25697 & ~n25698;
  assign n25700 = n24252 & ~n25699;
  assign n25701 = ~n25696 & ~n25700;
  assign n25702 = n24261 & ~n25701;
  assign n25703 = ~n24267 & ~n25702;
  assign n25704 = ~n20521 & ~n25703;
  assign n25705 = ~n24271 & ~n25704;
  assign n25706 = ~n20524 & ~n25705;
  assign po0332 = ~n25695 | n25706;
  assign n25708 = pi0063 & ~n20524;
  assign n25709 = n20521 & n25708;
  assign n25710 = pi0868 & n25691;
  assign n25711 = ~pi0868 & ~n24246;
  assign n25712 = ~n25710 & ~n25711;
  assign n25713 = n20524 & ~n25712;
  assign n25714 = ~n25709 & ~n25713;
  assign n25715 = pi0063 & ~n24252;
  assign n25716 = ~pi3245 & ~n12415;
  assign n25717 = pi3245 & ~n16676;
  assign n25718 = ~n25716 & ~n25717;
  assign n25719 = n24252 & ~n25718;
  assign n25720 = ~n25715 & ~n25719;
  assign n25721 = n24261 & ~n25720;
  assign n25722 = ~n24267 & ~n25721;
  assign n25723 = ~n20521 & ~n25722;
  assign n25724 = ~n24271 & ~n25723;
  assign n25725 = ~n20524 & ~n25724;
  assign po0333 = ~n25714 | n25725;
  assign n25727 = pi0064 & ~n24304;
  assign n25728 = n24302 & n25727;
  assign n25729 = n24304 & ~n25693;
  assign n25730 = ~n25728 & ~n25729;
  assign n25731 = pi0064 & ~n24310;
  assign n25732 = n24310 & ~n25699;
  assign n25733 = ~n25731 & ~n25732;
  assign n25734 = n24316 & ~n25733;
  assign n25735 = ~n24319 & ~n25734;
  assign n25736 = ~n24302 & ~n25735;
  assign n25737 = ~n24323 & ~n25736;
  assign n25738 = ~n24304 & ~n25737;
  assign po0334 = ~n25730 | n25738;
  assign n25740 = pi0065 & ~n24304;
  assign n25741 = n24302 & n25740;
  assign n25742 = n24304 & ~n25712;
  assign n25743 = ~n25741 & ~n25742;
  assign n25744 = pi0065 & ~n24310;
  assign n25745 = n24310 & ~n25718;
  assign n25746 = ~n25744 & ~n25745;
  assign n25747 = n24316 & ~n25746;
  assign n25748 = ~n24319 & ~n25747;
  assign n25749 = ~n24302 & ~n25748;
  assign n25750 = ~n24323 & ~n25749;
  assign n25751 = ~n24304 & ~n25750;
  assign po0335 = ~n25743 | n25751;
  assign n25753 = n20193 & n20379;
  assign n25754 = n20177 & n25753;
  assign n25755 = ~n20194 & ~n20234;
  assign n25756 = ~n20380 & n25755;
  assign n25757 = ~n25754 & ~n25756;
  assign n25758 = ~n20260 & ~n20334;
  assign n25759 = ~n25757 & ~n25758;
  assign n25760 = n25757 & n25758;
  assign n25761 = ~n25759 & ~n25760;
  assign n25762 = n24892 & ~n25761;
  assign n25763 = ~n11819 & ~n24905;
  assign n25764 = ~n25762 & ~n25763;
  assign n25765 = pi0343 & ~n12061;
  assign n25766 = ~n11929 & n25474;
  assign n25767 = ~n11933 & ~n25483;
  assign n25768 = ~n11929 & n25473;
  assign n25769 = ~n25767 & ~n25768;
  assign n25770 = ~n25491 & n25769;
  assign n25771 = ~n11947 & ~n25487;
  assign n25772 = n25770 & ~n25771;
  assign n25773 = ~n25479 & n25772;
  assign n25774 = ~n25471 & n25773;
  assign n25775 = ~n25766 & n25774;
  assign n25776 = ~pi0343 & ~n25775;
  assign n25777 = ~n25765 & ~n25776;
  assign n25778 = n25498 & ~n25777;
  assign n25779 = ~n16568 & n24913;
  assign n25780 = ~n12061 & n24916;
  assign n25781 = ~n25779 & ~n25780;
  assign n25782 = ~n25778 & n25781;
  assign n25783 = ~n24909 & n25782;
  assign n25784 = n25764 & n25783;
  assign n25785 = ~n11837 & n24922;
  assign n25786 = ~n11855 & n24925;
  assign n25787 = ~n25785 & ~n25786;
  assign n25788 = ~n11837 & n25462;
  assign n25789 = ~n11855 & n25465;
  assign n25790 = ~n25788 & ~n25789;
  assign n25791 = n25267 & n25323;
  assign n25792 = n25198 & n25320;
  assign n25793 = n25251 & n25317;
  assign n25794 = ~n25792 & ~n25793;
  assign n25795 = n25041 & n25209;
  assign n25796 = n25202 & n25276;
  assign n25797 = ~n25795 & ~n25796;
  assign n25798 = n24932 & n25215;
  assign n25799 = n25797 & ~n25798;
  assign n25800 = n25202 & n25207;
  assign n25801 = n25032 & n25220;
  assign n25802 = ~n25800 & ~n25801;
  assign n25803 = n25122 & n25246;
  assign n25804 = n25127 & n25151;
  assign n25805 = ~n25803 & ~n25804;
  assign n25806 = n25110 & n25165;
  assign n25807 = n25114 & n25149;
  assign n25808 = ~n25806 & ~n25807;
  assign n25809 = n25103 & n25130;
  assign n25810 = n25808 & ~n25809;
  assign n25811 = ~n25119 & n25810;
  assign n25812 = n25805 & n25811;
  assign n25813 = n25103 & n25257;
  assign n25814 = n24932 & n25213;
  assign n25815 = ~n25813 & ~n25814;
  assign n25816 = ~n25279 & ~n25285;
  assign n25817 = n25032 & n25224;
  assign n25818 = n25816 & ~n25817;
  assign n25819 = n25815 & n25818;
  assign n25820 = n25812 & n25819;
  assign n25821 = n25142 & n25230;
  assign n25822 = n25177 & n25198;
  assign n25823 = ~n25821 & ~n25822;
  assign n25824 = n25091 & n25149;
  assign n25825 = n25070 & n25230;
  assign n25826 = ~n25824 & ~n25825;
  assign n25827 = n25084 & n25158;
  assign n25828 = n25086 & n25165;
  assign n25829 = ~n25827 & ~n25828;
  assign n25830 = n25064 & n25290;
  assign n25831 = n25041 & n25078;
  assign n25832 = ~n25830 & ~n25831;
  assign n25833 = n25076 & n25290;
  assign n25834 = n25832 & ~n25833;
  assign n25835 = n25829 & n25834;
  assign n25836 = n25826 & n25835;
  assign n25837 = n25823 & n25836;
  assign n25838 = n25246 & n25329;
  assign n25839 = n25251 & n25327;
  assign n25840 = ~n25838 & ~n25839;
  assign n25841 = n25158 & n25179;
  assign n25842 = n25151 & n25182;
  assign n25843 = ~n25841 & ~n25842;
  assign n25844 = n25840 & n25843;
  assign n25845 = ~n25139 & n25844;
  assign n25846 = n25837 & n25845;
  assign n25847 = n25389 & n25846;
  assign n25848 = n25820 & n25847;
  assign n25849 = n25802 & n25848;
  assign n25850 = n25799 & n25849;
  assign n25851 = pi3516 & ~n11837;
  assign n25852 = n25850 & ~n25851;
  assign n25853 = n25237 & n25312;
  assign n25854 = n25267 & n25314;
  assign n25855 = ~n25853 & ~n25854;
  assign n25856 = n25852 & n25855;
  assign n25857 = n25794 & n25856;
  assign n25858 = ~n25791 & n25857;
  assign n25859 = n25443 & ~n25858;
  assign n25860 = n25097 & n25237;
  assign n25861 = n25100 & n25158;
  assign n25862 = ~n25860 & ~n25861;
  assign n25863 = n25189 & n25290;
  assign n25864 = n25144 & ~n25863;
  assign n25865 = n24932 & n25146;
  assign n25866 = n25153 & n25246;
  assign n25867 = ~n25865 & ~n25866;
  assign n25868 = n25267 & n25306;
  assign n25869 = n25251 & n25309;
  assign n25870 = ~n25868 & ~n25869;
  assign n25871 = n25349 & n25870;
  assign n25872 = n25867 & n25871;
  assign n25873 = n25864 & n25872;
  assign n25874 = n25158 & n25184;
  assign n25875 = n25181 & ~n25874;
  assign n25876 = n25028 & n25198;
  assign n25877 = n25036 & n25237;
  assign n25878 = ~n25876 & ~n25877;
  assign n25879 = n25049 & n25290;
  assign n25880 = n25878 & ~n25879;
  assign n25881 = n25094 & n25880;
  assign n25882 = ~n25183 & n25881;
  assign n25883 = n25875 & n25882;
  assign n25884 = n25873 & n25883;
  assign n25885 = n25202 & n25264;
  assign n25886 = n25032 & n25248;
  assign n25887 = ~n25885 & ~n25886;
  assign n25888 = n25243 & n25251;
  assign n25889 = n25887 & ~n25888;
  assign n25890 = n25041 & n25261;
  assign n25891 = n25202 & n25292;
  assign n25892 = ~n25890 & ~n25891;
  assign n25893 = n25151 & n25254;
  assign n25894 = n25230 & n25270;
  assign n25895 = ~n25893 & ~n25894;
  assign n25896 = n25892 & n25895;
  assign n25897 = ~n25258 & n25896;
  assign n25898 = n25889 & n25897;
  assign n25899 = n25160 & n25165;
  assign n25900 = n25149 & n25162;
  assign n25901 = ~n25899 & ~n25900;
  assign n25902 = n25151 & n25172;
  assign n25903 = n25169 & n25246;
  assign n25904 = ~n25902 & ~n25903;
  assign n25905 = n25195 & n25267;
  assign n25906 = n25204 & n25230;
  assign n25907 = ~n25905 & ~n25906;
  assign n25908 = n25904 & n25907;
  assign n25909 = n25211 & n25908;
  assign n25910 = n25901 & n25909;
  assign n25911 = n25898 & n25910;
  assign n25912 = n25103 & n25281;
  assign n25913 = n25280 & ~n25912;
  assign n25914 = n25041 & n25231;
  assign n25915 = n25227 & ~n25914;
  assign n25916 = n25103 & n25234;
  assign n25917 = n25165 & n25239;
  assign n25918 = ~n25916 & ~n25917;
  assign n25919 = n25915 & n25918;
  assign n25920 = ~n25285 & n25919;
  assign n25921 = n25913 & n25920;
  assign n25922 = n25911 & n25921;
  assign n25923 = n25884 & n25922;
  assign n25924 = n25862 & n25923;
  assign n25925 = n25134 & n25924;
  assign n25926 = n25032 & n25352;
  assign n25927 = n25149 & n25355;
  assign n25928 = ~n25926 & ~n25927;
  assign n25929 = n24932 & n25358;
  assign n25930 = n25198 & n25360;
  assign n25931 = ~n25929 & ~n25930;
  assign n25932 = n25326 & n25931;
  assign n25933 = n25928 & n25932;
  assign n25934 = n25925 & n25933;
  assign n25935 = pi3516 & ~n11855;
  assign n25936 = n25934 & ~n25935;
  assign n25937 = n25371 & ~n25936;
  assign n25938 = ~n25859 & ~n25937;
  assign n25939 = ~n16568 & n25508;
  assign n25940 = ~n12061 & n25512;
  assign n25941 = ~n25939 & ~n25940;
  assign n25942 = n25938 & n25941;
  assign n25943 = n25790 & n25942;
  assign n25944 = n25787 & n25943;
  assign n25945 = n25784 & n25944;
  assign n25946 = ~n16568 & n25449;
  assign n25947 = ~n25452 & ~n25946;
  assign n25948 = ~pi0342 & ~n25947;
  assign n25949 = pi0343 & ~n16568;
  assign n25950 = ~pi0343 & ~n12061;
  assign n25951 = ~n25949 & ~n25950;
  assign n25952 = n25458 & ~n25951;
  assign n25953 = ~n25948 & ~n25952;
  assign n25954 = n25945 & n25953;
  assign n25955 = n25544 & ~n25954;
  assign n25956 = pi0066 & n25533;
  assign n25957 = ~pi0213 & pi0979;
  assign n25958 = ~pi0214 & ~pi0979;
  assign n25959 = ~n25957 & ~n25958;
  assign n25960 = n25571 & ~n25959;
  assign n25961 = ~n11951 & ~n25582;
  assign n25962 = ~n11955 & n25582;
  assign n25963 = ~n25961 & ~n25962;
  assign n25964 = n25580 & ~n25963;
  assign n25965 = pi0066 & n25532;
  assign n25966 = ~n25964 & ~n25965;
  assign n25967 = n11938 & ~n25594;
  assign n25968 = n11942 & n25594;
  assign n25969 = ~n25967 & ~n25968;
  assign n25970 = n25591 & n25969;
  assign n25971 = n25966 & ~n25970;
  assign n25972 = ~n25960 & n25971;
  assign n25973 = n25606 & ~n25972;
  assign n25974 = ~n12061 & ~n25606;
  assign n25975 = ~n25973 & ~n25974;
  assign n25976 = n25564 & ~n25975;
  assign n25977 = ~n16568 & n25606;
  assign n25978 = ~n25606 & ~n25972;
  assign n25979 = ~n25977 & ~n25978;
  assign n25980 = ~n25564 & ~n25979;
  assign n25981 = ~n25976 & ~n25980;
  assign n25982 = ~n25533 & ~n25981;
  assign n25983 = ~n25956 & ~n25982;
  assign n25984 = ~n25544 & ~n25983;
  assign po0336 = n25955 | n25984;
  assign n25986 = n25620 & ~n25954;
  assign n25987 = pi0067 & ~n25625;
  assign n25988 = n25558 & ~n25963;
  assign n25989 = ~n24446 & ~n25558;
  assign n25990 = ~n25988 & ~n25989;
  assign n25991 = n25625 & ~n25990;
  assign n25992 = ~n25987 & ~n25991;
  assign n25993 = ~n25620 & ~n25992;
  assign po0337 = n25986 | n25993;
  assign n25995 = pi0068 & n20518;
  assign n25996 = pi0068 & ~n24259;
  assign n25997 = ~pi3245 & ~n14403;
  assign n25998 = pi3245 & ~n16891;
  assign n25999 = ~n25997 & ~n25998;
  assign n26000 = n24259 & ~n25999;
  assign n26001 = ~n25996 & ~n26000;
  assign n26002 = ~n20518 & ~n24260;
  assign n26003 = ~n26001 & n26002;
  assign n26004 = ~n25995 & ~n26003;
  assign n26005 = ~pi0051 & n24260;
  assign n26006 = ~n20518 & n26005;
  assign n26007 = n26004 & ~n26006;
  assign n26008 = ~n25637 & ~n26007;
  assign n26009 = ~n24091 & n24096;
  assign n26010 = n23286 & ~n26009;
  assign n26011 = n22762 & ~n26010;
  assign n26012 = n23300 & ~n26011;
  assign n26013 = n22109 & ~n26012;
  assign n26014 = ~n22104 & ~n26013;
  assign n26015 = ~n22105 & n26014;
  assign n26016 = ~n21675 & ~n21815;
  assign n26017 = ~n26015 & ~n26016;
  assign n26018 = n21675 & n21815;
  assign n26019 = ~n26017 & ~n26018;
  assign n26020 = n21680 & n21683;
  assign n26021 = ~n21680 & ~n21683;
  assign n26022 = ~n26020 & ~n26021;
  assign n26023 = n26019 & n26022;
  assign n26024 = ~n26019 & ~n26022;
  assign n26025 = ~n26023 & ~n26024;
  assign n26026 = pi0868 & n26025;
  assign n26027 = n21675 & ~n21815;
  assign n26028 = ~n21675 & n21815;
  assign n26029 = ~n26027 & ~n26028;
  assign n26030 = n26015 & ~n26029;
  assign n26031 = ~n26015 & n26029;
  assign n26032 = ~n26030 & ~n26031;
  assign n26033 = ~pi0868 & ~n26032;
  assign n26034 = ~n26026 & ~n26033;
  assign n26035 = n25637 & ~n26034;
  assign po0338 = n26008 | n26035;
  assign n26037 = pi0069 & n24300;
  assign n26038 = pi0069 & ~n24314;
  assign n26039 = n24314 & ~n25999;
  assign n26040 = ~n26038 & ~n26039;
  assign n26041 = ~n24300 & ~n24315;
  assign n26042 = ~n26040 & n26041;
  assign n26043 = ~n26037 & ~n26042;
  assign n26044 = ~pi0053 & n24315;
  assign n26045 = ~n24300 & n26044;
  assign n26046 = n26043 & ~n26045;
  assign n26047 = ~n25663 & ~n26046;
  assign n26048 = n25663 & ~n26034;
  assign po0339 = n26047 | n26048;
  assign n26050 = pi0979 & n20522;
  assign n26051 = ~pi1667 & n26050;
  assign n26052 = ~pi0070 & ~n26051;
  assign n26053 = ~n26034 & n26051;
  assign po0340 = n26052 | n26053;
  assign n26055 = ~pi1667 & n20522;
  assign n26056 = ~pi0979 & n26055;
  assign n26057 = ~pi0071 & ~n26056;
  assign n26058 = ~n26034 & n26056;
  assign po0341 = n26057 | n26058;
  assign n26060 = ~pi0734 & n9365;
  assign po3570 = pi3427 | n26060;
  assign n26062 = ~pi2555 & ~po3570;
  assign n26063 = ~pi2555 & ~n14816;
  assign n26064 = ~pi0072 & ~pi0330;
  assign n26065 = ~pi0073 & ~pi0127;
  assign n26066 = ~pi0128 & n26065;
  assign n26067 = ~pi0314 & ~pi0368;
  assign n26068 = n26066 & n26067;
  assign n26069 = n26064 & n26068;
  assign n26070 = ~pi1741 & ~pi1867;
  assign n26071 = ~pi1742 & ~pi1745;
  assign n26072 = n26070 & n26071;
  assign n26073 = n26069 & n26072;
  assign n26074 = pi1714 & ~n26073;
  assign n26075 = ~pi1714 & n26073;
  assign n26076 = ~n26074 & ~n26075;
  assign n26077 = pi1897 & n26076;
  assign n26078 = pi1714 & ~pi1897;
  assign n26079 = ~n26077 & ~n26078;
  assign n26080 = ~pi1741 & ~pi1742;
  assign n26081 = ~pi0368 & ~pi1867;
  assign n26082 = n26080 & n26081;
  assign n26083 = ~pi0072 & ~pi0127;
  assign n26084 = ~pi0073 & ~pi0128;
  assign n26085 = ~pi0314 & ~pi0330;
  assign n26086 = n26084 & n26085;
  assign n26087 = n26083 & n26086;
  assign n26088 = n26082 & n26087;
  assign n26089 = pi1745 & ~n26088;
  assign n26090 = ~pi1745 & n26088;
  assign n26091 = ~n26089 & ~n26090;
  assign n26092 = pi1897 & n26091;
  assign n26093 = pi1745 & ~pi1897;
  assign n26094 = ~n26092 & ~n26093;
  assign n26095 = n26064 & n26065;
  assign n26096 = n26067 & n26070;
  assign n26097 = n26095 & n26096;
  assign n26098 = ~pi0128 & n26097;
  assign n26099 = ~pi1742 & n26098;
  assign n26100 = pi1742 & ~n26098;
  assign n26101 = ~n26099 & ~n26100;
  assign n26102 = pi1897 & n26101;
  assign n26103 = pi1742 & ~pi1897;
  assign n26104 = ~n26102 & ~n26103;
  assign n26105 = ~n26094 & ~n26104;
  assign n26106 = ~pi1867 & n26069;
  assign n26107 = pi1867 & ~n26069;
  assign n26108 = ~n26106 & ~n26107;
  assign n26109 = pi1897 & n26108;
  assign n26110 = pi1867 & ~pi1897;
  assign n26111 = ~n26109 & ~n26110;
  assign n26112 = n26083 & n26084;
  assign n26113 = n26081 & n26085;
  assign n26114 = n26112 & n26113;
  assign n26115 = ~pi1741 & n26114;
  assign n26116 = pi1741 & ~n26114;
  assign n26117 = ~n26115 & ~n26116;
  assign n26118 = pi1897 & n26117;
  assign n26119 = pi1741 & ~pi1897;
  assign n26120 = ~n26118 & ~n26119;
  assign n26121 = ~n26111 & ~n26120;
  assign n26122 = pi0072 & ~n26066;
  assign n26123 = ~pi0072 & n26066;
  assign n26124 = ~n26122 & ~n26123;
  assign n26125 = pi1897 & n26124;
  assign n26126 = pi0072 & ~pi1897;
  assign n26127 = ~n26125 & ~n26126;
  assign n26128 = pi0330 & ~n26112;
  assign n26129 = ~pi0330 & n26112;
  assign n26130 = ~n26128 & ~n26129;
  assign n26131 = pi1897 & n26130;
  assign n26132 = pi0330 & ~pi1897;
  assign n26133 = ~n26131 & ~n26132;
  assign n26134 = ~n26127 & ~n26133;
  assign n26135 = pi0128 & ~pi1017;
  assign n26136 = pi0127 & ~n26084;
  assign n26137 = ~pi0127 & n26084;
  assign n26138 = ~n26136 & ~n26137;
  assign n26139 = pi1897 & n26138;
  assign n26140 = pi0127 & ~pi1897;
  assign n26141 = ~n26139 & ~n26140;
  assign n26142 = ~pi0073 & pi0128;
  assign n26143 = pi0073 & ~pi0128;
  assign n26144 = ~n26142 & ~n26143;
  assign n26145 = pi1897 & ~n26144;
  assign n26146 = pi0073 & ~pi1897;
  assign n26147 = ~n26145 & ~n26146;
  assign n26148 = ~n26141 & ~n26147;
  assign n26149 = n26135 & n26148;
  assign n26150 = n26134 & n26149;
  assign n26151 = ~pi0128 & n26095;
  assign n26152 = pi0314 & ~n26151;
  assign n26153 = ~pi0314 & n26151;
  assign n26154 = ~n26152 & ~n26153;
  assign n26155 = pi1897 & n26154;
  assign n26156 = pi0314 & ~pi1897;
  assign n26157 = ~n26155 & ~n26156;
  assign n26158 = pi1017 & n26157;
  assign n26159 = ~pi0368 & n26087;
  assign n26160 = pi0368 & ~n26087;
  assign n26161 = ~n26159 & ~n26160;
  assign n26162 = pi1897 & n26161;
  assign n26163 = pi0368 & ~pi1897;
  assign n26164 = ~n26162 & ~n26163;
  assign n26165 = ~n26158 & ~n26164;
  assign n26166 = n26150 & n26165;
  assign n26167 = ~pi1017 & ~n26157;
  assign n26168 = ~n26164 & n26167;
  assign n26169 = ~n26166 & ~n26168;
  assign n26170 = n26121 & ~n26169;
  assign n26171 = ~pi1714 & ~pi1745;
  assign n26172 = n26080 & n26171;
  assign n26173 = n26114 & n26172;
  assign n26174 = pi1744 & ~n26173;
  assign n26175 = ~pi1744 & n26173;
  assign n26176 = ~n26174 & ~n26175;
  assign n26177 = pi1897 & n26176;
  assign n26178 = pi1744 & ~pi1897;
  assign n26179 = ~n26177 & ~n26178;
  assign n26180 = n26170 & ~n26179;
  assign n26181 = n26105 & n26180;
  assign n26182 = ~n26079 & n26181;
  assign n26183 = ~n26094 & ~n26120;
  assign n26184 = ~n26111 & ~n26164;
  assign n26185 = n26135 & ~n26147;
  assign n26186 = ~n26141 & n26185;
  assign n26187 = ~n26127 & n26186;
  assign n26188 = ~n26133 & n26187;
  assign n26189 = ~n26158 & n26188;
  assign n26190 = ~n26167 & ~n26189;
  assign n26191 = n26184 & ~n26190;
  assign n26192 = ~n26104 & n26191;
  assign n26193 = ~n26079 & n26192;
  assign n26194 = n26183 & n26193;
  assign n26195 = ~n26179 & n26194;
  assign n26196 = n26179 & ~n26194;
  assign n26197 = ~n26195 & ~n26196;
  assign n26198 = pi1017 & n26197;
  assign n26199 = ~n26182 & ~n26198;
  assign n26200 = ~pi1714 & ~pi1744;
  assign n26201 = n26071 & n26096;
  assign n26202 = n26151 & n26201;
  assign n26203 = n26200 & n26202;
  assign n26204 = ~pi1743 & n26203;
  assign n26205 = pi1743 & ~n26203;
  assign n26206 = ~n26204 & ~n26205;
  assign n26207 = pi1897 & n26206;
  assign n26208 = pi1743 & ~pi1897;
  assign n26209 = ~n26207 & ~n26208;
  assign n26210 = ~pi1743 & ~pi1744;
  assign n26211 = n26082 & n26171;
  assign n26212 = n26087 & n26211;
  assign n26213 = n26210 & n26212;
  assign n26214 = ~pi1866 & n26213;
  assign n26215 = pi1866 & ~n26213;
  assign n26216 = ~n26214 & ~n26215;
  assign n26217 = pi1897 & n26216;
  assign n26218 = pi1866 & ~pi1897;
  assign n26219 = ~n26217 & ~n26218;
  assign n26220 = n26094 & n26104;
  assign n26221 = n26111 & n26120;
  assign n26222 = n26179 & n26219;
  assign n26223 = n26079 & n26209;
  assign n26224 = n26222 & n26223;
  assign n26225 = n26221 & n26224;
  assign n26226 = n26220 & n26225;
  assign n26227 = n26141 & n26147;
  assign n26228 = ~pi0128 & pi1897;
  assign n26229 = n26157 & n26164;
  assign n26230 = n26127 & n26133;
  assign n26231 = n26229 & n26230;
  assign n26232 = n26228 & n26231;
  assign n26233 = n26227 & n26232;
  assign n26234 = n26226 & n26233;
  assign n26235 = n26219 & ~n26234;
  assign n26236 = n26209 & n26235;
  assign n26237 = n26199 & n26236;
  assign n26238 = n26134 & ~n26141;
  assign n26239 = n26185 & n26238;
  assign n26240 = ~n26158 & n26239;
  assign n26241 = ~n26167 & ~n26240;
  assign n26242 = ~n26104 & ~n26241;
  assign n26243 = n26184 & n26242;
  assign n26244 = ~n26120 & n26243;
  assign n26245 = ~n26094 & n26244;
  assign n26246 = n26094 & ~n26244;
  assign n26247 = ~n26245 & ~n26246;
  assign n26248 = pi1017 & n26247;
  assign n26249 = n26105 & n26168;
  assign n26250 = n26121 & n26249;
  assign n26251 = n26105 & n26121;
  assign n26252 = n26165 & n26251;
  assign n26253 = n26134 & n26186;
  assign n26254 = n26252 & n26253;
  assign n26255 = ~n26250 & ~n26254;
  assign n26256 = n26079 & ~n26255;
  assign n26257 = ~n26079 & n26255;
  assign n26258 = ~n26256 & ~n26257;
  assign n26259 = ~pi1017 & ~n26258;
  assign n26260 = ~n26248 & ~n26259;
  assign n26261 = n26237 & n26260;
  assign n26262 = n26134 & n26165;
  assign n26263 = n26186 & n26262;
  assign n26264 = ~n26168 & ~n26263;
  assign n26265 = ~n26111 & n26264;
  assign n26266 = n26111 & ~n26264;
  assign n26267 = ~n26265 & ~n26266;
  assign n26268 = ~pi1017 & ~n26267;
  assign n26269 = n26164 & n26241;
  assign n26270 = ~n26164 & ~n26241;
  assign n26271 = ~n26269 & ~n26270;
  assign n26272 = pi1017 & n26271;
  assign n26273 = ~n26268 & ~n26272;
  assign n26274 = n26237 & n26273;
  assign n26275 = ~n26120 & ~n26191;
  assign n26276 = n26120 & n26191;
  assign n26277 = ~n26275 & ~n26276;
  assign n26278 = ~pi1017 & ~n26277;
  assign n26279 = pi1017 & ~n26267;
  assign n26280 = ~n26278 & ~n26279;
  assign n26281 = n26237 & n26280;
  assign n26282 = ~pi1017 & n26197;
  assign n26283 = pi1017 & ~n26258;
  assign n26284 = ~n26282 & ~n26283;
  assign n26285 = n26237 & n26284;
  assign n26286 = n26261 & n26285;
  assign n26287 = ~pi1017 & n26247;
  assign n26288 = n26104 & ~n26170;
  assign n26289 = ~n26104 & n26170;
  assign n26290 = ~n26288 & ~n26289;
  assign n26291 = pi1017 & n26290;
  assign n26292 = ~n26287 & ~n26291;
  assign n26293 = n26237 & n26292;
  assign n26294 = pi1017 & ~n26277;
  assign n26295 = ~pi1017 & n26290;
  assign n26296 = ~n26294 & ~n26295;
  assign n26297 = n26237 & n26296;
  assign n26298 = n26293 & n26297;
  assign n26299 = n26286 & n26298;
  assign n26300 = n26281 & n26299;
  assign n26301 = n26274 & n26300;
  assign n26302 = n26286 & ~n26299;
  assign n26303 = ~n26301 & ~n26302;
  assign n26304 = ~n26158 & ~n26167;
  assign n26305 = n26150 & n26304;
  assign n26306 = ~n26150 & ~n26304;
  assign n26307 = ~n26305 & ~n26306;
  assign n26308 = pi1017 & n26307;
  assign n26309 = ~pi1017 & n26271;
  assign n26310 = ~n26308 & ~n26309;
  assign n26311 = n26237 & ~n26310;
  assign n26312 = n26133 & ~n26187;
  assign n26313 = ~n26188 & ~n26312;
  assign n26314 = pi1017 & n26313;
  assign n26315 = ~pi1017 & n26307;
  assign n26316 = ~n26314 & ~n26315;
  assign n26317 = n26237 & ~n26316;
  assign n26318 = ~n26311 & ~n26317;
  assign n26319 = n26281 & n26318;
  assign n26320 = n26274 & n26319;
  assign n26321 = n26299 & n26320;
  assign n26322 = n26303 & ~n26321;
  assign n26323 = n26293 & ~n26297;
  assign n26324 = n26286 & n26323;
  assign n26325 = ~n26261 & n26285;
  assign n26326 = ~n26324 & ~n26325;
  assign n26327 = ~n26299 & ~n26326;
  assign n26328 = ~n26311 & n26317;
  assign n26329 = n26274 & ~n26328;
  assign n26330 = n26300 & ~n26329;
  assign n26331 = ~n26327 & ~n26330;
  assign n26332 = ~n26321 & n26331;
  assign n26333 = ~n26299 & n26332;
  assign n26334 = n26322 & n26333;
  assign n26335 = pi1017 & n26299;
  assign n26336 = ~n26322 & ~n26332;
  assign n26337 = ~n26320 & ~n26336;
  assign n26338 = n26335 & ~n26337;
  assign n26339 = n26334 & ~n26338;
  assign n26340 = n26261 & n26339;
  assign n26341 = ~n26317 & n26338;
  assign n26342 = ~n26340 & ~n26341;
  assign n26343 = ~n26299 & ~n26332;
  assign n26344 = n26322 & n26343;
  assign n26345 = ~n26334 & n26344;
  assign n26346 = n26293 & n26345;
  assign n26347 = ~n26322 & n26333;
  assign n26348 = n26297 & n26347;
  assign n26349 = ~n26322 & n26343;
  assign n26350 = n26281 & n26349;
  assign n26351 = n26299 & n26332;
  assign n26352 = n26322 & n26351;
  assign n26353 = n26274 & n26352;
  assign n26354 = n26299 & n26322;
  assign n26355 = ~n26332 & n26354;
  assign n26356 = ~n26311 & n26355;
  assign n26357 = ~n26322 & n26351;
  assign n26358 = ~n26317 & n26357;
  assign n26359 = n26127 & ~n26186;
  assign n26360 = ~n26187 & ~n26359;
  assign n26361 = pi1017 & n26360;
  assign n26362 = ~pi1017 & n26313;
  assign n26363 = ~n26361 & ~n26362;
  assign n26364 = n26237 & ~n26363;
  assign n26365 = ~n26357 & ~n26364;
  assign n26366 = ~n26358 & ~n26365;
  assign n26367 = ~n26355 & ~n26366;
  assign n26368 = ~n26356 & ~n26367;
  assign n26369 = ~n26352 & ~n26368;
  assign n26370 = ~n26353 & ~n26369;
  assign n26371 = ~n26349 & ~n26370;
  assign n26372 = ~n26350 & ~n26371;
  assign n26373 = ~n26347 & ~n26372;
  assign n26374 = ~n26348 & ~n26373;
  assign n26375 = ~n26334 & ~n26344;
  assign n26376 = ~n26374 & n26375;
  assign n26377 = ~n26346 & ~n26376;
  assign n26378 = ~n26338 & ~n26377;
  assign n26379 = n26342 & ~n26378;
  assign n26380 = pi1017 & n26379;
  assign n26381 = ~pi1017 & ~n26379;
  assign n26382 = ~n26380 & ~n26381;
  assign n26383 = pi2555 & ~n26382;
  assign n26384 = ~n26063 & ~n26383;
  assign n26385 = ~n26062 & ~n26384;
  assign n26386 = pi0072 & n26062;
  assign po0342 = n26385 | n26386;
  assign n26388 = ~pi2555 & ~n12061;
  assign n26389 = n26297 & n26339;
  assign n26390 = n26141 & ~n26185;
  assign n26391 = ~n26186 & ~n26390;
  assign n26392 = pi1017 & n26391;
  assign n26393 = ~pi1017 & n26360;
  assign n26394 = ~n26392 & ~n26393;
  assign n26395 = n26237 & ~n26394;
  assign n26396 = n26338 & ~n26395;
  assign n26397 = ~n26389 & ~n26396;
  assign n26398 = n26281 & n26345;
  assign n26399 = n26274 & n26347;
  assign n26400 = ~n26311 & n26349;
  assign n26401 = ~n26317 & n26352;
  assign n26402 = n26355 & ~n26364;
  assign n26403 = n26357 & ~n26395;
  assign n26404 = ~n26135 & n26147;
  assign n26405 = ~n26185 & ~n26404;
  assign n26406 = pi1017 & n26405;
  assign n26407 = ~pi1017 & n26391;
  assign n26408 = ~n26406 & ~n26407;
  assign n26409 = n26237 & ~n26408;
  assign n26410 = ~n26357 & ~n26409;
  assign n26411 = ~n26403 & ~n26410;
  assign n26412 = ~n26355 & ~n26411;
  assign n26413 = ~n26402 & ~n26412;
  assign n26414 = ~n26352 & ~n26413;
  assign n26415 = ~n26401 & ~n26414;
  assign n26416 = ~n26349 & ~n26415;
  assign n26417 = ~n26400 & ~n26416;
  assign n26418 = ~n26347 & ~n26417;
  assign n26419 = ~n26399 & ~n26418;
  assign n26420 = n26375 & ~n26419;
  assign n26421 = ~n26398 & ~n26420;
  assign n26422 = ~n26338 & ~n26421;
  assign n26423 = n26397 & ~n26422;
  assign n26424 = pi1017 & n26423;
  assign n26425 = ~pi1017 & ~n26423;
  assign n26426 = ~n26424 & ~n26425;
  assign n26427 = pi2555 & ~n26426;
  assign n26428 = ~n26388 & ~n26427;
  assign n26429 = ~n26062 & ~n26428;
  assign n26430 = pi0073 & n26062;
  assign po0343 = n26429 | n26430;
  assign n26432 = n24932 & n25231;
  assign n26433 = n25227 & ~n26432;
  assign n26434 = n25151 & n25234;
  assign n26435 = n25239 & n25251;
  assign n26436 = ~n26434 & ~n26435;
  assign n26437 = n25044 & n25218;
  assign n26438 = ~n24940 & n26437;
  assign n26439 = n25230 & n26438;
  assign n26440 = n25103 & n25360;
  assign n26441 = ~n26439 & ~n26440;
  assign n26442 = n25032 & n25355;
  assign n26443 = n25237 & n25358;
  assign n26444 = ~n26442 & ~n26443;
  assign n26445 = n25146 & n25237;
  assign n26446 = n25181 & ~n26445;
  assign n26447 = ~n25183 & n26446;
  assign n26448 = n24940 & n26437;
  assign n26449 = n25041 & n26448;
  assign n26450 = n26447 & ~n26449;
  assign n26451 = n25189 & n25198;
  assign n26452 = n25034 & n25074;
  assign n26453 = ~n24940 & n26452;
  assign n26454 = n25290 & n26453;
  assign n26455 = ~n26451 & ~n26454;
  assign n26456 = n25074 & n25222;
  assign n26457 = ~n24940 & n26456;
  assign n26458 = n25230 & n26457;
  assign n26459 = n24940 & n25286;
  assign n26460 = n25202 & n26459;
  assign n26461 = ~n26458 & ~n26460;
  assign n26462 = n24940 & n26456;
  assign n26463 = n25041 & n26462;
  assign n26464 = n26461 & ~n26463;
  assign n26465 = n25036 & n25060;
  assign n26466 = ~n25092 & ~n26465;
  assign n26467 = n25080 & n26466;
  assign n26468 = n26464 & n26467;
  assign n26469 = n26455 & n26468;
  assign n26470 = n26450 & n26469;
  assign n26471 = ~n25071 & ~n25087;
  assign n26472 = n25060 & n25153;
  assign n26473 = n26471 & ~n26472;
  assign n26474 = ~n25085 & n26473;
  assign n26475 = n26470 & n26474;
  assign n26476 = n25060 & n25352;
  assign n26477 = ~n25324 & ~n26476;
  assign n26478 = n25322 & n26477;
  assign n26479 = ~n25315 & n26478;
  assign n26480 = ~n25313 & n26479;
  assign n26481 = n25060 & n25309;
  assign n26482 = n25348 & ~n26481;
  assign n26483 = n25158 & n25306;
  assign n26484 = n26482 & ~n26483;
  assign n26485 = n25060 & n25097;
  assign n26486 = n25133 & ~n26485;
  assign n26487 = n25116 & n26486;
  assign n26488 = n25100 & n25246;
  assign n26489 = n26487 & ~n26488;
  assign n26490 = n25343 & n26489;
  assign n26491 = n26484 & n26490;
  assign n26492 = n26480 & n26491;
  assign n26493 = n26475 & n26492;
  assign n26494 = n26444 & n26493;
  assign n26495 = n26441 & n26494;
  assign n26496 = n25184 & n25246;
  assign n26497 = n25049 & n25198;
  assign n26498 = n25028 & n25103;
  assign n26499 = ~n26497 & ~n26498;
  assign n26500 = ~n25065 & n25144;
  assign n26501 = n26499 & n26500;
  assign n26502 = ~n26496 & n26501;
  assign n26503 = n26495 & n26502;
  assign n26504 = pi3516 & ~n13293;
  assign n26505 = n26503 & ~n26504;
  assign n26506 = n25060 & n25169;
  assign n26507 = ~n25173 & ~n26506;
  assign n26508 = n25149 & n25204;
  assign n26509 = n25211 & ~n26508;
  assign n26510 = n26507 & n26509;
  assign n26511 = n25158 & n25195;
  assign n26512 = n26510 & ~n26511;
  assign n26513 = n25160 & n25251;
  assign n26514 = n25032 & n25162;
  assign n26515 = ~n26513 & ~n26514;
  assign n26516 = n25165 & n25264;
  assign n26517 = n25149 & n25270;
  assign n26518 = ~n26516 & ~n26517;
  assign n26519 = n24940 & n25295;
  assign n26520 = n25202 & n26519;
  assign n26521 = n24932 & n25261;
  assign n26522 = ~n26520 & ~n26521;
  assign n26523 = n26518 & n26522;
  assign n26524 = n25060 & n25248;
  assign n26525 = ~n25258 & ~n26524;
  assign n26526 = n25060 & n25243;
  assign n26527 = ~n25255 & ~n26526;
  assign n26528 = n26525 & n26527;
  assign n26529 = n26523 & n26528;
  assign n26530 = n26515 & n26529;
  assign n26531 = n26512 & n26530;
  assign n26532 = n26505 & n26531;
  assign n26533 = n25151 & n25281;
  assign n26534 = n25237 & n25278;
  assign n26535 = ~n26533 & ~n26534;
  assign n26536 = ~n25277 & ~n25285;
  assign n26537 = n25044 & n25095;
  assign n26538 = ~n24940 & n26537;
  assign n26539 = n25290 & n26538;
  assign n26540 = n25267 & n25296;
  assign n26541 = ~n26539 & ~n26540;
  assign n26542 = n25267 & n25287;
  assign n26543 = n25165 & n25292;
  assign n26544 = ~n26542 & ~n26543;
  assign n26545 = n26541 & n26544;
  assign n26546 = n26536 & n26545;
  assign n26547 = n26535 & n26546;
  assign n26548 = n26532 & n26547;
  assign n26549 = n26436 & n26548;
  assign n26550 = n26433 & n26549;
  assign n26551 = n25371 & ~n26550;
  assign n26552 = n25153 & n25202;
  assign n26553 = n25142 & n25149;
  assign n26554 = ~n26552 & ~n26553;
  assign n26555 = n25103 & n25177;
  assign n26556 = n26554 & ~n26555;
  assign n26557 = n25179 & n25246;
  assign n26558 = n26556 & ~n26557;
  assign n26559 = n25110 & n25251;
  assign n26560 = n25032 & n25114;
  assign n26561 = ~n26559 & ~n26560;
  assign n26562 = n25124 & ~n25128;
  assign n26563 = pi3516 & ~n13297;
  assign n26564 = n25097 & n25290;
  assign n26565 = n25130 & n25151;
  assign n26566 = ~n26564 & ~n26565;
  assign n26567 = ~n26563 & n26566;
  assign n26568 = n26562 & n26567;
  assign n26569 = n26561 & n26568;
  assign n26570 = n25215 & n25237;
  assign n26571 = n24932 & n25209;
  assign n26572 = ~n26570 & ~n26571;
  assign n26573 = n25172 & n25267;
  assign n26574 = n25169 & n25202;
  assign n26575 = ~n26573 & ~n26574;
  assign n26576 = n25165 & n25207;
  assign n26577 = n25213 & n25237;
  assign n26578 = ~n26576 & ~n26577;
  assign n26579 = n26575 & n26578;
  assign n26580 = n25226 & n26579;
  assign n26581 = n26572 & n26580;
  assign n26582 = n25151 & n25257;
  assign n26583 = n25165 & n25276;
  assign n26584 = ~n26582 & ~n26583;
  assign n26585 = n25230 & n25243;
  assign n26586 = n25041 & n25248;
  assign n26587 = ~n26585 & ~n26586;
  assign n26588 = n25254 & n25267;
  assign n26589 = n26587 & ~n26588;
  assign n26590 = n25816 & n26589;
  assign n26591 = n26584 & n26590;
  assign n26592 = n26581 & n26591;
  assign n26593 = n25041 & n25352;
  assign n26594 = n25158 & n25314;
  assign n26595 = ~n26593 & ~n26594;
  assign n26596 = n25158 & n25323;
  assign n26597 = n25103 & n25320;
  assign n26598 = ~n26596 & ~n26597;
  assign n26599 = ~n25313 & ~n25318;
  assign n26600 = n26598 & n26599;
  assign n26601 = n26595 & n26600;
  assign n26602 = n26592 & n26601;
  assign n26603 = n25230 & n25309;
  assign n26604 = n26602 & ~n26603;
  assign n26605 = n25343 & n26604;
  assign n26606 = n25348 & n26605;
  assign n26607 = n26569 & n26606;
  assign n26608 = n25064 & n25198;
  assign n26609 = n25036 & n25290;
  assign n26610 = ~n26608 & ~n26609;
  assign n26611 = n25084 & n25246;
  assign n26612 = n25086 & n25251;
  assign n26613 = ~n26611 & ~n26612;
  assign n26614 = n25076 & n25198;
  assign n26615 = n24932 & n25078;
  assign n26616 = ~n26614 & ~n26615;
  assign n26617 = n25032 & n25091;
  assign n26618 = n25070 & n25149;
  assign n26619 = ~n26617 & ~n26618;
  assign n26620 = n26616 & n26619;
  assign n26621 = n26613 & n26620;
  assign n26622 = n26610 & n26621;
  assign n26623 = n26607 & n26622;
  assign n26624 = n25411 & n26623;
  assign n26625 = n26558 & n26624;
  assign n26626 = n25443 & ~n26625;
  assign n26627 = ~n26551 & ~n26626;
  assign n26628 = ~n16748 & n25508;
  assign n26629 = ~n13398 & n25512;
  assign n26630 = ~n26628 & ~n26629;
  assign n26631 = n26627 & n26630;
  assign n26632 = ~n13297 & n24922;
  assign n26633 = ~n13293 & n24925;
  assign n26634 = ~n26632 & ~n26633;
  assign n26635 = ~n13297 & n25462;
  assign n26636 = ~n13293 & n25465;
  assign n26637 = ~n26635 & ~n26636;
  assign n26638 = n26634 & n26637;
  assign n26639 = ~n16748 & n25449;
  assign n26640 = ~n25452 & ~n26639;
  assign n26641 = ~pi0342 & ~n26640;
  assign n26642 = pi0343 & ~n16748;
  assign n26643 = ~pi0343 & ~n13398;
  assign n26644 = ~n26642 & ~n26643;
  assign n26645 = n25458 & ~n26644;
  assign n26646 = ~n26641 & ~n26645;
  assign n26647 = ~n20316 & ~n20334;
  assign n26648 = n20318 & n20379;
  assign n26649 = ~n20030 & ~n20318;
  assign n26650 = ~n20380 & n26649;
  assign n26651 = ~n26648 & ~n26650;
  assign n26652 = n26647 & n26651;
  assign n26653 = ~n26647 & ~n26651;
  assign n26654 = ~n26652 & ~n26653;
  assign n26655 = n24892 & ~n26654;
  assign n26656 = ~n13173 & ~n24905;
  assign n26657 = ~n16748 & n24913;
  assign n26658 = ~n13398 & n24916;
  assign n26659 = ~n26657 & ~n26658;
  assign n26660 = ~n24909 & n26659;
  assign n26661 = ~n26656 & n26660;
  assign n26662 = ~n26655 & n26661;
  assign n26663 = ~n13204 & n25474;
  assign n26664 = ~n13208 & ~n25483;
  assign n26665 = ~n26663 & ~n26664;
  assign n26666 = ~n25479 & n26665;
  assign n26667 = ~n25491 & n26666;
  assign n26668 = ~n25471 & n26667;
  assign n26669 = ~n13182 & ~n25487;
  assign n26670 = ~n13204 & n25473;
  assign n26671 = ~n26669 & ~n26670;
  assign n26672 = n26668 & n26671;
  assign n26673 = ~pi0343 & ~n26672;
  assign n26674 = pi0343 & ~n13398;
  assign n26675 = ~n26673 & ~n26674;
  assign n26676 = n25498 & ~n26675;
  assign n26677 = n26662 & ~n26676;
  assign n26678 = n26646 & n26677;
  assign n26679 = n26638 & n26678;
  assign n26680 = n26631 & n26679;
  assign n26681 = n25544 & ~n26680;
  assign n26682 = ~pi0074 & n25533;
  assign n26683 = ~pi0132 & pi0979;
  assign n26684 = ~pi0133 & ~pi0979;
  assign n26685 = ~n26683 & ~n26684;
  assign n26686 = n25571 & ~n26685;
  assign n26687 = ~n13186 & ~n25582;
  assign n26688 = ~n13190 & n25582;
  assign n26689 = ~n26687 & ~n26688;
  assign n26690 = n25580 & ~n26689;
  assign n26691 = ~pi0074 & n25532;
  assign n26692 = ~n26690 & ~n26691;
  assign n26693 = n13195 & ~n25594;
  assign n26694 = n13199 & n25594;
  assign n26695 = ~n26693 & ~n26694;
  assign n26696 = n25591 & n26695;
  assign n26697 = n26692 & ~n26696;
  assign n26698 = ~n26686 & n26697;
  assign n26699 = n25606 & ~n26698;
  assign n26700 = ~n13398 & ~n25606;
  assign n26701 = ~n26699 & ~n26700;
  assign n26702 = n25564 & ~n26701;
  assign n26703 = ~n16748 & n25606;
  assign n26704 = ~n25606 & ~n26698;
  assign n26705 = ~n26703 & ~n26704;
  assign n26706 = ~n25564 & ~n26705;
  assign n26707 = ~n26702 & ~n26706;
  assign n26708 = ~n25533 & ~n26707;
  assign n26709 = ~n26682 & ~n26708;
  assign n26710 = ~n25544 & ~n26709;
  assign po0344 = n26681 | n26710;
  assign n26712 = n25230 & n26519;
  assign n26713 = n25198 & n25261;
  assign n26714 = ~n26712 & ~n26713;
  assign n26715 = n25149 & n25264;
  assign n26716 = n24932 & n25270;
  assign n26717 = ~n26715 & ~n26716;
  assign n26718 = ~n25287 & ~n25296;
  assign n26719 = n25202 & ~n26718;
  assign n26720 = n25149 & n25292;
  assign n26721 = ~n26719 & ~n26720;
  assign n26722 = n25165 & n25306;
  assign n26723 = n25343 & ~n26722;
  assign n26724 = n26482 & n26723;
  assign n26725 = n26528 & n26724;
  assign n26726 = n26721 & n26725;
  assign n26727 = n26717 & n26726;
  assign n26728 = n26714 & n26727;
  assign n26729 = n25097 & n25151;
  assign n26730 = n25100 & n25251;
  assign n26731 = ~n26729 & ~n26730;
  assign n26732 = n24932 & n25204;
  assign n26733 = n25211 & ~n26732;
  assign n26734 = n26507 & n26733;
  assign n26735 = n25165 & n25195;
  assign n26736 = n26734 & ~n26735;
  assign n26737 = n25032 & n25160;
  assign n26738 = n25162 & n25237;
  assign n26739 = ~n26737 & ~n26738;
  assign n26740 = n25041 & n26438;
  assign n26741 = n25158 & n25360;
  assign n26742 = ~n26740 & ~n26741;
  assign n26743 = n25237 & n25355;
  assign n26744 = n25103 & n25358;
  assign n26745 = ~n26743 & ~n26744;
  assign n26746 = n26742 & n26745;
  assign n26747 = n26739 & n26746;
  assign n26748 = n26736 & n26747;
  assign n26749 = ~n25183 & ~n26472;
  assign n26750 = n25184 & n25251;
  assign n26751 = n26749 & ~n26750;
  assign n26752 = n25181 & n26751;
  assign n26753 = n25290 & n26448;
  assign n26754 = n26752 & ~n26753;
  assign n26755 = n25036 & n25151;
  assign n26756 = n25080 & ~n26755;
  assign n26757 = n25049 & n25267;
  assign n26758 = n25290 & n26462;
  assign n26759 = ~n26757 & ~n26758;
  assign n26760 = n25230 & n26459;
  assign n26761 = n25041 & n26457;
  assign n26762 = ~n26760 & ~n26761;
  assign n26763 = n26759 & n26762;
  assign n26764 = ~n25092 & n26763;
  assign n26765 = n26756 & n26764;
  assign n26766 = n25189 & n25267;
  assign n26767 = n25103 & n25146;
  assign n26768 = ~n26766 & ~n26767;
  assign n26769 = n25144 & n26768;
  assign n26770 = n26765 & n26769;
  assign n26771 = n26754 & n26770;
  assign n26772 = n25028 & n25158;
  assign n26773 = n26771 & ~n26772;
  assign n26774 = n25072 & n25088;
  assign n26775 = n26773 & n26774;
  assign n26776 = n26480 & n26775;
  assign n26777 = n26748 & n26776;
  assign n26778 = n26731 & n26777;
  assign n26779 = n25134 & n26778;
  assign n26780 = pi3516 & ~n13790;
  assign n26781 = n25198 & n25231;
  assign n26782 = n25227 & ~n26781;
  assign n26783 = n25234 & n25246;
  assign n26784 = n25032 & n25239;
  assign n26785 = ~n26783 & ~n26784;
  assign n26786 = n25246 & n25281;
  assign n26787 = n25103 & n25278;
  assign n26788 = ~n26786 & ~n26787;
  assign n26789 = n26536 & n26788;
  assign n26790 = n26785 & n26789;
  assign n26791 = n26782 & n26790;
  assign n26792 = ~n26780 & n26791;
  assign n26793 = n26779 & n26792;
  assign n26794 = n26728 & n26793;
  assign n26795 = n25371 & ~n26794;
  assign n26796 = n25158 & n25320;
  assign n26797 = n25151 & n25312;
  assign n26798 = ~n26796 & ~n26797;
  assign n26799 = n25267 & ~n25385;
  assign n26800 = n25078 & n25198;
  assign n26801 = ~n26799 & ~n26800;
  assign n26802 = ~n25314 & ~n25323;
  assign n26803 = n25165 & ~n26802;
  assign n26804 = n25290 & n25352;
  assign n26805 = ~n26803 & ~n26804;
  assign n26806 = n26801 & n26805;
  assign n26807 = ~n25318 & n26806;
  assign n26808 = n26798 & n26807;
  assign n26809 = n25149 & n25207;
  assign n26810 = n25103 & n25213;
  assign n26811 = ~n26809 & ~n26810;
  assign n26812 = n25172 & n25202;
  assign n26813 = n25169 & n25230;
  assign n26814 = ~n26812 & ~n26813;
  assign n26815 = n25153 & n25230;
  assign n26816 = n25158 & n25177;
  assign n26817 = ~n26815 & ~n26816;
  assign n26818 = n24932 & n25142;
  assign n26819 = n26817 & ~n26818;
  assign n26820 = n25179 & n25251;
  assign n26821 = n26819 & ~n26820;
  assign n26822 = n26814 & n26821;
  assign n26823 = n25411 & n26822;
  assign n26824 = n25041 & n25309;
  assign n26825 = n25348 & ~n26824;
  assign n26826 = n25114 & n25237;
  assign n26827 = n25032 & n25110;
  assign n26828 = ~n26826 & ~n26827;
  assign n26829 = n25342 & n26828;
  assign n26830 = n25331 & n26829;
  assign n26831 = n26825 & n26830;
  assign n26832 = n25130 & n25246;
  assign n26833 = n26831 & ~n26832;
  assign n26834 = n26562 & n26833;
  assign n26835 = n26823 & n26834;
  assign n26836 = n25198 & n25209;
  assign n26837 = n25103 & n25215;
  assign n26838 = ~n26836 & ~n26837;
  assign n26839 = n26835 & n26838;
  assign n26840 = n25226 & n26839;
  assign n26841 = n26811 & n26840;
  assign n26842 = pi3516 & ~n13794;
  assign n26843 = n25246 & n25257;
  assign n26844 = n25149 & n25276;
  assign n26845 = ~n26843 & ~n26844;
  assign n26846 = n25816 & n26845;
  assign n26847 = n25202 & n25254;
  assign n26848 = n26846 & ~n26847;
  assign n26849 = n25041 & n25243;
  assign n26850 = n25248 & n25290;
  assign n26851 = ~n26849 & ~n26850;
  assign n26852 = n25084 & n25251;
  assign n26853 = n25032 & n25086;
  assign n26854 = ~n26852 & ~n26853;
  assign n26855 = n25091 & n25237;
  assign n26856 = n24932 & n25070;
  assign n26857 = ~n26855 & ~n26856;
  assign n26858 = n26854 & n26857;
  assign n26859 = n26851 & n26858;
  assign n26860 = n26848 & n26859;
  assign n26861 = ~n26842 & n26860;
  assign n26862 = n26841 & n26861;
  assign n26863 = n26808 & n26862;
  assign n26864 = n25443 & ~n26863;
  assign n26865 = ~n26795 & ~n26864;
  assign n26866 = ~n16712 & n25508;
  assign n26867 = ~n13988 & n25512;
  assign n26868 = ~n26866 & ~n26867;
  assign n26869 = n26865 & n26868;
  assign n26870 = ~n13794 & n24922;
  assign n26871 = ~n13790 & n24925;
  assign n26872 = ~n26870 & ~n26871;
  assign n26873 = ~n13794 & n25462;
  assign n26874 = ~n13790 & n25465;
  assign n26875 = ~n26873 & ~n26874;
  assign n26876 = n26872 & n26875;
  assign n26877 = ~n16712 & n25449;
  assign n26878 = ~n25452 & ~n26877;
  assign n26879 = ~pi0342 & ~n26878;
  assign n26880 = pi0343 & ~n16712;
  assign n26881 = ~pi0343 & ~n13988;
  assign n26882 = ~n26880 & ~n26881;
  assign n26883 = n25458 & ~n26882;
  assign n26884 = ~n26879 & ~n26883;
  assign n26885 = ~n20087 & n20379;
  assign n26886 = ~n20110 & n26885;
  assign n26887 = ~n20111 & ~n20312;
  assign n26888 = ~n20380 & n26887;
  assign n26889 = ~n26886 & ~n26888;
  assign n26890 = n20287 & ~n20304;
  assign n26891 = ~n20265 & ~n26890;
  assign n26892 = ~n20313 & ~n26891;
  assign n26893 = ~n20334 & ~n26892;
  assign n26894 = ~n26889 & n26893;
  assign n26895 = n26889 & ~n26893;
  assign n26896 = ~n26894 & ~n26895;
  assign n26897 = n24892 & n26896;
  assign n26898 = ~n13821 & ~n24905;
  assign n26899 = ~n16712 & n24913;
  assign n26900 = ~n13988 & n24916;
  assign n26901 = ~n26899 & ~n26900;
  assign n26902 = ~n24909 & n26901;
  assign n26903 = ~n26898 & n26902;
  assign n26904 = ~n26897 & n26903;
  assign n26905 = ~n13839 & ~n25475;
  assign n26906 = ~n25471 & ~n26905;
  assign n26907 = ~n13848 & ~n25487;
  assign n26908 = ~n13843 & ~n25483;
  assign n26909 = ~n26907 & ~n26908;
  assign n26910 = ~n25491 & n26909;
  assign n26911 = ~n25479 & n26910;
  assign n26912 = n26906 & n26911;
  assign n26913 = ~pi0343 & ~n26912;
  assign n26914 = pi0343 & ~n13988;
  assign n26915 = ~n26913 & ~n26914;
  assign n26916 = n25498 & ~n26915;
  assign n26917 = n26904 & ~n26916;
  assign n26918 = n26884 & n26917;
  assign n26919 = n26876 & n26918;
  assign n26920 = n26869 & n26919;
  assign n26921 = n25544 & ~n26920;
  assign n26922 = ~pi0075 & n25533;
  assign n26923 = ~pi0194 & pi0979;
  assign n26924 = ~pi0195 & ~pi0979;
  assign n26925 = ~n26923 & ~n26924;
  assign n26926 = n25571 & ~n26925;
  assign n26927 = ~n13852 & ~n25582;
  assign n26928 = ~n13856 & n25582;
  assign n26929 = ~n26927 & ~n26928;
  assign n26930 = n25580 & ~n26929;
  assign n26931 = ~pi0075 & n25532;
  assign n26932 = ~n26930 & ~n26931;
  assign n26933 = n13830 & ~n25594;
  assign n26934 = n13834 & n25594;
  assign n26935 = ~n26933 & ~n26934;
  assign n26936 = n25591 & n26935;
  assign n26937 = n26932 & ~n26936;
  assign n26938 = ~n26926 & n26937;
  assign n26939 = n25606 & ~n26938;
  assign n26940 = ~n13988 & ~n25606;
  assign n26941 = ~n26939 & ~n26940;
  assign n26942 = n25564 & ~n26941;
  assign n26943 = ~n16712 & n25606;
  assign n26944 = ~n25606 & ~n26938;
  assign n26945 = ~n26943 & ~n26944;
  assign n26946 = ~n25564 & ~n26945;
  assign n26947 = ~n26942 & ~n26946;
  assign n26948 = ~n25533 & ~n26947;
  assign n26949 = ~n26922 & ~n26948;
  assign n26950 = ~n25544 & ~n26949;
  assign po0345 = n26921 | n26950;
  assign n26952 = ~n12221 & n24922;
  assign n26953 = ~n12217 & n24925;
  assign n26954 = ~n26952 & ~n26953;
  assign n26955 = ~n12221 & n25462;
  assign n26956 = ~n12217 & n25465;
  assign n26957 = ~n26955 & ~n26956;
  assign n26958 = n25097 & n25246;
  assign n26959 = n25032 & n25100;
  assign n26960 = ~n26958 & ~n26959;
  assign n26961 = n25198 & n25204;
  assign n26962 = n26507 & ~n26961;
  assign n26963 = n25160 & n25237;
  assign n26964 = n25103 & n25162;
  assign n26965 = ~n26963 & ~n26964;
  assign n26966 = n25149 & n25195;
  assign n26967 = n26965 & ~n26966;
  assign n26968 = n25211 & n26967;
  assign n26969 = n26962 & n26968;
  assign n26970 = n25189 & n25202;
  assign n26971 = n26969 & ~n26970;
  assign n26972 = n25181 & n26749;
  assign n26973 = n25032 & n25184;
  assign n26974 = n25146 & n25158;
  assign n26975 = ~n26973 & ~n26974;
  assign n26976 = n25144 & n26975;
  assign n26977 = n26972 & n26976;
  assign n26978 = n26971 & n26977;
  assign n26979 = ~n25071 & ~n25092;
  assign n26980 = n25088 & n26979;
  assign n26981 = n25028 & n25165;
  assign n26982 = n25049 & n25202;
  assign n26983 = ~n26981 & ~n26982;
  assign n26984 = n25036 & n25246;
  assign n26985 = n26983 & ~n26984;
  assign n26986 = ~n25065 & n26985;
  assign n26987 = n25041 & n26459;
  assign n26988 = n25290 & n26457;
  assign n26989 = ~n26987 & ~n26988;
  assign n26990 = n26986 & n26989;
  assign n26991 = n25080 & n26990;
  assign n26992 = n26980 & n26991;
  assign n26993 = n26978 & n26992;
  assign n26994 = n25251 & n25281;
  assign n26995 = n25280 & ~n26994;
  assign n26996 = n25103 & n25355;
  assign n26997 = n25158 & n25358;
  assign n26998 = ~n26996 & ~n26997;
  assign n26999 = n25290 & n26438;
  assign n27000 = n25165 & n25360;
  assign n27001 = ~n26999 & ~n27000;
  assign n27002 = n25230 & n25296;
  assign n27003 = n25149 & n25306;
  assign n27004 = n26482 & ~n27003;
  assign n27005 = n25151 & n25352;
  assign n27006 = n25325 & ~n27005;
  assign n27007 = n25316 & n27006;
  assign n27008 = n25343 & n27007;
  assign n27009 = n27004 & n27008;
  assign n27010 = ~n27002 & n27009;
  assign n27011 = n27001 & n27010;
  assign n27012 = n26998 & n27011;
  assign n27013 = n24932 & n25264;
  assign n27014 = n25198 & n25270;
  assign n27015 = ~n27013 & ~n27014;
  assign n27016 = n25151 & n25248;
  assign n27017 = ~n25255 & ~n27016;
  assign n27018 = ~n26526 & n27017;
  assign n27019 = ~n25258 & n27018;
  assign n27020 = n25234 & n25251;
  assign n27021 = n25237 & n25239;
  assign n27022 = ~n27020 & ~n27021;
  assign n27023 = n25231 & n25267;
  assign n27024 = n27022 & ~n27023;
  assign n27025 = n25227 & n27024;
  assign n27026 = n27019 & n27025;
  assign n27027 = n25041 & n26519;
  assign n27028 = n25261 & n25267;
  assign n27029 = ~n27027 & ~n27028;
  assign n27030 = n27026 & n27029;
  assign n27031 = n27015 & n27030;
  assign n27032 = n27012 & n27031;
  assign n27033 = n25230 & n25287;
  assign n27034 = n24932 & n25292;
  assign n27035 = ~n27033 & ~n27034;
  assign n27036 = n27032 & n27035;
  assign n27037 = ~n25285 & n27036;
  assign n27038 = n26995 & n27037;
  assign n27039 = pi3516 & ~n12217;
  assign n27040 = n27038 & ~n27039;
  assign n27041 = n26993 & n27040;
  assign n27042 = n26960 & n27041;
  assign n27043 = n25134 & n27042;
  assign n27044 = n25371 & ~n27043;
  assign n27045 = n25149 & n25323;
  assign n27046 = n25165 & n25320;
  assign n27047 = ~n27045 & ~n27046;
  assign n27048 = n25246 & n25312;
  assign n27049 = n27047 & ~n27048;
  assign n27050 = n25290 & n25309;
  assign n27051 = n25348 & ~n27050;
  assign n27052 = n25331 & n27051;
  assign n27053 = n25342 & n27052;
  assign n27054 = n25110 & n25237;
  assign n27055 = n25103 & n25114;
  assign n27056 = ~n27054 & ~n27055;
  assign n27057 = n25130 & n25251;
  assign n27058 = pi3516 & ~n12221;
  assign n27059 = ~n27057 & ~n27058;
  assign n27060 = n26562 & n27059;
  assign n27061 = n27056 & n27060;
  assign n27062 = n27053 & n27061;
  assign n27063 = n24932 & n25207;
  assign n27064 = n25158 & n25213;
  assign n27065 = ~n27063 & ~n27064;
  assign n27066 = n25151 & ~n25420;
  assign n27067 = n27065 & ~n27066;
  assign n27068 = n25158 & n25215;
  assign n27069 = n25209 & n25267;
  assign n27070 = ~n27068 & ~n27069;
  assign n27071 = n25230 & n25254;
  assign n27072 = n25251 & n25257;
  assign n27073 = ~n27071 & ~n27072;
  assign n27074 = n25243 & n25290;
  assign n27075 = n24932 & n25276;
  assign n27076 = ~n27074 & ~n27075;
  assign n27077 = n27073 & n27076;
  assign n27078 = n25816 & n27077;
  assign n27079 = n25149 & n25314;
  assign n27080 = n27078 & ~n27079;
  assign n27081 = n25172 & n25230;
  assign n27082 = n25041 & n25169;
  assign n27083 = ~n27081 & ~n27082;
  assign n27084 = n27080 & n27083;
  assign n27085 = n27070 & n27084;
  assign n27086 = n27067 & n27085;
  assign n27087 = n27062 & n27086;
  assign n27088 = n25142 & n25198;
  assign n27089 = n25165 & n25177;
  assign n27090 = ~n27088 & ~n27089;
  assign n27091 = n25202 & ~n25385;
  assign n27092 = n25078 & n25267;
  assign n27093 = ~n27091 & ~n27092;
  assign n27094 = n25041 & n25153;
  assign n27095 = n25032 & n25179;
  assign n27096 = ~n27094 & ~n27095;
  assign n27097 = n27093 & n27096;
  assign n27098 = n25411 & n27097;
  assign n27099 = n27090 & n27098;
  assign n27100 = n25086 & n25237;
  assign n27101 = n25032 & n25084;
  assign n27102 = ~n27100 & ~n27101;
  assign n27103 = n25091 & n25103;
  assign n27104 = n25070 & n25198;
  assign n27105 = ~n27103 & ~n27104;
  assign n27106 = n27102 & n27105;
  assign n27107 = n27099 & n27106;
  assign n27108 = n27087 & n27107;
  assign n27109 = ~n25318 & n27108;
  assign n27110 = n27049 & n27109;
  assign n27111 = n25443 & ~n27110;
  assign n27112 = ~n27044 & ~n27111;
  assign n27113 = ~n16676 & n25508;
  assign n27114 = ~n12415 & n25512;
  assign n27115 = ~n27113 & ~n27114;
  assign n27116 = n27112 & n27115;
  assign n27117 = n26957 & n27116;
  assign n27118 = n26954 & n27117;
  assign n27119 = ~n16676 & n25449;
  assign n27120 = ~n25452 & ~n27119;
  assign n27121 = ~pi0342 & ~n27120;
  assign n27122 = pi0343 & ~n16676;
  assign n27123 = ~pi0343 & ~n12415;
  assign n27124 = ~n27122 & ~n27123;
  assign n27125 = n25458 & ~n27124;
  assign n27126 = ~n27121 & ~n27125;
  assign n27127 = n20313 & n20379;
  assign n27128 = ~n20313 & ~n26890;
  assign n27129 = ~n20380 & n27128;
  assign n27130 = ~n27127 & ~n27129;
  assign n27131 = ~n20265 & ~n20334;
  assign n27132 = ~n27130 & ~n27131;
  assign n27133 = n27130 & n27131;
  assign n27134 = ~n27132 & ~n27133;
  assign n27135 = n24892 & ~n27134;
  assign n27136 = ~n12248 & ~n24905;
  assign n27137 = ~n16676 & n24913;
  assign n27138 = ~n12415 & n24916;
  assign n27139 = ~n27137 & ~n27138;
  assign n27140 = ~n24909 & n27139;
  assign n27141 = ~n27136 & n27140;
  assign n27142 = ~n27135 & n27141;
  assign n27143 = ~n12270 & ~n25475;
  assign n27144 = ~n25471 & ~n27143;
  assign n27145 = ~n12257 & ~n25487;
  assign n27146 = ~n12274 & ~n25483;
  assign n27147 = ~n27145 & ~n27146;
  assign n27148 = ~n25491 & n27147;
  assign n27149 = ~n25479 & n27148;
  assign n27150 = n27144 & n27149;
  assign n27151 = ~pi0343 & ~n27150;
  assign n27152 = pi0343 & ~n12415;
  assign n27153 = ~n27151 & ~n27152;
  assign n27154 = n25498 & ~n27153;
  assign n27155 = n27142 & ~n27154;
  assign n27156 = n27126 & n27155;
  assign n27157 = n27118 & n27156;
  assign n27158 = n25544 & ~n27157;
  assign n27159 = ~pi0076 & n25533;
  assign n27160 = ~pi0187 & pi0979;
  assign n27161 = ~pi0188 & ~pi0979;
  assign n27162 = ~n27160 & ~n27161;
  assign n27163 = n25571 & ~n27162;
  assign n27164 = ~n12261 & ~n25582;
  assign n27165 = ~n12265 & n25582;
  assign n27166 = ~n27164 & ~n27165;
  assign n27167 = n25580 & ~n27166;
  assign n27168 = ~pi0076 & n25532;
  assign n27169 = ~n27167 & ~n27168;
  assign n27170 = n12279 & ~n25594;
  assign n27171 = n12283 & n25594;
  assign n27172 = ~n27170 & ~n27171;
  assign n27173 = n25591 & n27172;
  assign n27174 = n27169 & ~n27173;
  assign n27175 = ~n27163 & n27174;
  assign n27176 = n25606 & ~n27175;
  assign n27177 = ~n12415 & ~n25606;
  assign n27178 = ~n27176 & ~n27177;
  assign n27179 = n25564 & ~n27178;
  assign n27180 = ~n16676 & n25606;
  assign n27181 = ~n25606 & ~n27175;
  assign n27182 = ~n27180 & ~n27181;
  assign n27183 = ~n25564 & ~n27182;
  assign n27184 = ~n27179 & ~n27183;
  assign n27185 = ~n25533 & ~n27184;
  assign n27186 = ~n27159 & ~n27185;
  assign n27187 = ~n25544 & ~n27186;
  assign po0346 = n27158 | n27187;
  assign n27189 = pi3516 & ~n17217;
  assign n27190 = n25331 & n25336;
  assign n27191 = n25348 & n27190;
  assign n27192 = n25074 & n25112;
  assign n27193 = ~n24940 & n27192;
  assign n27194 = n25198 & n27193;
  assign n27195 = n25074 & n25108;
  assign n27196 = n24940 & n27195;
  assign n27197 = n24932 & n27196;
  assign n27198 = ~n27194 & ~n27197;
  assign n27199 = n25144 & n27198;
  assign n27200 = ~n24940 & n27195;
  assign n27201 = n25149 & n27200;
  assign n27202 = n27199 & ~n27201;
  assign n27203 = n25060 & n25184;
  assign n27204 = ~n26472 & ~n27203;
  assign n27205 = n27202 & n27204;
  assign n27206 = n25189 & n25246;
  assign n27207 = n25158 & n26453;
  assign n27208 = ~n27206 & ~n27207;
  assign n27209 = n24940 & n26452;
  assign n27210 = n25165 & n27209;
  assign n27211 = n25103 & n26448;
  assign n27212 = ~n27210 & ~n27211;
  assign n27213 = n27208 & n27212;
  assign n27214 = n25060 & n25146;
  assign n27215 = n25181 & ~n27214;
  assign n27216 = ~n25183 & n27215;
  assign n27217 = n27213 & n27216;
  assign n27218 = n25074 & n25140;
  assign n27219 = ~n24940 & n27218;
  assign n27220 = n25041 & n27219;
  assign n27221 = n25116 & ~n27220;
  assign n27222 = n25060 & n25100;
  assign n27223 = ~n26485 & ~n27222;
  assign n27224 = n24940 & n25140;
  assign n27225 = n25074 & n27224;
  assign n27226 = n25290 & n27225;
  assign n27227 = n25133 & ~n27226;
  assign n27228 = n27223 & n27227;
  assign n27229 = n27221 & n27228;
  assign n27230 = n25032 & n26459;
  assign n27231 = n26466 & ~n27230;
  assign n27232 = n25237 & n26457;
  assign n27233 = n25103 & n26462;
  assign n27234 = ~n27232 & ~n27233;
  assign n27235 = n25044 & n25082;
  assign n27236 = n24940 & n27235;
  assign n27237 = n24932 & n27236;
  assign n27238 = n27234 & ~n27237;
  assign n27239 = n25080 & n27238;
  assign n27240 = n27231 & n27239;
  assign n27241 = n27229 & n27240;
  assign n27242 = n25044 & n25175;
  assign n27243 = ~n24940 & n27242;
  assign n27244 = n25202 & n27243;
  assign n27245 = n25044 & n25089;
  assign n27246 = n24940 & n27245;
  assign n27247 = n25267 & n27246;
  assign n27248 = n25049 & n25246;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = n24940 & n27192;
  assign n27251 = n25267 & n27250;
  assign n27252 = n25026 & n25074;
  assign n27253 = ~n24940 & n27252;
  assign n27254 = n25202 & n27253;
  assign n27255 = ~n27251 & ~n27254;
  assign n27256 = ~n24940 & n27245;
  assign n27257 = n25198 & n27256;
  assign n27258 = n27255 & ~n27257;
  assign n27259 = n25060 & n25306;
  assign n27260 = n25341 & ~n26481;
  assign n27261 = ~n27259 & n27260;
  assign n27262 = n27258 & n27261;
  assign n27263 = n25028 & n25060;
  assign n27264 = n26774 & ~n27263;
  assign n27265 = n27262 & n27264;
  assign n27266 = n27249 & n27265;
  assign n27267 = ~n27244 & n27266;
  assign n27268 = n27241 & n27267;
  assign n27269 = n27217 & n27268;
  assign n27270 = n27205 & n27269;
  assign n27271 = n27191 & n27270;
  assign n27272 = n25060 & n25360;
  assign n27273 = ~n25321 & ~n27272;
  assign n27274 = ~n25315 & n27273;
  assign n27275 = ~n25324 & n27274;
  assign n27276 = n24940 & n27242;
  assign n27277 = n25230 & n27276;
  assign n27278 = ~n24940 & n25044;
  assign n27279 = n25068 & n27278;
  assign n27280 = n25041 & n27279;
  assign n27281 = ~n27277 & ~n27280;
  assign n27282 = n27275 & n27281;
  assign n27283 = n24940 & n26537;
  assign n27284 = n25165 & n27283;
  assign n27285 = n25237 & n26438;
  assign n27286 = ~n27284 & ~n27285;
  assign n27287 = n27282 & n27286;
  assign n27288 = n24940 & n27252;
  assign n27289 = n25230 & n27288;
  assign n27290 = n27287 & ~n27289;
  assign n27291 = n25060 & n25355;
  assign n27292 = n25060 & n25358;
  assign n27293 = ~n27291 & ~n27292;
  assign n27294 = n25060 & n25160;
  assign n27295 = n25060 & n25162;
  assign n27296 = ~n27294 & ~n27295;
  assign n27297 = n25060 & n25204;
  assign n27298 = n27296 & ~n27297;
  assign n27299 = n25060 & n25195;
  assign n27300 = n25151 & n25261;
  assign n27301 = n25032 & n26519;
  assign n27302 = ~n27300 & ~n27301;
  assign n27303 = n25060 & n25270;
  assign n27304 = n27302 & ~n27303;
  assign n27305 = n25060 & n25264;
  assign n27306 = n25060 & n25281;
  assign n27307 = n25280 & ~n27306;
  assign n27308 = ~n25285 & n27307;
  assign n27309 = n26528 & n27308;
  assign n27310 = n25158 & n26538;
  assign n27311 = n25251 & n25296;
  assign n27312 = ~n27310 & ~n27311;
  assign n27313 = n25251 & n25287;
  assign n27314 = n27312 & ~n27313;
  assign n27315 = n25060 & n25292;
  assign n27316 = n27314 & ~n27315;
  assign n27317 = n27309 & n27316;
  assign n27318 = ~n27305 & n27317;
  assign n27319 = n27304 & n27318;
  assign n27320 = n25227 & n27319;
  assign n27321 = n25060 & n25234;
  assign n27322 = n25060 & n25239;
  assign n27323 = ~n27321 & ~n27322;
  assign n27324 = ~n24940 & n27235;
  assign n27325 = n25149 & n27324;
  assign n27326 = n25151 & n25231;
  assign n27327 = ~n27325 & ~n27326;
  assign n27328 = n27323 & n27327;
  assign n27329 = n27320 & n27328;
  assign n27330 = ~n27299 & n27329;
  assign n27331 = n27298 & n27330;
  assign n27332 = n25211 & n26507;
  assign n27333 = n27331 & n27332;
  assign n27334 = n24940 & n25044;
  assign n27335 = n25290 & n27334;
  assign n27336 = n25068 & n27335;
  assign n27337 = n27333 & ~n27336;
  assign n27338 = n27293 & n27337;
  assign n27339 = n27290 & n27338;
  assign n27340 = ~n26476 & n26599;
  assign n27341 = n27339 & n27340;
  assign n27342 = n27271 & n27341;
  assign n27343 = ~n27189 & n27342;
  assign n27344 = n25371 & ~n27343;
  assign n27345 = n25237 & n25243;
  assign n27346 = n25103 & n25248;
  assign n27347 = ~n27345 & ~n27346;
  assign n27348 = n25251 & n25254;
  assign n27349 = n25041 & n25264;
  assign n27350 = ~n27348 & ~n27349;
  assign n27351 = n25270 & n25290;
  assign n27352 = n27350 & ~n27351;
  assign n27353 = n27347 & n27352;
  assign n27354 = ~n25258 & n27353;
  assign n27355 = n25041 & n25292;
  assign n27356 = n25165 & n25234;
  assign n27357 = n24932 & n25239;
  assign n27358 = ~n27356 & ~n27357;
  assign n27359 = n25032 & n25169;
  assign n27360 = n25172 & n25251;
  assign n27361 = ~n27359 & ~n27360;
  assign n27362 = n25151 & n25209;
  assign n27363 = n27361 & ~n27362;
  assign n27364 = n24932 & n25160;
  assign n27365 = n25162 & n25198;
  assign n27366 = ~n27364 & ~n27365;
  assign n27367 = n25195 & n25230;
  assign n27368 = n25204 & n25290;
  assign n27369 = ~n27367 & ~n27368;
  assign n27370 = n27366 & n27369;
  assign n27371 = ~n25208 & n27370;
  assign n27372 = n27363 & n27371;
  assign n27373 = n25165 & n25281;
  assign n27374 = n27372 & ~n27373;
  assign n27375 = ~n25221 & n27374;
  assign n27376 = n27358 & n27375;
  assign n27377 = ~n27355 & n27376;
  assign n27378 = n27354 & n27377;
  assign n27379 = ~n25214 & ~n25277;
  assign n27380 = ~n25279 & n27379;
  assign n27381 = ~n25216 & n27380;
  assign n27382 = n27378 & n27381;
  assign n27383 = ~n25225 & n27382;
  assign n27384 = ~n25285 & n27383;
  assign n27385 = n25326 & n27384;
  assign n27386 = n25103 & n25352;
  assign n27387 = n25198 & n25355;
  assign n27388 = ~n27386 & ~n27387;
  assign n27389 = n25267 & n25358;
  assign n27390 = n25202 & n25360;
  assign n27391 = ~n27389 & ~n27390;
  assign n27392 = n27388 & n27391;
  assign n27393 = n25097 & n25158;
  assign n27394 = n25100 & n25149;
  assign n27395 = ~n27393 & ~n27394;
  assign n27396 = n25134 & n27395;
  assign n27397 = n27392 & n27396;
  assign n27398 = n27385 & n27397;
  assign n27399 = n25064 & n25246;
  assign n27400 = n25036 & n25158;
  assign n27401 = ~n27399 & ~n27400;
  assign n27402 = n25230 & n25306;
  assign n27403 = n25237 & n25309;
  assign n27404 = ~n27402 & ~n27403;
  assign n27405 = n25349 & n27404;
  assign n27406 = n25076 & n25246;
  assign n27407 = n27405 & ~n27406;
  assign n27408 = n25028 & n25202;
  assign n27409 = n25078 & n25151;
  assign n27410 = ~n27408 & ~n27409;
  assign n27411 = n27407 & n27410;
  assign n27412 = n26980 & n27411;
  assign n27413 = n27401 & n27412;
  assign n27414 = pi3516 & ~n17221;
  assign n27415 = n25149 & n25184;
  assign n27416 = n25181 & ~n27415;
  assign n27417 = n25146 & n25267;
  assign n27418 = n25032 & n25153;
  assign n27419 = ~n27417 & ~n27418;
  assign n27420 = n25144 & n27419;
  assign n27421 = ~n25183 & n27420;
  assign n27422 = n27416 & n27421;
  assign n27423 = ~n27414 & n27422;
  assign n27424 = n27413 & n27423;
  assign n27425 = n27398 & n27424;
  assign n27426 = n25443 & ~n27425;
  assign n27427 = ~n27344 & ~n27426;
  assign n27428 = ~n17397 & n25508;
  assign n27429 = ~n17368 & n25512;
  assign n27430 = ~n27428 & ~n27429;
  assign n27431 = n27427 & n27430;
  assign n27432 = ~n17221 & n24922;
  assign n27433 = ~n17217 & n24925;
  assign n27434 = ~n27432 & ~n27433;
  assign n27435 = ~n17221 & n25462;
  assign n27436 = ~n17217 & n25465;
  assign n27437 = ~n27435 & ~n27436;
  assign n27438 = n27434 & n27437;
  assign n27439 = ~n16784 & n25449;
  assign n27440 = ~n25452 & ~n27439;
  assign n27441 = ~pi0342 & ~n27440;
  assign n27442 = pi0343 & ~n17397;
  assign n27443 = ~pi0343 & ~n17368;
  assign n27444 = ~n27442 & ~n27443;
  assign n27445 = n25458 & ~n27444;
  assign n27446 = ~n27441 & ~n27445;
  assign n27447 = ~n17248 & ~n24905;
  assign n27448 = n20427 & n24908;
  assign n27449 = ~n17397 & n24913;
  assign n27450 = ~n17368 & n24916;
  assign n27451 = ~n27449 & ~n27450;
  assign n27452 = n20387 & n24892;
  assign n27453 = n27451 & ~n27452;
  assign n27454 = ~n27448 & n27453;
  assign n27455 = ~n27447 & n27454;
  assign n27456 = ~n9498 & ~n25487;
  assign n27457 = ~n25491 & ~n27456;
  assign n27458 = ~n17327 & n25474;
  assign n27459 = ~n17331 & ~n25483;
  assign n27460 = ~n27458 & ~n27459;
  assign n27461 = ~n17327 & n25473;
  assign n27462 = ~n9498 & n25478;
  assign n27463 = ~n27461 & ~n27462;
  assign n27464 = ~n25471 & n27463;
  assign n27465 = n27460 & n27464;
  assign n27466 = n27457 & n27465;
  assign n27467 = ~pi0341 & ~pi0343;
  assign n27468 = ~n27466 & n27467;
  assign n27469 = ~pi0341 & pi0343;
  assign n27470 = ~n13121 & n27469;
  assign n27471 = ~n27468 & ~n27470;
  assign n27472 = pi0342 & ~n27471;
  assign n27473 = n27455 & ~n27472;
  assign n27474 = n27446 & n27473;
  assign n27475 = n27438 & n27474;
  assign n27476 = n27431 & n27475;
  assign n27477 = n25544 & ~n27476;
  assign n27478 = ~pi0077 & n25533;
  assign n27479 = ~pi0089 & pi0979;
  assign n27480 = ~pi0092 & ~pi0979;
  assign n27481 = ~n27479 & ~n27480;
  assign n27482 = n25571 & ~n27481;
  assign n27483 = ~n17318 & ~n25582;
  assign n27484 = ~n17322 & n25582;
  assign n27485 = ~n27483 & ~n27484;
  assign n27486 = n25580 & ~n27485;
  assign n27487 = ~pi0077 & n25532;
  assign n27488 = ~n27486 & ~n27487;
  assign n27489 = n17309 & ~n25594;
  assign n27490 = n17313 & n25594;
  assign n27491 = ~n27489 & ~n27490;
  assign n27492 = n25591 & n27491;
  assign n27493 = n27488 & ~n27492;
  assign n27494 = ~n27482 & n27493;
  assign n27495 = n25606 & ~n27494;
  assign n27496 = ~n17368 & ~n25606;
  assign n27497 = ~n27495 & ~n27496;
  assign n27498 = n25564 & ~n27497;
  assign n27499 = ~n17397 & n25606;
  assign n27500 = ~n25606 & ~n27494;
  assign n27501 = ~n27499 & ~n27500;
  assign n27502 = ~n25564 & ~n27501;
  assign n27503 = ~n27498 & ~n27502;
  assign n27504 = ~n25533 & ~n27503;
  assign n27505 = ~n27478 & ~n27504;
  assign n27506 = ~n25544 & ~n27505;
  assign po0347 = n27477 | n27506;
  assign n27508 = n25620 & ~n26680;
  assign n27509 = pi0078 & ~n25625;
  assign n27510 = n25558 & ~n26689;
  assign n27511 = ~n24769 & ~n25558;
  assign n27512 = ~n27510 & ~n27511;
  assign n27513 = n25625 & ~n27512;
  assign n27514 = ~n27509 & ~n27513;
  assign n27515 = ~n25620 & ~n27514;
  assign po0348 = n27508 | n27515;
  assign n27517 = n25620 & ~n26920;
  assign n27518 = pi0079 & ~n25625;
  assign n27519 = n25558 & ~n26929;
  assign n27520 = ~n25558 & ~n25699;
  assign n27521 = ~n27519 & ~n27520;
  assign n27522 = n25625 & ~n27521;
  assign n27523 = ~n27518 & ~n27522;
  assign n27524 = ~n25620 & ~n27523;
  assign po0349 = n27517 | n27524;
  assign n27526 = n25620 & ~n27157;
  assign n27527 = pi0080 & ~n25625;
  assign n27528 = n25558 & ~n27166;
  assign n27529 = ~n25558 & ~n25718;
  assign n27530 = ~n27528 & ~n27529;
  assign n27531 = n25625 & ~n27530;
  assign n27532 = ~n27527 & ~n27531;
  assign n27533 = ~n25620 & ~n27532;
  assign po0350 = n27526 | n27533;
  assign n27535 = n25620 & ~n27476;
  assign n27536 = pi0081 & ~n25625;
  assign n27537 = n25558 & ~n27485;
  assign n27538 = ~n24265 & ~n25558;
  assign n27539 = ~n27537 & ~n27538;
  assign n27540 = n25625 & ~n27539;
  assign n27541 = ~n27536 & ~n27540;
  assign n27542 = ~n25620 & ~n27541;
  assign po0351 = n27535 | n27542;
  assign n27544 = n24340 & ~n25712;
  assign n27545 = pi0082 & ~n24340;
  assign po0352 = n27544 | n27545;
  assign n27547 = n24340 & ~n25693;
  assign n27548 = pi0083 & ~n24340;
  assign po0353 = n27547 | n27548;
  assign n27550 = pi0084 & ~n24340;
  assign n27551 = n24340 & ~n25651;
  assign po0354 = n27550 | n27551;
  assign n27553 = ~pi0868 & n26025;
  assign n27554 = ~n21519 & ~n21534;
  assign n27555 = n21519 & n21534;
  assign n27556 = ~n27554 & ~n27555;
  assign n27557 = n24099 & ~n27556;
  assign n27558 = n21519 & ~n21534;
  assign n27559 = ~n21519 & n21534;
  assign n27560 = ~n27558 & ~n27559;
  assign n27561 = ~n24099 & ~n27560;
  assign n27562 = ~n27557 & ~n27561;
  assign n27563 = pi0868 & n27562;
  assign n27564 = ~n27553 & ~n27563;
  assign n27565 = n25637 & ~n27564;
  assign n27566 = pi0085 & n20518;
  assign n27567 = pi0085 & ~n24259;
  assign n27568 = ~pi3245 & ~n15426;
  assign n27569 = pi3245 & ~n16927;
  assign n27570 = ~n27568 & ~n27569;
  assign n27571 = n24259 & ~n27570;
  assign n27572 = ~n27567 & ~n27571;
  assign n27573 = n26002 & ~n27572;
  assign n27574 = ~n27566 & ~n27573;
  assign n27575 = ~n26006 & n27574;
  assign n27576 = ~n25637 & ~n27575;
  assign po0355 = n27565 | n27576;
  assign n27578 = pi0086 & n20518;
  assign n27579 = pi0086 & ~n24259;
  assign n27580 = n24259 & ~n24488;
  assign n27581 = ~n27579 & ~n27580;
  assign n27582 = n26002 & ~n27581;
  assign n27583 = ~n27578 & ~n27582;
  assign n27584 = ~n26006 & n27583;
  assign n27585 = ~n25637 & ~n27584;
  assign n27586 = ~n23249 & n23270;
  assign n27587 = ~n24091 & ~n27586;
  assign n27588 = n23249 & ~n23270;
  assign n27589 = ~n27587 & ~n27588;
  assign n27590 = n23251 & n23275;
  assign n27591 = ~n23251 & ~n23275;
  assign n27592 = ~n27590 & ~n27591;
  assign n27593 = n27589 & n27592;
  assign n27594 = ~n27589 & ~n27592;
  assign n27595 = ~n27593 & ~n27594;
  assign n27596 = pi0868 & n27595;
  assign n27597 = n23249 & n23270;
  assign n27598 = ~n23249 & ~n23270;
  assign n27599 = ~n27597 & ~n27598;
  assign n27600 = n24091 & ~n27599;
  assign n27601 = ~n24091 & n27599;
  assign n27602 = ~n27600 & ~n27601;
  assign n27603 = ~pi0868 & ~n27602;
  assign n27604 = ~n27596 & ~n27603;
  assign n27605 = ~pi1789 & ~pi1932;
  assign n27606 = ~n27604 & ~n27605;
  assign n27607 = n23804 & n24080;
  assign n27608 = n23920 & ~n27607;
  assign n27609 = ~n23694 & ~n24084;
  assign n27610 = ~n27608 & n27609;
  assign n27611 = n27608 & ~n27609;
  assign n27612 = ~n27610 & ~n27611;
  assign n27613 = pi0868 & n27612;
  assign n27614 = n23915 & ~n24080;
  assign n27615 = ~n23802 & ~n27614;
  assign n27616 = ~n23918 & ~n27615;
  assign n27617 = n23787 & n23789;
  assign n27618 = ~n23787 & ~n23789;
  assign n27619 = ~n27617 & ~n27618;
  assign n27620 = n27616 & n27619;
  assign n27621 = ~n27616 & ~n27619;
  assign n27622 = ~n27620 & ~n27621;
  assign n27623 = ~pi0868 & n27622;
  assign n27624 = ~n27613 & ~n27623;
  assign n27625 = pi0868 & n27622;
  assign n27626 = ~n23914 & ~n24080;
  assign n27627 = ~n23913 & n27626;
  assign n27628 = ~n23793 & n23801;
  assign n27629 = n23793 & ~n23801;
  assign n27630 = ~n27628 & ~n27629;
  assign n27631 = n27627 & n27630;
  assign n27632 = ~n27627 & ~n27630;
  assign n27633 = ~n27631 & ~n27632;
  assign n27634 = ~pi0868 & n27633;
  assign n27635 = ~n27625 & ~n27634;
  assign n27636 = n27624 & n27635;
  assign n27637 = pi0868 & n27633;
  assign n27638 = n23799 & ~n23864;
  assign n27639 = ~n23799 & n23864;
  assign n27640 = ~n27638 & ~n27639;
  assign n27641 = ~n23923 & ~n24079;
  assign n27642 = ~n23912 & ~n27641;
  assign n27643 = ~n27640 & ~n27642;
  assign n27644 = n27640 & n27642;
  assign n27645 = ~n27643 & ~n27644;
  assign n27646 = ~pi0868 & n27645;
  assign n27647 = ~n27637 & ~n27646;
  assign n27648 = pi0868 & n27645;
  assign n27649 = ~n23912 & ~n23923;
  assign n27650 = n24079 & ~n27649;
  assign n27651 = ~n24079 & n27649;
  assign n27652 = ~n27650 & ~n27651;
  assign n27653 = ~pi0868 & n27652;
  assign n27654 = ~n27648 & ~n27653;
  assign n27655 = n27647 & n27654;
  assign n27656 = ~n23310 & ~n23422;
  assign n27657 = n23310 & n23422;
  assign n27658 = ~n27656 & ~n27657;
  assign n27659 = n23424 & ~n23514;
  assign n27660 = n23701 & ~n27608;
  assign n27661 = ~n24085 & ~n27660;
  assign n27662 = ~n24086 & n27661;
  assign n27663 = ~n27659 & ~n27662;
  assign n27664 = ~n23515 & ~n27663;
  assign n27665 = ~n27658 & ~n27664;
  assign n27666 = n27658 & n27664;
  assign n27667 = ~n27665 & ~n27666;
  assign n27668 = ~pi0868 & n27667;
  assign n27669 = pi0868 & ~n27602;
  assign n27670 = ~n27668 & ~n27669;
  assign n27671 = pi0868 & n27667;
  assign n27672 = ~n23515 & ~n27659;
  assign n27673 = n27662 & ~n27672;
  assign n27674 = ~n27662 & n27672;
  assign n27675 = ~n27673 & ~n27674;
  assign n27676 = ~pi0868 & n27675;
  assign n27677 = ~n27671 & ~n27676;
  assign n27678 = n27670 & n27677;
  assign n27679 = pi0868 & n27675;
  assign n27680 = ~n23700 & ~n24086;
  assign n27681 = ~n23694 & ~n27608;
  assign n27682 = ~n24084 & ~n27681;
  assign n27683 = ~n27680 & n27682;
  assign n27684 = n27680 & ~n27682;
  assign n27685 = ~n27683 & ~n27684;
  assign n27686 = ~pi0868 & n27685;
  assign n27687 = ~n27679 & ~n27686;
  assign n27688 = pi0868 & n27685;
  assign n27689 = ~pi0868 & n27612;
  assign n27690 = ~n27688 & ~n27689;
  assign n27691 = n27687 & n27690;
  assign n27692 = n27678 & n27691;
  assign n27693 = n27655 & n27692;
  assign n27694 = n27636 & n27693;
  assign n27695 = ~pi0868 & ~n10970;
  assign n27696 = pi1472 & n27695;
  assign n27697 = ~n24025 & ~n24029;
  assign n27698 = ~n24028 & ~n27697;
  assign n27699 = ~n20543 & ~n24024;
  assign n27700 = n20543 & n24024;
  assign n27701 = ~n27699 & ~n27700;
  assign n27702 = n24028 & ~n27701;
  assign n27703 = ~n27698 & ~n27702;
  assign n27704 = pi0868 & n27703;
  assign n27705 = ~n27696 & ~n27704;
  assign n27706 = ~n24019 & ~n24048;
  assign n27707 = ~n24049 & ~n27706;
  assign n27708 = pi0868 & n27707;
  assign n27709 = ~pi0868 & n24046;
  assign n27710 = ~n27708 & ~n27709;
  assign n27711 = n27705 & n27710;
  assign n27712 = pi0868 & n24046;
  assign n27713 = ~pi0868 & n24041;
  assign n27714 = ~n27712 & ~n27713;
  assign n27715 = pi0868 & n24041;
  assign n27716 = ~pi0868 & n27703;
  assign n27717 = ~n27715 & ~n27716;
  assign n27718 = n27714 & n27717;
  assign n27719 = pi0868 & n27652;
  assign n27720 = n24055 & ~n24070;
  assign n27721 = n24057 & n24064;
  assign n27722 = ~n27720 & ~n27721;
  assign n27723 = n23909 & ~n24066;
  assign n27724 = ~n24074 & ~n27723;
  assign n27725 = ~n27722 & n27724;
  assign n27726 = n27722 & ~n27724;
  assign n27727 = ~n27725 & ~n27726;
  assign n27728 = ~pi0868 & n27727;
  assign n27729 = ~n27719 & ~n27728;
  assign n27730 = pi0868 & n27727;
  assign n27731 = n24057 & ~n24064;
  assign n27732 = ~n24057 & n24064;
  assign n27733 = ~n27731 & ~n27732;
  assign n27734 = n24055 & ~n27733;
  assign n27735 = ~n24055 & n27733;
  assign n27736 = ~n27734 & ~n27735;
  assign n27737 = ~pi0868 & n27736;
  assign n27738 = ~n27730 & ~n27737;
  assign n27739 = n27729 & n27738;
  assign n27740 = pi0868 & n27736;
  assign n27741 = ~n24050 & ~n24053;
  assign n27742 = ~n24052 & ~n27741;
  assign n27743 = ~n24005 & n24049;
  assign n27744 = n24005 & ~n24049;
  assign n27745 = ~n27743 & ~n27744;
  assign n27746 = n24052 & ~n27745;
  assign n27747 = ~n27742 & ~n27746;
  assign n27748 = ~pi0868 & n27747;
  assign n27749 = ~n27740 & ~n27748;
  assign n27750 = pi0868 & n27747;
  assign n27751 = ~pi0868 & n27707;
  assign n27752 = ~n27750 & ~n27751;
  assign n27753 = n27749 & n27752;
  assign n27754 = n27739 & n27753;
  assign n27755 = n27718 & n27754;
  assign n27756 = n27711 & n27755;
  assign n27757 = n27694 & n27756;
  assign n27758 = ~n27604 & ~n27757;
  assign n27759 = ~n27606 & ~n27758;
  assign n27760 = n25637 & ~n27759;
  assign po0356 = n27585 | n27760;
  assign n27762 = n25663 & ~n27564;
  assign n27763 = pi0087 & n24300;
  assign n27764 = pi0087 & ~n24314;
  assign n27765 = n24314 & ~n27570;
  assign n27766 = ~n27764 & ~n27765;
  assign n27767 = n26041 & ~n27766;
  assign n27768 = ~n27763 & ~n27767;
  assign n27769 = ~n26045 & n27768;
  assign n27770 = ~n25663 & ~n27769;
  assign po0357 = n27762 | n27770;
  assign n27772 = pi0088 & n24300;
  assign n27773 = pi0088 & ~n24314;
  assign n27774 = n24314 & ~n24488;
  assign n27775 = ~n27773 & ~n27774;
  assign n27776 = n26041 & ~n27775;
  assign n27777 = ~n27772 & ~n27776;
  assign n27778 = ~n26045 & n27777;
  assign n27779 = ~n25663 & ~n27778;
  assign n27780 = n25663 & ~n27759;
  assign po0358 = n27779 | n27780;
  assign n27782 = ~pi0089 & ~n26051;
  assign n27783 = ~n25651 & n26051;
  assign po0359 = n27782 | n27783;
  assign n27785 = n26051 & ~n27564;
  assign n27786 = ~pi0090 & ~n26051;
  assign po0360 = n27785 | n27786;
  assign n27788 = ~pi0091 & ~n26051;
  assign n27789 = n26051 & ~n27759;
  assign po0361 = n27788 | n27789;
  assign n27791 = ~pi0092 & ~n26056;
  assign n27792 = ~n25651 & n26056;
  assign po0362 = n27791 | n27792;
  assign n27794 = n26056 & ~n27564;
  assign n27795 = ~pi0093 & ~n26056;
  assign po0363 = n27794 | n27795;
  assign n27797 = ~pi0094 & ~n26056;
  assign n27798 = n26056 & ~n27759;
  assign po0364 = n27797 | n27798;
  assign n27800 = pi0343 & ~n16819;
  assign n27801 = ~pi0343 & ~n13701;
  assign n27802 = ~n27800 & ~n27801;
  assign n27803 = n25458 & ~n27802;
  assign n27804 = ~n20322 & ~n20334;
  assign n27805 = n19832 & n19848;
  assign n27806 = ~n19832 & ~n19848;
  assign n27807 = ~n27805 & ~n27806;
  assign n27808 = ~n20380 & ~n27807;
  assign n27809 = n19849 & n20379;
  assign n27810 = ~n27808 & ~n27809;
  assign n27811 = ~n27804 & n27810;
  assign n27812 = n27804 & ~n27810;
  assign n27813 = ~n27811 & ~n27812;
  assign n27814 = n24892 & n27813;
  assign n27815 = ~n13583 & ~n24905;
  assign n27816 = ~n27814 & ~n27815;
  assign n27817 = ~n13534 & n25474;
  assign n27818 = ~n25471 & ~n27817;
  assign n27819 = ~n13538 & ~n25483;
  assign n27820 = ~n13534 & n25473;
  assign n27821 = ~n27819 & ~n27820;
  assign n27822 = n27457 & n27821;
  assign n27823 = ~n25479 & n27822;
  assign n27824 = n27818 & n27823;
  assign n27825 = n27467 & ~n27824;
  assign n27826 = ~n27470 & ~n27825;
  assign n27827 = pi0342 & ~n27826;
  assign n27828 = ~n13701 & n24916;
  assign n27829 = ~n16819 & n24913;
  assign n27830 = ~n27828 & ~n27829;
  assign n27831 = ~n27827 & n27830;
  assign n27832 = ~n24909 & n27831;
  assign n27833 = n27816 & n27832;
  assign n27834 = ~n13556 & n24922;
  assign n27835 = ~n13552 & n24925;
  assign n27836 = ~n27834 & ~n27835;
  assign n27837 = ~n13556 & n25462;
  assign n27838 = ~n13552 & n25465;
  assign n27839 = ~n27837 & ~n27838;
  assign n27840 = n25097 & n25230;
  assign n27841 = n25114 & n25246;
  assign n27842 = ~n27840 & ~n27841;
  assign n27843 = n25267 & n25309;
  assign n27844 = n24932 & n25254;
  assign n27845 = n25041 & n25281;
  assign n27846 = ~n27844 & ~n27845;
  assign n27847 = n25243 & n25267;
  assign n27848 = n25202 & n25248;
  assign n27849 = ~n27847 & ~n27848;
  assign n27850 = n25202 & n25352;
  assign n27851 = n25237 & n25314;
  assign n27852 = ~n27850 & ~n27851;
  assign n27853 = n25215 & n25251;
  assign n27854 = n25103 & n25207;
  assign n27855 = ~n27853 & ~n27854;
  assign n27856 = n25213 & n25251;
  assign n27857 = n27855 & ~n27856;
  assign n27858 = n24932 & n25172;
  assign n27859 = n25165 & n25209;
  assign n27860 = ~n27858 & ~n27859;
  assign n27861 = n25041 & n25234;
  assign n27862 = n25169 & n25198;
  assign n27863 = ~n27861 & ~n27862;
  assign n27864 = n27860 & n27863;
  assign n27865 = n25226 & n27864;
  assign n27866 = n27857 & n27865;
  assign n27867 = ~n25258 & ~n25279;
  assign n27868 = n25103 & n25276;
  assign n27869 = n27867 & ~n27868;
  assign n27870 = ~n25285 & n27869;
  assign n27871 = n27866 & n27870;
  assign n27872 = n27852 & n27871;
  assign n27873 = n27849 & n27872;
  assign n27874 = n27846 & n27873;
  assign n27875 = n25237 & n25323;
  assign n27876 = n25032 & n25320;
  assign n27877 = ~n27875 & ~n27876;
  assign n27878 = n26599 & n27877;
  assign n27879 = n27874 & n27878;
  assign n27880 = n25349 & n27879;
  assign n27881 = ~n27843 & n27880;
  assign n27882 = n25142 & n25158;
  assign n27883 = ~n25139 & ~n25180;
  assign n27884 = ~n27882 & n27883;
  assign n27885 = n25184 & n25290;
  assign n27886 = n25032 & n25177;
  assign n27887 = ~n27885 & ~n27886;
  assign n27888 = n25153 & n25198;
  assign n27889 = n27887 & ~n27888;
  assign n27890 = ~n25183 & n27889;
  assign n27891 = n27884 & n27890;
  assign n27892 = n27881 & n27891;
  assign n27893 = n25100 & n25290;
  assign n27894 = n25110 & n25151;
  assign n27895 = ~n27893 & ~n27894;
  assign n27896 = n27892 & n27895;
  assign n27897 = n25133 & n27896;
  assign n27898 = n27842 & n27897;
  assign n27899 = n25070 & n25158;
  assign n27900 = n25091 & n25246;
  assign n27901 = ~n27899 & ~n27900;
  assign n27902 = n25086 & n25151;
  assign n27903 = n27901 & ~n27902;
  assign n27904 = n25064 & n25149;
  assign n27905 = n25036 & n25230;
  assign n27906 = ~n27904 & ~n27905;
  assign n27907 = n25076 & n25149;
  assign n27908 = n25078 & n25165;
  assign n27909 = ~n27907 & ~n27908;
  assign n27910 = n27906 & n27909;
  assign n27911 = ~n25085 & n27910;
  assign n27912 = n27903 & n27911;
  assign n27913 = n27898 & n27912;
  assign n27914 = pi3516 & ~n13556;
  assign n27915 = n27913 & ~n27914;
  assign n27916 = n25443 & ~n27915;
  assign n27917 = n25267 & n26438;
  assign n27918 = n25032 & n25360;
  assign n27919 = ~n27917 & ~n27918;
  assign n27920 = n25246 & n25355;
  assign n27921 = n25251 & n25358;
  assign n27922 = ~n27920 & ~n27921;
  assign n27923 = n25316 & n27922;
  assign n27924 = n27919 & n27923;
  assign n27925 = n25041 & n27283;
  assign n27926 = n27924 & ~n27925;
  assign n27927 = n25103 & n25264;
  assign n27928 = n25158 & n25270;
  assign n27929 = ~n27927 & ~n27928;
  assign n27930 = n25198 & n26519;
  assign n27931 = n25165 & n25261;
  assign n27932 = ~n27930 & ~n27931;
  assign n27933 = n25290 & n27324;
  assign n27934 = n25165 & n25231;
  assign n27935 = ~n27933 & ~n27934;
  assign n27936 = n25251 & n25278;
  assign n27937 = ~n27306 & ~n27936;
  assign n27938 = n26536 & n27937;
  assign n27939 = n25151 & n25239;
  assign n27940 = n25227 & ~n27939;
  assign n27941 = n27938 & n27940;
  assign n27942 = ~n27321 & n27941;
  assign n27943 = n27935 & n27942;
  assign n27944 = n25230 & n26538;
  assign n27945 = n24932 & n25296;
  assign n27946 = ~n27944 & ~n27945;
  assign n27947 = n24932 & n25287;
  assign n27948 = n25103 & n25292;
  assign n27949 = ~n27947 & ~n27948;
  assign n27950 = n27946 & n27949;
  assign n27951 = n27943 & n27950;
  assign n27952 = n26528 & n27951;
  assign n27953 = n27932 & n27952;
  assign n27954 = n27929 & n27953;
  assign n27955 = n25158 & n25204;
  assign n27956 = n26507 & ~n27955;
  assign n27957 = n25151 & n25160;
  assign n27958 = n25162 & n25246;
  assign n27959 = ~n27957 & ~n27958;
  assign n27960 = n25195 & n25237;
  assign n27961 = n27959 & ~n27960;
  assign n27962 = n25211 & n27961;
  assign n27963 = n27956 & n27962;
  assign n27964 = n27954 & n27963;
  assign n27965 = n25237 & n25306;
  assign n27966 = n26482 & ~n27965;
  assign n27967 = ~n25077 & ~n26465;
  assign n27968 = ~n25092 & n27967;
  assign n27969 = ~n25079 & n27968;
  assign n27970 = n25198 & n26459;
  assign n27971 = n27969 & ~n27970;
  assign n27972 = n25267 & n26457;
  assign n27973 = n25202 & n26462;
  assign n27974 = ~n27972 & ~n27973;
  assign n27975 = n25049 & n25149;
  assign n27976 = n25144 & ~n27975;
  assign n27977 = n27974 & n27976;
  assign n27978 = n27971 & n27977;
  assign n27979 = n25028 & n25032;
  assign n27980 = n27978 & ~n27979;
  assign n27981 = n25146 & n25251;
  assign n27982 = n25181 & ~n27981;
  assign n27983 = n25149 & n25189;
  assign n27984 = n25230 & n26453;
  assign n27985 = ~n27983 & ~n27984;
  assign n27986 = n25041 & n27209;
  assign n27987 = n25202 & n26448;
  assign n27988 = ~n27986 & ~n27987;
  assign n27989 = n27985 & n27988;
  assign n27990 = ~n25183 & n27989;
  assign n27991 = n27982 & n27990;
  assign n27992 = n25290 & n27200;
  assign n27993 = n27991 & ~n27992;
  assign n27994 = ~n26472 & n27993;
  assign n27995 = ~n27203 & n27994;
  assign n27996 = n27980 & n27995;
  assign n27997 = n26774 & n27223;
  assign n27998 = n27996 & n27997;
  assign n27999 = n25134 & n27998;
  assign n28000 = n25343 & n27999;
  assign n28001 = n27966 & n28000;
  assign n28002 = pi3516 & ~n13552;
  assign n28003 = n28001 & ~n28002;
  assign n28004 = n27964 & n28003;
  assign n28005 = n26478 & n28004;
  assign n28006 = n27926 & n28005;
  assign n28007 = n25371 & ~n28006;
  assign n28008 = ~n27916 & ~n28007;
  assign n28009 = ~n13701 & n25512;
  assign n28010 = ~n16819 & n25508;
  assign n28011 = ~n28009 & ~n28010;
  assign n28012 = n28008 & n28011;
  assign n28013 = n27839 & n28012;
  assign n28014 = n27836 & n28013;
  assign n28015 = n27833 & n28014;
  assign n28016 = ~n27441 & n28015;
  assign n28017 = ~n27803 & n28016;
  assign n28018 = n25544 & ~n28017;
  assign n28019 = ~pi0095 & n25533;
  assign n28020 = ~pi0147 & pi0979;
  assign n28021 = ~pi0148 & ~pi0979;
  assign n28022 = ~n28020 & ~n28021;
  assign n28023 = n25571 & ~n28022;
  assign n28024 = ~n13525 & ~n25582;
  assign n28025 = ~n13529 & n25582;
  assign n28026 = ~n28024 & ~n28025;
  assign n28027 = n25580 & ~n28026;
  assign n28028 = ~pi0095 & n25532;
  assign n28029 = ~n28027 & ~n28028;
  assign n28030 = n13516 & ~n25594;
  assign n28031 = n13520 & n25594;
  assign n28032 = ~n28030 & ~n28031;
  assign n28033 = n25591 & n28032;
  assign n28034 = n28029 & ~n28033;
  assign n28035 = ~n28023 & n28034;
  assign n28036 = n25606 & n28035;
  assign n28037 = n13701 & ~n25606;
  assign n28038 = ~n28036 & ~n28037;
  assign n28039 = n25564 & n28038;
  assign n28040 = ~n16819 & n25606;
  assign n28041 = ~n25606 & ~n28035;
  assign n28042 = ~n28040 & ~n28041;
  assign n28043 = ~n25564 & ~n28042;
  assign n28044 = ~n28039 & ~n28043;
  assign n28045 = ~n25533 & ~n28044;
  assign n28046 = ~n28019 & ~n28045;
  assign n28047 = ~n25544 & ~n28046;
  assign po0365 = n28018 | n28047;
  assign n28049 = n25202 & n25309;
  assign n28050 = n25348 & ~n28049;
  assign n28051 = n25153 & n25267;
  assign n28052 = n25177 & n25237;
  assign n28053 = ~n28051 & ~n28052;
  assign n28054 = n25142 & n25165;
  assign n28055 = n28053 & ~n28054;
  assign n28056 = n25151 & n25179;
  assign n28057 = n28055 & ~n28056;
  assign n28058 = n25202 & n25243;
  assign n28059 = n25230 & n25248;
  assign n28060 = ~n28058 & ~n28059;
  assign n28061 = n25198 & n25254;
  assign n28062 = n25281 & n25290;
  assign n28063 = ~n28061 & ~n28062;
  assign n28064 = n25237 & n25320;
  assign n28065 = n25103 & n25323;
  assign n28066 = ~n28064 & ~n28065;
  assign n28067 = n25032 & n25215;
  assign n28068 = n25158 & n25207;
  assign n28069 = ~n28067 & ~n28068;
  assign n28070 = n25032 & n25213;
  assign n28071 = n28069 & ~n28070;
  assign n28072 = n25172 & n25198;
  assign n28073 = n25149 & n25209;
  assign n28074 = ~n28072 & ~n28073;
  assign n28075 = n25234 & n25290;
  assign n28076 = n25169 & n25267;
  assign n28077 = ~n28075 & ~n28076;
  assign n28078 = n28074 & n28077;
  assign n28079 = n25226 & n28078;
  assign n28080 = n28071 & n28079;
  assign n28081 = n25158 & n25276;
  assign n28082 = n27867 & ~n28081;
  assign n28083 = ~n25285 & n28082;
  assign n28084 = n28080 & n28083;
  assign n28085 = n28066 & n28084;
  assign n28086 = n28063 & n28085;
  assign n28087 = n28060 & n28086;
  assign n28088 = n25230 & n25352;
  assign n28089 = n25103 & n25314;
  assign n28090 = ~n28088 & ~n28089;
  assign n28091 = n26599 & n28090;
  assign n28092 = n28087 & n28091;
  assign n28093 = n24932 & n25064;
  assign n28094 = n25036 & n25041;
  assign n28095 = ~n28093 & ~n28094;
  assign n28096 = n28092 & n28095;
  assign n28097 = n25411 & n28096;
  assign n28098 = n28057 & n28097;
  assign n28099 = n24932 & n25076;
  assign n28100 = n25078 & n25149;
  assign n28101 = ~n28099 & ~n28100;
  assign n28102 = n25091 & n25251;
  assign n28103 = n25070 & n25165;
  assign n28104 = ~n28102 & ~n28103;
  assign n28105 = n25086 & n25246;
  assign n28106 = n25084 & n25151;
  assign n28107 = ~n28105 & ~n28106;
  assign n28108 = n28104 & n28107;
  assign n28109 = n28101 & n28108;
  assign n28110 = n28098 & n28109;
  assign n28111 = pi3516 & ~n12962;
  assign n28112 = n28110 & ~n28111;
  assign n28113 = n25041 & n25097;
  assign n28114 = n25110 & n25246;
  assign n28115 = ~n28113 & ~n28114;
  assign n28116 = n25114 & n25251;
  assign n28117 = n25133 & ~n28116;
  assign n28118 = n28115 & n28117;
  assign n28119 = n28112 & n28118;
  assign n28120 = n25342 & n28119;
  assign n28121 = n25331 & n28120;
  assign n28122 = n28050 & n28121;
  assign n28123 = n25443 & ~n28122;
  assign n28124 = n25290 & n27209;
  assign n28125 = n25230 & n26448;
  assign n28126 = ~n28124 & ~n28125;
  assign n28127 = n25165 & n25204;
  assign n28128 = n26507 & ~n28127;
  assign n28129 = n25149 & n25231;
  assign n28130 = n25103 & n25195;
  assign n28131 = ~n28129 & ~n28130;
  assign n28132 = n25160 & n25246;
  assign n28133 = n25162 & n25251;
  assign n28134 = ~n28132 & ~n28133;
  assign n28135 = n28131 & n28134;
  assign n28136 = n25211 & n28135;
  assign n28137 = n28128 & n28136;
  assign n28138 = n25239 & n25246;
  assign n28139 = n28137 & ~n28138;
  assign n28140 = n25103 & n25306;
  assign n28141 = n25343 & ~n28140;
  assign n28142 = n26482 & n28141;
  assign n28143 = n25100 & n25151;
  assign n28144 = n28142 & ~n28143;
  assign n28145 = n25116 & n28144;
  assign n28146 = ~n27321 & n28145;
  assign n28147 = n28139 & n28146;
  assign n28148 = n25227 & n26486;
  assign n28149 = n28147 & n28148;
  assign n28150 = n24932 & n25189;
  assign n28151 = n25041 & n26453;
  assign n28152 = ~n28150 & ~n28151;
  assign n28153 = n25032 & n25146;
  assign n28154 = n25181 & ~n28153;
  assign n28155 = n28152 & n28154;
  assign n28156 = ~n25183 & n28155;
  assign n28157 = n25267 & n26459;
  assign n28158 = n25202 & n26457;
  assign n28159 = ~n28157 & ~n28158;
  assign n28160 = n25230 & n26462;
  assign n28161 = n26467 & ~n28160;
  assign n28162 = n28159 & n28161;
  assign n28163 = n28156 & n28162;
  assign n28164 = n28149 & n28163;
  assign n28165 = n28126 & n28164;
  assign n28166 = n26474 & n28165;
  assign n28167 = n25151 & n25184;
  assign n28168 = n24932 & n25049;
  assign n28169 = n25028 & n25237;
  assign n28170 = ~n28168 & ~n28169;
  assign n28171 = ~n25065 & n28170;
  assign n28172 = n25144 & n28171;
  assign n28173 = ~n28167 & n28172;
  assign n28174 = pi3516 & ~n12958;
  assign n28175 = n25202 & n26438;
  assign n28176 = n25237 & n25360;
  assign n28177 = ~n28175 & ~n28176;
  assign n28178 = n25316 & n28177;
  assign n28179 = n25290 & n27283;
  assign n28180 = n28178 & ~n28179;
  assign n28181 = n25158 & n25264;
  assign n28182 = n25165 & n25270;
  assign n28183 = ~n28181 & ~n28182;
  assign n28184 = n25032 & n25278;
  assign n28185 = ~n27306 & ~n28184;
  assign n28186 = n26536 & n28185;
  assign n28187 = n25267 & n26519;
  assign n28188 = n25149 & n25261;
  assign n28189 = ~n28187 & ~n28188;
  assign n28190 = n28186 & n28189;
  assign n28191 = n28183 & n28190;
  assign n28192 = n26528 & n28191;
  assign n28193 = n25041 & n26538;
  assign n28194 = n25198 & n25296;
  assign n28195 = ~n28193 & ~n28194;
  assign n28196 = n25198 & n25287;
  assign n28197 = n25158 & n25292;
  assign n28198 = ~n28196 & ~n28197;
  assign n28199 = n28195 & n28198;
  assign n28200 = n28192 & n28199;
  assign n28201 = n25251 & n25355;
  assign n28202 = n25032 & n25358;
  assign n28203 = ~n28201 & ~n28202;
  assign n28204 = n26478 & n28203;
  assign n28205 = n28200 & n28204;
  assign n28206 = n28180 & n28205;
  assign n28207 = ~n28174 & n28206;
  assign n28208 = n28173 & n28207;
  assign n28209 = n28166 & n28208;
  assign n28210 = n25371 & ~n28209;
  assign n28211 = ~n28123 & ~n28210;
  assign n28212 = ~n16784 & n25508;
  assign n28213 = ~n13121 & n25512;
  assign n28214 = ~n28212 & ~n28213;
  assign n28215 = n28211 & n28214;
  assign n28216 = ~n12962 & n24922;
  assign n28217 = ~n12958 & n24925;
  assign n28218 = ~n28216 & ~n28217;
  assign n28219 = ~n12962 & n25462;
  assign n28220 = ~n12958 & n25465;
  assign n28221 = ~n28219 & ~n28220;
  assign n28222 = n28218 & n28221;
  assign n28223 = ~n20030 & ~n20316;
  assign n28224 = ~n20318 & ~n28223;
  assign n28225 = ~n20334 & ~n28224;
  assign n28226 = ~n19974 & n19990;
  assign n28227 = n19974 & ~n19990;
  assign n28228 = ~n28226 & ~n28227;
  assign n28229 = ~n20380 & ~n28228;
  assign n28230 = n20321 & n20379;
  assign n28231 = ~n28229 & ~n28230;
  assign n28232 = ~n28225 & n28231;
  assign n28233 = n28225 & ~n28231;
  assign n28234 = ~n28232 & ~n28233;
  assign n28235 = n24892 & n28234;
  assign n28236 = ~n12989 & ~n24905;
  assign n28237 = ~n16784 & n24913;
  assign n28238 = ~n13121 & n24916;
  assign n28239 = ~n28237 & ~n28238;
  assign n28240 = ~n24909 & n28239;
  assign n28241 = ~n28236 & n28240;
  assign n28242 = ~n28235 & n28241;
  assign n28243 = ~n12940 & n25474;
  assign n28244 = ~n25471 & ~n28243;
  assign n28245 = ~n12940 & n25473;
  assign n28246 = ~n12944 & ~n25483;
  assign n28247 = ~n28245 & ~n28246;
  assign n28248 = n27457 & n28247;
  assign n28249 = ~n25479 & n28248;
  assign n28250 = n28244 & n28249;
  assign n28251 = n27467 & ~n28250;
  assign n28252 = ~n27470 & ~n28251;
  assign n28253 = pi0342 & ~n28252;
  assign n28254 = n28242 & ~n28253;
  assign n28255 = pi0343 & ~n16784;
  assign n28256 = ~pi0343 & ~n13121;
  assign n28257 = ~n28255 & ~n28256;
  assign n28258 = n25458 & ~n28257;
  assign n28259 = ~n27441 & ~n28258;
  assign n28260 = n28254 & n28259;
  assign n28261 = n28222 & n28260;
  assign n28262 = n28215 & n28261;
  assign n28263 = n25544 & ~n28262;
  assign n28264 = ~pi0096 & n25533;
  assign n28265 = ~pi0140 & pi0979;
  assign n28266 = ~pi0142 & ~pi0979;
  assign n28267 = ~n28265 & ~n28266;
  assign n28268 = n25571 & ~n28267;
  assign n28269 = ~n12931 & ~n25582;
  assign n28270 = ~n12935 & n25582;
  assign n28271 = ~n28269 & ~n28270;
  assign n28272 = n25580 & ~n28271;
  assign n28273 = ~pi0096 & n25532;
  assign n28274 = ~n28272 & ~n28273;
  assign n28275 = n12922 & ~n25594;
  assign n28276 = n12926 & n25594;
  assign n28277 = ~n28275 & ~n28276;
  assign n28278 = n25591 & n28277;
  assign n28279 = n28274 & ~n28278;
  assign n28280 = ~n28268 & n28279;
  assign n28281 = n25606 & ~n28280;
  assign n28282 = ~n13121 & ~n25606;
  assign n28283 = ~n28281 & ~n28282;
  assign n28284 = n25564 & ~n28283;
  assign n28285 = ~n16784 & n25606;
  assign n28286 = ~n25606 & ~n28280;
  assign n28287 = ~n28285 & ~n28286;
  assign n28288 = ~n25564 & ~n28287;
  assign n28289 = ~n28284 & ~n28288;
  assign n28290 = ~n25533 & ~n28289;
  assign n28291 = ~n28264 & ~n28290;
  assign n28292 = ~n25544 & ~n28291;
  assign po0366 = n28263 | n28292;
  assign n28294 = ~n16640 & n25508;
  assign n28295 = ~n14816 & n25512;
  assign n28296 = ~n28294 & ~n28295;
  assign n28297 = ~n20047 & n20379;
  assign n28298 = ~n20070 & n28297;
  assign n28299 = ~n20071 & ~n20154;
  assign n28300 = ~n20380 & n28299;
  assign n28301 = ~n28298 & ~n28300;
  assign n28302 = ~n20153 & ~n20263;
  assign n28303 = ~n20150 & ~n28302;
  assign n28304 = ~n20334 & ~n28303;
  assign n28305 = ~n28301 & n28304;
  assign n28306 = n28301 & ~n28304;
  assign n28307 = ~n28305 & ~n28306;
  assign n28308 = n24892 & n28307;
  assign n28309 = ~n14649 & ~n24905;
  assign n28310 = ~n16640 & n24913;
  assign n28311 = ~n14816 & n24916;
  assign n28312 = ~n28310 & ~n28311;
  assign n28313 = ~n24909 & n28312;
  assign n28314 = ~n28309 & n28313;
  assign n28315 = ~n28308 & n28314;
  assign n28316 = ~n16640 & n25449;
  assign n28317 = ~n25452 & ~n28316;
  assign n28318 = ~pi0342 & ~n28317;
  assign n28319 = pi0343 & ~n16640;
  assign n28320 = ~pi0343 & ~n14816;
  assign n28321 = ~n28319 & ~n28320;
  assign n28322 = n25458 & ~n28321;
  assign n28323 = ~n28318 & ~n28322;
  assign n28324 = ~n14609 & n25462;
  assign n28325 = ~n14605 & n25465;
  assign n28326 = ~n28324 & ~n28325;
  assign n28327 = ~n14676 & n25474;
  assign n28328 = ~n25479 & ~n28327;
  assign n28329 = ~n25471 & n28328;
  assign n28330 = ~n14680 & ~n25483;
  assign n28331 = n28329 & ~n28330;
  assign n28332 = ~n14685 & ~n25487;
  assign n28333 = ~n14676 & n25473;
  assign n28334 = ~n28332 & ~n28333;
  assign n28335 = n28331 & n28334;
  assign n28336 = ~n25491 & n28335;
  assign n28337 = ~pi0343 & ~n28336;
  assign n28338 = pi0343 & ~n14816;
  assign n28339 = ~n28337 & ~n28338;
  assign n28340 = n25498 & ~n28339;
  assign n28341 = ~n14609 & n24922;
  assign n28342 = ~n14605 & n24925;
  assign n28343 = ~n28341 & ~n28342;
  assign n28344 = ~n28340 & n28343;
  assign n28345 = n28326 & n28344;
  assign n28346 = n28323 & n28345;
  assign n28347 = n28315 & n28346;
  assign n28348 = n25028 & n25149;
  assign n28349 = n25036 & n25251;
  assign n28350 = ~n28348 & ~n28349;
  assign n28351 = n25290 & n26459;
  assign n28352 = n28350 & ~n28351;
  assign n28353 = ~n25087 & ~n25092;
  assign n28354 = ~n25085 & n28353;
  assign n28355 = n28352 & n28354;
  assign n28356 = n25049 & n25230;
  assign n28357 = n28355 & ~n28356;
  assign n28358 = n25097 & n25251;
  assign n28359 = n25100 & n25237;
  assign n28360 = ~n28358 & ~n28359;
  assign n28361 = pi3516 & ~n14605;
  assign n28362 = n25134 & ~n28361;
  assign n28363 = n28360 & n28362;
  assign n28364 = n25204 & n25267;
  assign n28365 = n26507 & ~n28364;
  assign n28366 = n25103 & n25160;
  assign n28367 = n25158 & n25162;
  assign n28368 = ~n28366 & ~n28367;
  assign n28369 = n24932 & n25195;
  assign n28370 = n28368 & ~n28369;
  assign n28371 = n25211 & n28370;
  assign n28372 = n28365 & n28371;
  assign n28373 = n25189 & n25230;
  assign n28374 = n28372 & ~n28373;
  assign n28375 = n25184 & n25237;
  assign n28376 = n25146 & n25165;
  assign n28377 = ~n28375 & ~n28376;
  assign n28378 = n25144 & n28377;
  assign n28379 = n26972 & n28378;
  assign n28380 = n28374 & n28379;
  assign n28381 = n28363 & n28380;
  assign n28382 = n25202 & n25231;
  assign n28383 = n25227 & ~n28382;
  assign n28384 = n25032 & n25234;
  assign n28385 = n25103 & n25239;
  assign n28386 = ~n28384 & ~n28385;
  assign n28387 = n25198 & n25264;
  assign n28388 = n25267 & n25270;
  assign n28389 = ~n28387 & ~n28388;
  assign n28390 = n25290 & n26519;
  assign n28391 = n25202 & n25261;
  assign n28392 = ~n28390 & ~n28391;
  assign n28393 = n25151 & n25243;
  assign n28394 = n25246 & n25248;
  assign n28395 = ~n28393 & ~n28394;
  assign n28396 = n28392 & n28395;
  assign n28397 = n25259 & n28396;
  assign n28398 = n28389 & n28397;
  assign n28399 = n25032 & n25281;
  assign n28400 = n25280 & ~n28399;
  assign n28401 = n25041 & n25287;
  assign n28402 = n25198 & n25292;
  assign n28403 = ~n28401 & ~n28402;
  assign n28404 = n25041 & n25296;
  assign n28405 = n28403 & ~n28404;
  assign n28406 = ~n25285 & n28405;
  assign n28407 = n28400 & n28406;
  assign n28408 = n28398 & n28407;
  assign n28409 = n24932 & n25306;
  assign n28410 = n25151 & n25309;
  assign n28411 = ~n28409 & ~n28410;
  assign n28412 = n25350 & n28411;
  assign n28413 = n25165 & n25358;
  assign n28414 = n25149 & n25360;
  assign n28415 = ~n28413 & ~n28414;
  assign n28416 = n25246 & n25352;
  assign n28417 = n25158 & n25355;
  assign n28418 = ~n28416 & ~n28417;
  assign n28419 = n28415 & n28418;
  assign n28420 = n28412 & n28419;
  assign n28421 = n28408 & n28420;
  assign n28422 = n28386 & n28421;
  assign n28423 = n28383 & n28422;
  assign n28424 = n28381 & n28423;
  assign n28425 = n25081 & n28424;
  assign n28426 = n28357 & n28425;
  assign n28427 = n25371 & ~n28426;
  assign n28428 = n25336 & n25348;
  assign n28429 = ~n25128 & ~n25330;
  assign n28430 = ~n25119 & ~n25340;
  assign n28431 = n28429 & n28430;
  assign n28432 = n28428 & n28431;
  assign n28433 = n25103 & n25110;
  assign n28434 = n25114 & n25158;
  assign n28435 = ~n28433 & ~n28434;
  assign n28436 = n25032 & n25130;
  assign n28437 = n25151 & n25327;
  assign n28438 = ~n28436 & ~n28437;
  assign n28439 = n28435 & n28438;
  assign n28440 = ~n25123 & n28439;
  assign n28441 = ~n25338 & n28440;
  assign n28442 = n25251 & n25312;
  assign n28443 = n25041 & n25254;
  assign n28444 = ~n28442 & ~n28443;
  assign n28445 = n25032 & n25257;
  assign n28446 = n28444 & ~n28445;
  assign n28447 = ~n25279 & n28446;
  assign n28448 = pi3516 & ~n14609;
  assign n28449 = n28447 & ~n28448;
  assign n28450 = n25246 & ~n25420;
  assign n28451 = n25198 & n25207;
  assign n28452 = n25165 & n25213;
  assign n28453 = ~n28451 & ~n28452;
  assign n28454 = n25165 & n25215;
  assign n28455 = n25202 & n25209;
  assign n28456 = ~n28454 & ~n28455;
  assign n28457 = n25041 & n25172;
  assign n28458 = n25169 & n25290;
  assign n28459 = ~n28457 & ~n28458;
  assign n28460 = n28456 & n28459;
  assign n28461 = n28453 & n28460;
  assign n28462 = ~n28450 & n28461;
  assign n28463 = n25151 & n25317;
  assign n28464 = n28462 & ~n28463;
  assign n28465 = ~n25285 & n28464;
  assign n28466 = n25198 & n25276;
  assign n28467 = n24932 & n25314;
  assign n28468 = ~n28466 & ~n28467;
  assign n28469 = n25149 & n25320;
  assign n28470 = n24932 & n25323;
  assign n28471 = ~n28469 & ~n28470;
  assign n28472 = n28468 & n28471;
  assign n28473 = n28465 & n28472;
  assign n28474 = n28449 & n28473;
  assign n28475 = n25091 & n25158;
  assign n28476 = n25070 & n25267;
  assign n28477 = ~n28475 & ~n28476;
  assign n28478 = n25153 & n25290;
  assign n28479 = n25179 & n25237;
  assign n28480 = ~n28478 & ~n28479;
  assign n28481 = n25142 & n25267;
  assign n28482 = n25149 & n25177;
  assign n28483 = ~n28481 & ~n28482;
  assign n28484 = n28480 & n28483;
  assign n28485 = n25411 & n28484;
  assign n28486 = n25078 & n25202;
  assign n28487 = n25230 & ~n25385;
  assign n28488 = ~n28486 & ~n28487;
  assign n28489 = n28485 & n28488;
  assign n28490 = n25084 & n25237;
  assign n28491 = n25086 & n25103;
  assign n28492 = ~n28490 & ~n28491;
  assign n28493 = n28489 & n28492;
  assign n28494 = n28477 & n28493;
  assign n28495 = n28474 & n28494;
  assign n28496 = n28441 & n28495;
  assign n28497 = n28432 & n28496;
  assign n28498 = n25443 & ~n28497;
  assign n28499 = ~n28427 & ~n28498;
  assign n28500 = n28347 & n28499;
  assign n28501 = n28296 & n28500;
  assign n28502 = n25544 & ~n28501;
  assign n28503 = ~pi0097 & n25533;
  assign n28504 = ~pi0219 & pi0979;
  assign n28505 = ~pi0221 & ~pi0979;
  assign n28506 = ~n28504 & ~n28505;
  assign n28507 = n25571 & ~n28506;
  assign n28508 = ~n14667 & ~n25582;
  assign n28509 = ~n14671 & n25582;
  assign n28510 = ~n28508 & ~n28509;
  assign n28511 = n25580 & ~n28510;
  assign n28512 = ~pi0097 & n25532;
  assign n28513 = ~n28511 & ~n28512;
  assign n28514 = n14658 & ~n25594;
  assign n28515 = n14662 & n25594;
  assign n28516 = ~n28514 & ~n28515;
  assign n28517 = n25591 & n28516;
  assign n28518 = n28513 & ~n28517;
  assign n28519 = ~n28507 & n28518;
  assign n28520 = n25606 & ~n28519;
  assign n28521 = ~n14816 & ~n25606;
  assign n28522 = ~n28520 & ~n28521;
  assign n28523 = n25564 & ~n28522;
  assign n28524 = ~n16640 & n25606;
  assign n28525 = ~n25606 & ~n28519;
  assign n28526 = ~n28524 & ~n28525;
  assign n28527 = ~n25564 & ~n28526;
  assign n28528 = ~n28523 & ~n28527;
  assign n28529 = ~n25533 & ~n28528;
  assign n28530 = ~n28503 & ~n28529;
  assign n28531 = ~n25544 & ~n28530;
  assign po0367 = n28502 | n28531;
  assign n28533 = n25177 & n25251;
  assign n28534 = ~n25183 & ~n28533;
  assign n28535 = n27883 & n28534;
  assign n28536 = n24932 & n25153;
  assign n28537 = n28535 & ~n28536;
  assign n28538 = n25041 & n25184;
  assign n28539 = n25103 & n25142;
  assign n28540 = ~n28538 & ~n28539;
  assign n28541 = n25064 & n25165;
  assign n28542 = n25070 & n25103;
  assign n28543 = ~n28541 & ~n28542;
  assign n28544 = n25091 & n25151;
  assign n28545 = n25088 & ~n28544;
  assign n28546 = n28543 & n28545;
  assign n28547 = n25076 & n25165;
  assign n28548 = n28546 & ~n28547;
  assign n28549 = n25036 & n25202;
  assign n28550 = n25078 & n25158;
  assign n28551 = ~n28549 & ~n28550;
  assign n28552 = n28548 & n28551;
  assign n28553 = n28540 & n28552;
  assign n28554 = n28537 & n28553;
  assign n28555 = n25251 & n25320;
  assign n28556 = n25032 & n25323;
  assign n28557 = ~n28555 & ~n28556;
  assign n28558 = n25237 & n25276;
  assign n28559 = n27867 & ~n28558;
  assign n28560 = n25230 & n25234;
  assign n28561 = n25207 & n25237;
  assign n28562 = ~n28560 & ~n28561;
  assign n28563 = n25160 & n25290;
  assign n28564 = n28562 & ~n28563;
  assign n28565 = n25215 & n25246;
  assign n28566 = n25158 & n25209;
  assign n28567 = ~n28565 & ~n28566;
  assign n28568 = n25239 & n25290;
  assign n28569 = n25213 & n25246;
  assign n28570 = ~n28568 & ~n28569;
  assign n28571 = n25226 & n28570;
  assign n28572 = n28567 & n28571;
  assign n28573 = n28564 & n28572;
  assign n28574 = n25149 & n25172;
  assign n28575 = n24932 & n25169;
  assign n28576 = ~n28574 & ~n28575;
  assign n28577 = n28573 & n28576;
  assign n28578 = ~n25285 & n28577;
  assign n28579 = n28559 & n28578;
  assign n28580 = n25149 & n25254;
  assign n28581 = n25230 & n25281;
  assign n28582 = ~n28580 & ~n28581;
  assign n28583 = n25198 & n25243;
  assign n28584 = n25248 & n25267;
  assign n28585 = ~n28583 & ~n28584;
  assign n28586 = n28582 & n28585;
  assign n28587 = n28579 & n28586;
  assign n28588 = n25267 & n25352;
  assign n28589 = n25032 & n25314;
  assign n28590 = ~n28588 & ~n28589;
  assign n28591 = n28587 & n28590;
  assign n28592 = n26599 & n28591;
  assign n28593 = n28557 & n28592;
  assign n28594 = n25198 & n25309;
  assign n28595 = n28593 & ~n28594;
  assign n28596 = n25343 & n28595;
  assign n28597 = n25348 & n28596;
  assign n28598 = pi3516 & ~n12520;
  assign n28599 = n28597 & ~n28598;
  assign n28600 = n25114 & n25151;
  assign n28601 = n25097 & n25202;
  assign n28602 = ~n28600 & ~n28601;
  assign n28603 = n25041 & n25100;
  assign n28604 = n28602 & ~n28603;
  assign n28605 = n25124 & n28604;
  assign n28606 = n28599 & n28605;
  assign n28607 = n25132 & n28606;
  assign n28608 = ~n25111 & n28607;
  assign n28609 = n28554 & n28608;
  assign n28610 = n25443 & ~n28609;
  assign n28611 = n24932 & n26519;
  assign n28612 = n25158 & n25261;
  assign n28613 = ~n28611 & ~n28612;
  assign n28614 = n25237 & n25264;
  assign n28615 = n25103 & n25270;
  assign n28616 = ~n28614 & ~n28615;
  assign n28617 = n25149 & n25287;
  assign n28618 = n25237 & n25292;
  assign n28619 = ~n28617 & ~n28618;
  assign n28620 = n25202 & n26538;
  assign n28621 = n25149 & n25296;
  assign n28622 = ~n28620 & ~n28621;
  assign n28623 = n25032 & n25306;
  assign n28624 = n26482 & ~n28623;
  assign n28625 = n24932 & n26459;
  assign n28626 = n25198 & n26457;
  assign n28627 = ~n28625 & ~n28626;
  assign n28628 = n25146 & n25246;
  assign n28629 = n25181 & ~n28628;
  assign n28630 = n25230 & n27209;
  assign n28631 = n25267 & n26448;
  assign n28632 = ~n28630 & ~n28631;
  assign n28633 = n25165 & n25189;
  assign n28634 = n25202 & n26453;
  assign n28635 = ~n28633 & ~n28634;
  assign n28636 = n28632 & n28635;
  assign n28637 = ~n25183 & n28636;
  assign n28638 = n28629 & n28637;
  assign n28639 = n27969 & n28638;
  assign n28640 = n25267 & n26462;
  assign n28641 = n25290 & n27236;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = n28639 & n28642;
  assign n28644 = n28627 & n28643;
  assign n28645 = n25041 & n27200;
  assign n28646 = n28644 & ~n28645;
  assign n28647 = ~n25065 & ~n27203;
  assign n28648 = n26471 & n28647;
  assign n28649 = ~n26472 & n28648;
  assign n28650 = n28646 & n28649;
  assign n28651 = n25049 & n25165;
  assign n28652 = n25028 & n25251;
  assign n28653 = ~n28651 & ~n28652;
  assign n28654 = n25290 & n27196;
  assign n28655 = ~n25085 & ~n28654;
  assign n28656 = n28653 & n28655;
  assign n28657 = n28650 & n28656;
  assign n28658 = n25144 & n27223;
  assign n28659 = n28657 & n28658;
  assign n28660 = n25343 & n28659;
  assign n28661 = n28624 & n28660;
  assign n28662 = n25134 & n28661;
  assign n28663 = n25246 & n25278;
  assign n28664 = ~n27306 & ~n28663;
  assign n28665 = n25227 & n27323;
  assign n28666 = n25041 & n27324;
  assign n28667 = n25158 & n25231;
  assign n28668 = ~n28666 & ~n28667;
  assign n28669 = n28665 & n28668;
  assign n28670 = n26536 & n28669;
  assign n28671 = n28664 & n28670;
  assign n28672 = n28662 & n28671;
  assign n28673 = n28622 & n28672;
  assign n28674 = n28619 & n28673;
  assign n28675 = n25198 & n26438;
  assign n28676 = n25251 & n25360;
  assign n28677 = ~n28675 & ~n28676;
  assign n28678 = n25316 & n28677;
  assign n28679 = n25230 & n27283;
  assign n28680 = n28678 & ~n28679;
  assign n28681 = n25103 & n25204;
  assign n28682 = n25211 & ~n27294;
  assign n28683 = n26507 & n28682;
  assign n28684 = ~n28681 & n28683;
  assign n28685 = n25032 & n25195;
  assign n28686 = n25151 & n25162;
  assign n28687 = ~n28685 & ~n28686;
  assign n28688 = n28684 & n28687;
  assign n28689 = n25151 & n25355;
  assign n28690 = n25246 & n25358;
  assign n28691 = ~n28689 & ~n28690;
  assign n28692 = n26478 & n28691;
  assign n28693 = n28688 & n28692;
  assign n28694 = n28680 & n28693;
  assign n28695 = n28674 & n28694;
  assign n28696 = n26528 & n28695;
  assign n28697 = n28616 & n28696;
  assign n28698 = n28613 & n28697;
  assign n28699 = pi3516 & ~n12516;
  assign n28700 = n28698 & ~n28699;
  assign n28701 = n25371 & ~n28700;
  assign n28702 = ~n28610 & ~n28701;
  assign n28703 = ~n16855 & n25508;
  assign n28704 = ~n12726 & n25512;
  assign n28705 = ~n28703 & ~n28704;
  assign n28706 = n28702 & n28705;
  assign n28707 = ~n12520 & n24922;
  assign n28708 = ~n12516 & n24925;
  assign n28709 = ~n28707 & ~n28708;
  assign n28710 = ~n12520 & n25462;
  assign n28711 = ~n12516 & n25465;
  assign n28712 = ~n28710 & ~n28711;
  assign n28713 = n28709 & n28712;
  assign n28714 = n19768 & n20379;
  assign n28715 = ~n19752 & n28714;
  assign n28716 = ~n19769 & ~n19810;
  assign n28717 = ~n20380 & n28716;
  assign n28718 = ~n28715 & ~n28717;
  assign n28719 = n19832 & ~n19848;
  assign n28720 = ~n20322 & ~n28719;
  assign n28721 = ~n19849 & ~n28720;
  assign n28722 = ~n20334 & ~n28721;
  assign n28723 = ~n28718 & ~n28722;
  assign n28724 = n28718 & n28722;
  assign n28725 = ~n28723 & ~n28724;
  assign n28726 = n24892 & ~n28725;
  assign n28727 = ~n12547 & ~n24905;
  assign n28728 = ~n12726 & n24916;
  assign n28729 = ~n16855 & n24913;
  assign n28730 = ~n28728 & ~n28729;
  assign n28731 = ~n24909 & n28730;
  assign n28732 = ~n28727 & n28731;
  assign n28733 = ~n28726 & n28732;
  assign n28734 = ~n12609 & n25474;
  assign n28735 = ~n25471 & ~n28734;
  assign n28736 = ~n12613 & ~n25483;
  assign n28737 = ~n12609 & n25473;
  assign n28738 = ~n28736 & ~n28737;
  assign n28739 = n27457 & n28738;
  assign n28740 = ~n25479 & n28739;
  assign n28741 = n28735 & n28740;
  assign n28742 = n27467 & ~n28741;
  assign n28743 = ~n27470 & ~n28742;
  assign n28744 = pi0342 & ~n28743;
  assign n28745 = n28733 & ~n28744;
  assign n28746 = pi0343 & ~n16855;
  assign n28747 = ~pi0343 & ~n12726;
  assign n28748 = ~n28746 & ~n28747;
  assign n28749 = n25458 & ~n28748;
  assign n28750 = ~n27441 & ~n28749;
  assign n28751 = n28745 & n28750;
  assign n28752 = n28713 & n28751;
  assign n28753 = n28706 & n28752;
  assign n28754 = n25544 & ~n28753;
  assign n28755 = ~pi0098 & n25533;
  assign n28756 = ~pi0139 & pi0979;
  assign n28757 = ~pi0141 & ~pi0979;
  assign n28758 = ~n28756 & ~n28757;
  assign n28759 = n25571 & ~n28758;
  assign n28760 = ~n12618 & ~n25582;
  assign n28761 = ~n12622 & n25582;
  assign n28762 = ~n28760 & ~n28761;
  assign n28763 = n25580 & ~n28762;
  assign n28764 = ~pi0098 & n25532;
  assign n28765 = ~n28763 & ~n28764;
  assign n28766 = n12627 & ~n25594;
  assign n28767 = n12631 & n25594;
  assign n28768 = ~n28766 & ~n28767;
  assign n28769 = n25591 & n28768;
  assign n28770 = n28765 & ~n28769;
  assign n28771 = ~n28759 & n28770;
  assign n28772 = n25606 & n28771;
  assign n28773 = n12726 & ~n25606;
  assign n28774 = ~n28772 & ~n28773;
  assign n28775 = n25564 & n28774;
  assign n28776 = ~n25606 & ~n28771;
  assign n28777 = ~n16855 & n25606;
  assign n28778 = ~n28776 & ~n28777;
  assign n28779 = ~n25564 & ~n28778;
  assign n28780 = ~n28775 & ~n28779;
  assign n28781 = ~n25533 & ~n28780;
  assign n28782 = ~n28755 & ~n28781;
  assign n28783 = ~n25544 & ~n28782;
  assign po0368 = n28754 | n28783;
  assign n28785 = n25097 & n25165;
  assign n28786 = n24932 & n25100;
  assign n28787 = ~n28785 & ~n28786;
  assign n28788 = n25158 & n25352;
  assign n28789 = n25267 & n25355;
  assign n28790 = ~n28788 & ~n28789;
  assign n28791 = n25202 & n25358;
  assign n28792 = n25230 & n25360;
  assign n28793 = ~n28791 & ~n28792;
  assign n28794 = n25032 & n25172;
  assign n28795 = n25169 & n25237;
  assign n28796 = ~n28794 & ~n28795;
  assign n28797 = n25209 & n25246;
  assign n28798 = ~n25208 & ~n28797;
  assign n28799 = n28796 & n28798;
  assign n28800 = n25041 & n25195;
  assign n28801 = n28799 & ~n28800;
  assign n28802 = n25160 & n25198;
  assign n28803 = n25162 & n25267;
  assign n28804 = ~n28802 & ~n28803;
  assign n28805 = n25103 & n25243;
  assign n28806 = n27867 & ~n28805;
  assign n28807 = n26536 & n28806;
  assign n28808 = n28804 & n28807;
  assign n28809 = n28801 & n28808;
  assign n28810 = n25290 & n25292;
  assign n28811 = n25032 & n25254;
  assign n28812 = ~n28810 & ~n28811;
  assign n28813 = n25264 & n25290;
  assign n28814 = n28812 & ~n28813;
  assign n28815 = n25158 & n25248;
  assign n28816 = n25149 & n25281;
  assign n28817 = ~n28815 & ~n28816;
  assign n28818 = n25149 & n25234;
  assign n28819 = n25198 & n25239;
  assign n28820 = ~n28818 & ~n28819;
  assign n28821 = n25227 & n28820;
  assign n28822 = n28817 & n28821;
  assign n28823 = n28814 & n28822;
  assign n28824 = n28809 & n28823;
  assign n28825 = n25326 & n28824;
  assign n28826 = n28793 & n28825;
  assign n28827 = n28790 & n28826;
  assign n28828 = n24932 & n25184;
  assign n28829 = n25142 & n25151;
  assign n28830 = ~n28828 & ~n28829;
  assign n28831 = n25036 & n25165;
  assign n28832 = n25028 & n25230;
  assign n28833 = ~n28831 & ~n28832;
  assign n28834 = n25076 & n25251;
  assign n28835 = n25078 & n25246;
  assign n28836 = ~n28834 & ~n28835;
  assign n28837 = n25064 & n25251;
  assign n28838 = n25070 & n25151;
  assign n28839 = ~n28837 & ~n28838;
  assign n28840 = n28836 & n28839;
  assign n28841 = n25093 & n28840;
  assign n28842 = n28833 & n28841;
  assign n28843 = ~n25180 & ~n25183;
  assign n28844 = ~n25178 & n28843;
  assign n28845 = ~n25139 & n28844;
  assign n28846 = n28842 & n28845;
  assign n28847 = n25146 & n25202;
  assign n28848 = n25153 & n25237;
  assign n28849 = ~n28847 & ~n28848;
  assign n28850 = n28846 & n28849;
  assign n28851 = n28830 & n28850;
  assign n28852 = n28827 & n28851;
  assign n28853 = n25041 & n25306;
  assign n28854 = n25103 & n25309;
  assign n28855 = ~n28853 & ~n28854;
  assign n28856 = n25349 & n28855;
  assign n28857 = pi3516 & ~n17018;
  assign n28858 = n28856 & ~n28857;
  assign n28859 = n28852 & n28858;
  assign n28860 = n28787 & n28859;
  assign n28861 = n25134 & n28860;
  assign n28862 = n25443 & ~n28861;
  assign n28863 = n25151 & n25270;
  assign n28864 = n25246 & n25261;
  assign n28865 = ~n28863 & ~n28864;
  assign n28866 = n25237 & n26519;
  assign n28867 = ~n27305 & ~n28866;
  assign n28868 = n28865 & n28867;
  assign n28869 = n25041 & n27288;
  assign n28870 = n28868 & ~n28869;
  assign n28871 = n25230 & n27253;
  assign n28872 = n25202 & n27250;
  assign n28873 = ~n28871 & ~n28872;
  assign n28874 = n25267 & n27256;
  assign n28875 = n27261 & ~n28874;
  assign n28876 = n28873 & n28875;
  assign n28877 = n25290 & n27219;
  assign n28878 = n28876 & ~n28877;
  assign n28879 = n25133 & n27223;
  assign n28880 = n25116 & n28879;
  assign n28881 = n28878 & n28880;
  assign n28882 = n25189 & n25251;
  assign n28883 = n25165 & n26453;
  assign n28884 = ~n28882 & ~n28883;
  assign n28885 = n25267 & n27193;
  assign n28886 = n25198 & n27196;
  assign n28887 = ~n28885 & ~n28886;
  assign n28888 = n24932 & n27200;
  assign n28889 = n27204 & ~n28888;
  assign n28890 = n28887 & n28889;
  assign n28891 = n25144 & n28890;
  assign n28892 = n27216 & n28891;
  assign n28893 = n25149 & n27209;
  assign n28894 = n25158 & n26448;
  assign n28895 = ~n28893 & ~n28894;
  assign n28896 = n28892 & n28895;
  assign n28897 = n28884 & n28896;
  assign n28898 = n28881 & n28897;
  assign n28899 = n25237 & n26459;
  assign n28900 = n26466 & ~n28899;
  assign n28901 = n25103 & n26457;
  assign n28902 = n25158 & n26462;
  assign n28903 = ~n28901 & ~n28902;
  assign n28904 = n25198 & n27236;
  assign n28905 = n28903 & ~n28904;
  assign n28906 = n25080 & n28905;
  assign n28907 = n28900 & n28906;
  assign n28908 = n25202 & n27246;
  assign n28909 = n25049 & n25251;
  assign n28910 = ~n28908 & ~n28909;
  assign n28911 = n25230 & n27243;
  assign n28912 = n27264 & ~n28911;
  assign n28913 = n28910 & n28912;
  assign n28914 = n28907 & n28913;
  assign n28915 = pi3516 & ~n17014;
  assign n28916 = n27191 & ~n28915;
  assign n28917 = n28914 & n28916;
  assign n28918 = n28898 & n28917;
  assign n28919 = n24932 & n27324;
  assign n28920 = n25231 & n25246;
  assign n28921 = ~n28919 & ~n28920;
  assign n28922 = n28665 & n28921;
  assign n28923 = n25151 & n25204;
  assign n28924 = n28922 & ~n28923;
  assign n28925 = n25149 & n27283;
  assign n28926 = n25103 & n26438;
  assign n28927 = ~n28925 & ~n28926;
  assign n28928 = n25290 & n27279;
  assign n28929 = n25041 & n27276;
  assign n28930 = ~n28928 & ~n28929;
  assign n28931 = n25032 & ~n26718;
  assign n28932 = n25165 & n26538;
  assign n28933 = ~n28931 & ~n28932;
  assign n28934 = ~n27315 & n28933;
  assign n28935 = n27275 & n28934;
  assign n28936 = n27308 & n28935;
  assign n28937 = n28930 & n28936;
  assign n28938 = n28927 & n28937;
  assign n28939 = n26507 & n27296;
  assign n28940 = n25211 & n28939;
  assign n28941 = n28938 & n28940;
  assign n28942 = n27293 & n28941;
  assign n28943 = ~n27299 & n28942;
  assign n28944 = n28924 & n28943;
  assign n28945 = n28918 & n28944;
  assign n28946 = n27340 & n28945;
  assign n28947 = n26528 & n28946;
  assign n28948 = n28870 & n28947;
  assign n28949 = n25371 & ~n28948;
  assign n28950 = ~n28862 & ~n28949;
  assign n28951 = ~n17105 & n25508;
  assign n28952 = ~n17199 & n25512;
  assign n28953 = ~n28951 & ~n28952;
  assign n28954 = n28950 & n28953;
  assign n28955 = ~n17018 & n24922;
  assign n28956 = ~n17014 & n24925;
  assign n28957 = ~n28955 & ~n28956;
  assign n28958 = ~n17018 & n25462;
  assign n28959 = ~n17014 & n25465;
  assign n28960 = ~n28958 & ~n28959;
  assign n28961 = n28957 & n28960;
  assign n28962 = ~n20327 & ~n20334;
  assign n28963 = n19693 & n20379;
  assign n28964 = ~n19693 & ~n20328;
  assign n28965 = ~n20380 & n28964;
  assign n28966 = ~n28963 & ~n28965;
  assign n28967 = n28962 & n28966;
  assign n28968 = ~n28962 & ~n28966;
  assign n28969 = ~n28967 & ~n28968;
  assign n28970 = n24892 & ~n28969;
  assign n28971 = ~n17045 & ~n24905;
  assign n28972 = ~n17105 & n24913;
  assign n28973 = ~n17199 & n24916;
  assign n28974 = ~n28972 & ~n28973;
  assign n28975 = ~n24909 & n28974;
  assign n28976 = ~n28971 & n28975;
  assign n28977 = ~n28970 & n28976;
  assign n28978 = ~n17071 & n25474;
  assign n28979 = ~n25471 & ~n28978;
  assign n28980 = ~n17071 & n25473;
  assign n28981 = ~n17075 & ~n25483;
  assign n28982 = ~n28980 & ~n28981;
  assign n28983 = n27457 & n28982;
  assign n28984 = ~n25479 & n28983;
  assign n28985 = n28979 & n28984;
  assign n28986 = n27467 & ~n28985;
  assign n28987 = ~n27470 & ~n28986;
  assign n28988 = pi0342 & ~n28987;
  assign n28989 = n28977 & ~n28988;
  assign n28990 = ~pi0343 & ~n17199;
  assign n28991 = pi0343 & ~n17105;
  assign n28992 = ~n28990 & ~n28991;
  assign n28993 = n25458 & ~n28992;
  assign n28994 = ~n27441 & ~n28993;
  assign n28995 = n28989 & n28994;
  assign n28996 = n28961 & n28995;
  assign n28997 = n28954 & n28996;
  assign n28998 = n25544 & ~n28997;
  assign n28999 = ~pi0099 & n25533;
  assign n29000 = ~pi0123 & pi0979;
  assign n29001 = ~pi0124 & ~pi0979;
  assign n29002 = ~n29000 & ~n29001;
  assign n29003 = n25571 & ~n29002;
  assign n29004 = ~n17062 & ~n25582;
  assign n29005 = ~n17066 & n25582;
  assign n29006 = ~n29004 & ~n29005;
  assign n29007 = n25580 & ~n29006;
  assign n29008 = ~pi0099 & n25532;
  assign n29009 = ~n29007 & ~n29008;
  assign n29010 = n17053 & ~n25594;
  assign n29011 = n17057 & n25594;
  assign n29012 = ~n29010 & ~n29011;
  assign n29013 = n25591 & n29012;
  assign n29014 = n29009 & ~n29013;
  assign n29015 = ~n29003 & n29014;
  assign n29016 = n25606 & ~n29015;
  assign n29017 = ~n17199 & ~n25606;
  assign n29018 = ~n29016 & ~n29017;
  assign n29019 = n25564 & ~n29018;
  assign n29020 = ~n17105 & n25606;
  assign n29021 = ~n25606 & ~n29015;
  assign n29022 = ~n29020 & ~n29021;
  assign n29023 = ~n25564 & ~n29022;
  assign n29024 = ~n29019 & ~n29023;
  assign n29025 = ~n25533 & ~n29024;
  assign n29026 = ~n28999 & ~n29025;
  assign n29027 = ~n25544 & ~n29026;
  assign po0369 = n28998 | n29027;
  assign n29029 = pi3516 & ~n9542;
  assign n29030 = n25097 & n25149;
  assign n29031 = n25100 & n25198;
  assign n29032 = ~n29030 & ~n29031;
  assign n29033 = n25134 & n29032;
  assign n29034 = n25032 & n25076;
  assign n29035 = n25078 & n25251;
  assign n29036 = ~n29034 & ~n29035;
  assign n29037 = n25032 & n25064;
  assign n29038 = n25070 & n25246;
  assign n29039 = ~n29037 & ~n29038;
  assign n29040 = n25036 & n25149;
  assign n29041 = n25028 & n25041;
  assign n29042 = ~n29040 & ~n29041;
  assign n29043 = n29039 & n29042;
  assign n29044 = n25093 & n29043;
  assign n29045 = n29036 & n29044;
  assign n29046 = n25146 & n25230;
  assign n29047 = n25103 & n25153;
  assign n29048 = ~n29046 & ~n29047;
  assign n29049 = n25290 & n25306;
  assign n29050 = n25158 & n25309;
  assign n29051 = ~n29049 & ~n29050;
  assign n29052 = n25349 & n29051;
  assign n29053 = n28845 & n29052;
  assign n29054 = n25184 & n25198;
  assign n29055 = n25142 & n25246;
  assign n29056 = ~n29054 & ~n29055;
  assign n29057 = n29053 & n29056;
  assign n29058 = n29048 & n29057;
  assign n29059 = n29045 & n29058;
  assign n29060 = n25151 & n25276;
  assign n29061 = n27867 & ~n29060;
  assign n29062 = n25160 & n25267;
  assign n29063 = n25162 & n25202;
  assign n29064 = ~n29062 & ~n29063;
  assign n29065 = n25195 & n25290;
  assign n29066 = n29064 & ~n29065;
  assign n29067 = n25151 & n25207;
  assign n29068 = n25209 & n25251;
  assign n29069 = ~n29067 & ~n29068;
  assign n29070 = n29066 & n29069;
  assign n29071 = n25172 & n25237;
  assign n29072 = n25103 & n25169;
  assign n29073 = ~n29071 & ~n29072;
  assign n29074 = n29070 & n29073;
  assign n29075 = ~n25285 & n29074;
  assign n29076 = n29061 & n29075;
  assign n29077 = n25237 & n25254;
  assign n29078 = n24932 & n25281;
  assign n29079 = ~n29077 & ~n29078;
  assign n29080 = n25158 & n25243;
  assign n29081 = n25165 & n25248;
  assign n29082 = ~n29080 & ~n29081;
  assign n29083 = n29079 & n29082;
  assign n29084 = n29076 & n29083;
  assign n29085 = n24932 & n25234;
  assign n29086 = n25239 & n25267;
  assign n29087 = ~n29085 & ~n29086;
  assign n29088 = n25326 & n29087;
  assign n29089 = n25227 & n29088;
  assign n29090 = n29084 & n29089;
  assign n29091 = n25230 & n25358;
  assign n29092 = n25041 & n25360;
  assign n29093 = ~n29091 & ~n29092;
  assign n29094 = n25165 & n25352;
  assign n29095 = n25202 & n25355;
  assign n29096 = ~n29094 & ~n29095;
  assign n29097 = n29093 & n29096;
  assign n29098 = n29090 & n29097;
  assign n29099 = n29059 & n29098;
  assign n29100 = n29033 & n29099;
  assign n29101 = ~n29029 & n29100;
  assign n29102 = n25443 & ~n29101;
  assign n29103 = pi3516 & ~n9538;
  assign n29104 = n24932 & n27209;
  assign n29105 = n25165 & n26448;
  assign n29106 = ~n29104 & ~n29105;
  assign n29107 = n25032 & n25189;
  assign n29108 = n25149 & n26453;
  assign n29109 = ~n29107 & ~n29108;
  assign n29110 = n27216 & n29109;
  assign n29111 = n29106 & n29110;
  assign n29112 = n25198 & n27200;
  assign n29113 = n29111 & ~n29112;
  assign n29114 = n25202 & n27193;
  assign n29115 = n25267 & n27196;
  assign n29116 = ~n29114 & ~n29115;
  assign n29117 = n27204 & n29116;
  assign n29118 = n25144 & n29117;
  assign n29119 = n29113 & n29118;
  assign n29120 = n25041 & n27243;
  assign n29121 = n29119 & ~n29120;
  assign n29122 = n25202 & n27256;
  assign n29123 = n25041 & n27253;
  assign n29124 = ~n29122 & ~n29123;
  assign n29125 = n25230 & n27250;
  assign n29126 = n29124 & ~n29125;
  assign n29127 = n27260 & n28429;
  assign n29128 = n28428 & n29127;
  assign n29129 = ~n27259 & n29128;
  assign n29130 = n29126 & n29129;
  assign n29131 = n25116 & n27223;
  assign n29132 = ~n25131 & ~n25328;
  assign n29133 = n29131 & n29132;
  assign n29134 = n25124 & n29133;
  assign n29135 = n29130 & n29134;
  assign n29136 = n25198 & n27324;
  assign n29137 = n25231 & n25251;
  assign n29138 = ~n29136 & ~n29137;
  assign n29139 = n25204 & n25246;
  assign n29140 = ~n27299 & ~n29139;
  assign n29141 = n29138 & n29140;
  assign n29142 = n28665 & n29141;
  assign n29143 = n25149 & n26538;
  assign n29144 = n25237 & n25296;
  assign n29145 = ~n29143 & ~n29144;
  assign n29146 = n25290 & n27276;
  assign n29147 = n27275 & ~n29146;
  assign n29148 = n24932 & n27283;
  assign n29149 = n25158 & n26438;
  assign n29150 = ~n29148 & ~n29149;
  assign n29151 = n29147 & n29150;
  assign n29152 = n27308 & n29151;
  assign n29153 = n25237 & n25287;
  assign n29154 = n25151 & n25292;
  assign n29155 = ~n29153 & ~n29154;
  assign n29156 = n29152 & n29155;
  assign n29157 = n29145 & n29156;
  assign n29158 = n29142 & n29157;
  assign n29159 = n29135 & n29158;
  assign n29160 = n27293 & n29159;
  assign n29161 = n28940 & n29160;
  assign n29162 = n25103 & n26459;
  assign n29163 = n26466 & ~n29162;
  assign n29164 = n25080 & n29163;
  assign n29165 = n25267 & n27236;
  assign n29166 = n29164 & ~n29165;
  assign n29167 = n25158 & n26457;
  assign n29168 = n25165 & n26462;
  assign n29169 = ~n29167 & ~n29168;
  assign n29170 = n25151 & n25264;
  assign n29171 = n25246 & n25270;
  assign n29172 = ~n29170 & ~n29171;
  assign n29173 = n25103 & n26519;
  assign n29174 = n25251 & n25261;
  assign n29175 = ~n29173 & ~n29174;
  assign n29176 = n26528 & n29175;
  assign n29177 = n29172 & n29176;
  assign n29178 = n25290 & n27288;
  assign n29179 = n29177 & ~n29178;
  assign n29180 = n27340 & n29179;
  assign n29181 = n29169 & n29180;
  assign n29182 = n29166 & n29181;
  assign n29183 = n29161 & n29182;
  assign n29184 = n25230 & n27246;
  assign n29185 = n25032 & n25049;
  assign n29186 = ~n29184 & ~n29185;
  assign n29187 = n27264 & n29186;
  assign n29188 = n29183 & n29187;
  assign n29189 = n29121 & n29188;
  assign n29190 = ~n29103 & n29189;
  assign n29191 = n25371 & ~n29190;
  assign n29192 = ~n29102 & ~n29191;
  assign n29193 = ~n9825 & n25512;
  assign n29194 = ~n16999 & n25508;
  assign n29195 = ~n29193 & ~n29194;
  assign n29196 = n29192 & n29195;
  assign n29197 = ~n9542 & n24922;
  assign n29198 = ~n9538 & n24925;
  assign n29199 = ~n29197 & ~n29198;
  assign n29200 = ~n9542 & n25462;
  assign n29201 = ~n9538 & n25465;
  assign n29202 = ~n29200 & ~n29201;
  assign n29203 = n29199 & n29202;
  assign n29204 = n19855 & ~n20324;
  assign n29205 = ~n19935 & ~n29204;
  assign n29206 = ~n19943 & ~n29205;
  assign n29207 = ~n20334 & ~n29206;
  assign n29208 = n19945 & n20379;
  assign n29209 = ~n19878 & n19896;
  assign n29210 = n19878 & ~n19896;
  assign n29211 = ~n29209 & ~n29210;
  assign n29212 = ~n20380 & ~n29211;
  assign n29213 = ~n29208 & ~n29212;
  assign n29214 = n29207 & ~n29213;
  assign n29215 = ~n29207 & n29213;
  assign n29216 = ~n29214 & ~n29215;
  assign n29217 = n24892 & n29216;
  assign n29218 = ~n9570 & ~n24905;
  assign n29219 = ~n9825 & n24916;
  assign n29220 = ~n16999 & n24913;
  assign n29221 = ~n29219 & ~n29220;
  assign n29222 = ~n24909 & n29221;
  assign n29223 = ~n29218 & n29222;
  assign n29224 = ~n29217 & n29223;
  assign n29225 = ~n9511 & n25474;
  assign n29226 = ~n25471 & ~n29225;
  assign n29227 = ~n9511 & n25473;
  assign n29228 = ~n9515 & ~n25483;
  assign n29229 = ~n29227 & ~n29228;
  assign n29230 = n27457 & n29229;
  assign n29231 = ~n25479 & n29230;
  assign n29232 = n29226 & n29231;
  assign n29233 = n27467 & ~n29232;
  assign n29234 = ~n27470 & ~n29233;
  assign n29235 = pi0342 & ~n29234;
  assign n29236 = n29224 & ~n29235;
  assign n29237 = pi0343 & ~n16999;
  assign n29238 = ~pi0343 & ~n9825;
  assign n29239 = ~n29237 & ~n29238;
  assign n29240 = n25458 & ~n29239;
  assign n29241 = ~n27441 & ~n29240;
  assign n29242 = n29236 & n29241;
  assign n29243 = n29203 & n29242;
  assign n29244 = n29196 & n29243;
  assign n29245 = n25544 & ~n29244;
  assign n29246 = ~pi0100 & n25533;
  assign n29247 = ~pi0121 & pi0979;
  assign n29248 = ~pi0125 & ~pi0979;
  assign n29249 = ~n29247 & ~n29248;
  assign n29250 = n25571 & ~n29249;
  assign n29251 = ~n9502 & ~n25582;
  assign n29252 = ~n9506 & n25582;
  assign n29253 = ~n29251 & ~n29252;
  assign n29254 = n25580 & ~n29253;
  assign n29255 = ~pi0100 & n25532;
  assign n29256 = ~n29254 & ~n29255;
  assign n29257 = n9489 & ~n25594;
  assign n29258 = n9493 & n25594;
  assign n29259 = ~n29257 & ~n29258;
  assign n29260 = n25591 & n29259;
  assign n29261 = n29256 & ~n29260;
  assign n29262 = ~n29250 & n29261;
  assign n29263 = n25606 & n29262;
  assign n29264 = n9825 & ~n25606;
  assign n29265 = ~n29263 & ~n29264;
  assign n29266 = n25564 & n29265;
  assign n29267 = ~n16999 & n25606;
  assign n29268 = ~n25606 & ~n29262;
  assign n29269 = ~n29267 & ~n29268;
  assign n29270 = ~n25564 & ~n29269;
  assign n29271 = ~n29266 & ~n29270;
  assign n29272 = ~n25533 & ~n29271;
  assign n29273 = ~n29246 & ~n29272;
  assign n29274 = ~n25544 & ~n29273;
  assign po0370 = n29245 | n29274;
  assign n29276 = n25267 & n27324;
  assign n29277 = n25032 & n25231;
  assign n29278 = ~n29276 & ~n29277;
  assign n29279 = n24932 & n26538;
  assign n29280 = n25103 & n25296;
  assign n29281 = ~n29279 & ~n29280;
  assign n29282 = n25103 & n25287;
  assign n29283 = n25246 & n25292;
  assign n29284 = ~n29282 & ~n29283;
  assign n29285 = n25204 & n25251;
  assign n29286 = n25211 & n27296;
  assign n29287 = n26507 & n29286;
  assign n29288 = ~n29285 & n29287;
  assign n29289 = n25165 & n26438;
  assign n29290 = ~n27272 & ~n29289;
  assign n29291 = n26478 & n27293;
  assign n29292 = n25290 & n27243;
  assign n29293 = n25041 & n27246;
  assign n29294 = ~n29292 & ~n29293;
  assign n29295 = n25158 & n26459;
  assign n29296 = n26466 & ~n29295;
  assign n29297 = n25165 & n26457;
  assign n29298 = n25149 & n26462;
  assign n29299 = ~n29297 & ~n29298;
  assign n29300 = n25202 & n27236;
  assign n29301 = n29299 & ~n29300;
  assign n29302 = n25080 & n29301;
  assign n29303 = n29296 & n29302;
  assign n29304 = n25049 & n25237;
  assign n29305 = n29303 & ~n29304;
  assign n29306 = n27264 & n29305;
  assign n29307 = n29294 & n29306;
  assign n29308 = n25198 & n27283;
  assign n29309 = n29307 & ~n29308;
  assign n29310 = n29291 & n29309;
  assign n29311 = n29290 & n29310;
  assign n29312 = n25316 & n29311;
  assign n29313 = n25151 & n25195;
  assign n29314 = n29312 & ~n29313;
  assign n29315 = n25290 & n27253;
  assign n29316 = n25041 & n27250;
  assign n29317 = ~n29315 & ~n29316;
  assign n29318 = n25230 & n27256;
  assign n29319 = n29317 & ~n29318;
  assign n29320 = n25151 & n25306;
  assign n29321 = n29319 & ~n29320;
  assign n29322 = n25124 & n27260;
  assign n29323 = n28428 & n29322;
  assign n29324 = n29321 & n29323;
  assign n29325 = n29131 & n29324;
  assign n29326 = n29314 & n29325;
  assign n29327 = n29132 & n29326;
  assign n29328 = n28429 & n29327;
  assign n29329 = n29288 & n29328;
  assign n29330 = n25246 & n25264;
  assign n29331 = n25251 & n25270;
  assign n29332 = ~n29330 & ~n29331;
  assign n29333 = n25158 & n26519;
  assign n29334 = n25032 & n25261;
  assign n29335 = ~n29333 & ~n29334;
  assign n29336 = n26528 & n29335;
  assign n29337 = n29332 & n29336;
  assign n29338 = n27308 & n29337;
  assign n29339 = n29329 & n29338;
  assign n29340 = n29284 & n29339;
  assign n29341 = n29281 & n29340;
  assign n29342 = n25189 & n25237;
  assign n29343 = n24932 & n26453;
  assign n29344 = ~n29342 & ~n29343;
  assign n29345 = n25198 & n27209;
  assign n29346 = n25149 & n26448;
  assign n29347 = ~n29345 & ~n29346;
  assign n29348 = n27216 & n29347;
  assign n29349 = n29344 & n29348;
  assign n29350 = n25267 & n27200;
  assign n29351 = n29349 & ~n29350;
  assign n29352 = n25230 & n27193;
  assign n29353 = n25202 & n27196;
  assign n29354 = ~n29352 & ~n29353;
  assign n29355 = n27204 & n29354;
  assign n29356 = n25144 & n29355;
  assign n29357 = n29351 & n29356;
  assign n29358 = n29341 & n29357;
  assign n29359 = n25227 & n29358;
  assign n29360 = n27323 & n29359;
  assign n29361 = n29278 & n29360;
  assign n29362 = pi3516 & ~n10456;
  assign n29363 = n29361 & ~n29362;
  assign n29364 = n25371 & ~n29363;
  assign n29365 = n24932 & n25036;
  assign n29366 = n25028 & n25290;
  assign n29367 = ~n29365 & ~n29366;
  assign n29368 = n25041 & n25146;
  assign n29369 = n25153 & n25158;
  assign n29370 = ~n29368 & ~n29369;
  assign n29371 = n25184 & n25267;
  assign n29372 = n25142 & n25251;
  assign n29373 = ~n29371 & ~n29372;
  assign n29374 = n25064 & n25237;
  assign n29375 = n25070 & n25251;
  assign n29376 = ~n29374 & ~n29375;
  assign n29377 = n25151 & ~n26802;
  assign n29378 = n25322 & ~n29377;
  assign n29379 = n25041 & n25358;
  assign n29380 = n25290 & n25360;
  assign n29381 = ~n29379 & ~n29380;
  assign n29382 = n25149 & n25352;
  assign n29383 = n25230 & n25355;
  assign n29384 = ~n29382 & ~n29383;
  assign n29385 = n29381 & n29384;
  assign n29386 = ~n25313 & n29385;
  assign n29387 = n29378 & n29386;
  assign n29388 = n28845 & n29387;
  assign n29389 = n29376 & n29388;
  assign n29390 = n29373 & n29389;
  assign n29391 = n29370 & n29390;
  assign n29392 = n25198 & n25234;
  assign n29393 = n25202 & n25239;
  assign n29394 = ~n29392 & ~n29393;
  assign n29395 = n24932 & n25097;
  assign n29396 = n25100 & n25267;
  assign n29397 = ~n29395 & ~n29396;
  assign n29398 = n25134 & n29397;
  assign n29399 = n25246 & n25276;
  assign n29400 = n27867 & ~n29399;
  assign n29401 = n25103 & n25172;
  assign n29402 = n25207 & n25246;
  assign n29403 = ~n29401 & ~n29402;
  assign n29404 = n25032 & n25209;
  assign n29405 = n29403 & ~n29404;
  assign n29406 = n25162 & n25230;
  assign n29407 = n29405 & ~n29406;
  assign n29408 = n25158 & n25169;
  assign n29409 = n25160 & n25202;
  assign n29410 = ~n29408 & ~n29409;
  assign n29411 = n29407 & n29410;
  assign n29412 = ~n25285 & n29411;
  assign n29413 = n29400 & n29412;
  assign n29414 = n25103 & n25254;
  assign n29415 = n25198 & n25281;
  assign n29416 = ~n29414 & ~n29415;
  assign n29417 = n25165 & n25243;
  assign n29418 = n25149 & n25248;
  assign n29419 = ~n29417 & ~n29418;
  assign n29420 = n29416 & n29419;
  assign n29421 = n29413 & n29420;
  assign n29422 = n29398 & n29421;
  assign n29423 = n29394 & n29422;
  assign n29424 = n25227 & n29423;
  assign n29425 = n25165 & n25309;
  assign n29426 = n29424 & ~n29425;
  assign n29427 = n25343 & n29426;
  assign n29428 = n25348 & n29427;
  assign n29429 = n29391 & n29428;
  assign n29430 = n25076 & n25237;
  assign n29431 = n25032 & n25078;
  assign n29432 = ~n29430 & ~n29431;
  assign n29433 = n29429 & n29432;
  assign n29434 = n25093 & n29433;
  assign n29435 = n29367 & n29434;
  assign n29436 = pi3516 & ~n10460;
  assign n29437 = n29435 & ~n29436;
  assign n29438 = n25443 & ~n29437;
  assign n29439 = ~n29364 & ~n29438;
  assign n29440 = ~n16963 & n25508;
  assign n29441 = ~n10608 & n25512;
  assign n29442 = ~n29440 & ~n29441;
  assign n29443 = n29439 & n29442;
  assign n29444 = ~n10460 & n24922;
  assign n29445 = ~n10456 & n24925;
  assign n29446 = ~n29444 & ~n29445;
  assign n29447 = ~n10460 & n25462;
  assign n29448 = ~n10456 & n25465;
  assign n29449 = ~n29447 & ~n29448;
  assign n29450 = n29446 & n29449;
  assign n29451 = ~n20334 & ~n29204;
  assign n29452 = n19943 & n20379;
  assign n29453 = ~n19935 & ~n19943;
  assign n29454 = ~n20380 & n29453;
  assign n29455 = ~n29452 & ~n29454;
  assign n29456 = n29451 & n29455;
  assign n29457 = ~n29451 & ~n29455;
  assign n29458 = ~n29456 & ~n29457;
  assign n29459 = n24892 & ~n29458;
  assign n29460 = ~n10487 & ~n24905;
  assign n29461 = ~n16963 & n24913;
  assign n29462 = ~n10608 & n24916;
  assign n29463 = ~n29461 & ~n29462;
  assign n29464 = ~n24909 & n29463;
  assign n29465 = ~n29460 & n29464;
  assign n29466 = ~n29459 & n29465;
  assign n29467 = ~n10420 & n25474;
  assign n29468 = ~n25471 & ~n29467;
  assign n29469 = ~n10420 & n25473;
  assign n29470 = ~n10424 & ~n25483;
  assign n29471 = ~n29469 & ~n29470;
  assign n29472 = n27457 & n29471;
  assign n29473 = ~n25479 & n29472;
  assign n29474 = n29468 & n29473;
  assign n29475 = n27467 & ~n29474;
  assign n29476 = ~n27470 & ~n29475;
  assign n29477 = pi0342 & ~n29476;
  assign n29478 = n29466 & ~n29477;
  assign n29479 = pi0343 & ~n16963;
  assign n29480 = ~pi0343 & ~n10608;
  assign n29481 = ~n29479 & ~n29480;
  assign n29482 = n25458 & ~n29481;
  assign n29483 = ~n27441 & ~n29482;
  assign n29484 = n29478 & n29483;
  assign n29485 = n29450 & n29484;
  assign n29486 = n29443 & n29485;
  assign n29487 = n25544 & ~n29486;
  assign n29488 = ~pi0101 & n25533;
  assign n29489 = ~pi0122 & pi0979;
  assign n29490 = ~pi0126 & ~pi0979;
  assign n29491 = ~n29489 & ~n29490;
  assign n29492 = n25571 & ~n29491;
  assign n29493 = ~n10429 & ~n25582;
  assign n29494 = ~n10433 & n25582;
  assign n29495 = ~n29493 & ~n29494;
  assign n29496 = n25580 & ~n29495;
  assign n29497 = ~pi0101 & n25532;
  assign n29498 = ~n29496 & ~n29497;
  assign n29499 = n10438 & ~n25594;
  assign n29500 = n10442 & n25594;
  assign n29501 = ~n29499 & ~n29500;
  assign n29502 = n25591 & n29501;
  assign n29503 = n29498 & ~n29502;
  assign n29504 = ~n29492 & n29503;
  assign n29505 = n25606 & ~n29504;
  assign n29506 = ~n10608 & ~n25606;
  assign n29507 = ~n29505 & ~n29506;
  assign n29508 = n25564 & ~n29507;
  assign n29509 = ~n16963 & n25606;
  assign n29510 = ~n25606 & ~n29504;
  assign n29511 = ~n29509 & ~n29510;
  assign n29512 = ~n25564 & ~n29511;
  assign n29513 = ~n29508 & ~n29512;
  assign n29514 = ~n25533 & ~n29513;
  assign n29515 = ~n29488 & ~n29514;
  assign n29516 = ~n25544 & ~n29515;
  assign po0371 = n29487 | n29516;
  assign n29518 = n25195 & n25246;
  assign n29519 = n29287 & ~n29518;
  assign n29520 = n25202 & n27324;
  assign n29521 = n25231 & n25237;
  assign n29522 = ~n29520 & ~n29521;
  assign n29523 = n25165 & n26459;
  assign n29524 = n26466 & ~n29523;
  assign n29525 = n25080 & n29524;
  assign n29526 = n25230 & n27236;
  assign n29527 = n29525 & ~n29526;
  assign n29528 = n25149 & n26457;
  assign n29529 = n24932 & n26462;
  assign n29530 = ~n29528 & ~n29529;
  assign n29531 = n24932 & n26448;
  assign n29532 = n25198 & n26453;
  assign n29533 = n25267 & n27209;
  assign n29534 = ~n29532 & ~n29533;
  assign n29535 = n25133 & ~n27214;
  assign n29536 = n29534 & n29535;
  assign n29537 = ~n29531 & n29536;
  assign n29538 = n25103 & n25189;
  assign n29539 = n25181 & ~n29538;
  assign n29540 = ~n25183 & n29539;
  assign n29541 = n29537 & n29540;
  assign n29542 = n25290 & n27250;
  assign n29543 = n25246 & n25306;
  assign n29544 = ~n29542 & ~n29543;
  assign n29545 = ~n25332 & n29544;
  assign n29546 = ~n26481 & n29545;
  assign n29547 = n25041 & n27256;
  assign n29548 = n29546 & ~n29547;
  assign n29549 = ~n25335 & ~n25346;
  assign n29550 = ~n25328 & n29549;
  assign n29551 = n29548 & n29550;
  assign n29552 = n25341 & ~n25347;
  assign n29553 = ~n25330 & n29552;
  assign n29554 = n29551 & n29553;
  assign n29555 = n29541 & n29554;
  assign n29556 = n29530 & n29555;
  assign n29557 = n29527 & n29556;
  assign n29558 = n25290 & n27246;
  assign n29559 = n25049 & n25103;
  assign n29560 = ~n29558 & ~n29559;
  assign n29561 = n25028 & n25151;
  assign n29562 = n26774 & ~n29561;
  assign n29563 = n29560 & n29562;
  assign n29564 = n25202 & n27200;
  assign n29565 = n29563 & ~n29564;
  assign n29566 = n25041 & n27193;
  assign n29567 = n25230 & n27196;
  assign n29568 = ~n29566 & ~n29567;
  assign n29569 = n27204 & n29568;
  assign n29570 = n25144 & n29569;
  assign n29571 = n29565 & n29570;
  assign n29572 = n29557 & n29571;
  assign n29573 = n25149 & n26438;
  assign n29574 = n25151 & n25360;
  assign n29575 = ~n29573 & ~n29574;
  assign n29576 = n25316 & n29575;
  assign n29577 = n25267 & n27283;
  assign n29578 = n29576 & ~n29577;
  assign n29579 = n29291 & n29578;
  assign n29580 = n29131 & n29579;
  assign n29581 = n29572 & n29580;
  assign n29582 = n25032 & n25204;
  assign n29583 = n29581 & ~n29582;
  assign n29584 = n25158 & n25287;
  assign n29585 = n25251 & n25292;
  assign n29586 = ~n29584 & ~n29585;
  assign n29587 = n25165 & n26519;
  assign n29588 = n25237 & n25261;
  assign n29589 = ~n29587 & ~n29588;
  assign n29590 = n25251 & n25264;
  assign n29591 = n25032 & n25270;
  assign n29592 = ~n29590 & ~n29591;
  assign n29593 = n26528 & n29592;
  assign n29594 = n29589 & n29593;
  assign n29595 = n27308 & n29594;
  assign n29596 = n25198 & n26538;
  assign n29597 = n25158 & n25296;
  assign n29598 = ~n29596 & ~n29597;
  assign n29599 = n29595 & n29598;
  assign n29600 = n29586 & n29599;
  assign n29601 = n25227 & n29600;
  assign n29602 = n29583 & n29601;
  assign n29603 = n27323 & n29602;
  assign n29604 = n29522 & n29603;
  assign n29605 = n29519 & n29604;
  assign n29606 = pi3516 & ~n15277;
  assign n29607 = n29605 & ~n29606;
  assign n29608 = n25371 & ~n29607;
  assign n29609 = n25234 & n25267;
  assign n29610 = n25230 & n25239;
  assign n29611 = ~n29609 & ~n29610;
  assign n29612 = n25097 & n25198;
  assign n29613 = n25100 & n25202;
  assign n29614 = ~n29612 & ~n29613;
  assign n29615 = n25134 & n29614;
  assign n29616 = n25251 & n25276;
  assign n29617 = n27867 & ~n29616;
  assign n29618 = n25165 & n25169;
  assign n29619 = n25160 & n25230;
  assign n29620 = ~n29618 & ~n29619;
  assign n29621 = n25041 & n25162;
  assign n29622 = n29620 & ~n29621;
  assign n29623 = n25158 & n25172;
  assign n29624 = n29622 & ~n29623;
  assign n29625 = n25207 & n25251;
  assign n29626 = n25209 & n25237;
  assign n29627 = ~n29625 & ~n29626;
  assign n29628 = n29624 & n29627;
  assign n29629 = ~n25285 & n29628;
  assign n29630 = n29617 & n29629;
  assign n29631 = n25149 & n25243;
  assign n29632 = n24932 & n25248;
  assign n29633 = ~n29631 & ~n29632;
  assign n29634 = n25158 & n25254;
  assign n29635 = n25267 & n25281;
  assign n29636 = ~n29634 & ~n29635;
  assign n29637 = n29633 & n29636;
  assign n29638 = n29630 & n29637;
  assign n29639 = n29615 & n29638;
  assign n29640 = n29611 & n29639;
  assign n29641 = n25227 & n29640;
  assign n29642 = n25149 & n25309;
  assign n29643 = n29641 & ~n29642;
  assign n29644 = n25246 & n25323;
  assign n29645 = n25151 & n25320;
  assign n29646 = ~n29644 & ~n29645;
  assign n29647 = n25041 & n25355;
  assign n29648 = n25290 & n25358;
  assign n29649 = ~n29647 & ~n29648;
  assign n29650 = n24932 & n25352;
  assign n29651 = n25246 & n25314;
  assign n29652 = ~n29650 & ~n29651;
  assign n29653 = n29649 & n29652;
  assign n29654 = n26599 & n29653;
  assign n29655 = n29646 & n29654;
  assign n29656 = n25064 & n25103;
  assign n29657 = n25032 & n25070;
  assign n29658 = ~n29656 & ~n29657;
  assign n29659 = n25036 & n25198;
  assign n29660 = n25078 & n25237;
  assign n29661 = ~n29659 & ~n29660;
  assign n29662 = n25076 & n25103;
  assign n29663 = n29661 & ~n29662;
  assign n29664 = n25093 & n29663;
  assign n29665 = n29658 & n29664;
  assign n29666 = n29655 & n29665;
  assign n29667 = n25343 & n29666;
  assign n29668 = n25348 & n29667;
  assign n29669 = n29643 & n29668;
  assign n29670 = n25151 & n25177;
  assign n29671 = n27883 & ~n29670;
  assign n29672 = n25146 & n25290;
  assign n29673 = n25153 & n25165;
  assign n29674 = ~n29672 & ~n29673;
  assign n29675 = n25184 & n25202;
  assign n29676 = n25032 & n25142;
  assign n29677 = ~n29675 & ~n29676;
  assign n29678 = n29674 & n29677;
  assign n29679 = ~n25183 & n29678;
  assign n29680 = n29671 & n29679;
  assign n29681 = n29669 & n29680;
  assign n29682 = pi3516 & ~n15281;
  assign n29683 = n29681 & ~n29682;
  assign n29684 = n25443 & ~n29683;
  assign n29685 = ~n29608 & ~n29684;
  assign n29686 = ~n15426 & n25512;
  assign n29687 = ~n16927 & n25508;
  assign n29688 = ~n29686 & ~n29687;
  assign n29689 = n29685 & n29688;
  assign n29690 = ~n15281 & n24922;
  assign n29691 = ~n15277 & n24925;
  assign n29692 = ~n29690 & ~n29691;
  assign n29693 = ~n15281 & n25462;
  assign n29694 = ~n15277 & n25465;
  assign n29695 = ~n29693 & ~n29694;
  assign n29696 = n29692 & n29695;
  assign n29697 = n19730 & n20379;
  assign n29698 = n19714 & n29697;
  assign n29699 = ~n19731 & ~n19811;
  assign n29700 = ~n20380 & n29699;
  assign n29701 = ~n29698 & ~n29700;
  assign n29702 = n19851 & ~n20323;
  assign n29703 = ~n19852 & ~n29702;
  assign n29704 = ~n19807 & ~n29703;
  assign n29705 = ~n20334 & ~n29704;
  assign n29706 = ~n29701 & n29705;
  assign n29707 = n29701 & ~n29705;
  assign n29708 = ~n29706 & ~n29707;
  assign n29709 = n24892 & n29708;
  assign n29710 = ~n15308 & ~n24905;
  assign n29711 = ~n15426 & n24916;
  assign n29712 = ~n16927 & n24913;
  assign n29713 = ~n29711 & ~n29712;
  assign n29714 = ~n24909 & n29713;
  assign n29715 = ~n29710 & n29714;
  assign n29716 = ~n29709 & n29715;
  assign n29717 = ~n15259 & n25474;
  assign n29718 = ~n25471 & ~n29717;
  assign n29719 = ~n15259 & n25473;
  assign n29720 = ~n15263 & ~n25483;
  assign n29721 = ~n29719 & ~n29720;
  assign n29722 = n27457 & n29721;
  assign n29723 = ~n25479 & n29722;
  assign n29724 = n29718 & n29723;
  assign n29725 = n27467 & ~n29724;
  assign n29726 = ~n27470 & ~n29725;
  assign n29727 = pi0342 & ~n29726;
  assign n29728 = n29716 & ~n29727;
  assign n29729 = pi0343 & ~n16927;
  assign n29730 = ~pi0343 & ~n15426;
  assign n29731 = ~n29729 & ~n29730;
  assign n29732 = n25458 & ~n29731;
  assign n29733 = ~n27441 & ~n29732;
  assign n29734 = n29728 & n29733;
  assign n29735 = n29696 & n29734;
  assign n29736 = n29689 & n29735;
  assign n29737 = n25544 & ~n29736;
  assign n29738 = ~pi0102 & n25533;
  assign n29739 = ~pi0090 & pi0979;
  assign n29740 = ~pi0093 & ~pi0979;
  assign n29741 = ~n29739 & ~n29740;
  assign n29742 = n25571 & ~n29741;
  assign n29743 = ~n15250 & ~n25582;
  assign n29744 = ~n15254 & n25582;
  assign n29745 = ~n29743 & ~n29744;
  assign n29746 = n25580 & ~n29745;
  assign n29747 = ~pi0102 & n25532;
  assign n29748 = ~n29746 & ~n29747;
  assign n29749 = n15241 & ~n25594;
  assign n29750 = n15245 & n25594;
  assign n29751 = ~n29749 & ~n29750;
  assign n29752 = n25591 & n29751;
  assign n29753 = n29748 & ~n29752;
  assign n29754 = ~n29742 & n29753;
  assign n29755 = n25606 & n29754;
  assign n29756 = n15426 & ~n25606;
  assign n29757 = ~n29755 & ~n29756;
  assign n29758 = n25564 & n29757;
  assign n29759 = ~n16927 & n25606;
  assign n29760 = ~n25606 & ~n29754;
  assign n29761 = ~n29759 & ~n29760;
  assign n29762 = ~n25564 & ~n29761;
  assign n29763 = ~n29758 & ~n29762;
  assign n29764 = ~n25533 & ~n29763;
  assign n29765 = ~n29738 & ~n29764;
  assign n29766 = ~n25544 & ~n29765;
  assign po0372 = n29737 | n29766;
  assign n29768 = n25149 & n26519;
  assign n29769 = n26527 & ~n29768;
  assign n29770 = n25237 & n25270;
  assign n29771 = n25103 & n25261;
  assign n29772 = ~n29770 & ~n29771;
  assign n29773 = n25032 & n25264;
  assign n29774 = n29772 & ~n29773;
  assign n29775 = ~n25258 & n29774;
  assign n29776 = ~n26524 & n29775;
  assign n29777 = n29769 & n29776;
  assign n29778 = n25230 & n27324;
  assign n29779 = n25103 & n25231;
  assign n29780 = ~n29778 & ~n29779;
  assign n29781 = n25202 & n27283;
  assign n29782 = n26477 & ~n29781;
  assign n29783 = n25151 & n25358;
  assign n29784 = n25246 & n25360;
  assign n29785 = ~n29783 & ~n29784;
  assign n29786 = ~n27291 & n29785;
  assign n29787 = ~n25313 & n29786;
  assign n29788 = n24932 & n26438;
  assign n29789 = n29787 & ~n29788;
  assign n29790 = n25204 & n25237;
  assign n29791 = n27296 & ~n29790;
  assign n29792 = n26507 & n29791;
  assign n29793 = n25195 & n25251;
  assign n29794 = n29792 & ~n29793;
  assign n29795 = n25211 & n29794;
  assign n29796 = ~n25315 & n29795;
  assign n29797 = n29789 & n29796;
  assign n29798 = n25146 & n25151;
  assign n29799 = n25181 & ~n29798;
  assign n29800 = n25202 & n27209;
  assign n29801 = n25198 & n26448;
  assign n29802 = ~n29800 & ~n29801;
  assign n29803 = n25158 & n25189;
  assign n29804 = n25267 & n26453;
  assign n29805 = ~n29803 & ~n29804;
  assign n29806 = n29802 & n29805;
  assign n29807 = ~n25183 & n29806;
  assign n29808 = n29799 & n29807;
  assign n29809 = n25088 & n29808;
  assign n29810 = n25049 & n25158;
  assign n29811 = n25028 & n25246;
  assign n29812 = ~n29810 & ~n29811;
  assign n29813 = n29809 & n29812;
  assign n29814 = n25198 & n26462;
  assign n29815 = n24932 & n26457;
  assign n29816 = ~n29814 & ~n29815;
  assign n29817 = n25149 & n26459;
  assign n29818 = n29816 & ~n29817;
  assign n29819 = n25041 & n27236;
  assign n29820 = n25080 & ~n29819;
  assign n29821 = ~n26465 & n29820;
  assign n29822 = ~n25092 & n29821;
  assign n29823 = n29818 & n29822;
  assign n29824 = n25230 & n27200;
  assign n29825 = n25041 & n27196;
  assign n29826 = ~n29824 & ~n29825;
  assign n29827 = n25290 & n27193;
  assign n29828 = n29826 & ~n29827;
  assign n29829 = n29823 & n29828;
  assign n29830 = n25144 & n29829;
  assign n29831 = n27204 & n29830;
  assign n29832 = n25072 & n29831;
  assign n29833 = n29813 & n29832;
  assign n29834 = n25290 & n27256;
  assign n29835 = n25251 & n25306;
  assign n29836 = ~n29834 & ~n29835;
  assign n29837 = n26482 & n29836;
  assign n29838 = n29131 & n29837;
  assign n29839 = n29833 & n29838;
  assign n29840 = n25133 & n25343;
  assign n29841 = n29839 & n29840;
  assign n29842 = n29797 & n29841;
  assign n29843 = n25322 & n29842;
  assign n29844 = n29782 & n29843;
  assign n29845 = pi3516 & ~n14255;
  assign n29846 = n29844 & ~n29845;
  assign n29847 = n25165 & ~n26718;
  assign n29848 = n25267 & n26538;
  assign n29849 = ~n29847 & ~n29848;
  assign n29850 = n25032 & n25292;
  assign n29851 = n25151 & n25278;
  assign n29852 = ~n29850 & ~n29851;
  assign n29853 = n26536 & n29852;
  assign n29854 = ~n27306 & n29853;
  assign n29855 = n29849 & n29854;
  assign n29856 = n25227 & n29855;
  assign n29857 = n29846 & n29856;
  assign n29858 = n27323 & n29857;
  assign n29859 = n29780 & n29858;
  assign n29860 = n29777 & n29859;
  assign n29861 = n25371 & ~n29860;
  assign n29862 = n25177 & n25246;
  assign n29863 = ~n25183 & ~n29862;
  assign n29864 = n27883 & n29863;
  assign n29865 = n25149 & n25153;
  assign n29866 = n29864 & ~n29865;
  assign n29867 = n25184 & n25230;
  assign n29868 = n25142 & n25237;
  assign n29869 = ~n29867 & ~n29868;
  assign n29870 = n24932 & n25243;
  assign n29871 = n25198 & n25248;
  assign n29872 = ~n29870 & ~n29871;
  assign n29873 = n25165 & n25254;
  assign n29874 = n25202 & n25281;
  assign n29875 = ~n29873 & ~n29874;
  assign n29876 = n24932 & n25309;
  assign n29877 = n25348 & ~n29876;
  assign n29878 = n25097 & n25267;
  assign n29879 = n25100 & n25230;
  assign n29880 = ~n29878 & ~n29879;
  assign n29881 = n25134 & n29880;
  assign n29882 = n25331 & n29881;
  assign n29883 = n29877 & n29882;
  assign n29884 = n25036 & n25267;
  assign n29885 = n25078 & n25103;
  assign n29886 = ~n29884 & ~n29885;
  assign n29887 = n25064 & n25158;
  assign n29888 = n25070 & n25237;
  assign n29889 = ~n29887 & ~n29888;
  assign n29890 = n25093 & n29889;
  assign n29891 = n25076 & n25158;
  assign n29892 = n29890 & ~n29891;
  assign n29893 = n25342 & n29892;
  assign n29894 = n29886 & n29893;
  assign n29895 = n29883 & n29894;
  assign n29896 = n25032 & n25207;
  assign n29897 = n25165 & n25172;
  assign n29898 = ~n29896 & ~n29897;
  assign n29899 = n25103 & n25209;
  assign n29900 = n29898 & ~n29899;
  assign n29901 = n25162 & n25290;
  assign n29902 = n29900 & ~n29901;
  assign n29903 = n25149 & n25169;
  assign n29904 = n25041 & n25160;
  assign n29905 = ~n29903 & ~n29904;
  assign n29906 = n25202 & n25234;
  assign n29907 = n25041 & n25239;
  assign n29908 = ~n29906 & ~n29907;
  assign n29909 = ~n25213 & ~n25215;
  assign n29910 = n25151 & ~n29909;
  assign n29911 = n25226 & ~n29910;
  assign n29912 = n29908 & n29911;
  assign n29913 = n29905 & n29912;
  assign n29914 = n29902 & n29913;
  assign n29915 = n25032 & n25276;
  assign n29916 = n27867 & ~n29915;
  assign n29917 = ~n25285 & n29916;
  assign n29918 = n29914 & n29917;
  assign n29919 = n29895 & n29918;
  assign n29920 = n29875 & n29919;
  assign n29921 = n29872 & n29920;
  assign n29922 = n25198 & n25352;
  assign n29923 = n25290 & n25355;
  assign n29924 = ~n29922 & ~n29923;
  assign n29925 = n25251 & n25314;
  assign n29926 = n29924 & ~n29925;
  assign n29927 = n29921 & n29926;
  assign n29928 = n25246 & n25320;
  assign n29929 = n25251 & n25323;
  assign n29930 = ~n29928 & ~n29929;
  assign n29931 = n26599 & n29930;
  assign n29932 = n29927 & n29931;
  assign n29933 = n29869 & n29932;
  assign n29934 = n29866 & n29933;
  assign n29935 = pi3516 & ~n14259;
  assign n29936 = n29934 & ~n29935;
  assign n29937 = n25443 & ~n29936;
  assign n29938 = ~n29861 & ~n29937;
  assign n29939 = ~n16891 & n25508;
  assign n29940 = ~n14403 & n25512;
  assign n29941 = ~n29939 & ~n29940;
  assign n29942 = n29938 & n29941;
  assign n29943 = ~n14259 & n24922;
  assign n29944 = ~n14255 & n24925;
  assign n29945 = ~n29943 & ~n29944;
  assign n29946 = ~n14259 & n25462;
  assign n29947 = ~n14255 & n25465;
  assign n29948 = ~n29946 & ~n29947;
  assign n29949 = n29945 & n29948;
  assign n29950 = n19807 & n20379;
  assign n29951 = ~n19807 & ~n19852;
  assign n29952 = ~n20380 & n29951;
  assign n29953 = ~n29950 & ~n29952;
  assign n29954 = ~n19851 & ~n20334;
  assign n29955 = ~n19953 & n27804;
  assign n29956 = ~n29954 & ~n29955;
  assign n29957 = ~n29953 & ~n29956;
  assign n29958 = n29953 & n29956;
  assign n29959 = ~n29957 & ~n29958;
  assign n29960 = n24892 & n29959;
  assign n29961 = ~n14286 & ~n24905;
  assign n29962 = ~n14403 & n24916;
  assign n29963 = ~n16891 & n24913;
  assign n29964 = ~n29962 & ~n29963;
  assign n29965 = ~n24909 & n29964;
  assign n29966 = ~n29961 & n29965;
  assign n29967 = ~n29960 & n29966;
  assign n29968 = ~n14219 & n25473;
  assign n29969 = ~n25471 & ~n29968;
  assign n29970 = ~n14223 & ~n25483;
  assign n29971 = ~n14219 & n25474;
  assign n29972 = ~n29970 & ~n29971;
  assign n29973 = n27457 & n29972;
  assign n29974 = ~n25479 & n29973;
  assign n29975 = n29969 & n29974;
  assign n29976 = n27467 & ~n29975;
  assign n29977 = ~n27470 & ~n29976;
  assign n29978 = pi0342 & ~n29977;
  assign n29979 = n29967 & ~n29978;
  assign n29980 = pi0343 & ~n16891;
  assign n29981 = ~pi0343 & ~n14403;
  assign n29982 = ~n29980 & ~n29981;
  assign n29983 = n25458 & ~n29982;
  assign n29984 = ~n27441 & ~n29983;
  assign n29985 = n29979 & n29984;
  assign n29986 = n29949 & n29985;
  assign n29987 = n29942 & n29986;
  assign n29988 = n25544 & ~n29987;
  assign n29989 = ~pi0103 & n25533;
  assign n29990 = ~pi0070 & pi0979;
  assign n29991 = ~pi0071 & ~pi0979;
  assign n29992 = ~n29990 & ~n29991;
  assign n29993 = n25571 & ~n29992;
  assign n29994 = ~n14228 & ~n25582;
  assign n29995 = ~n14232 & n25582;
  assign n29996 = ~n29994 & ~n29995;
  assign n29997 = n25580 & ~n29996;
  assign n29998 = ~pi0103 & n25532;
  assign n29999 = ~n29997 & ~n29998;
  assign n30000 = n14237 & ~n25594;
  assign n30001 = n14241 & n25594;
  assign n30002 = ~n30000 & ~n30001;
  assign n30003 = n25591 & n30002;
  assign n30004 = n29999 & ~n30003;
  assign n30005 = ~n29993 & n30004;
  assign n30006 = n25606 & n30005;
  assign n30007 = n14403 & ~n25606;
  assign n30008 = ~n30006 & ~n30007;
  assign n30009 = n25564 & n30008;
  assign n30010 = ~n25606 & ~n30005;
  assign n30011 = ~n16891 & n25606;
  assign n30012 = ~n30010 & ~n30011;
  assign n30013 = ~n25564 & ~n30012;
  assign n30014 = ~n30009 & ~n30013;
  assign n30015 = ~n25533 & ~n30014;
  assign n30016 = ~n29989 & ~n30015;
  assign n30017 = ~n25544 & ~n30016;
  assign po0373 = n29988 | n30017;
  assign n30019 = ~n16529 & n24913;
  assign n30020 = ~n11181 & n24916;
  assign n30021 = ~n30019 & ~n30020;
  assign n30022 = ~n20258 & ~n20334;
  assign n30023 = ~n20216 & n20232;
  assign n30024 = n20216 & ~n20232;
  assign n30025 = ~n30023 & ~n30024;
  assign n30026 = ~n20380 & ~n30025;
  assign n30027 = n20233 & n20379;
  assign n30028 = ~n30026 & ~n30027;
  assign n30029 = ~n30022 & n30028;
  assign n30030 = n30022 & ~n30028;
  assign n30031 = ~n30029 & ~n30030;
  assign n30032 = n24892 & n30031;
  assign n30033 = ~n11011 & ~n24905;
  assign n30034 = ~n30032 & ~n30033;
  assign n30035 = ~n10966 & n25474;
  assign n30036 = ~n25479 & ~n30035;
  assign n30037 = ~n25471 & n30036;
  assign n30038 = ~n10970 & ~n25483;
  assign n30039 = n30037 & ~n30038;
  assign n30040 = ~n10975 & ~n25487;
  assign n30041 = ~n10966 & n25473;
  assign n30042 = ~n30040 & ~n30041;
  assign n30043 = n30039 & n30042;
  assign n30044 = ~n25491 & n30043;
  assign n30045 = ~pi0343 & ~n30044;
  assign n30046 = pi0343 & ~n11181;
  assign n30047 = ~n30045 & ~n30046;
  assign n30048 = n25498 & ~n30047;
  assign n30049 = n30034 & ~n30048;
  assign n30050 = ~n24909 & n30049;
  assign n30051 = n30021 & n30050;
  assign n30052 = ~n11038 & n24922;
  assign n30053 = ~n11020 & n24925;
  assign n30054 = ~n30052 & ~n30053;
  assign n30055 = ~n11038 & n25462;
  assign n30056 = ~n11020 & n25465;
  assign n30057 = ~n30055 & ~n30056;
  assign n30058 = n25097 & n25103;
  assign n30059 = n25116 & ~n30058;
  assign n30060 = n25237 & n25352;
  assign n30061 = n24932 & n25355;
  assign n30062 = ~n30060 & ~n30061;
  assign n30063 = n25198 & n25358;
  assign n30064 = n25267 & n25360;
  assign n30065 = ~n30063 & ~n30064;
  assign n30066 = n25100 & n25165;
  assign n30067 = n25237 & n25248;
  assign n30068 = n25032 & n25243;
  assign n30069 = ~n30067 & ~n30068;
  assign n30070 = n25230 & n25292;
  assign n30071 = n30069 & ~n30070;
  assign n30072 = n25041 & n25270;
  assign n30073 = n25261 & n25290;
  assign n30074 = ~n30072 & ~n30073;
  assign n30075 = n25230 & n25264;
  assign n30076 = n25246 & n25254;
  assign n30077 = ~n30075 & ~n30076;
  assign n30078 = ~n25258 & n30077;
  assign n30079 = n30074 & n30078;
  assign n30080 = n30071 & n30079;
  assign n30081 = n25158 & n25281;
  assign n30082 = n30080 & ~n30081;
  assign n30083 = n25172 & n25246;
  assign n30084 = n25169 & n25251;
  assign n30085 = ~n30083 & ~n30084;
  assign n30086 = n25149 & n25160;
  assign n30087 = n24932 & n25162;
  assign n30088 = ~n30086 & ~n30087;
  assign n30089 = n25195 & n25202;
  assign n30090 = n25041 & n25204;
  assign n30091 = ~n30089 & ~n30090;
  assign n30092 = n30088 & n30091;
  assign n30093 = n25211 & n30092;
  assign n30094 = n30085 & n30093;
  assign n30095 = n25231 & n25290;
  assign n30096 = n25158 & n25234;
  assign n30097 = n25149 & n25239;
  assign n30098 = ~n30096 & ~n30097;
  assign n30099 = ~n30095 & n30098;
  assign n30100 = ~n25214 & n30099;
  assign n30101 = ~n25221 & n30100;
  assign n30102 = ~n25216 & n30101;
  assign n30103 = ~n25225 & n30102;
  assign n30104 = n30094 & n30103;
  assign n30105 = n26536 & n30104;
  assign n30106 = ~n25279 & n30105;
  assign n30107 = n30082 & n30106;
  assign n30108 = n25326 & n30107;
  assign n30109 = ~n30066 & n30108;
  assign n30110 = n30065 & n30109;
  assign n30111 = n30062 & n30110;
  assign n30112 = n25202 & n25306;
  assign n30113 = n25348 & ~n30112;
  assign n30114 = n25331 & n30113;
  assign n30115 = n25032 & n25309;
  assign n30116 = n30114 & ~n30115;
  assign n30117 = n25064 & n25151;
  assign n30118 = n25036 & n25103;
  assign n30119 = ~n30117 & ~n30118;
  assign n30120 = n25028 & n25267;
  assign n30121 = n25076 & n25151;
  assign n30122 = ~n30120 & ~n30121;
  assign n30123 = n30119 & n30122;
  assign n30124 = n25342 & n30123;
  assign n30125 = n30116 & n30124;
  assign n30126 = ~n25079 & n25088;
  assign n30127 = n26979 & n30126;
  assign n30128 = n30125 & n30127;
  assign n30129 = n25153 & n25251;
  assign n30130 = n25165 & n25184;
  assign n30131 = n25146 & n25198;
  assign n30132 = ~n30130 & ~n30131;
  assign n30133 = ~n30129 & n30132;
  assign n30134 = ~n25178 & n30133;
  assign n30135 = n30128 & n30134;
  assign n30136 = n28843 & n30135;
  assign n30137 = n25144 & n30136;
  assign n30138 = n30111 & n30137;
  assign n30139 = n25132 & n30138;
  assign n30140 = n25124 & n30139;
  assign n30141 = n30059 & n30140;
  assign n30142 = pi3516 & ~n11020;
  assign n30143 = n30141 & ~n30142;
  assign n30144 = n25371 & ~n30143;
  assign n30145 = n25103 & n25312;
  assign n30146 = n25202 & n25314;
  assign n30147 = ~n30145 & ~n30146;
  assign n30148 = n25165 & n25179;
  assign n30149 = n25182 & n25246;
  assign n30150 = ~n30148 & ~n30149;
  assign n30151 = n25041 & n25142;
  assign n30152 = n30150 & ~n30151;
  assign n30153 = n25084 & n25165;
  assign n30154 = n25086 & n25149;
  assign n30155 = ~n30153 & ~n30154;
  assign n30156 = n25251 & n25329;
  assign n30157 = n25151 & n25345;
  assign n30158 = ~n30156 & ~n30157;
  assign n30159 = n25032 & n25327;
  assign n30160 = n25336 & n29552;
  assign n30161 = ~n30159 & n30160;
  assign n30162 = n30158 & n30161;
  assign n30163 = n24932 & n25091;
  assign n30164 = n25177 & n25267;
  assign n30165 = ~n30163 & ~n30164;
  assign n30166 = n25041 & n25070;
  assign n30167 = n25078 & n25290;
  assign n30168 = ~n25139 & ~n30167;
  assign n30169 = ~n30166 & n30168;
  assign n30170 = n30165 & n30169;
  assign n30171 = n30162 & n30170;
  assign n30172 = n25207 & n25230;
  assign n30173 = n25198 & n25213;
  assign n30174 = ~n30172 & ~n30173;
  assign n30175 = n25151 & n25284;
  assign n30176 = n25224 & n25237;
  assign n30177 = ~n30175 & ~n30176;
  assign n30178 = n25127 & n25246;
  assign n30179 = n25122 & n25251;
  assign n30180 = ~n30178 & ~n30179;
  assign n30181 = n25110 & n25149;
  assign n30182 = n30180 & ~n30181;
  assign n30183 = n25220 & n25237;
  assign n30184 = n25198 & n25215;
  assign n30185 = ~n30183 & ~n30184;
  assign n30186 = n25230 & n25276;
  assign n30187 = n25209 & n25290;
  assign n30188 = ~n25279 & ~n30187;
  assign n30189 = ~n30186 & n30188;
  assign n30190 = n30185 & n30189;
  assign n30191 = n25158 & n25257;
  assign n30192 = n30190 & ~n30191;
  assign n30193 = n30182 & n30192;
  assign n30194 = n30177 & n30193;
  assign n30195 = n30174 & n30194;
  assign n30196 = n24932 & n25114;
  assign n30197 = n25130 & n25158;
  assign n30198 = ~n30196 & ~n30197;
  assign n30199 = ~n25119 & n30198;
  assign n30200 = n30195 & n30199;
  assign n30201 = n30171 & n30200;
  assign n30202 = n30155 & n30201;
  assign n30203 = n30152 & n30202;
  assign n30204 = pi3516 & ~n11038;
  assign n30205 = n30203 & ~n30204;
  assign n30206 = n25267 & n25320;
  assign n30207 = n25032 & n25317;
  assign n30208 = ~n30206 & ~n30207;
  assign n30209 = n25202 & n25323;
  assign n30210 = n30208 & ~n30209;
  assign n30211 = n30205 & n30210;
  assign n30212 = n30147 & n30211;
  assign n30213 = n25443 & ~n30212;
  assign n30214 = ~n30144 & ~n30213;
  assign n30215 = ~n16529 & n25508;
  assign n30216 = ~n11181 & n25512;
  assign n30217 = ~n30215 & ~n30216;
  assign n30218 = n30214 & n30217;
  assign n30219 = n30057 & n30218;
  assign n30220 = n30054 & n30219;
  assign n30221 = n30051 & n30220;
  assign n30222 = ~n16529 & n25449;
  assign n30223 = ~n25452 & ~n30222;
  assign n30224 = ~pi0342 & ~n30223;
  assign n30225 = pi0343 & ~n16529;
  assign n30226 = ~pi0343 & ~n11181;
  assign n30227 = ~n30225 & ~n30226;
  assign n30228 = n25458 & ~n30227;
  assign n30229 = ~n30224 & ~n30228;
  assign n30230 = n30221 & n30229;
  assign n30231 = n25544 & ~n30230;
  assign n30232 = ~pi0104 & n25533;
  assign n30233 = ~pi0091 & pi0979;
  assign n30234 = ~pi0094 & ~pi0979;
  assign n30235 = ~n30233 & ~n30234;
  assign n30236 = n25571 & ~n30235;
  assign n30237 = ~n10979 & ~n25582;
  assign n30238 = ~n10983 & n25582;
  assign n30239 = ~n30237 & ~n30238;
  assign n30240 = n25580 & ~n30239;
  assign n30241 = ~pi0104 & n25532;
  assign n30242 = ~n30240 & ~n30241;
  assign n30243 = n10957 & ~n25594;
  assign n30244 = n10961 & n25594;
  assign n30245 = ~n30243 & ~n30244;
  assign n30246 = n25591 & n30245;
  assign n30247 = n30242 & ~n30246;
  assign n30248 = ~n30236 & n30247;
  assign n30249 = n25606 & ~n30248;
  assign n30250 = ~n11181 & ~n25606;
  assign n30251 = ~n30249 & ~n30250;
  assign n30252 = n25564 & ~n30251;
  assign n30253 = ~n16529 & n25606;
  assign n30254 = ~n25606 & ~n30248;
  assign n30255 = ~n30253 & ~n30254;
  assign n30256 = ~n25564 & ~n30255;
  assign n30257 = ~n30252 & ~n30256;
  assign n30258 = ~n25533 & ~n30257;
  assign n30259 = ~n30232 & ~n30258;
  assign n30260 = ~n25544 & ~n30259;
  assign po0374 = n30231 | n30260;
  assign n30262 = n25620 & ~n28753;
  assign n30263 = pi0105 & ~n25625;
  assign n30264 = n25558 & n28762;
  assign n30265 = ~pi3245 & ~n12726;
  assign n30266 = pi3245 & ~n16855;
  assign n30267 = ~n30265 & ~n30266;
  assign n30268 = ~n25558 & n30267;
  assign n30269 = ~n30264 & ~n30268;
  assign n30270 = n25625 & n30269;
  assign n30271 = ~n30263 & ~n30270;
  assign n30272 = ~n25620 & ~n30271;
  assign po0375 = n30262 | n30272;
  assign n30274 = n25620 & ~n28501;
  assign n30275 = pi0106 & ~n25625;
  assign n30276 = n25558 & ~n28510;
  assign n30277 = ~n24256 & ~n25558;
  assign n30278 = ~n30276 & ~n30277;
  assign n30279 = n25625 & ~n30278;
  assign n30280 = ~n30275 & ~n30279;
  assign n30281 = ~n25620 & ~n30280;
  assign po0376 = n30274 | n30281;
  assign n30283 = n25620 & ~n28017;
  assign n30284 = pi0107 & ~n25625;
  assign n30285 = n25558 & n28026;
  assign n30286 = ~pi3245 & ~n13701;
  assign n30287 = pi3245 & ~n16819;
  assign n30288 = ~n30286 & ~n30287;
  assign n30289 = ~n25558 & n30288;
  assign n30290 = ~n30285 & ~n30289;
  assign n30291 = n25625 & n30290;
  assign n30292 = ~n30284 & ~n30291;
  assign n30293 = ~n25620 & ~n30292;
  assign po0377 = n30283 | n30293;
  assign n30295 = n25620 & ~n28262;
  assign n30296 = pi0108 & ~n25625;
  assign n30297 = n25558 & ~n28271;
  assign n30298 = ~n24744 & ~n25558;
  assign n30299 = ~n30297 & ~n30298;
  assign n30300 = n25625 & ~n30299;
  assign n30301 = ~n30296 & ~n30300;
  assign n30302 = ~n25620 & ~n30301;
  assign po0378 = n30295 | n30302;
  assign n30304 = n25620 & ~n28997;
  assign n30305 = pi0109 & ~n25625;
  assign n30306 = n25558 & ~n29006;
  assign n30307 = ~pi3245 & ~n17199;
  assign n30308 = pi3245 & ~n17105;
  assign n30309 = ~n30307 & ~n30308;
  assign n30310 = ~n25558 & ~n30309;
  assign n30311 = ~n30306 & ~n30310;
  assign n30312 = n25625 & ~n30311;
  assign n30313 = ~n30305 & ~n30312;
  assign n30314 = ~n25620 & ~n30313;
  assign po0379 = n30304 | n30314;
  assign n30316 = n25620 & ~n29244;
  assign n30317 = pi0110 & ~n25625;
  assign n30318 = n25558 & n29253;
  assign n30319 = ~pi3245 & ~n9825;
  assign n30320 = pi3245 & ~n16999;
  assign n30321 = ~n30319 & ~n30320;
  assign n30322 = ~n25558 & n30321;
  assign n30323 = ~n30318 & ~n30322;
  assign n30324 = n25625 & n30323;
  assign n30325 = ~n30317 & ~n30324;
  assign n30326 = ~n25620 & ~n30325;
  assign po0380 = n30316 | n30326;
  assign n30328 = n25620 & ~n29486;
  assign n30329 = pi0111 & ~n25625;
  assign n30330 = n25558 & n29495;
  assign n30331 = ~pi3245 & ~n10608;
  assign n30332 = pi3245 & ~n16963;
  assign n30333 = ~n30331 & ~n30332;
  assign n30334 = ~n25558 & n30333;
  assign n30335 = ~n30330 & ~n30334;
  assign n30336 = n25625 & n30335;
  assign n30337 = ~n30329 & ~n30336;
  assign n30338 = ~n25620 & ~n30337;
  assign po0381 = n30328 | n30338;
  assign n30340 = n25620 & ~n29736;
  assign n30341 = pi0112 & ~n25625;
  assign n30342 = n25558 & n29745;
  assign n30343 = ~n25558 & n27570;
  assign n30344 = ~n30342 & ~n30343;
  assign n30345 = n25625 & n30344;
  assign n30346 = ~n30341 & ~n30345;
  assign n30347 = ~n25620 & ~n30346;
  assign po0382 = n30340 | n30347;
  assign n30349 = n25620 & ~n29987;
  assign n30350 = pi0113 & ~n25625;
  assign n30351 = n25558 & n29996;
  assign n30352 = ~n25558 & n25999;
  assign n30353 = ~n30351 & ~n30352;
  assign n30354 = n25625 & n30353;
  assign n30355 = ~n30350 & ~n30354;
  assign n30356 = ~n25620 & ~n30355;
  assign po0383 = n30349 | n30356;
  assign n30358 = n25620 & ~n30230;
  assign n30359 = pi0114 & ~n25625;
  assign n30360 = n25558 & ~n30239;
  assign n30361 = ~n24488 & ~n25558;
  assign n30362 = ~n30360 & ~n30361;
  assign n30363 = n25625 & ~n30362;
  assign n30364 = ~n30359 & ~n30363;
  assign n30365 = ~n25620 & ~n30364;
  assign po0384 = n30358 | n30365;
  assign n30367 = pi0868 & n25648;
  assign n30368 = ~n21552 & ~n25641;
  assign n30369 = n25643 & ~n30368;
  assign n30370 = ~n25643 & n30368;
  assign n30371 = ~n30369 & ~n30370;
  assign n30372 = ~pi0868 & n30371;
  assign n30373 = ~n30367 & ~n30372;
  assign n30374 = n25637 & ~n30373;
  assign n30375 = pi0115 & n20518;
  assign n30376 = pi0115 & ~n24259;
  assign n30377 = n24259 & ~n30309;
  assign n30378 = ~n30376 & ~n30377;
  assign n30379 = n26002 & ~n30378;
  assign n30380 = ~n30375 & ~n30379;
  assign n30381 = ~n26006 & n30380;
  assign n30382 = ~n25637 & ~n30381;
  assign po0385 = n30374 | n30382;
  assign n30384 = n24099 & ~n27555;
  assign n30385 = ~n27554 & ~n30384;
  assign n30386 = n21536 & n21542;
  assign n30387 = ~n21536 & ~n21542;
  assign n30388 = ~n30386 & ~n30387;
  assign n30389 = ~n30385 & n30388;
  assign n30390 = n30385 & ~n30388;
  assign n30391 = ~n30389 & ~n30390;
  assign n30392 = ~pi0868 & n30391;
  assign n30393 = pi0868 & n30371;
  assign n30394 = ~n30392 & ~n30393;
  assign n30395 = n25637 & ~n30394;
  assign n30396 = pi0116 & n20518;
  assign n30397 = pi0116 & ~n24259;
  assign n30398 = n24259 & ~n30321;
  assign n30399 = ~n30397 & ~n30398;
  assign n30400 = n26002 & ~n30399;
  assign n30401 = ~n30396 & ~n30400;
  assign n30402 = ~n26006 & n30401;
  assign n30403 = ~n25637 & ~n30402;
  assign po0386 = n30395 | n30403;
  assign n30405 = pi0868 & n30391;
  assign n30406 = ~pi0868 & n27562;
  assign n30407 = ~n30405 & ~n30406;
  assign n30408 = n25637 & ~n30407;
  assign n30409 = pi0117 & n20518;
  assign n30410 = pi0117 & ~n24259;
  assign n30411 = n24259 & ~n30333;
  assign n30412 = ~n30410 & ~n30411;
  assign n30413 = n26002 & ~n30412;
  assign n30414 = ~n30409 & ~n30413;
  assign n30415 = ~n26006 & n30414;
  assign n30416 = ~n25637 & ~n30415;
  assign po0387 = n30408 | n30416;
  assign n30418 = n25663 & ~n30394;
  assign n30419 = pi0118 & n24300;
  assign n30420 = pi0118 & ~n24314;
  assign n30421 = n24314 & ~n30321;
  assign n30422 = ~n30420 & ~n30421;
  assign n30423 = n26041 & ~n30422;
  assign n30424 = ~n30419 & ~n30423;
  assign n30425 = ~n26045 & n30424;
  assign n30426 = ~n25663 & ~n30425;
  assign po0388 = n30418 | n30426;
  assign n30428 = n25663 & ~n30373;
  assign n30429 = pi0119 & n24300;
  assign n30430 = pi0119 & ~n24314;
  assign n30431 = n24314 & ~n30309;
  assign n30432 = ~n30430 & ~n30431;
  assign n30433 = n26041 & ~n30432;
  assign n30434 = ~n30429 & ~n30433;
  assign n30435 = ~n26045 & n30434;
  assign n30436 = ~n25663 & ~n30435;
  assign po0389 = n30428 | n30436;
  assign n30438 = n25663 & ~n30407;
  assign n30439 = pi0120 & n24300;
  assign n30440 = pi0120 & ~n24314;
  assign n30441 = n24314 & ~n30333;
  assign n30442 = ~n30440 & ~n30441;
  assign n30443 = n26041 & ~n30442;
  assign n30444 = ~n30439 & ~n30443;
  assign n30445 = ~n26045 & n30444;
  assign n30446 = ~n25663 & ~n30445;
  assign po0390 = n30438 | n30446;
  assign n30448 = n26051 & ~n30394;
  assign n30449 = ~pi0121 & ~n26051;
  assign po0391 = n30448 | n30449;
  assign n30451 = n26051 & ~n30407;
  assign n30452 = ~pi0122 & ~n26051;
  assign po0392 = n30451 | n30452;
  assign n30454 = n26051 & ~n30373;
  assign n30455 = ~pi0123 & ~n26051;
  assign po0393 = n30454 | n30455;
  assign n30457 = n26056 & ~n30373;
  assign n30458 = ~pi0124 & ~n26056;
  assign po0394 = n30457 | n30458;
  assign n30460 = n26056 & ~n30394;
  assign n30461 = ~pi0125 & ~n26056;
  assign po0395 = n30460 | n30461;
  assign n30463 = n26056 & ~n30407;
  assign n30464 = ~pi0126 & ~n26056;
  assign po0396 = n30463 | n30464;
  assign n30466 = ~pi2555 & ~n26062;
  assign n30467 = ~n15115 & n30466;
  assign n30468 = n26293 & n26339;
  assign n30469 = ~n26344 & n26347;
  assign n30470 = n26281 & n30469;
  assign n30471 = n26274 & n26349;
  assign n30472 = ~n26311 & n26352;
  assign n30473 = ~n26317 & n26355;
  assign n30474 = n26357 & ~n26364;
  assign n30475 = ~n26357 & ~n26395;
  assign n30476 = ~n30474 & ~n30475;
  assign n30477 = ~n26355 & ~n30476;
  assign n30478 = ~n30473 & ~n30477;
  assign n30479 = ~n26352 & ~n30478;
  assign n30480 = ~n30472 & ~n30479;
  assign n30481 = ~n26349 & ~n30480;
  assign n30482 = ~n30471 & ~n30481;
  assign n30483 = ~n26344 & ~n26347;
  assign n30484 = ~n30482 & n30483;
  assign n30485 = ~n30470 & ~n30484;
  assign n30486 = ~n26334 & ~n30485;
  assign n30487 = n26297 & n26345;
  assign n30488 = ~n30486 & ~n30487;
  assign n30489 = ~n26338 & ~n30488;
  assign n30490 = ~n30468 & ~n30489;
  assign n30491 = pi2555 & ~n30490;
  assign n30492 = pi2555 & n26338;
  assign n30493 = ~n26364 & n30492;
  assign n30494 = ~n30491 & ~n30493;
  assign n30495 = ~n26062 & ~n30494;
  assign n30496 = pi0127 & n26062;
  assign n30497 = ~n30495 & ~n30496;
  assign po0397 = n30467 | ~n30497;
  assign n30499 = ~n11181 & n30466;
  assign n30500 = ~n26311 & n30469;
  assign n30501 = ~n26317 & n26349;
  assign n30502 = n26352 & ~n26364;
  assign n30503 = n26355 & ~n26395;
  assign n30504 = n26357 & ~n26409;
  assign n30505 = ~pi1017 & n26405;
  assign n30506 = ~pi0128 & ~pi1017;
  assign n30507 = ~pi0128 & ~n30506;
  assign n30508 = pi1017 & ~n30507;
  assign n30509 = ~n30505 & ~n30508;
  assign n30510 = n26237 & ~n30509;
  assign n30511 = ~n26357 & ~n30510;
  assign n30512 = ~n30504 & ~n30511;
  assign n30513 = ~n26355 & ~n30512;
  assign n30514 = ~n30503 & ~n30513;
  assign n30515 = ~n26352 & ~n30514;
  assign n30516 = ~n30502 & ~n30515;
  assign n30517 = ~n26349 & ~n30516;
  assign n30518 = ~n30501 & ~n30517;
  assign n30519 = n30483 & ~n30518;
  assign n30520 = ~n30500 & ~n30519;
  assign n30521 = ~n26334 & ~n30520;
  assign n30522 = n26274 & n26345;
  assign n30523 = ~n30521 & ~n30522;
  assign n30524 = ~n26338 & ~n30523;
  assign n30525 = n26281 & n26339;
  assign n30526 = ~n30524 & ~n30525;
  assign n30527 = pi2555 & ~n30526;
  assign n30528 = ~n26409 & n30492;
  assign n30529 = ~n30527 & ~n30528;
  assign n30530 = ~n26062 & ~n30529;
  assign n30531 = pi0128 & n26062;
  assign n30532 = ~n30530 & ~n30531;
  assign po0398 = n30499 | ~n30532;
  assign n30534 = pi0979 & n9365;
  assign n30535 = pi0599 & n19569;
  assign n30536 = n30534 & ~n30535;
  assign n30537 = ~pi3426 & ~n19569;
  assign n30538 = ~n11181 & n25547;
  assign n30539 = ~n16529 & ~n25547;
  assign n30540 = ~n30538 & ~n30539;
  assign n30541 = ~n30537 & ~n30540;
  assign n30542 = n19630 & n20387;
  assign n30543 = ~n19630 & ~n20387;
  assign n30544 = ~n30542 & ~n30543;
  assign n30545 = pi2758 & ~n30544;
  assign n30546 = ~n19599 & ~n19630;
  assign n30547 = n19599 & n19630;
  assign n30548 = ~n30546 & ~n30547;
  assign n30549 = ~pi2758 & ~n30548;
  assign n30550 = ~n30545 & ~n30549;
  assign n30551 = ~pi2758 & ~n30550;
  assign n30552 = pi2758 & n30550;
  assign n30553 = ~n30551 & ~n30552;
  assign n30554 = n30537 & ~n30553;
  assign n30555 = ~n30541 & ~n30554;
  assign n30556 = n30536 & ~n30555;
  assign n30557 = pi0129 & ~n30536;
  assign po0399 = n30556 | n30557;
  assign n30559 = pi0130 & n20518;
  assign n30560 = pi0130 & ~n24259;
  assign n30561 = n24259 & ~n24769;
  assign n30562 = ~n30560 & ~n30561;
  assign n30563 = n26002 & ~n30562;
  assign n30564 = ~n30559 & ~n30563;
  assign n30565 = ~n26006 & n30564;
  assign n30566 = ~n25637 & ~n30565;
  assign n30567 = n22761 & ~n26010;
  assign n30568 = n23296 & ~n30567;
  assign n30569 = ~n22258 & ~n22419;
  assign n30570 = ~n30568 & ~n30569;
  assign n30571 = n22258 & n22419;
  assign n30572 = ~n30570 & ~n30571;
  assign n30573 = n22255 & n22261;
  assign n30574 = ~n22255 & ~n22261;
  assign n30575 = ~n30573 & ~n30574;
  assign n30576 = n30572 & n30575;
  assign n30577 = ~n30572 & ~n30575;
  assign n30578 = ~n30576 & ~n30577;
  assign n30579 = pi0868 & n30578;
  assign n30580 = n22258 & ~n22419;
  assign n30581 = ~n22258 & n22419;
  assign n30582 = ~n30580 & ~n30581;
  assign n30583 = n30568 & ~n30582;
  assign n30584 = ~n30568 & n30582;
  assign n30585 = ~n30583 & ~n30584;
  assign n30586 = ~pi0868 & ~n30585;
  assign n30587 = ~n30579 & ~n30586;
  assign n30588 = n25637 & ~n30587;
  assign po0400 = n30566 | n30588;
  assign n30590 = pi0131 & n24300;
  assign n30591 = pi0131 & ~n24314;
  assign n30592 = n24314 & ~n24769;
  assign n30593 = ~n30591 & ~n30592;
  assign n30594 = n26041 & ~n30593;
  assign n30595 = ~n30590 & ~n30594;
  assign n30596 = ~n26045 & n30595;
  assign n30597 = ~n25663 & ~n30596;
  assign n30598 = n25663 & ~n30587;
  assign po0401 = n30597 | n30598;
  assign n30600 = ~pi0132 & ~n26051;
  assign n30601 = n26051 & ~n30587;
  assign po0402 = n30600 | n30601;
  assign n30603 = ~pi0133 & ~n26056;
  assign n30604 = n26056 & ~n30587;
  assign po0403 = n30603 | n30604;
  assign n30606 = ~pi0134 & n19557;
  assign n30607 = ~n19557 & n20408;
  assign n30608 = ~n30606 & ~n30607;
  assign n30609 = pi1909 & pi3586;
  assign po3882 = pi0936 & n30609;
  assign po3897 = ~po0493 | po3882;
  assign po0404 = n30608 & ~po3897;
  assign n30613 = pi0135 & n20518;
  assign n30614 = pi0135 & ~n24259;
  assign n30615 = n24259 & ~n30267;
  assign n30616 = ~n30614 & ~n30615;
  assign n30617 = n26002 & ~n30616;
  assign n30618 = ~n30613 & ~n30617;
  assign n30619 = ~n26006 & n30618;
  assign n30620 = ~n25637 & ~n30619;
  assign n30621 = pi0868 & ~n26032;
  assign n30622 = ~n21960 & ~n22105;
  assign n30623 = ~n22108 & ~n26012;
  assign n30624 = ~n22103 & ~n30623;
  assign n30625 = ~n30622 & ~n30624;
  assign n30626 = n30622 & n30624;
  assign n30627 = ~n30625 & ~n30626;
  assign n30628 = ~pi0868 & ~n30627;
  assign n30629 = ~n30621 & ~n30628;
  assign n30630 = n25637 & ~n30629;
  assign po0405 = n30620 | n30630;
  assign n30632 = ~pi0868 & n30578;
  assign n30633 = ~n22103 & ~n22108;
  assign n30634 = n26012 & ~n30633;
  assign n30635 = ~n26012 & n30633;
  assign n30636 = ~n30634 & ~n30635;
  assign n30637 = pi0868 & n30636;
  assign n30638 = ~n30632 & ~n30637;
  assign n30639 = n25637 & ~n30638;
  assign n30640 = pi0136 & n20518;
  assign n30641 = pi0136 & ~n24259;
  assign n30642 = n24259 & ~n24744;
  assign n30643 = ~n30641 & ~n30642;
  assign n30644 = n26002 & ~n30643;
  assign n30645 = ~n30640 & ~n30644;
  assign n30646 = ~n26006 & n30645;
  assign n30647 = ~n25637 & ~n30646;
  assign po0406 = n30639 | n30647;
  assign n30649 = pi0137 & n24300;
  assign n30650 = pi0137 & ~n24314;
  assign n30651 = n24314 & ~n30267;
  assign n30652 = ~n30650 & ~n30651;
  assign n30653 = n26041 & ~n30652;
  assign n30654 = ~n30649 & ~n30653;
  assign n30655 = ~n26045 & n30654;
  assign n30656 = ~n25663 & ~n30655;
  assign n30657 = n25663 & ~n30629;
  assign po0407 = n30656 | n30657;
  assign n30659 = n25663 & ~n30638;
  assign n30660 = pi0138 & n24300;
  assign n30661 = pi0138 & ~n24314;
  assign n30662 = n24314 & ~n24744;
  assign n30663 = ~n30661 & ~n30662;
  assign n30664 = n26041 & ~n30663;
  assign n30665 = ~n30660 & ~n30664;
  assign n30666 = ~n26045 & n30665;
  assign n30667 = ~n25663 & ~n30666;
  assign po0408 = n30659 | n30667;
  assign n30669 = ~pi0139 & ~n26051;
  assign n30670 = n26051 & ~n30629;
  assign po0409 = n30669 | n30670;
  assign n30672 = n26051 & ~n30638;
  assign n30673 = ~pi0140 & ~n26051;
  assign po0410 = n30672 | n30673;
  assign n30675 = ~pi0141 & ~n26056;
  assign n30676 = n26056 & ~n30629;
  assign po0411 = n30675 | n30676;
  assign n30678 = n26056 & ~n30638;
  assign n30679 = ~pi0142 & ~n26056;
  assign po0412 = n30678 | n30679;
  assign n30681 = ~n9352 & n30537;
  assign n30682 = ~n19551 & ~n30681;
  assign n30683 = ~n19543 & n30682;
  assign n30684 = pi0143 & ~po3897;
  assign n30685 = n30683 & n30684;
  assign n30686 = n30537 & ~n30550;
  assign n30687 = ~pi0835 & ~n13988;
  assign n30688 = ~n30686 & ~n30687;
  assign n30689 = ~pi1612 & n20345;
  assign n30690 = ~pi1533 & n20347;
  assign n30691 = ~n30689 & ~n30690;
  assign n30692 = ~pi1613 & n20350;
  assign n30693 = ~pi1568 & n20353;
  assign n30694 = ~pi1551 & n20356;
  assign n30695 = ~n30693 & ~n30694;
  assign n30696 = ~pi1497 & n20360;
  assign n30697 = ~pi1479 & n20363;
  assign n30698 = ~n30696 & ~n30697;
  assign n30699 = n30695 & n30698;
  assign n30700 = ~n30692 & n30699;
  assign n30701 = n30691 & n30700;
  assign n30702 = n19550 & ~n30701;
  assign n30703 = n30688 & ~n30702;
  assign n30704 = ~n30683 & ~n30703;
  assign n30705 = ~po3897 & n30704;
  assign po0413 = n30685 | n30705;
  assign n30707 = ~pi0979 & ~pi3426;
  assign n30708 = ~n30535 & n30707;
  assign n30709 = ~n9352 & n30708;
  assign n30710 = ~n30555 & n30709;
  assign n30711 = pi0144 & ~n30709;
  assign po0414 = n30710 | n30711;
  assign n30713 = pi0868 & ~n30627;
  assign n30714 = ~pi0868 & n30636;
  assign n30715 = ~n30713 & ~n30714;
  assign n30716 = n25637 & ~n30715;
  assign n30717 = pi0145 & n20518;
  assign n30718 = pi0145 & ~n24259;
  assign n30719 = n24259 & ~n30288;
  assign n30720 = ~n30718 & ~n30719;
  assign n30721 = n26002 & ~n30720;
  assign n30722 = ~n30717 & ~n30721;
  assign n30723 = ~n26006 & n30722;
  assign n30724 = ~n25637 & ~n30723;
  assign po0415 = n30716 | n30724;
  assign n30726 = n25663 & ~n30715;
  assign n30727 = pi0146 & n24300;
  assign n30728 = pi0146 & ~n24314;
  assign n30729 = n24314 & ~n30288;
  assign n30730 = ~n30728 & ~n30729;
  assign n30731 = n26041 & ~n30730;
  assign n30732 = ~n30727 & ~n30731;
  assign n30733 = ~n26045 & n30732;
  assign n30734 = ~n25663 & ~n30733;
  assign po0416 = n30726 | n30734;
  assign n30736 = n26051 & ~n30715;
  assign n30737 = ~pi0147 & ~n26051;
  assign po0417 = n30736 | n30737;
  assign n30739 = n26056 & ~n30715;
  assign n30740 = ~pi0148 & ~n26056;
  assign po0418 = n30739 | n30740;
  assign n30742 = ~pi0835 & ~n11181;
  assign n30743 = n24900 & ~n28307;
  assign n30744 = n19554 & ~n30031;
  assign n30745 = n28725 & ~n29708;
  assign n30746 = ~n27813 & n30745;
  assign n30747 = ~n29959 & n30746;
  assign n30748 = n26654 & ~n28234;
  assign n30749 = n27134 & n30748;
  assign n30750 = ~n26896 & n30749;
  assign n30751 = n30747 & n30750;
  assign n30752 = ~n20387 & ~n29216;
  assign n30753 = n29458 & n30752;
  assign n30754 = n28969 & n30753;
  assign n30755 = n30751 & n30754;
  assign n30756 = n25761 & n30755;
  assign n30757 = n30744 & n30756;
  assign n30758 = n30743 & n30757;
  assign n30759 = ~n30742 & ~n30758;
  assign n30760 = ~n19557 & ~n30759;
  assign n30761 = ~pi1511 & n20360;
  assign n30762 = ~pi1493 & n20363;
  assign n30763 = ~n30761 & ~n30762;
  assign n30764 = ~pi1580 & n20353;
  assign n30765 = ~pi1564 & n20356;
  assign n30766 = ~n30764 & ~n30765;
  assign n30767 = ~pi1420 & n20345;
  assign n30768 = ~pi1547 & n20347;
  assign n30769 = ~n30767 & ~n30768;
  assign n30770 = ~pi1414 & n20350;
  assign n30771 = n30769 & ~n30770;
  assign n30772 = n30766 & n30771;
  assign n30773 = n30763 & n30772;
  assign n30774 = n19550 & ~n30773;
  assign n30775 = ~n19557 & n30774;
  assign n30776 = ~n30760 & ~n30775;
  assign n30777 = ~po3897 & ~n30776;
  assign n30778 = pi0149 & ~po3897;
  assign n30779 = n19557 & n30778;
  assign po0419 = n30777 | n30779;
  assign n30781 = ~pi0715 & pi2020;
  assign n30782 = n26050 & ~n30781;
  assign n30783 = pi0150 & ~n30782;
  assign n30784 = n20388 & n20427;
  assign n30785 = ~n20389 & ~n30784;
  assign n30786 = ~pi0715 & ~n30785;
  assign n30787 = pi0715 & ~n24265;
  assign n30788 = ~n30786 & ~n30787;
  assign n30789 = n30782 & ~n30788;
  assign po0420 = n30783 | n30789;
  assign n30791 = ~pi0979 & n20522;
  assign n30792 = ~n30781 & n30791;
  assign n30793 = pi0151 & ~n30792;
  assign n30794 = ~n30788 & n30792;
  assign po0421 = n30793 | n30794;
  assign n30796 = pi0152 & n19557;
  assign n30797 = ~n19557 & ~n20370;
  assign n30798 = ~n30796 & ~n30797;
  assign po0422 = ~po3897 & ~n30798;
  assign n30800 = pi0153 & ~n30782;
  assign n30801 = ~pi0715 & ~n20388;
  assign n30802 = ~n28725 & n30801;
  assign n30803 = pi0715 & ~n30267;
  assign n30804 = ~n30802 & ~n30803;
  assign n30805 = ~pi0715 & n20388;
  assign n30806 = ~n20427 & n30805;
  assign n30807 = n30804 & ~n30806;
  assign n30808 = n30782 & ~n30807;
  assign po0423 = n30800 | n30808;
  assign n30810 = pi0154 & ~n30782;
  assign n30811 = n27813 & n30801;
  assign n30812 = pi0715 & ~n30288;
  assign n30813 = ~n30811 & ~n30812;
  assign n30814 = ~n30806 & n30813;
  assign n30815 = n30782 & ~n30814;
  assign po0424 = n30810 | n30815;
  assign n30817 = pi0155 & ~n30782;
  assign n30818 = n28234 & n30801;
  assign n30819 = pi0715 & ~n24744;
  assign n30820 = ~n30818 & ~n30819;
  assign n30821 = ~n30806 & n30820;
  assign n30822 = n30782 & ~n30821;
  assign po0425 = n30817 | n30822;
  assign n30824 = pi0156 & ~n30782;
  assign n30825 = ~n26654 & n30801;
  assign n30826 = pi0715 & ~n24769;
  assign n30827 = ~n30825 & ~n30826;
  assign n30828 = ~n30806 & n30827;
  assign n30829 = n30782 & ~n30828;
  assign po0426 = n30824 | n30829;
  assign n30831 = pi0157 & ~n30782;
  assign n30832 = n26896 & n30801;
  assign n30833 = pi0715 & ~n25699;
  assign n30834 = ~n30832 & ~n30833;
  assign n30835 = ~n30806 & n30834;
  assign n30836 = n30782 & ~n30835;
  assign po0427 = n30831 | n30836;
  assign n30838 = pi0158 & ~n30782;
  assign n30839 = ~n27134 & n30801;
  assign n30840 = pi0715 & ~n25718;
  assign n30841 = ~n30839 & ~n30840;
  assign n30842 = ~n30806 & n30841;
  assign n30843 = n30782 & ~n30842;
  assign po0428 = n30838 | n30843;
  assign n30845 = pi0159 & ~n30782;
  assign n30846 = n28307 & n30801;
  assign n30847 = pi0715 & ~n24256;
  assign n30848 = ~n30846 & ~n30847;
  assign n30849 = ~n30806 & n30848;
  assign n30850 = n30782 & ~n30849;
  assign po0429 = n30845 | n30850;
  assign n30852 = pi0160 & ~n30782;
  assign n30853 = ~n24900 & n30801;
  assign n30854 = pi0715 & ~n24289;
  assign n30855 = ~n30853 & ~n30854;
  assign n30856 = ~n30806 & n30855;
  assign n30857 = n30782 & ~n30856;
  assign po0430 = n30852 | n30857;
  assign n30859 = pi0161 & ~n30782;
  assign n30860 = ~n25761 & n30801;
  assign n30861 = pi0715 & ~n24446;
  assign n30862 = ~n30860 & ~n30861;
  assign n30863 = ~n30806 & n30862;
  assign n30864 = n30782 & ~n30863;
  assign po0431 = n30859 | n30864;
  assign n30866 = pi0162 & ~n30782;
  assign n30867 = ~n28969 & n30801;
  assign n30868 = pi0715 & ~n30309;
  assign n30869 = ~n30867 & ~n30868;
  assign n30870 = ~n30806 & n30869;
  assign n30871 = n30782 & ~n30870;
  assign po0432 = n30866 | n30871;
  assign n30873 = pi0163 & ~n30782;
  assign n30874 = n29216 & n30801;
  assign n30875 = pi0715 & ~n30321;
  assign n30876 = ~n30874 & ~n30875;
  assign n30877 = ~n30806 & n30876;
  assign n30878 = n30782 & ~n30877;
  assign po0433 = n30873 | n30878;
  assign n30880 = pi0164 & ~n30782;
  assign n30881 = ~n29458 & n30801;
  assign n30882 = pi0715 & ~n30333;
  assign n30883 = ~n30881 & ~n30882;
  assign n30884 = ~n30806 & n30883;
  assign n30885 = n30782 & ~n30884;
  assign po0434 = n30880 | n30885;
  assign n30887 = pi0165 & ~n30782;
  assign n30888 = n29708 & n30801;
  assign n30889 = pi0715 & ~n27570;
  assign n30890 = ~n30888 & ~n30889;
  assign n30891 = ~n30806 & n30890;
  assign n30892 = n30782 & ~n30891;
  assign po0435 = n30887 | n30892;
  assign n30894 = pi0166 & ~n30782;
  assign n30895 = n29959 & n30801;
  assign n30896 = pi0715 & ~n25999;
  assign n30897 = ~n30895 & ~n30896;
  assign n30898 = ~n30806 & n30897;
  assign n30899 = n30782 & ~n30898;
  assign po0436 = n30894 | n30899;
  assign n30901 = pi0167 & ~n30792;
  assign n30902 = n30792 & ~n30807;
  assign po0437 = n30901 | n30902;
  assign n30904 = pi0168 & ~n30792;
  assign n30905 = n30792 & ~n30814;
  assign po0438 = n30904 | n30905;
  assign n30907 = pi0169 & ~n30792;
  assign n30908 = n30792 & ~n30821;
  assign po0439 = n30907 | n30908;
  assign n30910 = pi0170 & ~n30792;
  assign n30911 = n30792 & ~n30828;
  assign po0440 = n30910 | n30911;
  assign n30913 = pi0171 & ~n30792;
  assign n30914 = n30792 & ~n30835;
  assign po0441 = n30913 | n30914;
  assign n30916 = pi0172 & ~n30792;
  assign n30917 = n30792 & ~n30842;
  assign po0442 = n30916 | n30917;
  assign n30919 = pi0173 & ~n30792;
  assign n30920 = n30792 & ~n30849;
  assign po0443 = n30919 | n30920;
  assign n30922 = pi0174 & ~n30782;
  assign n30923 = n30031 & n30801;
  assign n30924 = pi0715 & ~n24488;
  assign n30925 = ~n30923 & ~n30924;
  assign n30926 = ~n30806 & n30925;
  assign n30927 = n30782 & ~n30926;
  assign po0444 = n30922 | n30927;
  assign n30929 = pi0175 & ~n30792;
  assign n30930 = n30792 & ~n30856;
  assign po0445 = n30929 | n30930;
  assign n30932 = pi0176 & ~n30792;
  assign n30933 = n30792 & ~n30863;
  assign po0446 = n30932 | n30933;
  assign n30935 = pi0177 & ~n30792;
  assign n30936 = n30792 & ~n30870;
  assign po0447 = n30935 | n30936;
  assign n30938 = pi0178 & ~n30792;
  assign n30939 = n30792 & ~n30877;
  assign po0448 = n30938 | n30939;
  assign n30941 = pi0179 & ~n30792;
  assign n30942 = n30792 & ~n30884;
  assign po0449 = n30941 | n30942;
  assign n30944 = pi0180 & ~n30792;
  assign n30945 = n30792 & ~n30891;
  assign po0450 = n30944 | n30945;
  assign n30947 = pi0181 & ~n30792;
  assign n30948 = n30792 & ~n30898;
  assign po0451 = n30947 | n30948;
  assign n30950 = pi0182 & ~n30792;
  assign n30951 = n30792 & ~n30926;
  assign po0452 = n30950 | n30951;
  assign n30953 = pi0709 & n26050;
  assign n30954 = ~pi2140 & n26050;
  assign n30955 = ~n30953 & ~n30954;
  assign n30956 = ~pi0709 & ~n29363;
  assign n30957 = pi0709 & ~n30333;
  assign n30958 = ~n30956 & ~n30957;
  assign n30959 = ~n30955 & ~n30958;
  assign n30960 = pi0183 & n30955;
  assign po0453 = n30959 | n30960;
  assign n30962 = pi0709 & n20522;
  assign n30963 = ~pi0979 & n30962;
  assign n30964 = ~pi2140 & n20522;
  assign n30965 = ~pi0979 & n30964;
  assign n30966 = ~n30963 & ~n30965;
  assign n30967 = ~n30958 & ~n30966;
  assign n30968 = pi0184 & n30966;
  assign po0454 = n30967 | n30968;
  assign n30970 = n22754 & ~n22759;
  assign n30971 = ~n22754 & n22759;
  assign n30972 = ~n30970 & ~n30971;
  assign n30973 = ~n22751 & ~n26010;
  assign n30974 = ~n23291 & ~n30973;
  assign n30975 = ~n30972 & n30974;
  assign n30976 = n30972 & ~n30974;
  assign n30977 = ~n30975 & ~n30976;
  assign n30978 = pi0868 & ~n30977;
  assign n30979 = n22732 & n22750;
  assign n30980 = ~n22732 & ~n22750;
  assign n30981 = ~n30979 & ~n30980;
  assign n30982 = ~n26010 & ~n30981;
  assign n30983 = n26010 & n30981;
  assign n30984 = ~n30982 & ~n30983;
  assign n30985 = ~pi0868 & n30984;
  assign n30986 = ~n30978 & ~n30985;
  assign n30987 = n25637 & ~n30986;
  assign n30988 = pi0185 & n20518;
  assign n30989 = pi0185 & ~n24259;
  assign n30990 = n24259 & ~n25718;
  assign n30991 = ~n30989 & ~n30990;
  assign n30992 = n26002 & ~n30991;
  assign n30993 = ~n30988 & ~n30992;
  assign n30994 = ~n26006 & n30993;
  assign n30995 = ~n25637 & ~n30994;
  assign po0455 = n30987 | n30995;
  assign n30997 = n25663 & ~n30986;
  assign n30998 = pi0186 & n24300;
  assign n30999 = pi0186 & ~n24314;
  assign n31000 = n24314 & ~n25718;
  assign n31001 = ~n30999 & ~n31000;
  assign n31002 = n26041 & ~n31001;
  assign n31003 = ~n30998 & ~n31002;
  assign n31004 = ~n26045 & n31003;
  assign n31005 = ~n25663 & ~n31004;
  assign po0456 = n30997 | n31005;
  assign n31007 = n26051 & ~n30986;
  assign n31008 = ~pi0187 & ~n26051;
  assign po0457 = n31007 | n31008;
  assign n31010 = n26056 & ~n30986;
  assign n31011 = ~pi0188 & ~n26056;
  assign po0458 = n31010 | n31011;
  assign n31013 = ~pi0582 & pi3530;
  assign n31014 = ~pi0831 & n9365;
  assign po3448 = n31013 | n31014;
  assign n31016 = pi2599 & ~po3448;
  assign n31017 = ~pi0610 & n31013;
  assign n31018 = ~n31016 & ~n31017;
  assign n31019 = ~pi0189 & n31016;
  assign n31020 = ~n31018 & ~n31019;
  assign n31021 = ~pi2599 & ~n31013;
  assign n31022 = pi0189 & ~pi0955;
  assign n31023 = pi0955 & ~pi1017;
  assign n31024 = pi0278 & ~pi1017;
  assign n31025 = ~pi0278 & pi1017;
  assign n31026 = ~n31024 & ~n31025;
  assign n31027 = pi0248 & pi0329;
  assign n31028 = ~n31026 & n31027;
  assign n31029 = pi1017 & n31028;
  assign n31030 = ~pi0248 & ~pi0329;
  assign n31031 = n31026 & n31030;
  assign n31032 = ~n31026 & n31030;
  assign n31033 = ~pi0248 & pi0329;
  assign n31034 = n31026 & n31033;
  assign n31035 = n31032 & ~n31034;
  assign n31036 = pi0331 & ~pi1017;
  assign n31037 = ~pi0331 & pi1017;
  assign n31038 = ~n31036 & ~n31037;
  assign n31039 = n31034 & n31038;
  assign n31040 = ~n31035 & ~n31039;
  assign n31041 = ~n31031 & ~n31040;
  assign n31042 = ~pi0350 & n31031;
  assign n31043 = ~n31041 & ~n31042;
  assign n31044 = n31029 & n31043;
  assign n31045 = pi1017 & ~n31028;
  assign n31046 = ~n31043 & ~n31045;
  assign n31047 = ~n31031 & n31034;
  assign n31048 = n31031 & n31038;
  assign n31049 = ~n31047 & ~n31048;
  assign n31050 = n31045 & ~n31049;
  assign n31051 = ~n31046 & ~n31050;
  assign n31052 = ~n31029 & n31051;
  assign n31053 = ~n31044 & ~n31052;
  assign n31054 = pi0479 & n31032;
  assign n31055 = ~n31026 & n31033;
  assign n31056 = pi0248 & ~pi0329;
  assign n31057 = n31026 & n31056;
  assign n31058 = ~n31026 & n31056;
  assign n31059 = n31026 & n31027;
  assign n31060 = n31058 & ~n31059;
  assign n31061 = n31038 & n31059;
  assign n31062 = ~n31060 & ~n31061;
  assign n31063 = ~n31057 & ~n31062;
  assign n31064 = ~pi0350 & n31057;
  assign n31065 = ~n31063 & ~n31064;
  assign n31066 = ~n31055 & n31065;
  assign n31067 = pi0370 & ~pi1017;
  assign n31068 = ~pi0370 & pi1017;
  assign n31069 = ~n31067 & ~n31068;
  assign n31070 = n31055 & ~n31069;
  assign n31071 = ~n31066 & ~n31070;
  assign n31072 = ~n31032 & ~n31071;
  assign n31073 = ~n31054 & ~n31072;
  assign n31074 = ~n31031 & n31073;
  assign n31075 = ~n31047 & ~n31074;
  assign n31076 = ~n31045 & ~n31075;
  assign n31077 = n31032 & ~n31069;
  assign n31078 = n31038 & n31057;
  assign n31079 = ~n31057 & n31059;
  assign n31080 = ~n31078 & ~n31079;
  assign n31081 = ~n31055 & ~n31080;
  assign n31082 = ~pi0350 & n31055;
  assign n31083 = ~n31081 & ~n31082;
  assign n31084 = ~n31032 & n31083;
  assign n31085 = ~n31077 & ~n31084;
  assign n31086 = ~n31034 & ~n31085;
  assign n31087 = pi0479 & n31034;
  assign n31088 = ~n31086 & ~n31087;
  assign n31089 = ~n31031 & ~n31088;
  assign n31090 = n31045 & ~n31089;
  assign n31091 = ~n31076 & ~n31090;
  assign n31092 = ~n31029 & ~n31091;
  assign n31093 = n31029 & ~n31075;
  assign n31094 = ~n31092 & ~n31093;
  assign n31095 = pi0479 & n31055;
  assign n31096 = ~n31038 & n31060;
  assign n31097 = pi0350 & n31059;
  assign n31098 = ~n31096 & ~n31097;
  assign n31099 = ~n31057 & ~n31098;
  assign n31100 = n31057 & ~n31069;
  assign n31101 = ~n31099 & ~n31100;
  assign n31102 = ~n31055 & ~n31101;
  assign n31103 = ~n31095 & ~n31102;
  assign n31104 = ~n31034 & n31103;
  assign n31105 = ~n31035 & ~n31104;
  assign n31106 = ~n31031 & ~n31105;
  assign n31107 = ~n31045 & n31106;
  assign n31108 = n31045 & ~n31075;
  assign n31109 = ~n31107 & ~n31108;
  assign n31110 = ~n31029 & ~n31109;
  assign n31111 = ~n31031 & ~n31034;
  assign n31112 = ~n31032 & n31055;
  assign n31113 = ~pi0479 & n31057;
  assign n31114 = n31059 & ~n31069;
  assign n31115 = pi0350 & n31058;
  assign n31116 = ~n31038 & ~n31058;
  assign n31117 = ~n31115 & ~n31116;
  assign n31118 = ~n31059 & ~n31117;
  assign n31119 = ~n31114 & ~n31118;
  assign n31120 = ~n31057 & n31119;
  assign n31121 = ~n31113 & ~n31120;
  assign n31122 = ~n31032 & ~n31121;
  assign n31123 = ~n31112 & ~n31122;
  assign n31124 = n31111 & ~n31123;
  assign n31125 = ~n31045 & n31124;
  assign n31126 = n31045 & n31106;
  assign n31127 = ~n31125 & ~n31126;
  assign n31128 = ~n31029 & ~n31127;
  assign n31129 = n31029 & n31124;
  assign n31130 = ~n31128 & ~n31129;
  assign n31131 = ~n31055 & n31057;
  assign n31132 = pi0479 & n31059;
  assign n31133 = n31058 & n31069;
  assign n31134 = ~pi0350 & ~n31058;
  assign n31135 = ~n31133 & ~n31134;
  assign n31136 = ~n31059 & n31135;
  assign n31137 = ~n31132 & ~n31136;
  assign n31138 = ~n31055 & n31137;
  assign n31139 = ~n31131 & ~n31138;
  assign n31140 = ~n31032 & ~n31034;
  assign n31141 = ~n31031 & n31140;
  assign n31142 = ~n31139 & n31141;
  assign n31143 = n31029 & ~n31142;
  assign n31144 = ~n31045 & n31142;
  assign n31145 = n31045 & n31124;
  assign n31146 = ~n31144 & ~n31145;
  assign n31147 = ~n31029 & n31146;
  assign n31148 = ~n31143 & ~n31147;
  assign n31149 = pi0479 & n31058;
  assign n31150 = ~n31058 & ~n31069;
  assign n31151 = ~n31149 & ~n31150;
  assign n31152 = ~n31059 & ~n31151;
  assign n31153 = n31111 & ~n31152;
  assign n31154 = ~n31055 & ~n31057;
  assign n31155 = n31153 & n31154;
  assign n31156 = ~n31032 & n31155;
  assign n31157 = n31029 & ~n31156;
  assign n31158 = ~n31045 & ~n31156;
  assign n31159 = n31045 & ~n31142;
  assign n31160 = ~n31158 & ~n31159;
  assign n31161 = ~n31029 & ~n31160;
  assign n31162 = ~n31157 & ~n31161;
  assign n31163 = pi0479 & ~n31058;
  assign n31164 = n31154 & ~n31163;
  assign n31165 = ~n31032 & ~n31059;
  assign n31166 = n31111 & n31165;
  assign n31167 = n31164 & n31166;
  assign n31168 = n31029 & ~n31167;
  assign n31169 = ~n31045 & ~n31167;
  assign n31170 = n31045 & ~n31156;
  assign n31171 = ~n31169 & ~n31170;
  assign n31172 = ~n31029 & ~n31171;
  assign n31173 = ~n31168 & ~n31172;
  assign n31174 = ~n31055 & ~n31059;
  assign n31175 = ~n31032 & ~n31057;
  assign n31176 = n31111 & n31175;
  assign n31177 = ~n31058 & n31176;
  assign n31178 = n31174 & n31177;
  assign n31179 = ~n31045 & ~n31178;
  assign n31180 = n31045 & ~n31167;
  assign n31181 = ~n31179 & ~n31180;
  assign n31182 = ~n31029 & ~n31181;
  assign n31183 = n31029 & ~n31178;
  assign n31184 = ~n31182 & ~n31183;
  assign n31185 = ~n31173 & ~n31184;
  assign n31186 = ~n31162 & n31185;
  assign n31187 = ~n31148 & n31186;
  assign n31188 = n31130 & n31187;
  assign n31189 = n31110 & ~n31188;
  assign n31190 = n31094 & ~n31189;
  assign n31191 = n31029 & ~n31089;
  assign n31192 = ~n31045 & ~n31089;
  assign n31193 = pi0479 & n31031;
  assign n31194 = ~pi0350 & n31032;
  assign n31195 = n31038 & n31055;
  assign n31196 = ~n31131 & ~n31195;
  assign n31197 = ~n31032 & ~n31196;
  assign n31198 = ~n31194 & ~n31197;
  assign n31199 = ~n31034 & n31198;
  assign n31200 = n31034 & ~n31069;
  assign n31201 = ~n31199 & ~n31200;
  assign n31202 = ~n31031 & ~n31201;
  assign n31203 = ~n31193 & ~n31202;
  assign n31204 = n31045 & n31203;
  assign n31205 = ~n31192 & ~n31204;
  assign n31206 = ~n31029 & ~n31205;
  assign n31207 = ~n31191 & ~n31206;
  assign n31208 = n31190 & n31207;
  assign n31209 = n31029 & ~n31203;
  assign n31210 = ~n31045 & ~n31203;
  assign n31211 = n31031 & ~n31069;
  assign n31212 = n31032 & n31038;
  assign n31213 = ~n31112 & ~n31212;
  assign n31214 = ~n31034 & ~n31213;
  assign n31215 = ~pi0350 & n31034;
  assign n31216 = ~n31214 & ~n31215;
  assign n31217 = ~n31031 & n31216;
  assign n31218 = ~n31211 & ~n31217;
  assign n31219 = n31045 & ~n31218;
  assign n31220 = ~n31210 & ~n31219;
  assign n31221 = ~n31029 & ~n31220;
  assign n31222 = ~n31209 & ~n31221;
  assign n31223 = n31029 & ~n31218;
  assign n31224 = ~n31045 & ~n31218;
  assign n31225 = n31043 & n31045;
  assign n31226 = ~n31224 & ~n31225;
  assign n31227 = ~n31029 & ~n31226;
  assign n31228 = ~n31223 & ~n31227;
  assign n31229 = ~n31222 & ~n31228;
  assign n31230 = n31208 & n31229;
  assign n31231 = ~n31053 & n31230;
  assign n31232 = ~n31045 & ~n31049;
  assign n31233 = n31031 & n31045;
  assign n31234 = ~n31232 & ~n31233;
  assign n31235 = ~n31029 & ~n31234;
  assign n31236 = n31029 & ~n31049;
  assign n31237 = ~n31235 & ~n31236;
  assign n31238 = ~n31231 & ~n31237;
  assign n31239 = n31231 & n31237;
  assign n31240 = ~n31238 & ~n31239;
  assign n31241 = ~pi1017 & ~n31240;
  assign n31242 = pi1017 & ~n31237;
  assign n31243 = ~n31241 & ~n31242;
  assign n31244 = n31207 & ~n31222;
  assign n31245 = n31130 & ~n31148;
  assign n31246 = n31186 & n31245;
  assign n31247 = n31110 & ~n31246;
  assign n31248 = n31094 & ~n31247;
  assign n31249 = ~n31228 & n31248;
  assign n31250 = n31244 & n31249;
  assign n31251 = n31053 & n31250;
  assign n31252 = ~n31053 & ~n31250;
  assign n31253 = ~n31251 & ~n31252;
  assign n31254 = ~pi1017 & n31253;
  assign n31255 = pi1017 & n31053;
  assign n31256 = ~n31254 & ~n31255;
  assign n31257 = n31243 & n31256;
  assign n31258 = pi1017 & n31228;
  assign n31259 = ~n31162 & ~n31173;
  assign n31260 = n31245 & n31259;
  assign n31261 = n31110 & ~n31260;
  assign n31262 = n31094 & ~n31261;
  assign n31263 = n31110 & n31184;
  assign n31264 = n31244 & ~n31263;
  assign n31265 = n31262 & n31264;
  assign n31266 = n31228 & ~n31265;
  assign n31267 = ~n31228 & n31265;
  assign n31268 = ~n31266 & ~n31267;
  assign n31269 = ~pi1017 & ~n31268;
  assign n31270 = ~n31258 & ~n31269;
  assign n31271 = ~pi1017 & ~n31208;
  assign n31272 = ~pi1017 & ~n31271;
  assign n31273 = n31222 & ~n31272;
  assign n31274 = n31208 & ~n31222;
  assign n31275 = ~pi1017 & n31274;
  assign n31276 = ~n31273 & ~n31275;
  assign n31277 = ~pi1017 & ~n31190;
  assign n31278 = ~pi1017 & ~n31277;
  assign n31279 = ~n31207 & ~n31278;
  assign n31280 = ~pi1017 & n31208;
  assign n31281 = ~n31279 & ~n31280;
  assign n31282 = ~pi1017 & n31247;
  assign n31283 = ~pi1017 & ~n31282;
  assign n31284 = ~n31094 & ~n31283;
  assign n31285 = ~pi1017 & n31248;
  assign n31286 = ~n31284 & ~n31285;
  assign n31287 = pi1017 & n31110;
  assign n31288 = ~n31184 & n31260;
  assign n31289 = n31110 & ~n31288;
  assign n31290 = ~n31110 & n31288;
  assign n31291 = ~n31289 & ~n31290;
  assign n31292 = ~pi1017 & n31291;
  assign n31293 = ~n31287 & ~n31292;
  assign n31294 = ~pi1017 & ~n31186;
  assign n31295 = ~pi1017 & ~n31294;
  assign n31296 = n31148 & ~n31295;
  assign n31297 = ~pi1017 & n31187;
  assign n31298 = ~n31296 & ~n31297;
  assign n31299 = ~pi1017 & ~n31185;
  assign n31300 = ~pi1017 & ~n31299;
  assign n31301 = n31162 & ~n31300;
  assign n31302 = ~pi1017 & n31186;
  assign n31303 = ~n31301 & ~n31302;
  assign n31304 = ~pi1017 & n31184;
  assign n31305 = ~pi1017 & ~n31304;
  assign n31306 = n31173 & ~n31305;
  assign n31307 = ~pi1017 & n31185;
  assign n31308 = ~n31306 & ~n31307;
  assign n31309 = ~pi1017 & ~n31184;
  assign n31310 = pi1017 & n31184;
  assign n31311 = ~n31309 & ~n31310;
  assign n31312 = n31308 & n31311;
  assign n31313 = n31303 & n31312;
  assign n31314 = n31298 & n31313;
  assign n31315 = n31293 & n31314;
  assign n31316 = ~pi1017 & ~n31187;
  assign n31317 = ~pi1017 & ~n31316;
  assign n31318 = ~n31130 & ~n31317;
  assign n31319 = ~pi1017 & n31188;
  assign n31320 = ~n31318 & ~n31319;
  assign n31321 = n31315 & n31320;
  assign n31322 = n31286 & n31321;
  assign n31323 = n31281 & n31322;
  assign n31324 = n31276 & n31323;
  assign n31325 = n31270 & n31324;
  assign n31326 = n31257 & n31325;
  assign n31327 = ~n31029 & n31045;
  assign n31328 = n31031 & ~n31327;
  assign n31329 = ~n31053 & ~n31228;
  assign n31330 = n31274 & n31329;
  assign n31331 = n31237 & n31330;
  assign n31332 = ~n31328 & ~n31331;
  assign n31333 = n31328 & n31331;
  assign n31334 = ~n31332 & ~n31333;
  assign n31335 = ~pi1017 & n31334;
  assign n31336 = pi1017 & n31328;
  assign n31337 = ~n31335 & ~n31336;
  assign n31338 = ~n31326 & ~n31337;
  assign n31339 = n31326 & n31337;
  assign n31340 = ~n31338 & ~n31339;
  assign n31341 = ~pi0247 & n31340;
  assign n31342 = pi0247 & ~n31337;
  assign n31343 = ~n31341 & ~n31342;
  assign n31344 = n31023 & ~n31343;
  assign n31345 = ~n31022 & ~n31344;
  assign n31346 = ~pi0247 & pi0955;
  assign n31347 = pi1017 & n31346;
  assign n31348 = n31345 & ~n31347;
  assign n31349 = n31021 & ~n31348;
  assign n31350 = pi2599 & ~n31013;
  assign n31351 = ~n10608 & n31350;
  assign n31352 = ~n31349 & ~n31351;
  assign n31353 = ~n31016 & ~n31352;
  assign po0459 = n31020 | n31353;
  assign n31355 = pi0190 & n20518;
  assign n31356 = pi0190 & ~n24259;
  assign n31357 = n24259 & ~n25699;
  assign n31358 = ~n31356 & ~n31357;
  assign n31359 = n26002 & ~n31358;
  assign n31360 = ~n31355 & ~n31359;
  assign n31361 = ~n26006 & n31360;
  assign n31362 = ~n25637 & ~n31361;
  assign n31363 = ~pi0868 & ~n30977;
  assign n31364 = pi0868 & ~n30585;
  assign n31365 = ~n31363 & ~n31364;
  assign n31366 = n25637 & ~n31365;
  assign po0460 = n31362 | n31366;
  assign n31368 = pi0191 & n24300;
  assign n31369 = pi0191 & ~n24314;
  assign n31370 = n24314 & ~n25699;
  assign n31371 = ~n31369 & ~n31370;
  assign n31372 = n26041 & ~n31371;
  assign n31373 = ~n31368 & ~n31372;
  assign n31374 = ~n26045 & n31373;
  assign n31375 = ~n25663 & ~n31374;
  assign n31376 = n25663 & ~n31365;
  assign po0461 = n31375 | n31376;
  assign n31378 = pi0979 & n24865;
  assign n31379 = pi0979 & n20515;
  assign n31380 = ~n20512 & ~n31379;
  assign n31381 = ~n31378 & n31380;
  assign n31382 = n20523 & ~n31381;
  assign n31383 = pi0192 & n31381;
  assign n31384 = ~n9352 & n31378;
  assign n31385 = ~n24265 & n31384;
  assign n31386 = pi0192 & ~n31384;
  assign n31387 = ~n31385 & ~n31386;
  assign n31388 = ~n24260 & ~n31381;
  assign n31389 = ~n31387 & n31388;
  assign n31390 = ~n31383 & ~n31389;
  assign n31391 = n26005 & ~n31381;
  assign n31392 = n31390 & ~n31391;
  assign n31393 = ~n31382 & ~n31392;
  assign n31394 = ~n27670 & n31382;
  assign po0462 = n31393 | n31394;
  assign n31396 = ~pi0979 & n24865;
  assign n31397 = ~pi0979 & n20515;
  assign n31398 = ~n24298 & ~n31397;
  assign n31399 = ~n31396 & n31398;
  assign n31400 = n24303 & ~n31399;
  assign n31401 = pi0193 & n31399;
  assign n31402 = ~n9352 & n31396;
  assign n31403 = ~n24265 & n31402;
  assign n31404 = pi0193 & ~n31402;
  assign n31405 = ~n31403 & ~n31404;
  assign n31406 = ~n24315 & ~n31399;
  assign n31407 = ~n31405 & n31406;
  assign n31408 = ~n31401 & ~n31407;
  assign n31409 = n26044 & ~n31399;
  assign n31410 = n31408 & ~n31409;
  assign n31411 = ~n31400 & ~n31410;
  assign n31412 = ~n27670 & n31400;
  assign po0463 = n31411 | n31412;
  assign n31414 = ~pi0194 & ~n26051;
  assign n31415 = n26051 & ~n31365;
  assign po0464 = n31414 | n31415;
  assign n31417 = ~pi0195 & ~n26056;
  assign n31418 = n26056 & ~n31365;
  assign po0465 = n31417 | n31418;
  assign n31420 = pi0196 & n19557;
  assign n31421 = ~n19557 & ~n20445;
  assign n31422 = ~n31420 & ~n31421;
  assign po0466 = ~po3897 & ~n31422;
  assign n31424 = pi0709 & ~n30267;
  assign n31425 = ~pi0709 & ~n28700;
  assign n31426 = ~n31424 & ~n31425;
  assign n31427 = ~n30955 & ~n31426;
  assign n31428 = pi0197 & n30955;
  assign po0467 = n31427 | n31428;
  assign n31430 = ~n30966 & ~n31426;
  assign n31431 = pi0198 & n30966;
  assign po0468 = n31430 | n31431;
  assign n31433 = pi3516 & n24928;
  assign n31434 = pi3518 & n31433;
  assign n31435 = ~pi2021 & n24928;
  assign n31436 = pi3516 & ~pi3518;
  assign n31437 = pi0152 & n31436;
  assign n31438 = n31435 & n31437;
  assign n31439 = n19587 & n31435;
  assign n31440 = ~n25053 & n31435;
  assign n31441 = ~pi0586 & n31440;
  assign n31442 = pi0586 & ~n31440;
  assign n31443 = ~n31441 & ~n31442;
  assign n31444 = n31439 & ~n31443;
  assign n31445 = ~n31438 & n31444;
  assign n31446 = ~n25245 & n31435;
  assign n31447 = n31440 & n31446;
  assign n31448 = ~n31440 & ~n31446;
  assign n31449 = ~n31447 & ~n31448;
  assign n31450 = n31439 & n31449;
  assign n31451 = ~n31439 & ~n31449;
  assign n31452 = ~n31450 & ~n31451;
  assign n31453 = ~n31438 & ~n31452;
  assign n31454 = ~n31445 & ~n31453;
  assign n31455 = ~n9534 & n31454;
  assign n31456 = ~n31438 & ~n31449;
  assign n31457 = ~n25250 & n31435;
  assign n31458 = ~n31440 & n31457;
  assign n31459 = n31440 & ~n31457;
  assign n31460 = ~n31458 & ~n31459;
  assign n31461 = ~n25031 & n31435;
  assign n31462 = ~n31440 & n31461;
  assign n31463 = n31440 & ~n31461;
  assign n31464 = ~n31462 & ~n31463;
  assign n31465 = n31460 & n31464;
  assign n31466 = ~n24931 & n31435;
  assign n31467 = ~n31440 & ~n31466;
  assign n31468 = n31440 & n31466;
  assign n31469 = ~n31467 & ~n31468;
  assign n31470 = ~n25148 & n31435;
  assign n31471 = ~n31440 & n31470;
  assign n31472 = n31440 & ~n31470;
  assign n31473 = ~n31471 & ~n31472;
  assign n31474 = ~n31469 & n31473;
  assign n31475 = ~n25236 & n31435;
  assign n31476 = ~n31440 & n31475;
  assign n31477 = n31440 & ~n31475;
  assign n31478 = ~n31476 & ~n31477;
  assign n31479 = ~n25102 & n31435;
  assign n31480 = n31440 & n31479;
  assign n31481 = ~n31440 & ~n31479;
  assign n31482 = ~n31480 & ~n31481;
  assign n31483 = n31478 & ~n31482;
  assign n31484 = ~n25164 & n31435;
  assign n31485 = ~n31440 & n31484;
  assign n31486 = n31440 & ~n31484;
  assign n31487 = ~n31485 & ~n31486;
  assign n31488 = n31483 & n31487;
  assign n31489 = ~n25157 & n31435;
  assign n31490 = n31440 & n31489;
  assign n31491 = ~n31440 & ~n31489;
  assign n31492 = ~n31490 & ~n31491;
  assign n31493 = n31488 & ~n31492;
  assign n31494 = n31474 & n31493;
  assign n31495 = n31465 & n31494;
  assign n31496 = ~n31444 & ~n31495;
  assign n31497 = n31456 & n31496;
  assign n31498 = ~n25201 & n31435;
  assign n31499 = n31440 & ~n31498;
  assign n31500 = ~n31440 & n31498;
  assign n31501 = ~n31499 & ~n31500;
  assign n31502 = ~n25266 & n31435;
  assign n31503 = ~n31440 & n31502;
  assign n31504 = n31440 & ~n31502;
  assign n31505 = ~n31503 & ~n31504;
  assign n31506 = ~n25197 & n31435;
  assign n31507 = ~n31440 & ~n31506;
  assign n31508 = n31440 & n31506;
  assign n31509 = ~n31507 & ~n31508;
  assign n31510 = ~n25229 & n31435;
  assign n31511 = ~n31440 & n31510;
  assign n31512 = n31440 & ~n31510;
  assign n31513 = ~n31511 & ~n31512;
  assign n31514 = ~n31509 & n31513;
  assign n31515 = n31505 & n31514;
  assign n31516 = n31501 & n31515;
  assign n31517 = n31473 & n31487;
  assign n31518 = ~n31492 & n31517;
  assign n31519 = ~n31469 & n31518;
  assign n31520 = ~n31516 & n31519;
  assign n31521 = n31465 & n31478;
  assign n31522 = ~n31482 & n31521;
  assign n31523 = ~n31520 & n31522;
  assign n31524 = n31456 & ~n31523;
  assign n31525 = ~n31444 & n31524;
  assign n31526 = ~n31497 & ~n31525;
  assign n31527 = ~n14618 & ~n31525;
  assign n31528 = ~n31526 & ~n31527;
  assign n31529 = ~n15006 & ~n31528;
  assign n31530 = ~n14618 & ~n31497;
  assign n31531 = ~n31529 & ~n31530;
  assign n31532 = n14618 & n31497;
  assign n31533 = ~n15006 & ~n31532;
  assign n31534 = n31528 & ~n31533;
  assign n31535 = n31487 & ~n31492;
  assign n31536 = n31505 & ~n31509;
  assign n31537 = ~n25289 & n31435;
  assign n31538 = n31440 & ~n31537;
  assign n31539 = ~n31440 & n31537;
  assign n31540 = ~n31538 & ~n31539;
  assign n31541 = ~n25040 & n31435;
  assign n31542 = ~n31440 & ~n31541;
  assign n31543 = n31440 & n31541;
  assign n31544 = ~n31542 & ~n31543;
  assign n31545 = n31540 & ~n31544;
  assign n31546 = n31513 & ~n31545;
  assign n31547 = n31501 & n31546;
  assign n31548 = n31536 & ~n31547;
  assign n31549 = n31474 & ~n31548;
  assign n31550 = n31535 & ~n31549;
  assign n31551 = ~n31482 & ~n31550;
  assign n31552 = n31478 & n31551;
  assign n31553 = n31465 & ~n31552;
  assign n31554 = n31456 & ~n31553;
  assign n31555 = ~n31444 & n31554;
  assign n31556 = n11850 & n31555;
  assign n31557 = ~n31540 & ~n31544;
  assign n31558 = n31513 & ~n31557;
  assign n31559 = n31501 & ~n31558;
  assign n31560 = n31505 & ~n31559;
  assign n31561 = ~n31509 & ~n31560;
  assign n31562 = ~n31469 & ~n31561;
  assign n31563 = n31473 & ~n31562;
  assign n31564 = n31487 & ~n31563;
  assign n31565 = ~n31492 & ~n31564;
  assign n31566 = ~n31482 & ~n31565;
  assign n31567 = n31478 & ~n31566;
  assign n31568 = n31464 & ~n31567;
  assign n31569 = n31460 & ~n31568;
  assign n31570 = ~n31449 & ~n31569;
  assign n31571 = ~n31438 & ~n31570;
  assign n31572 = ~n31444 & n31571;
  assign n31573 = n11033 & ~n31572;
  assign n31574 = ~n11850 & ~n31555;
  assign n31575 = n31573 & ~n31574;
  assign n31576 = ~n31556 & ~n31575;
  assign n31577 = ~n31534 & n31576;
  assign n31578 = n31531 & ~n31577;
  assign n31579 = ~n9534 & ~n31454;
  assign n31580 = n9534 & n31454;
  assign n31581 = ~n31579 & ~n31580;
  assign n31582 = n31578 & ~n31581;
  assign n31583 = ~n31455 & ~n31582;
  assign n31584 = n31434 & ~n31583;
  assign n31585 = ~pi2021 & n31434;
  assign n31586 = n19553 & n31585;
  assign n31587 = n31584 & n31586;
  assign n31588 = pi0867 & ~pi3426;
  assign n31589 = ~n31587 & ~n31588;
  assign n31590 = n24251 & ~n31589;
  assign n31591 = pi0867 & ~n12415;
  assign n31592 = ~pi0867 & ~n31454;
  assign n31593 = ~n31591 & ~n31592;
  assign n31594 = n31590 & ~n31593;
  assign n31595 = pi0199 & ~n31590;
  assign po0469 = n31594 | n31595;
  assign n31597 = ~pi0867 & n31497;
  assign n31598 = pi0867 & ~n14816;
  assign n31599 = ~n31597 & ~n31598;
  assign n31600 = n31590 & ~n31599;
  assign n31601 = pi0200 & ~n31590;
  assign po0470 = n31600 | n31601;
  assign n31603 = pi0867 & ~n15115;
  assign n31604 = ~pi0867 & n31525;
  assign n31605 = ~n31603 & ~n31604;
  assign n31606 = n31590 & ~n31605;
  assign n31607 = pi0201 & ~n31590;
  assign po0471 = n31606 | n31607;
  assign n31609 = pi0867 & ~n12061;
  assign n31610 = ~pi0867 & n31555;
  assign n31611 = ~n31609 & ~n31610;
  assign n31612 = n31590 & ~n31611;
  assign n31613 = pi0202 & ~n31590;
  assign po0472 = n31612 | n31613;
  assign n31615 = n24309 & ~n31589;
  assign n31616 = ~n31593 & n31615;
  assign n31617 = pi0203 & ~n31615;
  assign po0473 = n31616 | n31617;
  assign n31619 = ~n31599 & n31615;
  assign n31620 = pi0204 & ~n31615;
  assign po0474 = n31619 | n31620;
  assign n31622 = ~pi0867 & ~n31572;
  assign n31623 = pi0867 & ~n11181;
  assign n31624 = ~n31622 & ~n31623;
  assign n31625 = n31590 & ~n31624;
  assign n31626 = pi0205 & ~n31590;
  assign po0475 = n31625 | n31626;
  assign n31628 = ~n31611 & n31615;
  assign n31629 = pi0206 & ~n31615;
  assign po0476 = n31628 | n31629;
  assign n31631 = ~n31605 & n31615;
  assign n31632 = pi0207 & ~n31615;
  assign po0477 = n31631 | n31632;
  assign n31634 = n31615 & ~n31624;
  assign n31635 = pi0208 & ~n31615;
  assign po0478 = n31634 | n31635;
  assign n31637 = ~n24091 & ~n24095;
  assign n31638 = n23280 & ~n31637;
  assign n31639 = ~n23020 & ~n23284;
  assign n31640 = ~n31638 & n31639;
  assign n31641 = n31638 & ~n31639;
  assign n31642 = ~n31640 & ~n31641;
  assign n31643 = pi0868 & n31642;
  assign n31644 = ~pi0868 & n27595;
  assign n31645 = ~n31643 & ~n31644;
  assign n31646 = n25637 & ~n31645;
  assign n31647 = pi0209 & n20518;
  assign n31648 = pi0209 & ~n24259;
  assign n31649 = n24259 & ~n24446;
  assign n31650 = ~n31648 & ~n31649;
  assign n31651 = n26002 & ~n31650;
  assign n31652 = ~n31647 & ~n31651;
  assign n31653 = ~n26006 & n31652;
  assign n31654 = ~n25637 & ~n31653;
  assign po0479 = n31646 | n31654;
  assign n31656 = n25663 & ~n31645;
  assign n31657 = pi0210 & n24300;
  assign n31658 = pi0210 & ~n24314;
  assign n31659 = n24314 & ~n24446;
  assign n31660 = ~n31658 & ~n31659;
  assign n31661 = n26041 & ~n31660;
  assign n31662 = ~n31657 & ~n31661;
  assign n31663 = ~n26045 & n31662;
  assign n31664 = ~n25663 & ~n31663;
  assign po0480 = n31656 | n31664;
  assign n31666 = ~n27677 & n31382;
  assign n31667 = pi0211 & n31381;
  assign n31668 = ~n30309 & n31384;
  assign n31669 = pi0211 & ~n31384;
  assign n31670 = ~n31668 & ~n31669;
  assign n31671 = n31388 & ~n31670;
  assign n31672 = ~n31667 & ~n31671;
  assign n31673 = ~n31391 & n31672;
  assign n31674 = ~n31382 & ~n31673;
  assign po0481 = n31666 | n31674;
  assign n31676 = ~n27677 & n31400;
  assign n31677 = pi0212 & n31399;
  assign n31678 = ~n30309 & n31402;
  assign n31679 = pi0212 & ~n31402;
  assign n31680 = ~n31678 & ~n31679;
  assign n31681 = n31406 & ~n31680;
  assign n31682 = ~n31677 & ~n31681;
  assign n31683 = ~n31409 & n31682;
  assign n31684 = ~n31400 & ~n31683;
  assign po0482 = n31676 | n31684;
  assign n31686 = n26051 & ~n31645;
  assign n31687 = ~pi0213 & ~n26051;
  assign po0483 = n31686 | n31687;
  assign n31689 = n26056 & ~n31645;
  assign n31690 = ~pi0214 & ~n26056;
  assign po0484 = n31689 | n31690;
  assign n31692 = pi0868 & n30984;
  assign n31693 = ~n23020 & ~n23280;
  assign n31694 = ~n23020 & n31637;
  assign n31695 = ~n23284 & ~n31694;
  assign n31696 = ~n31693 & n31695;
  assign n31697 = ~n22915 & ~n23282;
  assign n31698 = ~n31696 & n31697;
  assign n31699 = n31696 & ~n31697;
  assign n31700 = ~n31698 & ~n31699;
  assign n31701 = ~pi0868 & n31700;
  assign n31702 = ~n31692 & ~n31701;
  assign n31703 = n25637 & ~n31702;
  assign n31704 = pi0215 & n20518;
  assign n31705 = pi0215 & ~n24259;
  assign n31706 = ~n24256 & n24259;
  assign n31707 = ~n31705 & ~n31706;
  assign n31708 = n26002 & ~n31707;
  assign n31709 = ~n31704 & ~n31708;
  assign n31710 = ~n26006 & n31709;
  assign n31711 = ~n25637 & ~n31710;
  assign po0485 = n31703 | n31711;
  assign n31713 = ~pi0868 & n31642;
  assign n31714 = pi0868 & n31700;
  assign n31715 = ~n31713 & ~n31714;
  assign n31716 = n25637 & ~n31715;
  assign n31717 = pi0216 & n20518;
  assign n31718 = pi0216 & ~n24259;
  assign n31719 = n24259 & ~n24289;
  assign n31720 = ~n31718 & ~n31719;
  assign n31721 = n26002 & ~n31720;
  assign n31722 = ~n31717 & ~n31721;
  assign n31723 = ~n26006 & n31722;
  assign n31724 = ~n25637 & ~n31723;
  assign po0486 = n31716 | n31724;
  assign n31726 = n25663 & ~n31715;
  assign n31727 = pi0217 & n24300;
  assign n31728 = pi0217 & ~n24314;
  assign n31729 = ~n24289 & n24314;
  assign n31730 = ~n31728 & ~n31729;
  assign n31731 = n26041 & ~n31730;
  assign n31732 = ~n31727 & ~n31731;
  assign n31733 = ~n26045 & n31732;
  assign n31734 = ~n25663 & ~n31733;
  assign po0487 = n31726 | n31734;
  assign n31736 = n25663 & ~n31702;
  assign n31737 = pi0218 & n24300;
  assign n31738 = pi0218 & ~n24314;
  assign n31739 = ~n24256 & n24314;
  assign n31740 = ~n31738 & ~n31739;
  assign n31741 = n26041 & ~n31740;
  assign n31742 = ~n31737 & ~n31741;
  assign n31743 = ~n26045 & n31742;
  assign n31744 = ~n25663 & ~n31743;
  assign po0488 = n31736 | n31744;
  assign n31746 = n26051 & ~n31702;
  assign n31747 = ~pi0219 & ~n26051;
  assign po0489 = n31746 | n31747;
  assign n31749 = n26051 & ~n31715;
  assign n31750 = ~pi0220 & ~n26051;
  assign po0490 = n31749 | n31750;
  assign n31752 = n26056 & ~n31702;
  assign n31753 = ~pi0221 & ~n26056;
  assign po0491 = n31752 | n31753;
  assign n31755 = n26056 & ~n31715;
  assign n31756 = ~pi0222 & ~n26056;
  assign po0492 = n31755 | n31756;
  assign n31758 = ~pi1426 & ~po3853;
  assign n31759 = pi1426 & ~po1235;
  assign po0494 = n31758 | n31759;
  assign n31761 = pi0827 & ~pi3681;
  assign n31762 = ~pi0496 & ~pi0577;
  assign n31763 = ~pi0653 & ~pi0863;
  assign n31764 = ~pi0398 & ~pi0458;
  assign n31765 = ~pi0336 & ~pi0367;
  assign n31766 = ~pi0223 & ~pi0246;
  assign n31767 = ~pi0277 & ~pi0303;
  assign n31768 = n31766 & n31767;
  assign n31769 = n31765 & n31768;
  assign n31770 = n31764 & n31769;
  assign n31771 = ~pi0849 & n31770;
  assign n31772 = n31763 & n31771;
  assign n31773 = n31762 & n31772;
  assign n31774 = ~pi0822 & n31773;
  assign n31775 = ~pi0699 & n31774;
  assign n31776 = ~pi0728 & n31775;
  assign n31777 = n31761 & n31776;
  assign n31778 = ~pi3472 & ~pi3681;
  assign n31779 = ~pi3438 & n31778;
  assign n31780 = pi1722 & ~n31779;
  assign n31781 = n31777 & n31780;
  assign n31782 = ~pi2095 & n31779;
  assign n31783 = ~n31781 & ~n31782;
  assign n31784 = ~pi0728 & ~pi0822;
  assign n31785 = ~pi0699 & ~pi0849;
  assign n31786 = n31784 & n31785;
  assign n31787 = ~pi3681 & ~n31786;
  assign n31788 = pi0863 & n31787;
  assign n31789 = pi0653 & n31788;
  assign n31790 = pi0496 & n31789;
  assign n31791 = pi0577 & n31790;
  assign n31792 = pi0577 & n31789;
  assign n31793 = pi0496 & n31792;
  assign n31794 = ~pi0496 & ~n31792;
  assign n31795 = ~n31793 & ~n31794;
  assign n31796 = ~pi0577 & ~n31789;
  assign n31797 = ~n31792 & ~n31796;
  assign n31798 = ~pi0653 & ~n31788;
  assign n31799 = ~n31789 & ~n31798;
  assign n31800 = ~pi0863 & ~n31787;
  assign n31801 = ~n31788 & ~n31800;
  assign n31802 = ~n31799 & ~n31801;
  assign n31803 = ~n31797 & n31802;
  assign n31804 = ~n31795 & n31803;
  assign n31805 = ~n31791 & n31804;
  assign n31806 = n31791 & ~n31804;
  assign n31807 = ~n31805 & ~n31806;
  assign n31808 = ~pi3681 & n31807;
  assign n31809 = pi0458 & n31808;
  assign n31810 = pi0398 & n31809;
  assign n31811 = pi0336 & n31810;
  assign n31812 = pi0367 & n31811;
  assign n31813 = pi0367 & n31810;
  assign n31814 = pi0336 & n31813;
  assign n31815 = ~pi0336 & ~n31813;
  assign n31816 = ~n31814 & ~n31815;
  assign n31817 = ~pi0367 & ~n31810;
  assign n31818 = ~n31813 & ~n31817;
  assign n31819 = ~pi0398 & ~n31809;
  assign n31820 = ~n31810 & ~n31819;
  assign n31821 = ~pi0458 & ~n31808;
  assign n31822 = ~n31809 & ~n31821;
  assign n31823 = ~n31820 & ~n31822;
  assign n31824 = ~n31818 & n31823;
  assign n31825 = ~n31816 & n31824;
  assign n31826 = ~n31812 & n31825;
  assign n31827 = n31812 & ~n31825;
  assign n31828 = ~n31826 & ~n31827;
  assign n31829 = ~pi3681 & n31828;
  assign n31830 = pi0303 & n31829;
  assign n31831 = pi0277 & n31830;
  assign n31832 = pi0246 & n31831;
  assign n31833 = pi0223 & ~n31832;
  assign n31834 = ~pi0277 & ~n31830;
  assign n31835 = ~n31831 & ~n31834;
  assign n31836 = ~pi0303 & ~n31829;
  assign n31837 = ~n31830 & ~n31836;
  assign n31838 = ~n31835 & ~n31837;
  assign n31839 = n31833 & ~n31838;
  assign n31840 = ~pi0246 & ~n31831;
  assign n31841 = ~n31832 & ~n31840;
  assign n31842 = n31833 & n31841;
  assign n31843 = ~pi0223 & n31832;
  assign n31844 = n31838 & ~n31841;
  assign n31845 = n31843 & ~n31844;
  assign n31846 = ~n31842 & ~n31845;
  assign n31847 = ~n31839 & n31846;
  assign n31848 = pi3641 & ~n31847;
  assign n31849 = ~n31833 & ~n31843;
  assign n31850 = pi3641 & n31844;
  assign n31851 = n31849 & n31850;
  assign n31852 = ~n31848 & ~n31851;
  assign n31853 = pi0223 & ~pi3641;
  assign n31854 = n31852 & ~n31853;
  assign n31855 = ~n31777 & ~n31854;
  assign n31856 = ~pi0827 & ~pi3681;
  assign n31857 = pi0691 & pi1370;
  assign n31858 = pi1605 & pi1681;
  assign n31859 = pi1704 & n31858;
  assign n31860 = pi1606 & n31859;
  assign n31861 = pi0620 & n31860;
  assign n31862 = pi0619 & n31861;
  assign n31863 = n31857 & n31862;
  assign n31864 = ~pi3681 & ~n31863;
  assign n31865 = ~n31856 & ~n31864;
  assign n31866 = n31855 & n31865;
  assign n31867 = pi0223 & ~n31865;
  assign n31868 = ~n31777 & n31867;
  assign n31869 = ~n31866 & ~n31868;
  assign n31870 = ~n31779 & ~n31869;
  assign po0495 = ~n31783 | n31870;
  assign n31872 = ~pi0622 & n31013;
  assign n31873 = ~n31016 & ~n31872;
  assign n31874 = ~pi0224 & n31016;
  assign n31875 = ~n31873 & ~n31874;
  assign n31876 = ~n15426 & n31350;
  assign n31877 = n31276 & n31281;
  assign n31878 = n31256 & n31322;
  assign n31879 = n31877 & n31878;
  assign n31880 = n31270 & n31879;
  assign n31881 = ~n31243 & ~n31880;
  assign n31882 = n31243 & n31880;
  assign n31883 = ~n31881 & ~n31882;
  assign n31884 = ~pi0247 & n31883;
  assign n31885 = pi0247 & ~n31243;
  assign n31886 = ~n31884 & ~n31885;
  assign n31887 = pi0955 & ~pi2599;
  assign n31888 = ~n31886 & n31887;
  assign n31889 = ~pi0955 & ~pi2599;
  assign n31890 = pi0224 & n31889;
  assign n31891 = ~n31888 & ~n31890;
  assign n31892 = ~n31013 & ~n31891;
  assign n31893 = ~n31876 & ~n31892;
  assign n31894 = ~n31016 & ~n31893;
  assign po0496 = n31875 | n31894;
  assign n31896 = ~pi0621 & n31013;
  assign n31897 = ~n31016 & ~n31896;
  assign n31898 = ~pi0225 & n31016;
  assign n31899 = ~n31897 & ~n31898;
  assign n31900 = ~n14403 & n31350;
  assign n31901 = n31286 & n31877;
  assign n31902 = n31321 & n31901;
  assign n31903 = n31270 & n31902;
  assign n31904 = n31256 & n31903;
  assign n31905 = ~n31256 & ~n31903;
  assign n31906 = ~n31904 & ~n31905;
  assign n31907 = ~pi0247 & n31906;
  assign n31908 = pi0247 & ~n31256;
  assign n31909 = ~n31907 & ~n31908;
  assign n31910 = n31887 & ~n31909;
  assign n31911 = pi0225 & n31889;
  assign n31912 = ~n31910 & ~n31911;
  assign n31913 = ~n31013 & ~n31912;
  assign n31914 = ~n31900 & ~n31913;
  assign n31915 = ~n31016 & ~n31914;
  assign po0497 = n31899 | n31915;
  assign n31917 = pi0709 & ~n25999;
  assign n31918 = ~pi0709 & ~n29860;
  assign n31919 = ~n31917 & ~n31918;
  assign n31920 = ~n30955 & ~n31919;
  assign n31921 = pi0226 & n30955;
  assign po0498 = n31920 | n31921;
  assign n31923 = ~n30966 & ~n31919;
  assign n31924 = pi0227 & n30966;
  assign po0499 = n31923 | n31924;
  assign n31926 = ~n27687 & n31382;
  assign n31927 = pi0228 & n31381;
  assign n31928 = n30321 & n31384;
  assign n31929 = ~pi0228 & ~n31384;
  assign n31930 = ~n31928 & ~n31929;
  assign n31931 = n31388 & n31930;
  assign n31932 = ~n31927 & ~n31931;
  assign n31933 = ~n31391 & n31932;
  assign n31934 = ~n31382 & ~n31933;
  assign po0500 = n31926 | n31934;
  assign n31936 = ~n27687 & n31400;
  assign n31937 = pi0229 & n31399;
  assign n31938 = n30321 & n31402;
  assign n31939 = ~pi0229 & ~n31402;
  assign n31940 = ~n31938 & ~n31939;
  assign n31941 = n31406 & n31940;
  assign n31942 = ~n31937 & ~n31941;
  assign n31943 = ~n31409 & n31942;
  assign n31944 = ~n31400 & ~n31943;
  assign po0501 = n31936 | n31944;
  assign n31946 = pi1953 & n19569;
  assign n31947 = n20522 & ~n31946;
  assign n31948 = pi0979 & n31947;
  assign n31949 = ~pi0230 & ~n31948;
  assign n31950 = n20387 & ~n30537;
  assign n31951 = ~n28969 & n30537;
  assign n31952 = ~n31950 & ~n31951;
  assign n31953 = n31948 & ~n31952;
  assign po0502 = n31949 | n31953;
  assign n31955 = ~pi0979 & n31947;
  assign n31956 = ~pi0231 & ~n31955;
  assign n31957 = ~n31952 & n31955;
  assign po0503 = n31956 | n31957;
  assign n31959 = ~pi0631 & n31013;
  assign n31960 = ~n31016 & ~n31959;
  assign n31961 = ~pi0232 & n31016;
  assign n31962 = ~n31960 & ~n31961;
  assign n31963 = ~n13701 & n31350;
  assign n31964 = pi0247 & ~n31276;
  assign n31965 = ~n31276 & ~n31323;
  assign n31966 = ~n31324 & ~n31965;
  assign n31967 = ~pi0247 & n31966;
  assign n31968 = ~n31964 & ~n31967;
  assign n31969 = n31887 & ~n31968;
  assign n31970 = pi0232 & n31889;
  assign n31971 = ~n31969 & ~n31970;
  assign n31972 = ~n31013 & ~n31971;
  assign n31973 = ~n31963 & ~n31972;
  assign n31974 = ~n31016 & ~n31973;
  assign po0504 = n31962 | n31974;
  assign n31976 = ~pi0709 & ~n29607;
  assign n31977 = pi0709 & ~n27570;
  assign n31978 = ~n31976 & ~n31977;
  assign n31979 = ~n30955 & ~n31978;
  assign n31980 = pi0233 & n30955;
  assign po0505 = n31979 | n31980;
  assign n31982 = ~n30966 & ~n31978;
  assign n31983 = pi0234 & n30966;
  assign po0506 = n31982 | n31983;
  assign n31985 = pi0710 & n26050;
  assign n31986 = ~n30954 & ~n31985;
  assign n31987 = ~pi0710 & ~n27915;
  assign n31988 = pi0710 & ~n30288;
  assign n31989 = ~n31987 & ~n31988;
  assign n31990 = ~n31986 & ~n31989;
  assign n31991 = pi0235 & n31986;
  assign po0507 = n31990 | n31991;
  assign n31993 = pi0710 & n20522;
  assign n31994 = ~pi0979 & n31993;
  assign n31995 = ~n30965 & ~n31994;
  assign n31996 = ~n31989 & ~n31995;
  assign n31997 = pi0236 & n31995;
  assign po0508 = n31996 | n31997;
  assign n31999 = ~pi0608 & n31013;
  assign n32000 = ~n31016 & ~n31999;
  assign n32001 = ~pi0237 & n31016;
  assign n32002 = ~n32000 & ~n32001;
  assign n32003 = ~n12726 & n31350;
  assign n32004 = n31313 & n31320;
  assign n32005 = n31298 & n32004;
  assign n32006 = n31877 & n32005;
  assign n32007 = n31293 & n32006;
  assign n32008 = n31286 & n32007;
  assign n32009 = ~n31270 & ~n32008;
  assign n32010 = n31270 & n32008;
  assign n32011 = ~n32009 & ~n32010;
  assign n32012 = ~pi0247 & n32011;
  assign n32013 = pi0247 & ~n31270;
  assign n32014 = ~n32012 & ~n32013;
  assign n32015 = n31887 & ~n32014;
  assign n32016 = pi0237 & n31889;
  assign n32017 = ~n32015 & ~n32016;
  assign n32018 = ~n31013 & ~n32017;
  assign n32019 = ~n32003 & ~n32018;
  assign n32020 = ~n31016 & ~n32019;
  assign po0509 = n32002 | n32020;
  assign n32022 = ~pi0709 & ~n28006;
  assign n32023 = pi0709 & ~n30288;
  assign n32024 = ~n32022 & ~n32023;
  assign n32025 = ~n30955 & ~n32024;
  assign n32026 = pi0238 & n30955;
  assign po0510 = n32025 | n32026;
  assign n32028 = ~n30966 & ~n32024;
  assign n32029 = pi0239 & n30966;
  assign po0511 = n32028 | n32029;
  assign n32031 = ~n27690 & n31382;
  assign n32032 = pi0240 & n31381;
  assign n32033 = n30333 & n31384;
  assign n32034 = ~pi0240 & ~n31384;
  assign n32035 = ~n32033 & ~n32034;
  assign n32036 = n31388 & n32035;
  assign n32037 = ~n32032 & ~n32036;
  assign n32038 = ~n31391 & n32037;
  assign n32039 = ~n31382 & ~n32038;
  assign po0512 = n32031 | n32039;
  assign n32041 = ~n27690 & n31400;
  assign n32042 = pi0241 & n31399;
  assign n32043 = n30333 & n31402;
  assign n32044 = ~pi0241 & ~n31402;
  assign n32045 = ~n32043 & ~n32044;
  assign n32046 = n31406 & n32045;
  assign n32047 = ~n32042 & ~n32046;
  assign n32048 = ~n31409 & n32047;
  assign n32049 = ~n31400 & ~n32048;
  assign po0513 = n32041 | n32049;
  assign n32051 = ~n28969 & ~n30537;
  assign n32052 = n29216 & n30537;
  assign n32053 = ~n32051 & ~n32052;
  assign n32054 = n31948 & ~n32053;
  assign n32055 = ~pi0242 & ~n31948;
  assign po0514 = n32054 | n32055;
  assign n32057 = ~pi0243 & ~n31948;
  assign n32058 = n29216 & ~n30537;
  assign n32059 = ~n29458 & n30537;
  assign n32060 = ~n32058 & ~n32059;
  assign n32061 = n31948 & ~n32060;
  assign po0515 = n32057 | n32061;
  assign n32063 = n31955 & ~n32053;
  assign n32064 = ~pi0244 & ~n31955;
  assign po0516 = n32063 | n32064;
  assign n32066 = ~pi0245 & ~n31955;
  assign n32067 = n31955 & ~n32060;
  assign po0517 = n32066 | n32067;
  assign n32069 = ~n31838 & n31841;
  assign n32070 = ~n31844 & ~n32069;
  assign n32071 = n31865 & ~n32070;
  assign n32072 = pi3641 & n32071;
  assign n32073 = pi3641 & n31865;
  assign n32074 = pi0246 & ~n32073;
  assign n32075 = ~n32072 & ~n32074;
  assign n32076 = ~n31777 & ~n32075;
  assign n32077 = pi1723 & n31777;
  assign n32078 = ~n32076 & ~n32077;
  assign n32079 = ~n31779 & ~n32078;
  assign n32080 = ~pi2394 & n31779;
  assign po0518 = n32079 | n32080;
  assign n32082 = ~pi0630 & n31013;
  assign n32083 = ~n31016 & ~n32082;
  assign n32084 = ~pi0247 & n31016;
  assign n32085 = ~n32083 & ~n32084;
  assign n32086 = pi0247 & ~n31281;
  assign n32087 = ~n31281 & ~n31322;
  assign n32088 = ~n31323 & ~n32087;
  assign n32089 = ~pi0247 & n32088;
  assign n32090 = ~n32086 & ~n32089;
  assign n32091 = n31887 & ~n32090;
  assign n32092 = pi0247 & n31889;
  assign n32093 = ~n32091 & ~n32092;
  assign n32094 = ~n31013 & ~n32093;
  assign n32095 = ~n13121 & n31350;
  assign n32096 = ~n32094 & ~n32095;
  assign n32097 = ~n31016 & ~n32096;
  assign po0519 = n32085 | n32097;
  assign n32099 = ~pi0629 & n31013;
  assign n32100 = ~n31016 & ~n32099;
  assign n32101 = ~pi0248 & n31016;
  assign n32102 = ~n32100 & ~n32101;
  assign n32103 = ~n13398 & n31350;
  assign n32104 = pi0247 & ~n31286;
  assign n32105 = ~n31286 & ~n31321;
  assign n32106 = ~n31322 & ~n32105;
  assign n32107 = ~pi0247 & n32106;
  assign n32108 = ~n32104 & ~n32107;
  assign n32109 = n31887 & ~n32108;
  assign n32110 = pi0248 & n31889;
  assign n32111 = ~n32109 & ~n32110;
  assign n32112 = ~n31013 & ~n32111;
  assign n32113 = ~n32103 & ~n32112;
  assign n32114 = ~n31016 & ~n32113;
  assign po0520 = n32102 | n32114;
  assign n32116 = pi0710 & ~n30267;
  assign n32117 = ~pi0710 & ~n28609;
  assign n32118 = ~n32116 & ~n32117;
  assign n32119 = ~n31986 & ~n32118;
  assign n32120 = pi0249 & n31986;
  assign po0521 = n32119 | n32120;
  assign n32122 = ~pi0710 & ~n28122;
  assign n32123 = pi0710 & ~n24744;
  assign n32124 = ~n32122 & ~n32123;
  assign n32125 = ~n31986 & ~n32124;
  assign n32126 = pi0250 & n31986;
  assign po0522 = n32125 | n32126;
  assign n32128 = ~pi0710 & ~n27425;
  assign n32129 = pi0710 & ~n24265;
  assign n32130 = ~n32128 & ~n32129;
  assign n32131 = ~n31986 & ~n32130;
  assign n32132 = pi0251 & n31986;
  assign po0523 = n32131 | n32132;
  assign n32134 = ~n31995 & ~n32118;
  assign n32135 = pi0252 & n31995;
  assign po0524 = n32134 | n32135;
  assign n32137 = ~n31995 & ~n32124;
  assign n32138 = pi0253 & n31995;
  assign po0525 = n32137 | n32138;
  assign n32140 = ~n31995 & ~n32130;
  assign n32141 = pi0254 & n31995;
  assign po0526 = n32140 | n32141;
  assign n32143 = ~n27624 & n31382;
  assign n32144 = pi0255 & n31381;
  assign n32145 = n27570 & n31384;
  assign n32146 = ~pi0255 & ~n31384;
  assign n32147 = ~n32145 & ~n32146;
  assign n32148 = n31388 & n32147;
  assign n32149 = ~n32144 & ~n32148;
  assign n32150 = ~n31391 & n32149;
  assign n32151 = ~n31382 & ~n32150;
  assign po0527 = n32143 | n32151;
  assign n32153 = ~n27635 & n31382;
  assign n32154 = pi0256 & n31381;
  assign n32155 = n25999 & n31384;
  assign n32156 = ~pi0256 & ~n31384;
  assign n32157 = ~n32155 & ~n32156;
  assign n32158 = n31388 & n32157;
  assign n32159 = ~n32154 & ~n32158;
  assign n32160 = ~n31391 & n32159;
  assign n32161 = ~n31382 & ~n32160;
  assign po0528 = n32153 | n32161;
  assign n32163 = ~n27624 & n31400;
  assign n32164 = pi0257 & n31399;
  assign n32165 = n27570 & n31402;
  assign n32166 = ~pi0257 & ~n31402;
  assign n32167 = ~n32165 & ~n32166;
  assign n32168 = n31406 & n32167;
  assign n32169 = ~n32164 & ~n32168;
  assign n32170 = ~n31409 & n32169;
  assign n32171 = ~n31400 & ~n32170;
  assign po0529 = n32163 | n32171;
  assign n32173 = ~n27635 & n31400;
  assign n32174 = pi0258 & n31399;
  assign n32175 = n25999 & n31402;
  assign n32176 = ~pi0258 & ~n31402;
  assign n32177 = ~n32175 & ~n32176;
  assign n32178 = n31406 & n32177;
  assign n32179 = ~n32174 & ~n32178;
  assign n32180 = ~n31409 & n32179;
  assign n32181 = ~n31400 & ~n32180;
  assign po0530 = n32173 | n32181;
  assign n32183 = ~pi0709 & ~n26794;
  assign n32184 = pi0709 & ~n25699;
  assign n32185 = ~n32183 & ~n32184;
  assign n32186 = ~n30955 & ~n32185;
  assign n32187 = pi0259 & n30955;
  assign po0531 = n32186 | n32187;
  assign n32189 = ~pi0709 & ~n26550;
  assign n32190 = pi0709 & ~n24769;
  assign n32191 = ~n32189 & ~n32190;
  assign n32192 = ~n30955 & ~n32191;
  assign n32193 = pi0260 & n30955;
  assign po0532 = n32192 | n32193;
  assign n32195 = ~pi0709 & ~n29190;
  assign n32196 = pi0709 & ~n30321;
  assign n32197 = ~n32195 & ~n32196;
  assign n32198 = ~n30955 & ~n32197;
  assign n32199 = pi0261 & n30955;
  assign po0533 = n32198 | n32199;
  assign n32201 = pi0709 & ~n24488;
  assign n32202 = ~pi0709 & ~n30143;
  assign n32203 = ~n32201 & ~n32202;
  assign n32204 = ~n30955 & ~n32203;
  assign n32205 = pi0262 & n30955;
  assign po0534 = n32204 | n32205;
  assign n32207 = ~n30966 & ~n32185;
  assign n32208 = pi0263 & n30966;
  assign po0535 = n32207 | n32208;
  assign n32210 = ~n30966 & ~n32191;
  assign n32211 = pi0264 & n30966;
  assign po0536 = n32210 | n32211;
  assign n32213 = ~n30966 & ~n32197;
  assign n32214 = pi0265 & n30966;
  assign po0537 = n32213 | n32214;
  assign n32216 = ~n30966 & ~n32203;
  assign n32217 = pi0266 & n30966;
  assign po0538 = n32216 | n32217;
  assign n32219 = ~n27647 & n31382;
  assign n32220 = pi0267 & n31381;
  assign n32221 = n30267 & n31384;
  assign n32222 = ~pi0267 & ~n31384;
  assign n32223 = ~n32221 & ~n32222;
  assign n32224 = n31388 & n32223;
  assign n32225 = ~n32220 & ~n32224;
  assign n32226 = ~n31391 & n32225;
  assign n32227 = ~n31382 & ~n32226;
  assign po0539 = n32219 | n32227;
  assign n32229 = ~n27647 & n31400;
  assign n32230 = pi0268 & n31399;
  assign n32231 = n30267 & n31402;
  assign n32232 = ~pi0268 & ~n31402;
  assign n32233 = ~n32231 & ~n32232;
  assign n32234 = n31406 & n32233;
  assign n32235 = ~n32230 & ~n32234;
  assign n32236 = ~n31409 & n32235;
  assign n32237 = ~n31400 & ~n32236;
  assign po0540 = n32229 | n32237;
  assign n32239 = ~pi0709 & ~n27043;
  assign n32240 = pi0709 & ~n25718;
  assign n32241 = ~n32239 & ~n32240;
  assign n32242 = ~n30955 & ~n32241;
  assign n32243 = pi0269 & n30955;
  assign po0541 = n32242 | n32243;
  assign n32245 = ~n30966 & ~n32241;
  assign n32246 = pi0270 & n30966;
  assign po0542 = n32245 | n32246;
  assign n32248 = pi0710 & ~n30333;
  assign n32249 = ~pi0710 & ~n29437;
  assign n32250 = ~n32248 & ~n32249;
  assign n32251 = ~n31986 & ~n32250;
  assign n32252 = pi0271 & n31986;
  assign po0543 = n32251 | n32252;
  assign n32254 = ~n31995 & ~n32250;
  assign n32255 = pi0272 & n31995;
  assign po0544 = n32254 | n32255;
  assign n32257 = ~n29458 & ~n30537;
  assign n32258 = n29708 & n30537;
  assign n32259 = ~n32257 & ~n32258;
  assign n32260 = n31948 & ~n32259;
  assign n32261 = ~pi0273 & ~n31948;
  assign po0545 = n32260 | n32261;
  assign n32263 = ~pi0274 & ~n31948;
  assign n32264 = n29708 & ~n30537;
  assign n32265 = n29959 & n30537;
  assign n32266 = ~n32264 & ~n32265;
  assign n32267 = n31948 & ~n32266;
  assign po0546 = n32263 | n32267;
  assign n32269 = n31955 & ~n32259;
  assign n32270 = ~pi0275 & ~n31955;
  assign po0547 = n32269 | n32270;
  assign n32272 = ~pi0276 & ~n31955;
  assign n32273 = n31955 & ~n32266;
  assign po0548 = n32272 | n32273;
  assign n32275 = n31835 & n31837;
  assign n32276 = ~n31838 & ~n32275;
  assign n32277 = n31865 & ~n32276;
  assign n32278 = pi3641 & n32277;
  assign n32279 = pi0277 & ~n32073;
  assign n32280 = ~n32278 & ~n32279;
  assign n32281 = ~n31777 & ~n32280;
  assign n32282 = pi1879 & n31777;
  assign n32283 = ~n32281 & ~n32282;
  assign n32284 = ~n31779 & ~n32283;
  assign n32285 = ~pi2097 & n31779;
  assign po0549 = n32284 | n32285;
  assign n32287 = ~pi0611 & n31013;
  assign n32288 = ~n31016 & ~n32287;
  assign n32289 = ~pi0278 & n31016;
  assign n32290 = ~n32288 & ~n32289;
  assign n32291 = ~n13988 & n31350;
  assign n32292 = ~n31293 & n32005;
  assign n32293 = n31293 & ~n32005;
  assign n32294 = ~n32292 & ~n32293;
  assign n32295 = ~pi0247 & ~n32294;
  assign n32296 = pi0247 & ~n31293;
  assign n32297 = ~n32295 & ~n32296;
  assign n32298 = n31887 & ~n32297;
  assign n32299 = pi0278 & n31889;
  assign n32300 = ~n32298 & ~n32299;
  assign n32301 = ~n31013 & ~n32300;
  assign n32302 = ~n32291 & ~n32301;
  assign n32303 = ~n31016 & ~n32302;
  assign po0550 = n32290 | n32303;
  assign n32305 = ~pi0709 & ~n28209;
  assign n32306 = pi0709 & ~n24744;
  assign n32307 = ~n32305 & ~n32306;
  assign n32308 = ~n30955 & ~n32307;
  assign n32309 = pi0279 & n30955;
  assign po0551 = n32308 | n32309;
  assign n32311 = ~n30966 & ~n32307;
  assign n32312 = pi0280 & n30966;
  assign po0552 = n32311 | n32312;
  assign n32314 = ~pi0710 & ~n29683;
  assign n32315 = pi0710 & ~n27570;
  assign n32316 = ~n32314 & ~n32315;
  assign n32317 = ~n31986 & ~n32316;
  assign n32318 = pi0281 & n31986;
  assign po0553 = n32317 | n32318;
  assign n32320 = pi0710 & ~n25999;
  assign n32321 = ~pi0710 & ~n29936;
  assign n32322 = ~n32320 & ~n32321;
  assign n32323 = ~n31986 & ~n32322;
  assign n32324 = pi0282 & n31986;
  assign po0554 = n32323 | n32324;
  assign n32326 = ~n31995 & ~n32316;
  assign n32327 = pi0283 & n31995;
  assign po0555 = n32326 | n32327;
  assign n32329 = ~n31995 & ~n32322;
  assign n32330 = pi0284 & n31995;
  assign po0556 = n32329 | n32330;
  assign n32332 = ~pi0709 & ~n27343;
  assign n32333 = pi0709 & ~n24265;
  assign n32334 = ~n32332 & ~n32333;
  assign n32335 = ~n30955 & ~n32334;
  assign n32336 = pi0285 & n30955;
  assign po0557 = n32335 | n32336;
  assign n32338 = ~n30966 & ~n32334;
  assign n32339 = pi0286 & n30966;
  assign po0558 = n32338 | n32339;
  assign n32341 = ~pi0710 & ~n26625;
  assign n32342 = pi0710 & ~n24769;
  assign n32343 = ~n32341 & ~n32342;
  assign n32344 = ~n31986 & ~n32343;
  assign n32345 = pi0287 & n31986;
  assign po0559 = n32344 | n32345;
  assign n32347 = ~pi0710 & ~n26863;
  assign n32348 = pi0710 & ~n25699;
  assign n32349 = ~n32347 & ~n32348;
  assign n32350 = ~n31986 & ~n32349;
  assign n32351 = pi0288 & n31986;
  assign po0560 = n32350 | n32351;
  assign n32353 = ~pi0710 & ~n25858;
  assign n32354 = pi0710 & ~n24446;
  assign n32355 = ~n32353 & ~n32354;
  assign n32356 = ~n31986 & ~n32355;
  assign n32357 = pi0289 & n31986;
  assign po0561 = n32356 | n32357;
  assign n32359 = ~n31995 & ~n32343;
  assign n32360 = pi0290 & n31995;
  assign po0562 = n32359 | n32360;
  assign n32362 = ~n31995 & ~n32349;
  assign n32363 = pi0291 & n31995;
  assign po0563 = n32362 | n32363;
  assign n32365 = ~n31995 & ~n32355;
  assign n32366 = pi0292 & n31995;
  assign po0564 = n32365 | n32366;
  assign n32368 = ~n27654 & n31382;
  assign n32369 = pi0293 & n31381;
  assign n32370 = n30288 & n31384;
  assign n32371 = ~pi0293 & ~n31384;
  assign n32372 = ~n32370 & ~n32371;
  assign n32373 = n31388 & n32372;
  assign n32374 = ~n32369 & ~n32373;
  assign n32375 = ~n31391 & n32374;
  assign n32376 = ~n31382 & ~n32375;
  assign po0565 = n32368 | n32376;
  assign n32378 = ~n27654 & n31400;
  assign n32379 = pi0294 & n31399;
  assign n32380 = n30288 & n31402;
  assign n32381 = ~pi0294 & ~n31402;
  assign n32382 = ~n32380 & ~n32381;
  assign n32383 = n31406 & n32382;
  assign n32384 = ~n32379 & ~n32383;
  assign n32385 = ~n31409 & n32384;
  assign n32386 = ~n31400 & ~n32385;
  assign po0566 = n32378 | n32386;
  assign n32388 = ~pi0295 & ~n31948;
  assign n32389 = n29959 & ~n30537;
  assign n32390 = ~n28725 & n30537;
  assign n32391 = ~n32389 & ~n32390;
  assign n32392 = n31948 & ~n32391;
  assign po0567 = n32388 | n32392;
  assign n32394 = ~pi0296 & ~n31955;
  assign n32395 = n31955 & ~n32391;
  assign po0568 = n32394 | n32395;
  assign n32397 = ~pi0709 & ~n28948;
  assign n32398 = pi0709 & ~n30309;
  assign n32399 = ~n32397 & ~n32398;
  assign n32400 = ~n30955 & ~n32399;
  assign n32401 = pi0297 & n30955;
  assign po0569 = n32400 | n32401;
  assign n32403 = ~n30966 & ~n32399;
  assign n32404 = pi0298 & n30966;
  assign po0570 = n32403 | n32404;
  assign n32406 = ~pi0710 & ~n25441;
  assign n32407 = pi0710 & ~n24289;
  assign n32408 = ~n32406 & ~n32407;
  assign n32409 = ~n31986 & ~n32408;
  assign n32410 = pi0299 & n31986;
  assign po0571 = n32409 | n32410;
  assign n32412 = ~n31995 & ~n32408;
  assign n32413 = pi0300 & n31995;
  assign po0572 = n32412 | n32413;
  assign n32415 = ~n28725 & ~n30537;
  assign n32416 = n27813 & n30537;
  assign n32417 = ~n32415 & ~n32416;
  assign n32418 = n31948 & ~n32417;
  assign n32419 = ~pi0301 & ~n31948;
  assign po0573 = n32418 | n32419;
  assign n32421 = n31955 & ~n32417;
  assign n32422 = ~pi0302 & ~n31955;
  assign po0574 = n32421 | n32422;
  assign n32424 = pi3641 & ~n31837;
  assign n32425 = pi0303 & ~pi3641;
  assign n32426 = ~n32424 & ~n32425;
  assign n32427 = n31865 & ~n32426;
  assign n32428 = pi0303 & ~n31865;
  assign n32429 = ~n32427 & ~n32428;
  assign n32430 = ~n31777 & ~n32429;
  assign n32431 = pi1880 & n31777;
  assign n32432 = ~n32430 & ~n32431;
  assign n32433 = ~n31779 & ~n32432;
  assign n32434 = ~pi2096 & n31779;
  assign po0575 = n32433 | n32434;
  assign n32436 = ~pi0709 & ~n28426;
  assign n32437 = pi0709 & ~n24256;
  assign n32438 = ~n32436 & ~n32437;
  assign n32439 = ~n30955 & ~n32438;
  assign n32440 = pi0304 & n30955;
  assign po0576 = n32439 | n32440;
  assign n32442 = ~pi0709 & ~n25936;
  assign n32443 = pi0709 & ~n24446;
  assign n32444 = ~n32442 & ~n32443;
  assign n32445 = ~n30955 & ~n32444;
  assign n32446 = pi0305 & n30955;
  assign po0577 = n32445 | n32446;
  assign n32448 = ~n30966 & ~n32438;
  assign n32449 = pi0306 & n30966;
  assign po0578 = n32448 | n32449;
  assign n32451 = ~n30966 & ~n32444;
  assign n32452 = pi0307 & n30966;
  assign po0579 = n32451 | n32452;
  assign n32454 = ~pi0710 & ~n29101;
  assign n32455 = pi0710 & ~n30321;
  assign n32456 = ~n32454 & ~n32455;
  assign n32457 = ~n31986 & ~n32456;
  assign n32458 = pi0308 & n31986;
  assign po0580 = n32457 | n32458;
  assign n32460 = ~pi0710 & ~n30212;
  assign n32461 = pi0710 & ~n24488;
  assign n32462 = ~n32460 & ~n32461;
  assign n32463 = ~n31986 & ~n32462;
  assign n32464 = pi0309 & n31986;
  assign po0581 = n32463 | n32464;
  assign n32466 = ~n31995 & ~n32456;
  assign n32467 = pi0310 & n31995;
  assign po0582 = n32466 | n32467;
  assign n32469 = ~n31995 & ~n32462;
  assign n32470 = pi0311 & n31995;
  assign po0583 = n32469 | n32470;
  assign n32472 = ~n27729 & n31382;
  assign n32473 = pi0312 & n31381;
  assign n32474 = ~n24744 & n31384;
  assign n32475 = pi0312 & ~n31384;
  assign n32476 = ~n32474 & ~n32475;
  assign n32477 = n31388 & ~n32476;
  assign n32478 = ~n32473 & ~n32477;
  assign n32479 = ~n31391 & n32478;
  assign n32480 = ~n31382 & ~n32479;
  assign po0584 = n32472 | n32480;
  assign n32482 = ~n27729 & n31400;
  assign n32483 = pi0313 & n31399;
  assign n32484 = ~n24744 & n31402;
  assign n32485 = pi0313 & ~n31402;
  assign n32486 = ~n32484 & ~n32485;
  assign n32487 = n31406 & ~n32486;
  assign n32488 = ~n32483 & ~n32487;
  assign n32489 = ~n31409 & n32488;
  assign n32490 = ~n31400 & ~n32489;
  assign po0585 = n32482 | n32490;
  assign n32492 = pi1017 & n26322;
  assign n32493 = ~pi1017 & ~n26322;
  assign n32494 = ~n32492 & ~n32493;
  assign n32495 = pi2555 & ~n32494;
  assign n32496 = ~pi2555 & ~n13988;
  assign n32497 = ~n32495 & ~n32496;
  assign n32498 = ~n26062 & ~n32497;
  assign n32499 = pi0314 & n26062;
  assign po0586 = n32498 | n32499;
  assign n32501 = ~pi0709 & ~n25367;
  assign n32502 = pi0709 & ~n24289;
  assign n32503 = ~n32501 & ~n32502;
  assign n32504 = ~n30955 & ~n32503;
  assign n32505 = pi0315 & n30955;
  assign po0587 = n32504 | n32505;
  assign n32507 = ~n30966 & ~n32503;
  assign n32508 = pi0316 & n30966;
  assign po0588 = n32507 | n32508;
  assign n32510 = ~pi0710 & ~n27110;
  assign n32511 = pi0710 & ~n25718;
  assign n32512 = ~n32510 & ~n32511;
  assign n32513 = ~n31986 & ~n32512;
  assign n32514 = pi0317 & n31986;
  assign po0589 = n32513 | n32514;
  assign n32516 = ~pi0710 & ~n28861;
  assign n32517 = pi0710 & ~n30309;
  assign n32518 = ~n32516 & ~n32517;
  assign n32519 = ~n31986 & ~n32518;
  assign n32520 = pi0318 & n31986;
  assign po0590 = n32519 | n32520;
  assign n32522 = ~n31995 & ~n32512;
  assign n32523 = pi0319 & n31995;
  assign po0591 = n32522 | n32523;
  assign n32525 = ~n31995 & ~n32518;
  assign n32526 = pi0320 & n31995;
  assign po0592 = n32525 | n32526;
  assign n32528 = ~pi0321 & ~n31948;
  assign n32529 = n27813 & ~n30537;
  assign n32530 = n28234 & n30537;
  assign n32531 = ~n32529 & ~n32530;
  assign n32532 = n31948 & ~n32531;
  assign po0593 = n32528 | n32532;
  assign n32534 = ~pi0322 & ~n31955;
  assign n32535 = n31955 & ~n32531;
  assign po0594 = n32534 | n32535;
  assign n32537 = ~pi0710 & ~n28497;
  assign n32538 = pi0710 & ~n24256;
  assign n32539 = ~n32537 & ~n32538;
  assign n32540 = ~n31986 & ~n32539;
  assign n32541 = pi0323 & n31986;
  assign po0595 = n32540 | n32541;
  assign n32543 = ~n31995 & ~n32539;
  assign n32544 = pi0324 & n31995;
  assign po0596 = n32543 | n32544;
  assign n32546 = ~pi0325 & ~n31948;
  assign n32547 = n28234 & ~n30537;
  assign n32548 = ~n26654 & n30537;
  assign n32549 = ~n32547 & ~n32548;
  assign n32550 = n31948 & ~n32549;
  assign po0597 = n32546 | n32550;
  assign n32552 = ~pi0326 & ~n31955;
  assign n32553 = n31955 & ~n32549;
  assign po0598 = n32552 | n32553;
  assign n32555 = ~n27738 & n31382;
  assign n32556 = pi0327 & n31381;
  assign n32557 = ~n24769 & n31384;
  assign n32558 = pi0327 & ~n31384;
  assign n32559 = ~n32557 & ~n32558;
  assign n32560 = n31388 & ~n32559;
  assign n32561 = ~n32556 & ~n32560;
  assign n32562 = ~n31391 & n32561;
  assign n32563 = ~n31382 & ~n32562;
  assign po0599 = n32555 | n32563;
  assign n32565 = ~n27738 & n31400;
  assign n32566 = pi0328 & n31399;
  assign n32567 = ~n24769 & n31402;
  assign n32568 = pi0328 & ~n31402;
  assign n32569 = ~n32567 & ~n32568;
  assign n32570 = n31406 & ~n32569;
  assign n32571 = ~n32566 & ~n32570;
  assign n32572 = ~n31409 & n32571;
  assign n32573 = ~n31400 & ~n32572;
  assign po0600 = n32565 | n32573;
  assign n32575 = ~pi0628 & n31013;
  assign n32576 = ~n31016 & ~n32575;
  assign n32577 = ~pi0329 & n31016;
  assign n32578 = ~n32576 & ~n32577;
  assign n32579 = pi0247 & ~n31320;
  assign n32580 = n31314 & n31320;
  assign n32581 = ~n31314 & ~n31320;
  assign n32582 = ~n32580 & ~n32581;
  assign n32583 = ~pi0247 & n32582;
  assign n32584 = ~n32579 & ~n32583;
  assign n32585 = n31887 & ~n32584;
  assign n32586 = pi0329 & n31889;
  assign n32587 = ~n32585 & ~n32586;
  assign n32588 = ~n31013 & ~n32587;
  assign n32589 = ~n12415 & n31350;
  assign n32590 = ~n32588 & ~n32589;
  assign n32591 = ~n31016 & ~n32590;
  assign po0601 = n32578 | n32591;
  assign n32593 = pi2555 & ~n26332;
  assign n32594 = ~pi2555 & ~n12415;
  assign n32595 = ~n32593 & ~n32594;
  assign n32596 = ~n26062 & ~n32595;
  assign n32597 = pi0330 & n26062;
  assign po0602 = n32596 | n32597;
  assign n32599 = ~pi0627 & n31013;
  assign n32600 = ~n31016 & ~n32599;
  assign n32601 = ~pi0331 & n31016;
  assign n32602 = ~n32600 & ~n32601;
  assign n32603 = pi0247 & ~n31298;
  assign n32604 = ~n31298 & ~n31313;
  assign n32605 = ~n31314 & ~n32604;
  assign n32606 = ~pi0247 & n32605;
  assign n32607 = ~n32603 & ~n32606;
  assign n32608 = n31887 & ~n32607;
  assign n32609 = pi0331 & n31889;
  assign n32610 = ~n32608 & ~n32609;
  assign n32611 = ~n31013 & ~n32610;
  assign n32612 = ~n14816 & n31350;
  assign n32613 = ~n32611 & ~n32612;
  assign n32614 = ~n31016 & ~n32613;
  assign po0603 = n32602 | n32614;
  assign n32616 = ~n9530 & ~n13284;
  assign n32617 = ~n12208 & n32616;
  assign n32618 = ~n13781 & n32617;
  assign n32619 = n24995 & n32618;
  assign n32620 = n14623 & n15011;
  assign n32621 = n32619 & n32620;
  assign n32622 = n24928 & n32621;
  assign n32623 = ~pi2021 & n32622;
  assign n32624 = n19587 & n32623;
  assign n32625 = ~pi3518 & n31435;
  assign n32626 = ~n32624 & ~n32625;
  assign n32627 = pi0712 & n32626;
  assign n32628 = n26050 & ~n32627;
  assign n32629 = pi0712 & ~n31572;
  assign n32630 = ~pi0712 & ~n24488;
  assign n32631 = ~n32629 & ~n32630;
  assign n32632 = n32628 & ~n32631;
  assign n32633 = pi0332 & ~n32628;
  assign po0604 = n32632 | n32633;
  assign n32635 = n30791 & ~n32627;
  assign n32636 = ~n32631 & n32635;
  assign n32637 = pi0333 & ~n32635;
  assign po0605 = n32636 | n32637;
  assign n32639 = ~n27749 & n31382;
  assign n32640 = pi0334 & n31381;
  assign n32641 = ~n25699 & n31384;
  assign n32642 = pi0334 & ~n31384;
  assign n32643 = ~n32641 & ~n32642;
  assign n32644 = n31388 & ~n32643;
  assign n32645 = ~n32640 & ~n32644;
  assign n32646 = ~n31391 & n32645;
  assign n32647 = ~n31382 & ~n32646;
  assign po0606 = n32639 | n32647;
  assign n32649 = ~n27749 & n31400;
  assign n32650 = pi0335 & n31399;
  assign n32651 = ~n25699 & n31402;
  assign n32652 = pi0335 & ~n31402;
  assign n32653 = ~n32651 & ~n32652;
  assign n32654 = n31406 & ~n32653;
  assign n32655 = ~n32650 & ~n32654;
  assign n32656 = ~n31409 & n32655;
  assign n32657 = ~n31400 & ~n32656;
  assign po0607 = n32649 | n32657;
  assign n32659 = pi0336 & ~n31865;
  assign n32660 = n31816 & ~n31824;
  assign n32661 = ~n31825 & ~n32660;
  assign n32662 = pi3641 & ~n32661;
  assign n32663 = pi0336 & ~pi3641;
  assign n32664 = ~n32662 & ~n32663;
  assign n32665 = n31865 & ~n32664;
  assign n32666 = ~n32659 & ~n32665;
  assign n32667 = ~n31777 & ~n32666;
  assign n32668 = pi1724 & n31777;
  assign n32669 = ~n32667 & ~n32668;
  assign n32670 = ~n31779 & ~n32669;
  assign n32671 = ~pi1881 & n31779;
  assign po0608 = n32670 | n32671;
  assign n32673 = ~n26654 & ~n30537;
  assign n32674 = n26896 & n30537;
  assign n32675 = ~n32673 & ~n32674;
  assign n32676 = n31948 & ~n32675;
  assign n32677 = ~pi0337 & ~n31948;
  assign po0609 = n32676 | n32677;
  assign n32679 = ~pi0338 & ~n31948;
  assign n32680 = n26896 & ~n30537;
  assign n32681 = ~n27134 & n30537;
  assign n32682 = ~n32680 & ~n32681;
  assign n32683 = n31948 & ~n32682;
  assign po0610 = n32679 | n32683;
  assign n32685 = n31955 & ~n32675;
  assign n32686 = ~pi0339 & ~n31955;
  assign po0611 = n32685 | n32686;
  assign n32688 = ~pi0340 & ~n31955;
  assign n32689 = n31955 & ~n32682;
  assign po0612 = n32688 | n32689;
  assign n32691 = n20513 & n24870;
  assign n32692 = ~n24883 & ~n32691;
  assign n32693 = n24888 & ~n32692;
  assign n32694 = n25510 & n32693;
  assign n32695 = pi3245 & ~po3872;
  assign n32696 = n32693 & n32695;
  assign n32697 = ~po3872 & n20513;
  assign n32698 = n24874 & n24888;
  assign n32699 = n32697 & n32698;
  assign n32700 = n20519 & n32698;
  assign n32701 = n32695 & n32700;
  assign n32702 = n25510 & n32700;
  assign n32703 = ~n32701 & ~n32702;
  assign n32704 = ~n32699 & n32703;
  assign n32705 = ~n32696 & n32704;
  assign n32706 = n32694 & n32705;
  assign n32707 = ~n32694 & ~n32696;
  assign n32708 = ~n32699 & n32707;
  assign n32709 = ~n32701 & n32708;
  assign n32710 = ~n32702 & n32709;
  assign n32711 = n32702 & n32709;
  assign po0615 = n32710 | n32711;
  assign n32713 = n32699 & n32707;
  assign n32714 = n32703 & n32713;
  assign n32715 = n32701 & n32708;
  assign n32716 = ~n32702 & n32715;
  assign po0614 = n32714 | n32716;
  assign n32718 = ~po0615 & ~po0614;
  assign n32719 = ~n32694 & n32696;
  assign n32720 = n32704 & n32719;
  assign n32721 = n32718 & ~n32720;
  assign po0613 = n32706 | ~n32721;
  assign n32723 = ~n32706 & ~n32716;
  assign po0616 = n32710 | ~n32723;
  assign n32725 = ~n27752 & n31382;
  assign n32726 = pi0344 & n31381;
  assign n32727 = ~n25718 & n31384;
  assign n32728 = pi0344 & ~n31384;
  assign n32729 = ~n32727 & ~n32728;
  assign n32730 = n31388 & ~n32729;
  assign n32731 = ~n32726 & ~n32730;
  assign n32732 = ~n31391 & n32731;
  assign n32733 = ~n31382 & ~n32732;
  assign po0617 = n32725 | n32733;
  assign n32735 = ~n27752 & n31400;
  assign n32736 = pi0345 & n31399;
  assign n32737 = ~n25718 & n31402;
  assign n32738 = pi0345 & ~n31402;
  assign n32739 = ~n32737 & ~n32738;
  assign n32740 = n31406 & ~n32739;
  assign n32741 = ~n32736 & ~n32740;
  assign n32742 = ~n31409 & n32741;
  assign n32743 = ~n31400 & ~n32742;
  assign po0618 = n32735 | n32743;
  assign n32745 = ~n27134 & ~n30537;
  assign n32746 = n28307 & n30537;
  assign n32747 = ~n32745 & ~n32746;
  assign n32748 = n31948 & ~n32747;
  assign n32749 = ~pi0346 & ~n31948;
  assign po0619 = n32748 | n32749;
  assign n32751 = ~pi0347 & ~n31948;
  assign n32752 = n28307 & ~n30537;
  assign n32753 = ~n24900 & n30537;
  assign n32754 = ~n32752 & ~n32753;
  assign n32755 = n31948 & ~n32754;
  assign po0620 = n32751 | n32755;
  assign n32757 = n31955 & ~n32747;
  assign n32758 = ~pi0348 & ~n31955;
  assign po0621 = n32757 | n32758;
  assign n32760 = ~pi0349 & ~n31955;
  assign n32761 = n31955 & ~n32754;
  assign po0622 = n32760 | n32761;
  assign n32763 = ~pi0626 & n31013;
  assign n32764 = ~n31016 & ~n32763;
  assign n32765 = ~pi0350 & n31016;
  assign n32766 = ~n32764 & ~n32765;
  assign n32767 = pi0247 & ~n31303;
  assign n32768 = ~n31303 & ~n31312;
  assign n32769 = ~n31313 & ~n32768;
  assign n32770 = ~pi0247 & n32769;
  assign n32771 = ~n32767 & ~n32770;
  assign n32772 = n31887 & ~n32771;
  assign n32773 = pi0350 & n31889;
  assign n32774 = ~n32772 & ~n32773;
  assign n32775 = ~n31013 & ~n32774;
  assign n32776 = ~n15115 & n31350;
  assign n32777 = ~n32775 & ~n32776;
  assign n32778 = ~n31016 & ~n32777;
  assign po0623 = n32766 | n32778;
  assign n32780 = pi0975 & ~pi1422;
  assign n32781 = ~pi3147 & pi3580;
  assign n32782 = pi3578 & n32781;
  assign n32783 = pi1937 & n32780;
  assign n32784 = pi1770 & pi1855;
  assign n32785 = n32783 & n32784;
  assign n32786 = ~pi3428 & ~n32780;
  assign n32787 = ~n32785 & ~n32786;
  assign n32788 = pi2515 & ~n32787;
  assign n32789 = ~n32782 & ~n32788;
  assign n32790 = ~n32780 & ~n32789;
  assign n32791 = pi0351 & ~n32790;
  assign n32792 = ~n8591 & n8592;
  assign n32793 = ~pi3445 & ~n32792;
  assign n32794 = pi3560 & pi3566;
  assign n32795 = pi3553 & pi3565;
  assign n32796 = pi3563 & pi3564;
  assign n32797 = n32795 & n32796;
  assign n32798 = pi3577 & n32797;
  assign n32799 = pi3574 & n32798;
  assign n32800 = ~pi3567 & n32799;
  assign n32801 = n32794 & n32800;
  assign n32802 = pi4168 & n32801;
  assign n32803 = pi3567 & n32799;
  assign n32804 = pi3560 & ~pi3566;
  assign n32805 = n32803 & n32804;
  assign n32806 = pi4144 & n32805;
  assign n32807 = ~n32802 & ~n32806;
  assign n32808 = pi3567 & pi3574;
  assign n32809 = n32794 & n32808;
  assign n32810 = pi3565 & pi3577;
  assign n32811 = pi3553 & n32810;
  assign n32812 = n32809 & n32811;
  assign n32813 = ~pi3563 & pi3564;
  assign n32814 = n32812 & n32813;
  assign n32815 = pi4096 & n32814;
  assign n32816 = n32796 & n32809;
  assign n32817 = pi3553 & n32816;
  assign n32818 = ~pi3565 & pi3577;
  assign n32819 = n32817 & n32818;
  assign n32820 = pi4048 & n32819;
  assign n32821 = ~n32815 & ~n32820;
  assign n32822 = n32810 & n32816;
  assign n32823 = ~pi3553 & n32822;
  assign n32824 = pi3563 & ~pi3564;
  assign n32825 = n32812 & n32824;
  assign n32826 = pi3566 & pi3567;
  assign n32827 = n32798 & n32826;
  assign n32828 = pi3560 & ~pi3574;
  assign n32829 = n32827 & n32828;
  assign n32830 = ~pi3577 & n32797;
  assign n32831 = n32809 & n32830;
  assign n32832 = ~n32829 & ~n32831;
  assign n32833 = ~n32823 & n32832;
  assign n32834 = ~pi3560 & n32826;
  assign n32835 = n32799 & n32834;
  assign n32836 = ~n32801 & ~n32835;
  assign n32837 = ~n32805 & n32836;
  assign n32838 = n32833 & n32837;
  assign n32839 = ~n32814 & n32838;
  assign n32840 = ~n32819 & n32839;
  assign n32841 = ~n32825 & n32840;
  assign n32842 = ~n32823 & ~n32841;
  assign n32843 = pi4024 & ~n32842;
  assign n32844 = pi4072 & n32825;
  assign n32845 = ~n32843 & ~n32844;
  assign n32846 = n32821 & n32845;
  assign n32847 = n32807 & n32846;
  assign n32848 = pi4120 & n32835;
  assign n32849 = n32847 & ~n32848;
  assign n32850 = pi4192 & n32829;
  assign n32851 = pi4216 & n32831;
  assign n32852 = ~n32850 & ~n32851;
  assign n32853 = n32849 & n32852;
  assign n32854 = n32792 & ~n32853;
  assign n32855 = ~n32793 & ~n32854;
  assign n32856 = ~n8593 & ~n32855;
  assign n32857 = n8593 & ~n16855;
  assign n32858 = ~n32856 & ~n32857;
  assign n32859 = ~n10768 & ~n32858;
  assign n32860 = n10768 & ~n12726;
  assign n32861 = ~n32859 & ~n32860;
  assign n32862 = n32790 & ~n32861;
  assign po0624 = n32791 | n32862;
  assign n32864 = pi0352 & ~n32790;
  assign n32865 = ~pi3474 & ~n32792;
  assign n32866 = pi4167 & n32801;
  assign n32867 = pi4143 & n32805;
  assign n32868 = ~n32866 & ~n32867;
  assign n32869 = pi4095 & n32814;
  assign n32870 = pi4047 & n32819;
  assign n32871 = ~n32869 & ~n32870;
  assign n32872 = pi4023 & ~n32842;
  assign n32873 = pi4071 & n32825;
  assign n32874 = ~n32872 & ~n32873;
  assign n32875 = n32871 & n32874;
  assign n32876 = n32868 & n32875;
  assign n32877 = pi4119 & n32835;
  assign n32878 = n32876 & ~n32877;
  assign n32879 = pi4191 & n32829;
  assign n32880 = pi4215 & n32831;
  assign n32881 = ~n32879 & ~n32880;
  assign n32882 = n32878 & n32881;
  assign n32883 = n32792 & ~n32882;
  assign n32884 = ~n32865 & ~n32883;
  assign n32885 = ~n8593 & ~n32884;
  assign n32886 = n8593 & ~n16819;
  assign n32887 = ~n32885 & ~n32886;
  assign n32888 = ~n10768 & ~n32887;
  assign n32889 = n10768 & ~n13701;
  assign n32890 = ~n32888 & ~n32889;
  assign n32891 = n32790 & ~n32890;
  assign po0625 = n32864 | n32891;
  assign n32893 = pi0353 & ~n32790;
  assign n32894 = n10768 & ~n13121;
  assign n32895 = pi4166 & n32801;
  assign n32896 = pi4142 & n32805;
  assign n32897 = ~n32895 & ~n32896;
  assign n32898 = pi4094 & n32814;
  assign n32899 = pi4046 & n32819;
  assign n32900 = ~n32898 & ~n32899;
  assign n32901 = pi4022 & ~n32842;
  assign n32902 = pi4070 & n32825;
  assign n32903 = ~n32901 & ~n32902;
  assign n32904 = n32900 & n32903;
  assign n32905 = n32897 & n32904;
  assign n32906 = pi4118 & n32835;
  assign n32907 = n32905 & ~n32906;
  assign n32908 = pi4190 & n32829;
  assign n32909 = pi4214 & n32831;
  assign n32910 = ~n32908 & ~n32909;
  assign n32911 = n32907 & n32910;
  assign n32912 = n32792 & ~n32911;
  assign n32913 = ~pi3477 & ~n32792;
  assign n32914 = ~n32912 & ~n32913;
  assign n32915 = ~n8593 & ~n32914;
  assign n32916 = n8593 & ~n16784;
  assign n32917 = ~n32915 & ~n32916;
  assign n32918 = ~n10768 & ~n32917;
  assign n32919 = ~n32894 & ~n32918;
  assign n32920 = n32790 & ~n32919;
  assign po0626 = n32893 | n32920;
  assign n32922 = pi0354 & ~n32790;
  assign n32923 = n10768 & ~n13398;
  assign n32924 = pi4165 & n32801;
  assign n32925 = pi4141 & n32805;
  assign n32926 = ~n32924 & ~n32925;
  assign n32927 = pi4093 & n32814;
  assign n32928 = pi4045 & n32819;
  assign n32929 = ~n32927 & ~n32928;
  assign n32930 = pi4021 & ~n32842;
  assign n32931 = pi4069 & n32825;
  assign n32932 = ~n32930 & ~n32931;
  assign n32933 = n32929 & n32932;
  assign n32934 = n32926 & n32933;
  assign n32935 = pi4117 & n32835;
  assign n32936 = n32934 & ~n32935;
  assign n32937 = pi4189 & n32829;
  assign n32938 = pi4213 & n32831;
  assign n32939 = ~n32937 & ~n32938;
  assign n32940 = n32936 & n32939;
  assign n32941 = n32792 & ~n32940;
  assign n32942 = ~pi3476 & ~n32792;
  assign n32943 = ~n32941 & ~n32942;
  assign n32944 = ~n8593 & ~n32943;
  assign n32945 = n8593 & ~n16748;
  assign n32946 = ~n32944 & ~n32945;
  assign n32947 = ~n10768 & ~n32946;
  assign n32948 = ~n32923 & ~n32947;
  assign n32949 = n32790 & ~n32948;
  assign po0627 = n32922 | n32949;
  assign n32951 = pi0355 & ~n32790;
  assign n32952 = n10768 & ~n13988;
  assign n32953 = pi4164 & n32801;
  assign n32954 = pi4140 & n32805;
  assign n32955 = ~n32953 & ~n32954;
  assign n32956 = pi4092 & n32814;
  assign n32957 = pi4044 & n32819;
  assign n32958 = ~n32956 & ~n32957;
  assign n32959 = pi4020 & ~n32842;
  assign n32960 = pi4068 & n32825;
  assign n32961 = ~n32959 & ~n32960;
  assign n32962 = n32958 & n32961;
  assign n32963 = n32955 & n32962;
  assign n32964 = pi4116 & n32835;
  assign n32965 = n32963 & ~n32964;
  assign n32966 = pi4188 & n32829;
  assign n32967 = pi4212 & n32831;
  assign n32968 = ~n32966 & ~n32967;
  assign n32969 = n32965 & n32968;
  assign n32970 = n32792 & ~n32969;
  assign n32971 = ~pi3475 & ~n32792;
  assign n32972 = ~n32970 & ~n32971;
  assign n32973 = ~n8593 & ~n32972;
  assign n32974 = n8593 & ~n16712;
  assign n32975 = ~n32973 & ~n32974;
  assign n32976 = ~n10768 & ~n32975;
  assign n32977 = ~n32952 & ~n32976;
  assign n32978 = n32790 & ~n32977;
  assign po0628 = n32951 | n32978;
  assign n32980 = pi0356 & ~n32790;
  assign n32981 = n10768 & ~n12415;
  assign n32982 = pi4163 & n32801;
  assign n32983 = pi4139 & n32805;
  assign n32984 = ~n32982 & ~n32983;
  assign n32985 = pi4091 & n32814;
  assign n32986 = pi4043 & n32819;
  assign n32987 = ~n32985 & ~n32986;
  assign n32988 = pi4019 & ~n32842;
  assign n32989 = pi4067 & n32825;
  assign n32990 = ~n32988 & ~n32989;
  assign n32991 = n32987 & n32990;
  assign n32992 = n32984 & n32991;
  assign n32993 = pi4115 & n32835;
  assign n32994 = n32992 & ~n32993;
  assign n32995 = pi4187 & n32829;
  assign n32996 = pi4211 & n32831;
  assign n32997 = ~n32995 & ~n32996;
  assign n32998 = n32994 & n32997;
  assign n32999 = n32792 & ~n32998;
  assign n33000 = ~pi3470 & ~n32792;
  assign n33001 = ~n32999 & ~n33000;
  assign n33002 = ~n8593 & ~n33001;
  assign n33003 = n8593 & ~n16676;
  assign n33004 = ~n33002 & ~n33003;
  assign n33005 = ~n10768 & ~n33004;
  assign n33006 = ~n32981 & ~n33005;
  assign n33007 = n32790 & ~n33006;
  assign po0629 = n32980 | n33007;
  assign n33009 = pi0357 & ~n32790;
  assign n33010 = n10768 & ~n14816;
  assign n33011 = pi4162 & n32801;
  assign n33012 = pi4138 & n32805;
  assign n33013 = ~n33011 & ~n33012;
  assign n33014 = pi4090 & n32814;
  assign n33015 = pi4042 & n32819;
  assign n33016 = ~n33014 & ~n33015;
  assign n33017 = pi4018 & ~n32842;
  assign n33018 = pi4066 & n32825;
  assign n33019 = ~n33017 & ~n33018;
  assign n33020 = n33016 & n33019;
  assign n33021 = n33013 & n33020;
  assign n33022 = pi4114 & n32835;
  assign n33023 = n33021 & ~n33022;
  assign n33024 = pi4186 & n32829;
  assign n33025 = pi4210 & n32831;
  assign n33026 = ~n33024 & ~n33025;
  assign n33027 = n33023 & n33026;
  assign n33028 = n32792 & ~n33027;
  assign n33029 = ~pi3446 & ~n32792;
  assign n33030 = ~n33028 & ~n33029;
  assign n33031 = ~n8593 & ~n33030;
  assign n33032 = n8593 & ~n16640;
  assign n33033 = ~n33031 & ~n33032;
  assign n33034 = ~n10768 & ~n33033;
  assign n33035 = ~n33010 & ~n33034;
  assign n33036 = n32790 & ~n33035;
  assign po0630 = n33009 | n33036;
  assign n33038 = pi0358 & ~n32790;
  assign n33039 = n10768 & ~n15115;
  assign n33040 = pi4161 & n32801;
  assign n33041 = pi4137 & n32805;
  assign n33042 = ~n33040 & ~n33041;
  assign n33043 = pi4089 & n32814;
  assign n33044 = pi4041 & n32819;
  assign n33045 = ~n33043 & ~n33044;
  assign n33046 = pi4017 & ~n32842;
  assign n33047 = pi4065 & n32825;
  assign n33048 = ~n33046 & ~n33047;
  assign n33049 = n33045 & n33048;
  assign n33050 = n33042 & n33049;
  assign n33051 = pi4113 & n32835;
  assign n33052 = n33050 & ~n33051;
  assign n33053 = pi4185 & n32829;
  assign n33054 = pi4209 & n32831;
  assign n33055 = ~n33053 & ~n33054;
  assign n33056 = n33052 & n33055;
  assign n33057 = n32792 & ~n33056;
  assign n33058 = ~pi3462 & ~n32792;
  assign n33059 = ~n33057 & ~n33058;
  assign n33060 = ~n8593 & ~n33059;
  assign n33061 = n8593 & ~n16604;
  assign n33062 = ~n33060 & ~n33061;
  assign n33063 = ~n10768 & ~n33062;
  assign n33064 = ~n33039 & ~n33063;
  assign n33065 = n32790 & ~n33064;
  assign po0631 = n33038 | n33065;
  assign n33067 = pi0359 & ~n32790;
  assign n33068 = n10768 & ~n12061;
  assign n33069 = pi4160 & n32801;
  assign n33070 = pi4136 & n32805;
  assign n33071 = ~n33069 & ~n33070;
  assign n33072 = pi4088 & n32814;
  assign n33073 = pi4040 & n32819;
  assign n33074 = ~n33072 & ~n33073;
  assign n33075 = pi4016 & ~n32842;
  assign n33076 = pi4064 & n32825;
  assign n33077 = ~n33075 & ~n33076;
  assign n33078 = n33074 & n33077;
  assign n33079 = n33071 & n33078;
  assign n33080 = pi4112 & n32835;
  assign n33081 = n33079 & ~n33080;
  assign n33082 = pi4184 & n32829;
  assign n33083 = pi4208 & n32831;
  assign n33084 = ~n33082 & ~n33083;
  assign n33085 = n33081 & n33084;
  assign n33086 = n32792 & ~n33085;
  assign n33087 = ~pi3468 & ~n32792;
  assign n33088 = ~n33086 & ~n33087;
  assign n33089 = ~n8593 & ~n33088;
  assign n33090 = n8593 & ~n16568;
  assign n33091 = ~n33089 & ~n33090;
  assign n33092 = ~n10768 & ~n33091;
  assign n33093 = ~n33068 & ~n33092;
  assign n33094 = n32790 & ~n33093;
  assign po0632 = n33067 | n33094;
  assign n33096 = pi0360 & ~n32790;
  assign n33097 = n10768 & ~n17368;
  assign n33098 = ~pi3467 & ~n32792;
  assign n33099 = pi4174 & n32801;
  assign n33100 = pi4150 & n32805;
  assign n33101 = ~n33099 & ~n33100;
  assign n33102 = pi4102 & n32814;
  assign n33103 = pi4054 & n32819;
  assign n33104 = ~n33102 & ~n33103;
  assign n33105 = pi4030 & ~n32842;
  assign n33106 = pi4078 & n32825;
  assign n33107 = ~n33105 & ~n33106;
  assign n33108 = n33104 & n33107;
  assign n33109 = n33101 & n33108;
  assign n33110 = pi4126 & n32835;
  assign n33111 = n33109 & ~n33110;
  assign n33112 = pi4198 & n32829;
  assign n33113 = pi4222 & n32831;
  assign n33114 = ~n33112 & ~n33113;
  assign n33115 = n33111 & n33114;
  assign n33116 = n32792 & ~n33115;
  assign n33117 = ~n33098 & ~n33116;
  assign n33118 = ~n8593 & ~n33117;
  assign n33119 = n8593 & ~n17397;
  assign n33120 = ~n33118 & ~n33119;
  assign n33121 = ~n10768 & ~n33120;
  assign n33122 = ~n33097 & ~n33121;
  assign n33123 = n32790 & ~n33122;
  assign po0633 = n33096 | n33123;
  assign n33125 = pi0361 & ~n32790;
  assign n33126 = n10768 & ~n17199;
  assign n33127 = ~pi3465 & ~n32792;
  assign n33128 = pi4173 & n32801;
  assign n33129 = pi4149 & n32805;
  assign n33130 = ~n33128 & ~n33129;
  assign n33131 = pi4101 & n32814;
  assign n33132 = pi4053 & n32819;
  assign n33133 = ~n33131 & ~n33132;
  assign n33134 = pi4029 & ~n32842;
  assign n33135 = pi4077 & n32825;
  assign n33136 = ~n33134 & ~n33135;
  assign n33137 = n33133 & n33136;
  assign n33138 = n33130 & n33137;
  assign n33139 = pi4125 & n32835;
  assign n33140 = n33138 & ~n33139;
  assign n33141 = pi4197 & n32829;
  assign n33142 = pi4221 & n32831;
  assign n33143 = ~n33141 & ~n33142;
  assign n33144 = n33140 & n33143;
  assign n33145 = n32792 & ~n33144;
  assign n33146 = ~n33127 & ~n33145;
  assign n33147 = ~n8593 & ~n33146;
  assign n33148 = n8593 & ~n17105;
  assign n33149 = ~n33147 & ~n33148;
  assign n33150 = ~n10768 & ~n33149;
  assign n33151 = ~n33126 & ~n33150;
  assign n33152 = n32790 & ~n33151;
  assign po0634 = n33125 | n33152;
  assign n33154 = pi0362 & ~n32790;
  assign n33155 = ~pi3466 & ~n32792;
  assign n33156 = pi4172 & n32801;
  assign n33157 = pi4148 & n32805;
  assign n33158 = ~n33156 & ~n33157;
  assign n33159 = pi4100 & n32814;
  assign n33160 = pi4052 & n32819;
  assign n33161 = ~n33159 & ~n33160;
  assign n33162 = pi4028 & ~n32842;
  assign n33163 = pi4076 & n32825;
  assign n33164 = ~n33162 & ~n33163;
  assign n33165 = n33161 & n33164;
  assign n33166 = n33158 & n33165;
  assign n33167 = pi4124 & n32835;
  assign n33168 = n33166 & ~n33167;
  assign n33169 = pi4196 & n32829;
  assign n33170 = pi4220 & n32831;
  assign n33171 = ~n33169 & ~n33170;
  assign n33172 = n33168 & n33171;
  assign n33173 = n32792 & ~n33172;
  assign n33174 = ~n33155 & ~n33173;
  assign n33175 = ~n8593 & ~n33174;
  assign n33176 = n8593 & ~n16999;
  assign n33177 = ~n33175 & ~n33176;
  assign n33178 = ~n10768 & ~n33177;
  assign n33179 = ~n9825 & n10768;
  assign n33180 = ~n33178 & ~n33179;
  assign n33181 = n32790 & ~n33180;
  assign po0635 = n33154 | n33181;
  assign n33183 = pi0363 & ~n32790;
  assign n33184 = ~pi3447 & ~n32792;
  assign n33185 = pi4171 & n32801;
  assign n33186 = pi4147 & n32805;
  assign n33187 = ~n33185 & ~n33186;
  assign n33188 = pi4099 & n32814;
  assign n33189 = pi4051 & n32819;
  assign n33190 = ~n33188 & ~n33189;
  assign n33191 = pi4027 & ~n32842;
  assign n33192 = pi4075 & n32825;
  assign n33193 = ~n33191 & ~n33192;
  assign n33194 = n33190 & n33193;
  assign n33195 = n33187 & n33194;
  assign n33196 = pi4123 & n32835;
  assign n33197 = n33195 & ~n33196;
  assign n33198 = pi4195 & n32829;
  assign n33199 = pi4219 & n32831;
  assign n33200 = ~n33198 & ~n33199;
  assign n33201 = n33197 & n33200;
  assign n33202 = n32792 & ~n33201;
  assign n33203 = ~n33184 & ~n33202;
  assign n33204 = ~n8593 & ~n33203;
  assign n33205 = n8593 & ~n16963;
  assign n33206 = ~n33204 & ~n33205;
  assign n33207 = ~n10768 & ~n33206;
  assign n33208 = ~n10608 & n10768;
  assign n33209 = ~n33207 & ~n33208;
  assign n33210 = n32790 & ~n33209;
  assign po0636 = n33183 | n33210;
  assign n33212 = pi0364 & ~n32790;
  assign n33213 = ~pi3463 & ~n32792;
  assign n33214 = pi4170 & n32801;
  assign n33215 = pi4146 & n32805;
  assign n33216 = ~n33214 & ~n33215;
  assign n33217 = pi4098 & n32814;
  assign n33218 = pi4050 & n32819;
  assign n33219 = ~n33217 & ~n33218;
  assign n33220 = pi4026 & ~n32842;
  assign n33221 = pi4074 & n32825;
  assign n33222 = ~n33220 & ~n33221;
  assign n33223 = n33219 & n33222;
  assign n33224 = n33216 & n33223;
  assign n33225 = pi4122 & n32835;
  assign n33226 = n33224 & ~n33225;
  assign n33227 = pi4194 & n32829;
  assign n33228 = pi4218 & n32831;
  assign n33229 = ~n33227 & ~n33228;
  assign n33230 = n33226 & n33229;
  assign n33231 = n32792 & ~n33230;
  assign n33232 = ~n33213 & ~n33231;
  assign n33233 = ~n8593 & ~n33232;
  assign n33234 = n8593 & ~n16927;
  assign n33235 = ~n33233 & ~n33234;
  assign n33236 = ~n10768 & ~n33235;
  assign n33237 = n10768 & ~n15426;
  assign n33238 = ~n33236 & ~n33237;
  assign n33239 = n32790 & ~n33238;
  assign po0637 = n33212 | n33239;
  assign n33241 = pi0365 & ~n32790;
  assign n33242 = ~pi3448 & ~n32792;
  assign n33243 = pi4169 & n32801;
  assign n33244 = pi4145 & n32805;
  assign n33245 = ~n33243 & ~n33244;
  assign n33246 = pi4097 & n32814;
  assign n33247 = pi4049 & n32819;
  assign n33248 = ~n33246 & ~n33247;
  assign n33249 = pi4025 & ~n32842;
  assign n33250 = pi4073 & n32825;
  assign n33251 = ~n33249 & ~n33250;
  assign n33252 = n33248 & n33251;
  assign n33253 = n33245 & n33252;
  assign n33254 = pi4121 & n32835;
  assign n33255 = n33253 & ~n33254;
  assign n33256 = pi4193 & n32829;
  assign n33257 = pi4217 & n32831;
  assign n33258 = ~n33256 & ~n33257;
  assign n33259 = n33255 & n33258;
  assign n33260 = n32792 & ~n33259;
  assign n33261 = ~n33242 & ~n33260;
  assign n33262 = ~n8593 & ~n33261;
  assign n33263 = n8593 & ~n16891;
  assign n33264 = ~n33262 & ~n33263;
  assign n33265 = ~n10768 & ~n33264;
  assign n33266 = n10768 & ~n14403;
  assign n33267 = ~n33265 & ~n33266;
  assign n33268 = n32790 & ~n33267;
  assign po0638 = n33241 | n33268;
  assign n33270 = pi0366 & ~n32790;
  assign n33271 = n10768 & ~n11181;
  assign n33272 = pi4159 & n32801;
  assign n33273 = pi4135 & n32805;
  assign n33274 = ~n33272 & ~n33273;
  assign n33275 = pi4087 & n32814;
  assign n33276 = pi4039 & n32819;
  assign n33277 = ~n33275 & ~n33276;
  assign n33278 = pi4015 & ~n32842;
  assign n33279 = pi4063 & n32825;
  assign n33280 = ~n33278 & ~n33279;
  assign n33281 = n33277 & n33280;
  assign n33282 = n33274 & n33281;
  assign n33283 = pi4111 & n32835;
  assign n33284 = n33282 & ~n33283;
  assign n33285 = pi4183 & n32829;
  assign n33286 = pi4207 & n32831;
  assign n33287 = ~n33285 & ~n33286;
  assign n33288 = n33284 & n33287;
  assign n33289 = n32792 & ~n33288;
  assign n33290 = ~pi3464 & ~n32792;
  assign n33291 = ~n33289 & ~n33290;
  assign n33292 = ~n8593 & ~n33291;
  assign n33293 = n8593 & ~n16529;
  assign n33294 = ~n33292 & ~n33293;
  assign n33295 = ~n10768 & ~n33294;
  assign n33296 = ~n33271 & ~n33295;
  assign n33297 = n32790 & ~n33296;
  assign po0639 = n33270 | n33297;
  assign n33299 = n31818 & ~n31823;
  assign n33300 = ~n31824 & ~n33299;
  assign n33301 = n31865 & ~n33300;
  assign n33302 = pi3641 & n33301;
  assign n33303 = pi0367 & ~n32073;
  assign n33304 = ~n33302 & ~n33303;
  assign n33305 = ~n31777 & ~n33304;
  assign n33306 = pi1725 & n31777;
  assign n33307 = ~n33305 & ~n33306;
  assign n33308 = ~n31779 & ~n33307;
  assign n33309 = ~pi2395 & n31779;
  assign po0640 = n33308 | n33309;
  assign n33311 = pi2555 & n26299;
  assign n33312 = ~pi2555 & ~n13398;
  assign n33313 = ~n33311 & ~n33312;
  assign n33314 = ~n26062 & ~n33313;
  assign n33315 = pi0368 & n26062;
  assign po0641 = n33314 | n33315;
  assign n33317 = ~pi2567 & pi3142;
  assign n33318 = ~pi3246 & n33317;
  assign n33319 = ~pi3255 & ~pi3271;
  assign n33320 = pi3266 & n33319;
  assign n33321 = n33318 & n33320;
  assign n33322 = pi0785 & n33321;
  assign n33323 = ~pi3682 & ~n33172;
  assign n33324 = ~pi3261 & pi3682;
  assign n33325 = ~n33323 & ~n33324;
  assign n33326 = pi3305 & ~n33325;
  assign n33327 = ~n33322 & ~n33326;
  assign n33328 = pi3305 & ~n9352;
  assign n33329 = ~n33321 & ~n33328;
  assign n33330 = ~pi1008 & ~pi3426;
  assign n33331 = ~pi3305 & ~n33330;
  assign n33332 = pi3142 & n33331;
  assign n33333 = pi2567 & n33332;
  assign n33334 = ~n33329 & ~n33333;
  assign n33335 = ~n9352 & n33330;
  assign n33336 = ~n33333 & n33335;
  assign n33337 = ~n33334 & ~n33336;
  assign n33338 = ~n33327 & ~n33337;
  assign n33339 = pi0369 & n33337;
  assign po0642 = n33338 | n33339;
  assign n33341 = ~pi0694 & n31013;
  assign n33342 = ~n31016 & ~n33341;
  assign n33343 = ~pi0370 & n31016;
  assign n33344 = ~n33342 & ~n33343;
  assign n33345 = ~n12061 & n31350;
  assign n33346 = pi0247 & ~n31308;
  assign n33347 = ~n31308 & ~n31311;
  assign n33348 = ~n31312 & ~n33347;
  assign n33349 = ~pi0247 & n33348;
  assign n33350 = ~n33346 & ~n33349;
  assign n33351 = n31887 & ~n33350;
  assign n33352 = pi0370 & n31889;
  assign n33353 = ~n33351 & ~n33352;
  assign n33354 = ~n31013 & ~n33353;
  assign n33355 = ~n33345 & ~n33354;
  assign n33356 = ~n31016 & ~n33355;
  assign po0643 = n33344 | n33356;
  assign n33358 = pi0825 & n33321;
  assign n33359 = ~pi3682 & ~n33201;
  assign n33360 = ~pi3283 & pi3682;
  assign n33361 = ~n33359 & ~n33360;
  assign n33362 = pi3305 & ~n33361;
  assign n33363 = ~n33358 & ~n33362;
  assign n33364 = ~n33337 & ~n33363;
  assign n33365 = pi0371 & n33337;
  assign po0644 = n33364 | n33365;
  assign n33367 = pi0855 & n33321;
  assign n33368 = ~pi3682 & ~n33230;
  assign n33369 = ~pi3273 & pi3682;
  assign n33370 = ~n33368 & ~n33369;
  assign n33371 = pi3305 & ~n33370;
  assign n33372 = ~n33367 & ~n33371;
  assign n33373 = ~n33337 & ~n33372;
  assign n33374 = pi0372 & n33337;
  assign po0645 = n33373 | n33374;
  assign n33376 = pi0856 & n33321;
  assign n33377 = ~pi3682 & ~n33259;
  assign n33378 = ~pi3263 & pi3682;
  assign n33379 = ~n33377 & ~n33378;
  assign n33380 = pi3305 & ~n33379;
  assign n33381 = ~n33376 & ~n33380;
  assign n33382 = ~n33337 & ~n33381;
  assign n33383 = pi0373 & n33337;
  assign po0646 = n33382 | n33383;
  assign n33385 = pi0857 & n33321;
  assign n33386 = ~pi3682 & ~n32853;
  assign n33387 = ~pi3282 & pi3682;
  assign n33388 = ~n33386 & ~n33387;
  assign n33389 = pi3305 & ~n33388;
  assign n33390 = ~n33385 & ~n33389;
  assign n33391 = ~n33337 & ~n33390;
  assign n33392 = pi0374 & n33337;
  assign po0647 = n33391 | n33392;
  assign n33394 = pi0858 & n33321;
  assign n33395 = ~pi3682 & ~n32882;
  assign n33396 = ~pi3264 & pi3682;
  assign n33397 = ~n33395 & ~n33396;
  assign n33398 = pi3305 & ~n33397;
  assign n33399 = ~n33394 & ~n33398;
  assign n33400 = ~n33337 & ~n33399;
  assign n33401 = pi0375 & n33337;
  assign po0648 = n33400 | n33401;
  assign n33403 = ~n17368 & n33330;
  assign n33404 = ~n33337 & ~n33403;
  assign n33405 = ~pi0376 & n33337;
  assign n33406 = ~n33404 & ~n33405;
  assign n33407 = ~pi3682 & ~n32911;
  assign n33408 = ~pi3274 & pi3682;
  assign n33409 = ~n33407 & ~n33408;
  assign n33410 = pi3305 & ~n33409;
  assign n33411 = pi0824 & n33321;
  assign n33412 = ~n33410 & ~n33411;
  assign n33413 = ~n33337 & ~n33412;
  assign po0649 = n33406 | n33413;
  assign n33415 = ~n17199 & n33330;
  assign n33416 = ~n33337 & ~n33415;
  assign n33417 = ~pi0377 & n33337;
  assign n33418 = ~n33416 & ~n33417;
  assign n33419 = ~pi3682 & ~n32940;
  assign n33420 = ~pi3280 & pi3682;
  assign n33421 = ~n33419 & ~n33420;
  assign n33422 = pi3305 & ~n33421;
  assign n33423 = pi0823 & n33321;
  assign n33424 = ~n33422 & ~n33423;
  assign n33425 = ~n33337 & ~n33424;
  assign po0650 = n33418 | n33425;
  assign n33427 = ~n9825 & n33330;
  assign n33428 = ~n33337 & ~n33427;
  assign n33429 = ~pi0378 & n33337;
  assign n33430 = ~n33428 & ~n33429;
  assign n33431 = ~pi3682 & ~n32969;
  assign n33432 = ~pi3279 & pi3682;
  assign n33433 = ~n33431 & ~n33432;
  assign n33434 = pi3305 & ~n33433;
  assign n33435 = pi0859 & n33321;
  assign n33436 = ~n33434 & ~n33435;
  assign n33437 = ~n33337 & ~n33436;
  assign po0651 = n33430 | n33437;
  assign n33439 = pi0853 & n33321;
  assign n33440 = ~pi3682 & ~n33115;
  assign n33441 = ~pi3253 & pi3682;
  assign n33442 = ~n33440 & ~n33441;
  assign n33443 = pi3305 & ~n33442;
  assign n33444 = ~n33439 & ~n33443;
  assign n33445 = ~n33337 & ~n33444;
  assign n33446 = pi0379 & n33337;
  assign po0652 = n33445 | n33446;
  assign n33448 = pi0854 & n33321;
  assign n33449 = ~pi3682 & ~n33144;
  assign n33450 = ~pi3272 & pi3682;
  assign n33451 = ~n33449 & ~n33450;
  assign n33452 = pi3305 & ~n33451;
  assign n33453 = ~n33448 & ~n33452;
  assign n33454 = ~n33337 & ~n33453;
  assign n33455 = pi0380 & n33337;
  assign po0653 = n33454 | n33455;
  assign n33457 = ~n10608 & n33330;
  assign n33458 = ~n33337 & ~n33457;
  assign n33459 = ~pi0381 & n33337;
  assign n33460 = ~n33458 & ~n33459;
  assign n33461 = ~pi3682 & ~n32998;
  assign n33462 = ~pi3275 & pi3682;
  assign n33463 = ~n33461 & ~n33462;
  assign n33464 = pi3305 & ~n33463;
  assign n33465 = pi0730 & n33321;
  assign n33466 = ~n33464 & ~n33465;
  assign n33467 = ~n33337 & ~n33466;
  assign po0654 = n33460 | n33467;
  assign n33469 = ~n12726 & n33330;
  assign n33470 = ~n33337 & ~n33469;
  assign n33471 = ~pi0382 & n33337;
  assign n33472 = ~n33470 & ~n33471;
  assign n33473 = ~pi3682 & ~n33085;
  assign n33474 = ~pi3258 & pi3682;
  assign n33475 = ~n33473 & ~n33474;
  assign n33476 = pi3305 & ~n33475;
  assign n33477 = pi0851 & n33321;
  assign n33478 = ~n33476 & ~n33477;
  assign n33479 = ~n33337 & ~n33478;
  assign po0655 = n33472 | n33479;
  assign n33481 = ~n13701 & n33330;
  assign n33482 = ~n33337 & ~n33481;
  assign n33483 = ~pi0383 & n33337;
  assign n33484 = ~n33482 & ~n33483;
  assign n33485 = ~pi3682 & ~n33288;
  assign n33486 = ~pi3259 & pi3682;
  assign n33487 = ~n33485 & ~n33486;
  assign n33488 = pi3305 & ~n33487;
  assign n33489 = pi0860 & n33321;
  assign n33490 = ~n33488 & ~n33489;
  assign n33491 = ~n33337 & ~n33490;
  assign po0656 = n33484 | n33491;
  assign n33493 = ~n13121 & n33330;
  assign n33494 = ~n33337 & ~n33493;
  assign n33495 = ~pi0384 & n33337;
  assign n33496 = ~n33494 & ~n33495;
  assign n33497 = pi4158 & n32801;
  assign n33498 = pi4134 & n32805;
  assign n33499 = ~n33497 & ~n33498;
  assign n33500 = pi4086 & n32814;
  assign n33501 = pi4038 & n32819;
  assign n33502 = ~n33500 & ~n33501;
  assign n33503 = pi4014 & ~n32842;
  assign n33504 = pi4062 & n32825;
  assign n33505 = ~n33503 & ~n33504;
  assign n33506 = n33502 & n33505;
  assign n33507 = n33499 & n33506;
  assign n33508 = pi4110 & n32835;
  assign n33509 = n33507 & ~n33508;
  assign n33510 = pi4182 & n32829;
  assign n33511 = pi4206 & n32831;
  assign n33512 = ~n33510 & ~n33511;
  assign n33513 = n33509 & n33512;
  assign n33514 = ~pi3682 & ~n33513;
  assign n33515 = ~pi3286 & pi3682;
  assign n33516 = ~n33514 & ~n33515;
  assign n33517 = pi3305 & ~n33516;
  assign n33518 = pi0852 & n33321;
  assign n33519 = ~n33517 & ~n33518;
  assign n33520 = ~n33337 & ~n33519;
  assign po0657 = n33496 | n33520;
  assign n33522 = ~n13398 & n33330;
  assign n33523 = ~n33337 & ~n33522;
  assign n33524 = ~pi0385 & n33337;
  assign n33525 = ~n33523 & ~n33524;
  assign n33526 = pi4157 & n32801;
  assign n33527 = pi4133 & n32805;
  assign n33528 = ~n33526 & ~n33527;
  assign n33529 = pi4085 & n32814;
  assign n33530 = pi4037 & n32819;
  assign n33531 = ~n33529 & ~n33530;
  assign n33532 = pi4013 & ~n32842;
  assign n33533 = pi4061 & n32825;
  assign n33534 = ~n33532 & ~n33533;
  assign n33535 = n33531 & n33534;
  assign n33536 = n33528 & n33535;
  assign n33537 = pi4109 & n32835;
  assign n33538 = n33536 & ~n33537;
  assign n33539 = pi4181 & n32829;
  assign n33540 = pi4205 & n32831;
  assign n33541 = ~n33539 & ~n33540;
  assign n33542 = n33538 & n33541;
  assign n33543 = ~pi3682 & ~n33542;
  assign n33544 = ~pi3287 & pi3682;
  assign n33545 = ~n33543 & ~n33544;
  assign n33546 = pi3305 & ~n33545;
  assign n33547 = pi0821 & n33321;
  assign n33548 = ~n33546 & ~n33547;
  assign n33549 = ~n33337 & ~n33548;
  assign po0658 = n33525 | n33549;
  assign n33551 = ~n13988 & n33330;
  assign n33552 = ~n33337 & ~n33551;
  assign n33553 = ~pi0386 & n33337;
  assign n33554 = ~n33552 & ~n33553;
  assign n33555 = pi4156 & n32801;
  assign n33556 = pi4132 & n32805;
  assign n33557 = ~n33555 & ~n33556;
  assign n33558 = pi4084 & n32814;
  assign n33559 = pi4036 & n32819;
  assign n33560 = ~n33558 & ~n33559;
  assign n33561 = pi4012 & ~n32842;
  assign n33562 = pi4060 & n32825;
  assign n33563 = ~n33561 & ~n33562;
  assign n33564 = n33560 & n33563;
  assign n33565 = n33557 & n33564;
  assign n33566 = pi4108 & n32835;
  assign n33567 = n33565 & ~n33566;
  assign n33568 = pi4180 & n32829;
  assign n33569 = pi4204 & n32831;
  assign n33570 = ~n33568 & ~n33569;
  assign n33571 = n33567 & n33570;
  assign n33572 = ~pi3682 & ~n33571;
  assign n33573 = ~pi3289 & pi3682;
  assign n33574 = ~n33572 & ~n33573;
  assign n33575 = pi3305 & ~n33574;
  assign n33576 = ~pi0937 & n33321;
  assign n33577 = ~n33575 & ~n33576;
  assign n33578 = ~n33337 & ~n33577;
  assign po0659 = n33554 | n33578;
  assign n33580 = ~n12415 & n33330;
  assign n33581 = ~n33337 & ~n33580;
  assign n33582 = ~pi0387 & n33337;
  assign n33583 = ~n33581 & ~n33582;
  assign n33584 = pi4155 & n32801;
  assign n33585 = pi4131 & n32805;
  assign n33586 = ~n33584 & ~n33585;
  assign n33587 = pi4083 & n32814;
  assign n33588 = pi4035 & n32819;
  assign n33589 = ~n33587 & ~n33588;
  assign n33590 = pi4011 & ~n32842;
  assign n33591 = pi4059 & n32825;
  assign n33592 = ~n33590 & ~n33591;
  assign n33593 = n33589 & n33592;
  assign n33594 = n33586 & n33593;
  assign n33595 = pi4107 & n32835;
  assign n33596 = n33594 & ~n33595;
  assign n33597 = pi4179 & n32829;
  assign n33598 = pi4203 & n32831;
  assign n33599 = ~n33597 & ~n33598;
  assign n33600 = n33596 & n33599;
  assign n33601 = ~pi3682 & ~n33600;
  assign n33602 = ~pi3288 & pi3682;
  assign n33603 = ~n33601 & ~n33602;
  assign n33604 = pi3305 & ~n33603;
  assign n33605 = ~pi1045 & n33321;
  assign n33606 = ~n33604 & ~n33605;
  assign n33607 = ~n33337 & ~n33606;
  assign po0660 = n33583 | n33607;
  assign n33609 = ~n14816 & n33330;
  assign n33610 = ~n33337 & ~n33609;
  assign n33611 = ~pi0388 & n33337;
  assign n33612 = ~n33610 & ~n33611;
  assign n33613 = pi4154 & n32801;
  assign n33614 = pi4130 & n32805;
  assign n33615 = ~n33613 & ~n33614;
  assign n33616 = pi4082 & n32814;
  assign n33617 = pi4034 & n32819;
  assign n33618 = ~n33616 & ~n33617;
  assign n33619 = pi4010 & ~n32842;
  assign n33620 = pi4058 & n32825;
  assign n33621 = ~n33619 & ~n33620;
  assign n33622 = n33618 & n33621;
  assign n33623 = n33615 & n33622;
  assign n33624 = pi4106 & n32835;
  assign n33625 = n33623 & ~n33624;
  assign n33626 = pi4178 & n32829;
  assign n33627 = pi4202 & n32831;
  assign n33628 = ~n33626 & ~n33627;
  assign n33629 = n33625 & n33628;
  assign n33630 = ~pi3682 & ~n33629;
  assign n33631 = ~pi3260 & pi3682;
  assign n33632 = ~n33630 & ~n33631;
  assign n33633 = pi3305 & ~n33632;
  assign n33634 = ~pi1082 & n33321;
  assign n33635 = ~n33633 & ~n33634;
  assign n33636 = ~n33337 & ~n33635;
  assign po0661 = n33612 | n33636;
  assign n33638 = ~n15115 & n33330;
  assign n33639 = ~n33337 & ~n33638;
  assign n33640 = ~pi0389 & n33337;
  assign n33641 = ~n33639 & ~n33640;
  assign n33642 = pi4153 & n32801;
  assign n33643 = pi4129 & n32805;
  assign n33644 = ~n33642 & ~n33643;
  assign n33645 = pi4081 & n32814;
  assign n33646 = pi4033 & n32819;
  assign n33647 = ~n33645 & ~n33646;
  assign n33648 = pi4009 & ~n32842;
  assign n33649 = pi4057 & n32825;
  assign n33650 = ~n33648 & ~n33649;
  assign n33651 = n33647 & n33650;
  assign n33652 = n33644 & n33651;
  assign n33653 = pi4105 & n32835;
  assign n33654 = n33652 & ~n33653;
  assign n33655 = pi4177 & n32829;
  assign n33656 = pi4201 & n32831;
  assign n33657 = ~n33655 & ~n33656;
  assign n33658 = n33654 & n33657;
  assign n33659 = ~pi3682 & ~n33658;
  assign n33660 = ~pi3284 & pi3682;
  assign n33661 = ~n33659 & ~n33660;
  assign n33662 = pi3305 & ~n33661;
  assign n33663 = ~pi1080 & n33321;
  assign n33664 = ~n33662 & ~n33663;
  assign n33665 = ~n33337 & ~n33664;
  assign po0662 = n33641 | n33665;
  assign n33667 = ~n12061 & n33330;
  assign n33668 = ~n33337 & ~n33667;
  assign n33669 = ~pi0390 & n33337;
  assign n33670 = ~n33668 & ~n33669;
  assign n33671 = pi4152 & n32801;
  assign n33672 = pi4128 & n32805;
  assign n33673 = ~n33671 & ~n33672;
  assign n33674 = pi4080 & n32814;
  assign n33675 = pi4032 & n32819;
  assign n33676 = ~n33674 & ~n33675;
  assign n33677 = pi4008 & ~n32842;
  assign n33678 = pi4056 & n32825;
  assign n33679 = ~n33677 & ~n33678;
  assign n33680 = n33676 & n33679;
  assign n33681 = n33673 & n33680;
  assign n33682 = pi4104 & n32835;
  assign n33683 = n33681 & ~n33682;
  assign n33684 = pi4176 & n32829;
  assign n33685 = pi4200 & n32831;
  assign n33686 = ~n33684 & ~n33685;
  assign n33687 = n33683 & n33686;
  assign n33688 = ~pi3682 & ~n33687;
  assign n33689 = ~pi3262 & pi3682;
  assign n33690 = ~n33688 & ~n33689;
  assign n33691 = pi3305 & ~n33690;
  assign n33692 = ~pi1052 & n33321;
  assign n33693 = ~n33691 & ~n33692;
  assign n33694 = ~n33337 & ~n33693;
  assign po0663 = n33670 | n33694;
  assign n33696 = ~n15426 & n33330;
  assign n33697 = ~n33337 & ~n33696;
  assign n33698 = ~pi0391 & n33337;
  assign n33699 = ~n33697 & ~n33698;
  assign n33700 = ~pi3682 & ~n33027;
  assign n33701 = ~pi3276 & pi3682;
  assign n33702 = ~n33700 & ~n33701;
  assign n33703 = pi3305 & ~n33702;
  assign n33704 = pi0731 & n33321;
  assign n33705 = ~n33703 & ~n33704;
  assign n33706 = ~n33337 & ~n33705;
  assign po0664 = n33699 | n33706;
  assign n33708 = ~n14403 & n33330;
  assign n33709 = ~n33337 & ~n33708;
  assign n33710 = ~pi0392 & n33337;
  assign n33711 = ~n33709 & ~n33710;
  assign n33712 = ~pi3682 & ~n33056;
  assign n33713 = ~pi3265 & pi3682;
  assign n33714 = ~n33712 & ~n33713;
  assign n33715 = pi3305 & ~n33714;
  assign n33716 = pi0938 & n33321;
  assign n33717 = ~n33715 & ~n33716;
  assign n33718 = ~n33337 & ~n33717;
  assign po0665 = n33711 | n33718;
  assign n33720 = ~n11181 & n33330;
  assign n33721 = ~n33337 & ~n33720;
  assign n33722 = ~pi0393 & n33337;
  assign n33723 = ~n33721 & ~n33722;
  assign n33724 = pi4151 & n32801;
  assign n33725 = pi4127 & n32805;
  assign n33726 = ~n33724 & ~n33725;
  assign n33727 = pi4079 & n32814;
  assign n33728 = pi4031 & n32819;
  assign n33729 = ~n33727 & ~n33728;
  assign n33730 = pi4007 & ~n32842;
  assign n33731 = pi4055 & n32825;
  assign n33732 = ~n33730 & ~n33731;
  assign n33733 = n33729 & n33732;
  assign n33734 = n33726 & n33733;
  assign n33735 = pi4103 & n32835;
  assign n33736 = n33734 & ~n33735;
  assign n33737 = pi4175 & n32829;
  assign n33738 = pi4199 & n32831;
  assign n33739 = ~n33737 & ~n33738;
  assign n33740 = n33736 & n33739;
  assign n33741 = ~pi3682 & ~n33740;
  assign n33742 = ~pi3277 & pi3682;
  assign n33743 = ~n33741 & ~n33742;
  assign n33744 = pi3305 & ~n33743;
  assign n33745 = ~pi0911 & n33321;
  assign n33746 = ~n33744 & ~n33745;
  assign n33747 = ~n33337 & ~n33746;
  assign po0666 = n33723 | n33747;
  assign n33749 = ~pi0712 & ~n24446;
  assign n33750 = pi0712 & n31555;
  assign n33751 = ~n33749 & ~n33750;
  assign n33752 = n32628 & ~n33751;
  assign n33753 = pi0394 & ~n32628;
  assign po0667 = n33752 | n33753;
  assign n33755 = n32635 & ~n33751;
  assign n33756 = pi0395 & ~n32635;
  assign po0668 = n33755 | n33756;
  assign n33758 = ~n27710 & n31382;
  assign n33759 = pi0396 & n31381;
  assign n33760 = ~n24256 & n31384;
  assign n33761 = pi0396 & ~n31384;
  assign n33762 = ~n33760 & ~n33761;
  assign n33763 = n31388 & ~n33762;
  assign n33764 = ~n33759 & ~n33763;
  assign n33765 = ~n31391 & n33764;
  assign n33766 = ~n31382 & ~n33765;
  assign po0669 = n33758 | n33766;
  assign n33768 = ~n27710 & n31400;
  assign n33769 = pi0397 & n31399;
  assign n33770 = ~n24256 & n31402;
  assign n33771 = pi0397 & ~n31402;
  assign n33772 = ~n33770 & ~n33771;
  assign n33773 = n31406 & ~n33772;
  assign n33774 = ~n33769 & ~n33773;
  assign n33775 = ~n31409 & n33774;
  assign n33776 = ~n31400 & ~n33775;
  assign po0670 = n33768 | n33776;
  assign n33778 = n31820 & n31822;
  assign n33779 = ~n31823 & ~n33778;
  assign n33780 = n31865 & ~n33779;
  assign n33781 = pi3641 & n33780;
  assign n33782 = pi0398 & ~n32073;
  assign n33783 = ~n33781 & ~n33782;
  assign n33784 = ~n31777 & ~n33783;
  assign n33785 = pi1877 & n31777;
  assign n33786 = ~n33784 & ~n33785;
  assign n33787 = ~n31779 & ~n33786;
  assign n33788 = ~pi2090 & n31779;
  assign po0671 = n33787 | n33788;
  assign n33790 = ~pi0712 & ~n24289;
  assign n33791 = pi0712 & n31525;
  assign n33792 = ~n33790 & ~n33791;
  assign n33793 = n32628 & ~n33792;
  assign n33794 = pi0399 & ~n32628;
  assign po0672 = n33793 | n33794;
  assign n33796 = n32635 & ~n33792;
  assign n33797 = pi0400 & ~n32635;
  assign po0673 = n33796 | n33797;
  assign n33799 = ~n24900 & ~n30537;
  assign n33800 = ~n25761 & n30537;
  assign n33801 = ~n33799 & ~n33800;
  assign n33802 = n31948 & ~n33801;
  assign n33803 = ~pi0401 & ~n31948;
  assign po0674 = n33802 | n33803;
  assign n33805 = n31955 & ~n33801;
  assign n33806 = ~pi0402 & ~n31955;
  assign po0675 = n33805 | n33806;
  assign n33808 = pi3362 & n8563;
  assign n33809 = ~pi0565 & n33808;
  assign n33810 = ~pi3589 & n33809;
  assign n33811 = pi2813 & ~pi3552;
  assign po3685 = n33810 | n33811;
  assign n33813 = ~po3831 & ~po3685;
  assign n33814 = ~n33325 & ~n33813;
  assign n33815 = n33317 & n33320;
  assign n33816 = pi3246 & n33815;
  assign n33817 = pi0785 & n33816;
  assign n33818 = pi0403 & ~n33816;
  assign n33819 = ~n33817 & ~n33818;
  assign n33820 = n33813 & ~n33819;
  assign po0677 = n33814 | n33820;
  assign n33822 = ~po3873 & ~po3948;
  assign n33823 = ~po3848 & n33822;
  assign n33824 = pi0404 & n33823;
  assign n33825 = po0767 & n33824;
  assign n33826 = ~pi0404 & po0767;
  assign n33827 = n9345 & n33823;
  assign n33828 = ~pi2479 & pi2900;
  assign n33829 = pi2900 & pi3056;
  assign n33830 = ~n33828 & ~n33829;
  assign n33831 = n33828 & n33829;
  assign n33832 = ~n33830 & ~n33831;
  assign n33833 = ~pi2480 & pi3072;
  assign n33834 = pi3072 & pi3108;
  assign n33835 = ~n33833 & ~n33834;
  assign n33836 = n33833 & n33834;
  assign n33837 = ~n33835 & ~n33836;
  assign n33838 = ~pi2477 & pi2955;
  assign n33839 = pi2955 & pi3095;
  assign n33840 = ~n33838 & ~n33839;
  assign n33841 = n33838 & n33839;
  assign n33842 = ~n33840 & ~n33841;
  assign n33843 = ~pi2478 & pi2995;
  assign n33844 = pi2995 & pi3011;
  assign n33845 = ~n33843 & ~n33844;
  assign n33846 = n33843 & n33844;
  assign n33847 = ~n33845 & ~n33846;
  assign n33848 = ~n33842 & ~n33847;
  assign n33849 = ~n33837 & n33848;
  assign n33850 = ~n33832 & n33849;
  assign n33851 = ~pi2483 & pi2907;
  assign n33852 = pi2907 & pi2977;
  assign n33853 = ~n33851 & ~n33852;
  assign n33854 = n33851 & n33852;
  assign n33855 = ~n33853 & ~n33854;
  assign n33856 = ~pi2516 & pi3001;
  assign n33857 = pi3001 & pi3016;
  assign n33858 = ~n33856 & ~n33857;
  assign n33859 = n33856 & n33857;
  assign n33860 = ~n33858 & ~n33859;
  assign n33861 = ~pi2481 & pi3067;
  assign n33862 = pi2991 & pi3067;
  assign n33863 = ~n33861 & ~n33862;
  assign n33864 = n33861 & n33862;
  assign n33865 = ~n33863 & ~n33864;
  assign n33866 = ~pi2482 & pi3073;
  assign n33867 = pi3012 & pi3073;
  assign n33868 = ~n33866 & ~n33867;
  assign n33869 = n33866 & n33867;
  assign n33870 = ~n33868 & ~n33869;
  assign n33871 = ~n33865 & ~n33870;
  assign n33872 = ~n33860 & n33871;
  assign n33873 = ~n33855 & n33872;
  assign n33874 = n33850 & n33873;
  assign n33875 = ~pi2475 & pi2954;
  assign n33876 = pi2954 & pi3009;
  assign n33877 = ~n33875 & ~n33876;
  assign n33878 = n33875 & n33876;
  assign n33879 = ~n33877 & ~n33878;
  assign n33880 = ~pi2476 & pi2994;
  assign n33881 = pi2994 & pi3010;
  assign n33882 = ~n33880 & ~n33881;
  assign n33883 = n33880 & n33881;
  assign n33884 = ~n33882 & ~n33883;
  assign n33885 = ~pi2518 & pi2999;
  assign n33886 = pi2959 & pi2999;
  assign n33887 = ~n33885 & ~n33886;
  assign n33888 = n33885 & n33886;
  assign n33889 = ~n33887 & ~n33888;
  assign n33890 = ~pi2517 & pi3000;
  assign n33891 = pi2786 & pi3000;
  assign n33892 = ~n33890 & ~n33891;
  assign n33893 = n33890 & n33891;
  assign n33894 = ~n33892 & ~n33893;
  assign n33895 = ~n33889 & ~n33894;
  assign n33896 = ~n33884 & n33895;
  assign n33897 = ~n33879 & n33896;
  assign n33898 = ~pi2514 & pi2908;
  assign n33899 = pi2908 & pi2984;
  assign n33900 = n33898 & ~n33899;
  assign n33901 = ~n33898 & n33899;
  assign n33902 = ~n33900 & ~n33901;
  assign n33903 = n33897 & n33902;
  assign n33904 = pi2485 & pi2886;
  assign n33905 = ~pi2485 & ~pi2886;
  assign n33906 = ~n33904 & ~n33905;
  assign n33907 = pi2901 & ~n33906;
  assign n33908 = pi2408 & pi2972;
  assign n33909 = ~pi2408 & ~pi2972;
  assign n33910 = ~n33908 & ~n33909;
  assign n33911 = pi2887 & ~n33910;
  assign n33912 = ~n33907 & ~n33911;
  assign n33913 = pi2484 & pi3015;
  assign n33914 = ~pi2484 & ~pi3015;
  assign n33915 = ~n33913 & ~n33914;
  assign n33916 = pi2998 & ~n33915;
  assign n33917 = ~pi2400 & pi3014;
  assign n33918 = pi2400 & ~pi3014;
  assign n33919 = ~n33917 & ~n33918;
  assign n33920 = pi2997 & n33919;
  assign n33921 = ~n33916 & ~n33920;
  assign n33922 = n33912 & n33921;
  assign n33923 = ~pi2996 & n33922;
  assign n33924 = ~pi2643 & n33923;
  assign n33925 = ~pi2472 & pi3013;
  assign n33926 = pi2472 & ~pi3013;
  assign n33927 = ~n33925 & ~n33926;
  assign n33928 = n33924 & ~n33927;
  assign n33929 = n33903 & n33928;
  assign n33930 = n33874 & n33929;
  assign n33931 = ~pi2475 & pi2880;
  assign n33932 = pi2815 & pi2880;
  assign n33933 = ~n33931 & ~n33932;
  assign n33934 = n33931 & n33932;
  assign n33935 = ~n33933 & ~n33934;
  assign n33936 = ~pi2476 & pi3002;
  assign n33937 = pi3002 & pi3017;
  assign n33938 = ~n33936 & ~n33937;
  assign n33939 = n33936 & n33937;
  assign n33940 = ~n33938 & ~n33939;
  assign n33941 = ~pi2518 & pi3077;
  assign n33942 = pi3023 & pi3077;
  assign n33943 = ~n33941 & ~n33942;
  assign n33944 = n33941 & n33942;
  assign n33945 = ~n33943 & ~n33944;
  assign n33946 = ~pi2517 & pi3085;
  assign n33947 = pi3024 & pi3085;
  assign n33948 = ~n33946 & ~n33947;
  assign n33949 = n33946 & n33947;
  assign n33950 = ~n33948 & ~n33949;
  assign n33951 = ~n33945 & ~n33950;
  assign n33952 = ~n33940 & n33951;
  assign n33953 = ~n33935 & n33952;
  assign n33954 = ~pi2479 & pi2884;
  assign n33955 = pi2884 & pi2956;
  assign n33956 = ~n33954 & ~n33955;
  assign n33957 = n33954 & n33955;
  assign n33958 = ~n33956 & ~n33957;
  assign n33959 = ~pi2480 & pi2821;
  assign n33960 = pi2821 & pi3019;
  assign n33961 = ~n33959 & ~n33960;
  assign n33962 = n33959 & n33960;
  assign n33963 = ~n33961 & ~n33962;
  assign n33964 = ~pi2477 & pi3003;
  assign n33965 = pi3003 & pi3066;
  assign n33966 = ~n33964 & ~n33965;
  assign n33967 = n33964 & n33965;
  assign n33968 = ~n33966 & ~n33967;
  assign n33969 = ~pi2478 & pi3004;
  assign n33970 = pi3004 & pi3018;
  assign n33971 = ~n33969 & ~n33970;
  assign n33972 = n33969 & n33970;
  assign n33973 = ~n33971 & ~n33972;
  assign n33974 = ~n33968 & ~n33973;
  assign n33975 = ~n33963 & n33974;
  assign n33976 = ~n33958 & n33975;
  assign n33977 = n33953 & n33976;
  assign n33978 = ~pi2483 & pi2838;
  assign n33979 = pi2838 & pi3021;
  assign n33980 = ~n33978 & ~n33979;
  assign n33981 = n33978 & n33979;
  assign n33982 = ~n33980 & ~n33981;
  assign n33983 = ~pi2516 & pi3008;
  assign n33984 = pi3008 & pi3025;
  assign n33985 = ~n33983 & ~n33984;
  assign n33986 = n33983 & n33984;
  assign n33987 = ~n33985 & ~n33986;
  assign n33988 = ~pi2481 & pi2822;
  assign n33989 = pi2790 & pi2822;
  assign n33990 = ~n33988 & ~n33989;
  assign n33991 = n33988 & n33989;
  assign n33992 = ~n33990 & ~n33991;
  assign n33993 = ~pi2482 & pi2839;
  assign n33994 = pi2839 & pi3020;
  assign n33995 = ~n33993 & ~n33994;
  assign n33996 = n33993 & n33994;
  assign n33997 = ~n33995 & ~n33996;
  assign n33998 = ~n33992 & ~n33997;
  assign n33999 = ~n33987 & n33998;
  assign n34000 = ~n33982 & n33999;
  assign n34001 = ~pi2514 & pi2858;
  assign n34002 = pi2858 & pi2909;
  assign n34003 = n34001 & ~n34002;
  assign n34004 = ~n34001 & n34002;
  assign n34005 = ~n34003 & ~n34004;
  assign n34006 = n34000 & n34005;
  assign n34007 = ~pi2472 & pi3022;
  assign n34008 = pi2472 & ~pi3022;
  assign n34009 = ~n34007 & ~n34008;
  assign n34010 = pi2484 & pi2906;
  assign n34011 = ~pi2484 & ~pi2906;
  assign n34012 = ~n34010 & ~n34011;
  assign n34013 = pi3007 & ~n34012;
  assign n34014 = pi2485 & pi2885;
  assign n34015 = ~pi2485 & ~pi2885;
  assign n34016 = ~n34014 & ~n34015;
  assign n34017 = pi3094 & ~n34016;
  assign n34018 = ~n34013 & ~n34017;
  assign n34019 = pi2408 & pi2910;
  assign n34020 = ~pi2408 & ~pi2910;
  assign n34021 = ~n34019 & ~n34020;
  assign n34022 = pi2857 & ~n34021;
  assign n34023 = ~pi2400 & pi2837;
  assign n34024 = pi2400 & ~pi2837;
  assign n34025 = ~n34023 & ~n34024;
  assign n34026 = pi3006 & n34025;
  assign n34027 = ~n34022 & ~n34026;
  assign n34028 = n34018 & n34027;
  assign n34029 = ~pi3005 & n34028;
  assign n34030 = ~pi2643 & n34029;
  assign n34031 = ~n34009 & n34030;
  assign n34032 = n34006 & n34031;
  assign n34033 = n33977 & n34032;
  assign n34034 = pi2800 & ~pi3644;
  assign n34035 = ~pi3362 & n34034;
  assign n34036 = ~pi3643 & n34035;
  assign n34037 = pi0408 & ~pi2762;
  assign n34038 = n8607 & n9373;
  assign n34039 = ~pi0405 & ~pi0421;
  assign n34040 = n34038 & n34039;
  assign n34041 = n34037 & n34040;
  assign n34042 = ~pi2417 & ~pi3426;
  assign n34043 = pi3026 & pi3040;
  assign n34044 = ~pi1028 & pi3026;
  assign n34045 = ~n34043 & ~n34044;
  assign n34046 = n34043 & n34044;
  assign n34047 = ~n34045 & ~n34046;
  assign n34048 = pi3081 & pi3103;
  assign n34049 = ~pi1029 & pi3081;
  assign n34050 = ~n34048 & ~n34049;
  assign n34051 = n34048 & n34049;
  assign n34052 = ~n34050 & ~n34051;
  assign n34053 = pi3046 & pi3078;
  assign n34054 = ~pi1037 & pi3078;
  assign n34055 = ~n34053 & ~n34054;
  assign n34056 = n34053 & n34054;
  assign n34057 = ~n34055 & ~n34056;
  assign n34058 = pi3031 & pi3061;
  assign n34059 = ~pi1038 & pi3031;
  assign n34060 = ~n34058 & ~n34059;
  assign n34061 = n34058 & n34059;
  assign n34062 = ~n34060 & ~n34061;
  assign n34063 = ~n34057 & ~n34062;
  assign n34064 = ~n34052 & n34063;
  assign n34065 = ~n34047 & n34064;
  assign n34066 = pi2806 & pi3029;
  assign n34067 = ~pi2979 & pi3029;
  assign n34068 = ~n34066 & n34067;
  assign n34069 = n34066 & ~n34067;
  assign n34070 = ~n34068 & ~n34069;
  assign n34071 = pi3028 & pi3042;
  assign n34072 = ~pi1012 & pi3028;
  assign n34073 = ~n34071 & ~n34072;
  assign n34074 = n34071 & n34072;
  assign n34075 = ~n34073 & ~n34074;
  assign n34076 = pi3032 & pi3047;
  assign n34077 = ~pi1039 & pi3032;
  assign n34078 = ~n34076 & ~n34077;
  assign n34079 = n34076 & n34077;
  assign n34080 = ~n34078 & ~n34079;
  assign n34081 = pi3041 & pi3060;
  assign n34082 = ~pi1033 & pi3060;
  assign n34083 = ~n34081 & ~n34082;
  assign n34084 = n34081 & n34082;
  assign n34085 = ~n34083 & ~n34084;
  assign n34086 = pi2811 & pi2859;
  assign n34087 = ~pi1034 & pi2859;
  assign n34088 = ~n34086 & ~n34087;
  assign n34089 = n34086 & n34087;
  assign n34090 = ~n34088 & ~n34089;
  assign n34091 = ~n34085 & ~n34090;
  assign n34092 = ~n34080 & n34091;
  assign n34093 = ~n34075 & n34092;
  assign n34094 = pi2791 & pi3027;
  assign n34095 = ~pi1013 & pi3027;
  assign n34096 = ~n34094 & ~n34095;
  assign n34097 = n34094 & n34095;
  assign n34098 = ~n34096 & ~n34097;
  assign n34099 = pi2970 & pi3062;
  assign n34100 = ~pi1032 & pi3062;
  assign n34101 = ~n34099 & ~n34100;
  assign n34102 = n34099 & n34100;
  assign n34103 = ~n34101 & ~n34102;
  assign n34104 = pi2898 & pi3087;
  assign n34105 = ~pi1030 & pi3087;
  assign n34106 = ~n34104 & ~n34105;
  assign n34107 = n34104 & n34105;
  assign n34108 = ~n34106 & ~n34107;
  assign n34109 = pi3090 & pi3092;
  assign n34110 = ~pi1031 & pi3090;
  assign n34111 = ~n34109 & ~n34110;
  assign n34112 = n34109 & n34110;
  assign n34113 = ~n34111 & ~n34112;
  assign n34114 = ~n34108 & ~n34113;
  assign n34115 = ~n34103 & n34114;
  assign n34116 = ~n34098 & n34115;
  assign n34117 = n34093 & n34116;
  assign n34118 = n34070 & n34117;
  assign n34119 = n34065 & n34118;
  assign n34120 = pi3045 & pi3070;
  assign n34121 = ~pi1035 & pi3070;
  assign n34122 = ~n34120 & n34121;
  assign n34123 = n34120 & ~n34121;
  assign n34124 = ~n34122 & ~n34123;
  assign n34125 = n34119 & n34124;
  assign n34126 = pi3030 & pi3088;
  assign n34127 = ~pi1036 & pi3030;
  assign n34128 = ~n34126 & ~n34127;
  assign n34129 = n34126 & n34127;
  assign n34130 = ~n34128 & ~n34129;
  assign n34131 = pi2904 & pi3058;
  assign n34132 = ~pi2981 & pi3058;
  assign n34133 = ~n34131 & ~n34132;
  assign n34134 = n34131 & n34132;
  assign n34135 = ~n34133 & ~n34134;
  assign n34136 = pi3044 & pi3057;
  assign n34137 = ~pi2980 & pi3057;
  assign n34138 = ~n34136 & ~n34137;
  assign n34139 = n34136 & n34137;
  assign n34140 = ~n34138 & ~n34139;
  assign n34141 = ~n34135 & ~n34140;
  assign n34142 = ~n34130 & n34141;
  assign n34143 = n34125 & n34142;
  assign n34144 = n34042 & n34143;
  assign n34145 = ~pi2978 & pi3043;
  assign n34146 = pi2978 & ~pi3043;
  assign n34147 = ~n34145 & ~n34146;
  assign n34148 = ~pi2902 & ~pi3083;
  assign n34149 = ~n34147 & n34148;
  assign n34150 = n34144 & n34149;
  assign n34151 = ~pi2409 & pi3043;
  assign n34152 = pi2409 & ~pi3043;
  assign n34153 = ~n34151 & ~n34152;
  assign n34154 = ~pi2644 & pi3087;
  assign n34155 = ~n34104 & n34154;
  assign n34156 = n34104 & ~n34154;
  assign n34157 = ~n34155 & ~n34156;
  assign n34158 = ~pi2797 & pi3090;
  assign n34159 = ~n34109 & n34158;
  assign n34160 = n34109 & ~n34158;
  assign n34161 = ~n34159 & ~n34160;
  assign n34162 = n34157 & n34161;
  assign n34163 = ~pi2645 & pi3027;
  assign n34164 = ~n34094 & n34163;
  assign n34165 = n34094 & ~n34163;
  assign n34166 = ~n34164 & ~n34165;
  assign n34167 = ~pi2553 & pi3062;
  assign n34168 = ~n34099 & n34167;
  assign n34169 = n34099 & ~n34167;
  assign n34170 = ~n34168 & ~n34169;
  assign n34171 = n34166 & n34170;
  assign n34172 = ~pi2549 & pi3028;
  assign n34173 = ~n34071 & ~n34172;
  assign n34174 = n34071 & n34172;
  assign n34175 = ~n34173 & ~n34174;
  assign n34176 = ~pi2540 & pi3032;
  assign n34177 = ~n34076 & ~n34176;
  assign n34178 = n34076 & n34176;
  assign n34179 = ~n34177 & ~n34178;
  assign n34180 = ~pi2551 & pi3060;
  assign n34181 = ~n34081 & ~n34180;
  assign n34182 = n34081 & n34180;
  assign n34183 = ~n34181 & ~n34182;
  assign n34184 = ~pi2646 & pi2859;
  assign n34185 = ~n34086 & ~n34184;
  assign n34186 = n34086 & n34184;
  assign n34187 = ~n34185 & ~n34186;
  assign n34188 = ~n34183 & ~n34187;
  assign n34189 = ~n34179 & n34188;
  assign n34190 = ~n34175 & n34189;
  assign n34191 = ~pi2794 & pi3026;
  assign n34192 = ~n34043 & ~n34191;
  assign n34193 = n34043 & n34191;
  assign n34194 = ~n34192 & ~n34193;
  assign n34195 = ~pi2796 & pi3081;
  assign n34196 = ~n34048 & ~n34195;
  assign n34197 = n34048 & n34195;
  assign n34198 = ~n34196 & ~n34197;
  assign n34199 = ~pi2953 & pi3078;
  assign n34200 = ~n34053 & ~n34199;
  assign n34201 = n34053 & n34199;
  assign n34202 = ~n34200 & ~n34201;
  assign n34203 = ~pi2788 & pi3031;
  assign n34204 = ~n34058 & ~n34203;
  assign n34205 = n34058 & n34203;
  assign n34206 = ~n34204 & ~n34205;
  assign n34207 = ~n34202 & ~n34206;
  assign n34208 = ~n34198 & n34207;
  assign n34209 = ~n34194 & n34208;
  assign n34210 = n34190 & n34209;
  assign n34211 = ~pi2473 & pi3029;
  assign n34212 = ~n34066 & ~n34211;
  assign n34213 = n34066 & n34211;
  assign n34214 = ~n34212 & ~n34213;
  assign n34215 = n34210 & ~n34214;
  assign n34216 = n34171 & n34215;
  assign n34217 = n34162 & n34216;
  assign n34218 = ~pi2647 & pi3070;
  assign n34219 = ~n34120 & n34218;
  assign n34220 = n34120 & ~n34218;
  assign n34221 = ~n34219 & ~n34220;
  assign n34222 = n34217 & n34221;
  assign n34223 = ~pi2529 & pi3030;
  assign n34224 = ~n34126 & ~n34223;
  assign n34225 = n34126 & n34223;
  assign n34226 = ~n34224 & ~n34225;
  assign n34227 = ~pi2405 & pi3058;
  assign n34228 = ~n34131 & ~n34227;
  assign n34229 = n34131 & n34227;
  assign n34230 = ~n34228 & ~n34229;
  assign n34231 = ~pi2404 & pi3057;
  assign n34232 = ~n34136 & ~n34231;
  assign n34233 = n34136 & n34231;
  assign n34234 = ~n34232 & ~n34233;
  assign n34235 = ~n34230 & ~n34234;
  assign n34236 = ~n34226 & n34235;
  assign n34237 = n34222 & n34236;
  assign n34238 = pi2902 & n34237;
  assign n34239 = ~pi3083 & n34238;
  assign n34240 = ~n34153 & n34239;
  assign n34241 = ~pi2409 & pi3052;
  assign n34242 = pi2409 & ~pi3052;
  assign n34243 = ~n34241 & ~n34242;
  assign n34244 = pi2823 & ~pi2953;
  assign n34245 = pi2823 & pi3069;
  assign n34246 = n34244 & ~n34245;
  assign n34247 = ~n34244 & n34245;
  assign n34248 = ~n34246 & ~n34247;
  assign n34249 = ~pi2788 & pi2883;
  assign n34250 = pi2775 & pi2883;
  assign n34251 = n34249 & ~n34250;
  assign n34252 = ~n34249 & n34250;
  assign n34253 = ~n34251 & ~n34252;
  assign n34254 = n34248 & n34253;
  assign n34255 = ~pi2794 & pi3033;
  assign n34256 = pi2899 & pi3033;
  assign n34257 = n34255 & ~n34256;
  assign n34258 = ~n34255 & n34256;
  assign n34259 = ~n34257 & ~n34258;
  assign n34260 = pi2792 & ~pi2796;
  assign n34261 = pi2792 & pi3048;
  assign n34262 = n34260 & ~n34261;
  assign n34263 = ~n34260 & n34261;
  assign n34264 = ~n34262 & ~n34263;
  assign n34265 = n34259 & n34264;
  assign n34266 = ~pi2549 & pi3037;
  assign n34267 = pi2818 & pi3037;
  assign n34268 = ~n34266 & ~n34267;
  assign n34269 = n34266 & n34267;
  assign n34270 = ~n34268 & ~n34269;
  assign n34271 = ~pi2540 & pi2973;
  assign n34272 = pi2882 & pi2973;
  assign n34273 = ~n34271 & ~n34272;
  assign n34274 = n34271 & n34272;
  assign n34275 = ~n34273 & ~n34274;
  assign n34276 = ~pi2551 & pi3036;
  assign n34277 = pi2957 & pi3036;
  assign n34278 = ~n34276 & ~n34277;
  assign n34279 = n34276 & n34277;
  assign n34280 = ~n34278 & ~n34279;
  assign n34281 = ~pi2646 & pi2905;
  assign n34282 = pi2905 & pi2958;
  assign n34283 = ~n34281 & ~n34282;
  assign n34284 = n34281 & n34282;
  assign n34285 = ~n34283 & ~n34284;
  assign n34286 = ~n34280 & ~n34285;
  assign n34287 = ~n34275 & n34286;
  assign n34288 = ~n34270 & n34287;
  assign n34289 = ~pi2645 & pi3035;
  assign n34290 = pi3035 & pi3110;
  assign n34291 = ~n34289 & ~n34290;
  assign n34292 = n34289 & n34290;
  assign n34293 = ~n34291 & ~n34292;
  assign n34294 = ~pi2553 & pi2903;
  assign n34295 = pi2903 & pi2971;
  assign n34296 = ~n34294 & ~n34295;
  assign n34297 = n34294 & n34295;
  assign n34298 = ~n34296 & ~n34297;
  assign n34299 = ~pi2644 & pi3034;
  assign n34300 = pi3034 & pi3049;
  assign n34301 = ~n34299 & ~n34300;
  assign n34302 = n34299 & n34300;
  assign n34303 = ~n34301 & ~n34302;
  assign n34304 = ~pi2797 & pi2881;
  assign n34305 = pi2881 & pi3050;
  assign n34306 = ~n34304 & ~n34305;
  assign n34307 = n34304 & n34305;
  assign n34308 = ~n34306 & ~n34307;
  assign n34309 = ~n34303 & ~n34308;
  assign n34310 = ~n34298 & n34309;
  assign n34311 = ~n34293 & n34310;
  assign n34312 = n34288 & n34311;
  assign n34313 = ~pi2473 & pi3038;
  assign n34314 = pi3038 & pi3053;
  assign n34315 = ~n34313 & ~n34314;
  assign n34316 = n34313 & n34314;
  assign n34317 = ~n34315 & ~n34316;
  assign n34318 = n34312 & ~n34317;
  assign n34319 = n34265 & n34318;
  assign n34320 = n34254 & n34319;
  assign n34321 = ~pi2647 & pi3064;
  assign n34322 = pi3064 & pi3080;
  assign n34323 = n34321 & ~n34322;
  assign n34324 = ~n34321 & n34322;
  assign n34325 = ~n34323 & ~n34324;
  assign n34326 = n34320 & n34325;
  assign n34327 = ~pi2529 & pi3071;
  assign n34328 = pi2915 & pi3071;
  assign n34329 = ~n34327 & ~n34328;
  assign n34330 = n34327 & n34328;
  assign n34331 = ~n34329 & ~n34330;
  assign n34332 = ~pi2405 & pi3039;
  assign n34333 = pi3039 & pi3054;
  assign n34334 = ~n34332 & ~n34333;
  assign n34335 = n34332 & n34333;
  assign n34336 = ~n34334 & ~n34335;
  assign n34337 = ~pi2404 & pi3089;
  assign n34338 = pi2930 & pi3089;
  assign n34339 = ~n34337 & ~n34338;
  assign n34340 = n34337 & n34338;
  assign n34341 = ~n34339 & ~n34340;
  assign n34342 = ~n34336 & ~n34341;
  assign n34343 = ~n34331 & n34342;
  assign n34344 = n34326 & n34343;
  assign n34345 = pi3051 & n34344;
  assign n34346 = ~pi3082 & n34345;
  assign n34347 = ~n34243 & n34346;
  assign n34348 = ~n34240 & ~n34347;
  assign n34349 = ~pi2802 & ~n34348;
  assign n34350 = ~pi3426 & n34349;
  assign n34351 = ~pi1028 & pi3033;
  assign n34352 = ~n34256 & ~n34351;
  assign n34353 = n34256 & n34351;
  assign n34354 = ~n34352 & ~n34353;
  assign n34355 = ~pi1029 & pi2792;
  assign n34356 = ~n34261 & ~n34355;
  assign n34357 = n34261 & n34355;
  assign n34358 = ~n34356 & ~n34357;
  assign n34359 = ~pi1037 & pi2823;
  assign n34360 = ~n34245 & ~n34359;
  assign n34361 = n34245 & n34359;
  assign n34362 = ~n34360 & ~n34361;
  assign n34363 = ~pi1038 & pi2883;
  assign n34364 = ~n34250 & ~n34363;
  assign n34365 = n34250 & n34363;
  assign n34366 = ~n34364 & ~n34365;
  assign n34367 = ~n34362 & ~n34366;
  assign n34368 = ~n34358 & n34367;
  assign n34369 = ~n34354 & n34368;
  assign n34370 = ~pi2979 & pi3038;
  assign n34371 = ~n34314 & n34370;
  assign n34372 = n34314 & ~n34370;
  assign n34373 = ~n34371 & ~n34372;
  assign n34374 = ~pi1012 & pi3037;
  assign n34375 = ~n34267 & ~n34374;
  assign n34376 = n34267 & n34374;
  assign n34377 = ~n34375 & ~n34376;
  assign n34378 = ~pi1039 & pi2973;
  assign n34379 = ~n34272 & ~n34378;
  assign n34380 = n34272 & n34378;
  assign n34381 = ~n34379 & ~n34380;
  assign n34382 = ~pi1033 & pi3036;
  assign n34383 = ~n34277 & ~n34382;
  assign n34384 = n34277 & n34382;
  assign n34385 = ~n34383 & ~n34384;
  assign n34386 = ~pi1034 & pi2905;
  assign n34387 = ~n34282 & ~n34386;
  assign n34388 = n34282 & n34386;
  assign n34389 = ~n34387 & ~n34388;
  assign n34390 = ~n34385 & ~n34389;
  assign n34391 = ~n34381 & n34390;
  assign n34392 = ~n34377 & n34391;
  assign n34393 = ~pi1013 & pi3035;
  assign n34394 = ~n34290 & ~n34393;
  assign n34395 = n34290 & n34393;
  assign n34396 = ~n34394 & ~n34395;
  assign n34397 = ~pi1032 & pi2903;
  assign n34398 = ~n34295 & ~n34397;
  assign n34399 = n34295 & n34397;
  assign n34400 = ~n34398 & ~n34399;
  assign n34401 = ~pi1030 & pi3034;
  assign n34402 = ~n34300 & ~n34401;
  assign n34403 = n34300 & n34401;
  assign n34404 = ~n34402 & ~n34403;
  assign n34405 = ~pi1031 & pi2881;
  assign n34406 = ~n34305 & ~n34405;
  assign n34407 = n34305 & n34405;
  assign n34408 = ~n34406 & ~n34407;
  assign n34409 = ~n34404 & ~n34408;
  assign n34410 = ~n34400 & n34409;
  assign n34411 = ~n34396 & n34410;
  assign n34412 = n34392 & n34411;
  assign n34413 = n34373 & n34412;
  assign n34414 = n34369 & n34413;
  assign n34415 = ~pi1035 & pi3064;
  assign n34416 = ~n34322 & n34415;
  assign n34417 = n34322 & ~n34415;
  assign n34418 = ~n34416 & ~n34417;
  assign n34419 = n34414 & n34418;
  assign n34420 = ~pi1036 & pi3071;
  assign n34421 = ~n34328 & ~n34420;
  assign n34422 = n34328 & n34420;
  assign n34423 = ~n34421 & ~n34422;
  assign n34424 = ~pi2981 & pi3039;
  assign n34425 = ~n34333 & ~n34424;
  assign n34426 = n34333 & n34424;
  assign n34427 = ~n34425 & ~n34426;
  assign n34428 = ~pi2980 & pi3089;
  assign n34429 = ~n34338 & ~n34428;
  assign n34430 = n34338 & n34428;
  assign n34431 = ~n34429 & ~n34430;
  assign n34432 = ~n34427 & ~n34431;
  assign n34433 = ~n34423 & n34432;
  assign n34434 = n34419 & n34433;
  assign n34435 = n34042 & n34434;
  assign n34436 = ~pi2978 & pi3052;
  assign n34437 = pi2978 & ~pi3052;
  assign n34438 = ~n34436 & ~n34437;
  assign n34439 = ~pi3051 & ~pi3082;
  assign n34440 = ~n34438 & n34439;
  assign n34441 = n34435 & n34440;
  assign n34442 = ~n34350 & ~n34441;
  assign n34443 = ~n34150 & n34442;
  assign n34444 = ~pi2761 & ~n34443;
  assign n34445 = ~n34041 & ~n34444;
  assign n34446 = ~n34036 & n34445;
  assign n34447 = ~n34033 & n34446;
  assign n34448 = ~n33930 & n34447;
  assign n34449 = n33827 & ~n34448;
  assign n34450 = po3831 & n34449;
  assign n34451 = n33826 & n34450;
  assign po0678 = n33825 | n34451;
  assign n34453 = ~n33397 & ~n33813;
  assign n34454 = pi0858 & n33816;
  assign n34455 = pi0405 & ~n33816;
  assign n34456 = ~n34454 & ~n34455;
  assign n34457 = n33813 & ~n34456;
  assign po0679 = n34453 | n34457;
  assign n34459 = ~n33463 & ~n33813;
  assign n34460 = pi0730 & n33816;
  assign n34461 = pi0406 & ~n33816;
  assign n34462 = ~n34460 & ~n34461;
  assign n34463 = n33813 & ~n34462;
  assign po0680 = n34459 | n34463;
  assign n34465 = ~n33690 & ~n33813;
  assign n34466 = ~pi1052 & n33816;
  assign n34467 = ~pi0407 & ~n33816;
  assign n34468 = ~n34466 & ~n34467;
  assign n34469 = n33813 & ~n34468;
  assign po0681 = n34465 | n34469;
  assign n34471 = ~n33603 & ~n33813;
  assign n34472 = ~pi1045 & n33816;
  assign n34473 = pi0408 & ~n33816;
  assign n34474 = ~n34472 & ~n34473;
  assign n34475 = n33813 & ~n34474;
  assign po0682 = n34471 | n34475;
  assign n34477 = ~n33475 & ~n33813;
  assign n34478 = pi0851 & n33816;
  assign n34479 = pi0409 & ~n33816;
  assign n34480 = ~n34478 & ~n34479;
  assign n34481 = n33813 & ~n34480;
  assign po0683 = n34477 | n34481;
  assign n34483 = ~n33487 & ~n33813;
  assign n34484 = pi0860 & n33816;
  assign n34485 = pi0410 & ~n33816;
  assign n34486 = ~n34484 & ~n34485;
  assign n34487 = n33813 & ~n34486;
  assign po0684 = n34483 | n34487;
  assign n34489 = ~n33516 & ~n33813;
  assign n34490 = pi0852 & n33816;
  assign n34491 = pi0411 & ~n33816;
  assign n34492 = ~n34490 & ~n34491;
  assign n34493 = n33813 & ~n34492;
  assign po0685 = n34489 | n34493;
  assign n34495 = ~n33545 & ~n33813;
  assign n34496 = pi0821 & n33816;
  assign n34497 = pi0412 & ~n33816;
  assign n34498 = ~n34496 & ~n34497;
  assign n34499 = n33813 & ~n34498;
  assign po0686 = n34495 | n34499;
  assign n34501 = ~n33574 & ~n33813;
  assign n34502 = ~pi0937 & n33816;
  assign n34503 = pi0413 & ~n33816;
  assign n34504 = ~n34502 & ~n34503;
  assign n34505 = n33813 & ~n34504;
  assign po0687 = n34501 | n34505;
  assign n34507 = ~n33632 & ~n33813;
  assign n34508 = ~pi1082 & n33816;
  assign n34509 = pi0414 & ~n33816;
  assign n34510 = ~n34508 & ~n34509;
  assign n34511 = n33813 & ~n34510;
  assign po0688 = n34507 | n34511;
  assign n34513 = ~n33661 & ~n33813;
  assign n34514 = ~pi1080 & n33816;
  assign n34515 = pi0415 & ~n33816;
  assign n34516 = ~n34514 & ~n34515;
  assign n34517 = n33813 & ~n34516;
  assign po0689 = n34513 | n34517;
  assign n34519 = ~n33442 & ~n33813;
  assign n34520 = pi0853 & n33816;
  assign n34521 = pi0416 & ~n33816;
  assign n34522 = ~n34520 & ~n34521;
  assign n34523 = n33813 & ~n34522;
  assign po0690 = n34519 | n34523;
  assign n34525 = ~n33451 & ~n33813;
  assign n34526 = pi0854 & n33816;
  assign n34527 = pi0417 & ~n33816;
  assign n34528 = ~n34526 & ~n34527;
  assign n34529 = n33813 & ~n34528;
  assign po0691 = n34525 | n34529;
  assign n34531 = ~n33361 & ~n33813;
  assign n34532 = pi0825 & n33816;
  assign n34533 = pi0418 & ~n33816;
  assign n34534 = ~n34532 & ~n34533;
  assign n34535 = n33813 & ~n34534;
  assign po0692 = n34531 | n34535;
  assign n34537 = ~n33370 & ~n33813;
  assign n34538 = pi0855 & n33816;
  assign n34539 = pi0419 & ~n33816;
  assign n34540 = ~n34538 & ~n34539;
  assign n34541 = n33813 & ~n34540;
  assign po0693 = n34537 | n34541;
  assign n34543 = ~n33379 & ~n33813;
  assign n34544 = pi0856 & n33816;
  assign n34545 = pi0420 & ~n33816;
  assign n34546 = ~n34544 & ~n34545;
  assign n34547 = n33813 & ~n34546;
  assign po0694 = n34543 | n34547;
  assign n34549 = ~n33388 & ~n33813;
  assign n34550 = pi0857 & n33816;
  assign n34551 = pi0421 & ~n33816;
  assign n34552 = ~n34550 & ~n34551;
  assign n34553 = n33813 & ~n34552;
  assign po0695 = n34549 | n34553;
  assign n34555 = ~n33409 & ~n33813;
  assign n34556 = pi0824 & n33816;
  assign n34557 = pi0422 & ~n33816;
  assign n34558 = ~n34556 & ~n34557;
  assign n34559 = n33813 & ~n34558;
  assign po0696 = n34555 | n34559;
  assign n34561 = ~n33421 & ~n33813;
  assign n34562 = pi0823 & n33816;
  assign n34563 = pi0423 & ~n33816;
  assign n34564 = ~n34562 & ~n34563;
  assign n34565 = n33813 & ~n34564;
  assign po0697 = n34561 | n34565;
  assign n34567 = ~n33433 & ~n33813;
  assign n34568 = pi0859 & n33816;
  assign n34569 = pi0424 & ~n33816;
  assign n34570 = ~n34568 & ~n34569;
  assign n34571 = n33813 & ~n34570;
  assign po0698 = n34567 | n34571;
  assign n34573 = ~n33702 & ~n33813;
  assign n34574 = pi0731 & n33816;
  assign n34575 = pi0425 & ~n33816;
  assign n34576 = ~n34574 & ~n34575;
  assign n34577 = n33813 & ~n34576;
  assign po0699 = n34573 | n34577;
  assign n34579 = ~n33714 & ~n33813;
  assign n34580 = pi0938 & n33816;
  assign n34581 = pi0426 & ~n33816;
  assign n34582 = ~n34580 & ~n34581;
  assign n34583 = n33813 & ~n34582;
  assign po0700 = n34579 | n34583;
  assign n34585 = ~n33743 & ~n33813;
  assign n34586 = ~pi0911 & n33816;
  assign n34587 = ~pi0427 & ~n33816;
  assign n34588 = ~n34586 & ~n34587;
  assign n34589 = n33813 & ~n34588;
  assign po0701 = n34585 | n34589;
  assign n34591 = pi0975 & ~n32782;
  assign n34592 = ~pi0975 & ~n32788;
  assign n34593 = ~n34591 & ~n34592;
  assign n34594 = ~pi1771 & ~pi3580;
  assign n34595 = pi3581 & n34594;
  assign n34596 = n34593 & ~n34595;
  assign n34597 = ~pi1422 & n34596;
  assign n34598 = pi0428 & ~n34597;
  assign n34599 = n32792 & ~n33542;
  assign n34600 = ~n32942 & ~n34599;
  assign n34601 = ~n8593 & n34597;
  assign n34602 = ~n34600 & n34601;
  assign po0702 = n34598 | n34602;
  assign n34604 = pi0429 & ~n34597;
  assign n34605 = n32792 & ~n33571;
  assign n34606 = ~n32971 & ~n34605;
  assign n34607 = n34601 & ~n34606;
  assign po0703 = n34604 | n34607;
  assign n34609 = pi0430 & ~n34597;
  assign n34610 = n32792 & ~n33600;
  assign n34611 = ~n33000 & ~n34610;
  assign n34612 = n34601 & ~n34611;
  assign po0704 = n34609 | n34612;
  assign n34614 = pi0431 & ~n34597;
  assign n34615 = n32792 & ~n33629;
  assign n34616 = ~n33029 & ~n34615;
  assign n34617 = n34601 & ~n34616;
  assign po0705 = n34614 | n34617;
  assign n34619 = pi0432 & ~n34597;
  assign n34620 = n32792 & ~n33658;
  assign n34621 = ~n33058 & ~n34620;
  assign n34622 = n34601 & ~n34621;
  assign po0706 = n34619 | n34622;
  assign n34624 = pi0433 & ~n34597;
  assign n34625 = n32792 & ~n33687;
  assign n34626 = ~n33087 & ~n34625;
  assign n34627 = n34601 & ~n34626;
  assign po0707 = n34624 | n34627;
  assign n34629 = pi0434 & ~n34597;
  assign n34630 = n32792 & ~n33740;
  assign n34631 = ~n33290 & ~n34630;
  assign n34632 = n34601 & ~n34631;
  assign po0708 = n34629 | n34632;
  assign n34634 = pi0435 & ~n34597;
  assign n34635 = n32792 & ~n33513;
  assign n34636 = ~n32913 & ~n34635;
  assign n34637 = n34601 & ~n34636;
  assign po0709 = n34634 | n34637;
  assign n34639 = ~n25761 & ~n30537;
  assign n34640 = n30031 & n30537;
  assign n34641 = ~n34639 & ~n34640;
  assign n34642 = n31948 & ~n34641;
  assign n34643 = ~pi0436 & ~n31948;
  assign po0710 = n34642 | n34643;
  assign n34645 = n31955 & ~n34641;
  assign n34646 = ~pi0437 & ~n31955;
  assign po0711 = n34645 | n34646;
  assign n34648 = pi3419 & ~n12726;
  assign n34649 = n10773 & n34648;
  assign n34650 = ~pi0438 & ~pi3419;
  assign n34651 = ~n34649 & ~n34650;
  assign n34652 = n8586 & ~n16568;
  assign n34653 = pi3099 & n16211;
  assign n34654 = n8578 & n34653;
  assign n34655 = ~n33085 & n34654;
  assign n34656 = ~n34652 & ~n34655;
  assign n34657 = pi3419 & ~n34656;
  assign po0712 = ~n34651 | n34657;
  assign n34659 = pi3419 & ~n13701;
  assign n34660 = n10773 & n34659;
  assign n34661 = ~pi0439 & ~pi3419;
  assign n34662 = ~n34660 & ~n34661;
  assign n34663 = n8586 & ~n16529;
  assign n34664 = ~n33288 & n34654;
  assign n34665 = ~n34663 & ~n34664;
  assign n34666 = pi3419 & ~n34665;
  assign po0713 = ~n34662 | n34666;
  assign n34668 = ~n33513 & n34654;
  assign n34669 = n10773 & ~n13121;
  assign n34670 = ~n34668 & ~n34669;
  assign n34671 = pi3419 & ~n34670;
  assign n34672 = ~pi0440 & ~pi3419;
  assign po0714 = n34671 | n34672;
  assign n34674 = ~n33542 & n34654;
  assign n34675 = n10773 & ~n13398;
  assign n34676 = ~n34674 & ~n34675;
  assign n34677 = pi3419 & ~n34676;
  assign n34678 = ~pi0441 & ~pi3419;
  assign po0715 = n34677 | n34678;
  assign n34680 = ~n33571 & n34654;
  assign n34681 = n10773 & ~n13988;
  assign n34682 = ~n34680 & ~n34681;
  assign n34683 = pi3419 & ~n34682;
  assign n34684 = ~pi0442 & ~pi3419;
  assign po0716 = n34683 | n34684;
  assign n34686 = ~n33600 & n34654;
  assign n34687 = n10773 & ~n12415;
  assign n34688 = ~n34686 & ~n34687;
  assign n34689 = pi3419 & ~n34688;
  assign n34690 = ~pi0443 & ~pi3419;
  assign po0717 = n34689 | n34690;
  assign n34692 = ~n33629 & n34654;
  assign n34693 = n10773 & ~n14816;
  assign n34694 = ~n34692 & ~n34693;
  assign n34695 = pi3419 & ~n34694;
  assign n34696 = ~pi0444 & ~pi3419;
  assign po0718 = n34695 | n34696;
  assign n34698 = ~n33115 & n34654;
  assign n34699 = n8586 & ~n17397;
  assign n34700 = ~n34698 & ~n34699;
  assign n34701 = pi3419 & ~n34700;
  assign n34702 = ~pi0445 & ~pi3419;
  assign po0719 = n34701 | n34702;
  assign n34704 = ~n33144 & n34654;
  assign n34705 = n8586 & ~n17105;
  assign n34706 = ~n34704 & ~n34705;
  assign n34707 = pi3419 & ~n34706;
  assign n34708 = ~pi0446 & ~pi3419;
  assign po0720 = n34707 | n34708;
  assign n34710 = ~n33172 & n34654;
  assign n34711 = n8586 & ~n16999;
  assign n34712 = ~n34710 & ~n34711;
  assign n34713 = pi3419 & ~n34712;
  assign n34714 = ~pi0447 & ~pi3419;
  assign po0721 = n34713 | n34714;
  assign n34716 = ~n33201 & n34654;
  assign n34717 = n8586 & ~n16963;
  assign n34718 = ~n34716 & ~n34717;
  assign n34719 = pi3419 & ~n34718;
  assign n34720 = ~pi0448 & ~pi3419;
  assign po0722 = n34719 | n34720;
  assign n34722 = ~n33687 & n34654;
  assign n34723 = n10773 & ~n12061;
  assign n34724 = ~n34722 & ~n34723;
  assign n34725 = pi3419 & ~n34724;
  assign n34726 = ~pi0449 & ~pi3419;
  assign po0723 = n34725 | n34726;
  assign n34728 = ~n33230 & n34654;
  assign n34729 = n8586 & ~n16927;
  assign n34730 = ~n34728 & ~n34729;
  assign n34731 = pi3419 & ~n34730;
  assign n34732 = ~pi0450 & ~pi3419;
  assign po0724 = n34731 | n34732;
  assign n34734 = ~n33259 & n34654;
  assign n34735 = n8586 & ~n16891;
  assign n34736 = ~n34734 & ~n34735;
  assign n34737 = pi3419 & ~n34736;
  assign n34738 = ~pi0451 & ~pi3419;
  assign po0725 = n34737 | n34738;
  assign n34740 = ~n32882 & n34654;
  assign n34741 = n8586 & ~n16819;
  assign n34742 = ~n34740 & ~n34741;
  assign n34743 = pi3419 & ~n34742;
  assign n34744 = ~pi0452 & ~pi3419;
  assign po0726 = n34743 | n34744;
  assign n34746 = pi3419 & ~n17368;
  assign n34747 = n10773 & n34746;
  assign n34748 = ~pi0453 & ~pi3419;
  assign n34749 = ~n34747 & ~n34748;
  assign n34750 = n8586 & ~n16784;
  assign n34751 = ~n32911 & n34654;
  assign n34752 = ~n34750 & ~n34751;
  assign n34753 = pi3419 & ~n34752;
  assign po0727 = ~n34749 | n34753;
  assign n34755 = pi3419 & ~n17199;
  assign n34756 = n10773 & n34755;
  assign n34757 = ~pi0454 & ~pi3419;
  assign n34758 = ~n34756 & ~n34757;
  assign n34759 = n8586 & ~n16748;
  assign n34760 = ~n32940 & n34654;
  assign n34761 = ~n34759 & ~n34760;
  assign n34762 = pi3419 & ~n34761;
  assign po0728 = ~n34758 | n34762;
  assign n34764 = pi3419 & ~n10608;
  assign n34765 = n10773 & n34764;
  assign n34766 = ~pi0455 & ~pi3419;
  assign n34767 = ~n34765 & ~n34766;
  assign n34768 = n8586 & ~n16676;
  assign n34769 = ~n32998 & n34654;
  assign n34770 = ~n34768 & ~n34769;
  assign n34771 = pi3419 & ~n34770;
  assign po0729 = ~n34767 | n34771;
  assign n34773 = pi3419 & ~n15426;
  assign n34774 = n10773 & n34773;
  assign n34775 = ~pi0456 & ~pi3419;
  assign n34776 = ~n34774 & ~n34775;
  assign n34777 = n8586 & ~n16640;
  assign n34778 = ~n33027 & n34654;
  assign n34779 = ~n34777 & ~n34778;
  assign n34780 = pi3419 & ~n34779;
  assign po0730 = ~n34776 | n34780;
  assign n34782 = pi3419 & ~n14403;
  assign n34783 = n10773 & n34782;
  assign n34784 = ~pi0457 & ~pi3419;
  assign n34785 = ~n34783 & ~n34784;
  assign n34786 = n8586 & ~n16604;
  assign n34787 = ~n33056 & n34654;
  assign n34788 = ~n34786 & ~n34787;
  assign n34789 = pi3419 & ~n34788;
  assign po0731 = ~n34785 | n34789;
  assign n34791 = pi3641 & ~n31822;
  assign n34792 = pi0458 & ~pi3641;
  assign n34793 = ~n34791 & ~n34792;
  assign n34794 = n31865 & ~n34793;
  assign n34795 = pi0458 & ~n31865;
  assign n34796 = ~n34794 & ~n34795;
  assign n34797 = ~n31777 & ~n34796;
  assign n34798 = pi1878 & n31777;
  assign n34799 = ~n34797 & ~n34798;
  assign n34800 = ~n31779 & ~n34799;
  assign n34801 = ~pi2091 & n31779;
  assign po0732 = n34800 | n34801;
  assign n34803 = ~n33658 & n34654;
  assign n34804 = n10773 & ~n15115;
  assign n34805 = ~n34803 & ~n34804;
  assign n34806 = pi3419 & ~n34805;
  assign n34807 = ~pi0459 & ~pi3419;
  assign po0733 = n34806 | n34807;
  assign n34809 = ~n33740 & n34654;
  assign n34810 = n10773 & ~n11181;
  assign n34811 = ~n34809 & ~n34810;
  assign n34812 = pi3419 & ~n34811;
  assign n34813 = ~pi0460 & ~pi3419;
  assign po0734 = n34812 | n34813;
  assign n34815 = pi3419 & ~n9825;
  assign n34816 = n10773 & n34815;
  assign n34817 = ~pi0461 & ~pi3419;
  assign n34818 = ~n34816 & ~n34817;
  assign n34819 = n8586 & ~n16712;
  assign n34820 = ~n32969 & n34654;
  assign n34821 = ~n34819 & ~n34820;
  assign n34822 = pi3419 & ~n34821;
  assign po0735 = ~n34818 | n34822;
  assign n34824 = ~n32853 & n34654;
  assign n34825 = n8586 & ~n16855;
  assign n34826 = ~n34824 & ~n34825;
  assign n34827 = pi3419 & ~n34826;
  assign n34828 = ~pi0462 & ~pi3419;
  assign po0736 = n34827 | n34828;
  assign n34830 = ~pi0463 & ~n31948;
  assign n34831 = ~n30031 & ~n30537;
  assign n34832 = n17234 & n30537;
  assign n34833 = ~n34831 & ~n34832;
  assign n34834 = n31948 & n34833;
  assign po0737 = n34830 | n34834;
  assign n34836 = ~pi0464 & ~n31955;
  assign n34837 = n31955 & n34833;
  assign po0738 = n34836 | n34837;
  assign n34839 = pi0887 & pi1739;
  assign n34840 = ~pi0888 & pi3667;
  assign n34841 = pi0888 & ~pi3667;
  assign n34842 = ~n34840 & ~n34841;
  assign n34843 = ~pi0887 & ~n34842;
  assign po0739 = ~n34839 & ~n34843;
  assign n34845 = pi0525 & pi0527;
  assign n34846 = pi0526 & n34845;
  assign n34847 = pi0554 & n34846;
  assign n34848 = pi0531 & n34847;
  assign n34849 = ~pi0791 & ~pi0889;
  assign n34850 = pi3249 & pi3647;
  assign n34851 = ~pi0790 & pi3670;
  assign n34852 = pi0790 & po0036;
  assign n34853 = ~n34851 & ~n34852;
  assign n34854 = pi0881 & ~n34853;
  assign n34855 = ~pi0881 & n34853;
  assign po3569 = ~n34854 & ~n34855;
  assign po2701 = n34850 & po3569;
  assign n34858 = n34849 & po2701;
  assign n34859 = pi0791 & ~pi0889;
  assign n34860 = ~pi2387 & n34859;
  assign n34861 = ~pi0791 & pi0889;
  assign n34862 = pi3550 & n34861;
  assign n34863 = pi3493 & ~n34861;
  assign n34864 = ~n34862 & ~n34863;
  assign n34865 = ~n34859 & ~n34864;
  assign n34866 = ~n34860 & ~n34865;
  assign n34867 = ~n34849 & ~n34866;
  assign n34868 = ~n34858 & ~n34867;
  assign n34869 = ~pi0654 & n34868;
  assign n34870 = ~n34848 & ~n34869;
  assign n34871 = ~pi0474 & n34870;
  assign n34872 = pi0543 & n34871;
  assign n34873 = ~pi0882 & ~pi0883;
  assign n34874 = ~pi0543 & ~pi0696;
  assign n34875 = n34870 & n34874;
  assign n34876 = ~n34873 & n34875;
  assign n34877 = ~pi0465 & ~n34870;
  assign n34878 = ~n34876 & ~n34877;
  assign po0740 = n34872 | ~n34878;
  assign n34880 = pi0543 & n34870;
  assign n34881 = ~pi0478 & n34880;
  assign n34882 = ~pi0466 & ~n34870;
  assign n34883 = ~n34876 & ~n34882;
  assign po0741 = n34881 | ~n34883;
  assign n34885 = ~pi0466 & n34870;
  assign n34886 = pi0543 & n34885;
  assign n34887 = ~pi0467 & ~n34870;
  assign n34888 = ~n34876 & ~n34887;
  assign po0742 = n34886 | ~n34888;
  assign n34890 = ~pi0467 & n34870;
  assign n34891 = pi0543 & n34890;
  assign n34892 = ~pi0468 & ~n34870;
  assign n34893 = ~n34876 & ~n34892;
  assign po0743 = n34891 | ~n34893;
  assign n34895 = ~pi0468 & n34870;
  assign n34896 = pi0543 & n34895;
  assign n34897 = ~pi0469 & ~n34870;
  assign n34898 = ~n34876 & ~n34897;
  assign po0744 = n34896 | ~n34898;
  assign n34900 = ~pi0469 & n34870;
  assign n34901 = pi0543 & n34900;
  assign n34902 = ~pi0470 & ~n34870;
  assign n34903 = ~n34876 & ~n34902;
  assign po0745 = n34901 | ~n34903;
  assign n34905 = ~pi0470 & n34870;
  assign n34906 = pi0543 & n34905;
  assign n34907 = ~pi0471 & ~n34870;
  assign n34908 = ~n34876 & ~n34907;
  assign po0746 = n34906 | ~n34908;
  assign n34910 = ~pi0697 & n34870;
  assign n34911 = pi0543 & n34910;
  assign n34912 = ~pi0472 & ~n34870;
  assign n34913 = ~n34876 & ~n34912;
  assign po0747 = n34911 | ~n34913;
  assign n34915 = ~pi0472 & n34870;
  assign n34916 = pi0543 & n34915;
  assign n34917 = ~pi0473 & ~n34870;
  assign n34918 = ~n34876 & ~n34917;
  assign po0748 = n34916 | ~n34918;
  assign n34920 = ~pi0473 & n34870;
  assign n34921 = pi0543 & n34920;
  assign n34922 = ~pi0474 & ~n34870;
  assign n34923 = ~n34876 & ~n34922;
  assign po0749 = n34921 | ~n34923;
  assign n34925 = ~pi0465 & n34870;
  assign n34926 = pi0543 & n34925;
  assign n34927 = ~pi0475 & ~n34870;
  assign n34928 = ~n34876 & ~n34927;
  assign po0750 = n34926 | ~n34928;
  assign n34930 = ~pi0475 & n34870;
  assign n34931 = pi0543 & n34930;
  assign n34932 = ~pi0476 & ~n34870;
  assign n34933 = ~n34876 & ~n34932;
  assign po0751 = n34931 | ~n34933;
  assign n34935 = ~pi0476 & n34870;
  assign n34936 = pi0543 & n34935;
  assign n34937 = ~pi0477 & ~n34870;
  assign n34938 = ~n34876 & ~n34937;
  assign po0752 = n34936 | ~n34938;
  assign n34940 = ~pi0477 & n34880;
  assign n34941 = ~pi0478 & ~n34870;
  assign n34942 = ~n34876 & ~n34941;
  assign po0753 = n34940 | ~n34942;
  assign n34944 = pi0479 & n31016;
  assign n34945 = pi2599 & ~n11181;
  assign n34946 = pi0955 & ~n31311;
  assign n34947 = pi0479 & ~pi0955;
  assign n34948 = ~n34946 & ~n34947;
  assign n34949 = ~pi2599 & ~n34948;
  assign n34950 = ~n34945 & ~n34949;
  assign n34951 = ~n31013 & ~n34950;
  assign n34952 = ~pi0693 & n31013;
  assign n34953 = ~n34951 & ~n34952;
  assign n34954 = ~n31016 & ~n34953;
  assign po0754 = n34944 | n34954;
  assign n34956 = pi0712 & n31497;
  assign n34957 = ~pi0712 & ~n24256;
  assign n34958 = ~n34956 & ~n34957;
  assign n34959 = n32628 & ~n34958;
  assign n34960 = pi0480 & ~n32628;
  assign po0755 = n34959 | n34960;
  assign n34962 = n32635 & ~n34958;
  assign n34963 = pi0481 & ~n32635;
  assign po0756 = n34962 | n34963;
  assign n34965 = pi0832 & pi0921;
  assign n34966 = pi2763 & pi3394;
  assign n34967 = ~pi3330 & n34966;
  assign n34968 = pi3398 & n34967;
  assign n34969 = pi3392 & n34968;
  assign n34970 = pi0482 & n34969;
  assign n34971 = n24380 & n24391;
  assign n34972 = n16000 & n34971;
  assign n34973 = ~n34970 & ~n34972;
  assign n34974 = ~pi2487 & pi3392;
  assign n34975 = n34973 & ~n34974;
  assign n34976 = pi0615 & ~n34975;
  assign n34977 = pi0616 & pi0647;
  assign n34978 = ~pi1821 & n34977;
  assign n34979 = ~pi0616 & ~pi0647;
  assign n34980 = ~pi1810 & n34979;
  assign n34981 = ~n34978 & ~n34980;
  assign n34982 = ~pi0616 & pi0647;
  assign n34983 = ~pi1665 & n34982;
  assign n34984 = pi0616 & ~pi0647;
  assign n34985 = ~pi1657 & n34984;
  assign n34986 = ~n34983 & ~n34985;
  assign n34987 = n34981 & n34986;
  assign n34988 = n34976 & ~n34987;
  assign n34989 = ~pi0585 & ~n34976;
  assign n34990 = ~n34988 & ~n34989;
  assign n34991 = n34965 & ~n34990;
  assign n34992 = ~n11181 & ~n34965;
  assign n34993 = ~n34991 & ~n34992;
  assign n34994 = n34965 & ~n34974;
  assign n34995 = n15555 & n34971;
  assign n34996 = ~n34969 & ~n34995;
  assign n34997 = n34994 & n34996;
  assign n34998 = ~n9352 & ~n34997;
  assign n34999 = ~n34993 & n34998;
  assign n35000 = ~pi0585 & ~pi0632;
  assign n35001 = pi0585 & pi0632;
  assign n35002 = ~n35000 & ~n35001;
  assign n35003 = ~n34976 & ~n35002;
  assign n35004 = ~pi1817 & n34977;
  assign n35005 = ~pi1711 & n34979;
  assign n35006 = ~n35004 & ~n35005;
  assign n35007 = ~pi1630 & n34982;
  assign n35008 = ~pi1638 & n34984;
  assign n35009 = ~n35007 & ~n35008;
  assign n35010 = n35006 & n35009;
  assign n35011 = n34976 & ~n35010;
  assign n35012 = ~n35003 & ~n35011;
  assign n35013 = n34965 & ~n35012;
  assign n35014 = ~n12061 & ~n34965;
  assign n35015 = ~n35013 & ~n35014;
  assign n35016 = ~pi0592 & n35000;
  assign n35017 = pi0592 & ~n35000;
  assign n35018 = ~n35016 & ~n35017;
  assign n35019 = ~n34976 & ~n35018;
  assign n35020 = ~pi1816 & n34977;
  assign n35021 = ~pi1806 & n34979;
  assign n35022 = ~n35020 & ~n35021;
  assign n35023 = ~pi1662 & n34982;
  assign n35024 = ~pi1654 & n34984;
  assign n35025 = ~n35023 & ~n35024;
  assign n35026 = n35022 & n35025;
  assign n35027 = n34976 & ~n35026;
  assign n35028 = ~n35019 & ~n35027;
  assign n35029 = n34965 & ~n35028;
  assign n35030 = ~n15115 & ~n34965;
  assign n35031 = ~n35029 & ~n35030;
  assign n35032 = n9825 & ~n34965;
  assign n35033 = ~pi0594 & ~pi0595;
  assign n35034 = ~pi0590 & ~pi0593;
  assign n35035 = ~pi0591 & ~pi0603;
  assign n35036 = n35016 & n35035;
  assign n35037 = ~pi0578 & n35036;
  assign n35038 = ~pi0572 & n35037;
  assign n35039 = ~pi0571 & ~pi0602;
  assign n35040 = n35038 & n35039;
  assign n35041 = n35034 & n35040;
  assign n35042 = n35033 & n35041;
  assign n35043 = pi0573 & n35042;
  assign n35044 = ~pi0573 & ~n35042;
  assign n35045 = ~n35043 & ~n35044;
  assign n35046 = ~n34976 & ~n35045;
  assign n35047 = ~pi1818 & n34977;
  assign n35048 = ~pi1807 & n34979;
  assign n35049 = ~n35047 & ~n35048;
  assign n35050 = ~pi1655 & n34984;
  assign n35051 = n35049 & ~n35050;
  assign n35052 = ~pi1663 & n34982;
  assign n35053 = n35051 & ~n35052;
  assign n35054 = n34976 & n35053;
  assign n35055 = ~n35046 & ~n35054;
  assign n35056 = n34965 & ~n35055;
  assign n35057 = ~n35032 & ~n35056;
  assign n35058 = n15426 & ~n34965;
  assign n35059 = ~pi0590 & ~pi0602;
  assign n35060 = ~pi0571 & ~pi0594;
  assign n35061 = ~pi0603 & n35016;
  assign n35062 = ~pi0591 & n35061;
  assign n35063 = ~pi0572 & ~pi0578;
  assign n35064 = n35062 & n35063;
  assign n35065 = n35060 & n35064;
  assign n35066 = n35059 & n35065;
  assign n35067 = pi0595 & n35066;
  assign n35068 = ~pi0595 & ~n35066;
  assign n35069 = ~n35067 & ~n35068;
  assign n35070 = ~n34976 & ~n35069;
  assign n35071 = ~pi1819 & n34977;
  assign n35072 = ~pi1809 & n34979;
  assign n35073 = ~n35071 & ~n35072;
  assign n35074 = ~pi1656 & n34984;
  assign n35075 = n35073 & ~n35074;
  assign n35076 = ~pi1664 & n34982;
  assign n35077 = n35075 & ~n35076;
  assign n35078 = n34976 & n35077;
  assign n35079 = ~n35070 & ~n35078;
  assign n35080 = n34965 & ~n35079;
  assign n35081 = ~n35058 & ~n35080;
  assign n35082 = pi0591 & ~n35061;
  assign n35083 = ~n35062 & ~n35082;
  assign n35084 = ~n34976 & ~n35083;
  assign n35085 = ~pi1815 & n34977;
  assign n35086 = ~pi1804 & n34979;
  assign n35087 = ~n35085 & ~n35086;
  assign n35088 = ~pi1660 & n34982;
  assign n35089 = ~pi1653 & n34984;
  assign n35090 = ~n35088 & ~n35089;
  assign n35091 = n35087 & n35090;
  assign n35092 = n34976 & ~n35091;
  assign n35093 = ~n35084 & ~n35092;
  assign n35094 = n34965 & ~n35093;
  assign n35095 = ~n12415 & ~n34965;
  assign n35096 = ~n35094 & ~n35095;
  assign n35097 = ~pi0571 & ~pi0572;
  assign n35098 = ~pi0578 & n35061;
  assign n35099 = ~pi0591 & n35098;
  assign n35100 = n35059 & n35099;
  assign n35101 = n35097 & n35100;
  assign n35102 = pi0594 & n35101;
  assign n35103 = ~pi0594 & ~n35101;
  assign n35104 = ~n35102 & ~n35103;
  assign n35105 = ~n34976 & ~n35104;
  assign n35106 = ~pi1820 & n34977;
  assign n35107 = ~pi1710 & n34979;
  assign n35108 = ~n35106 & ~n35107;
  assign n35109 = ~pi1634 & n34984;
  assign n35110 = n35108 & ~n35109;
  assign n35111 = ~pi1632 & n34982;
  assign n35112 = n35110 & ~n35111;
  assign n35113 = n34976 & n35112;
  assign n35114 = ~n35105 & ~n35113;
  assign n35115 = n34965 & n35114;
  assign n35116 = ~n14403 & ~n34965;
  assign n35117 = ~n35115 & ~n35116;
  assign n35118 = ~n10608 & ~n34965;
  assign n35119 = ~pi1631 & n34982;
  assign n35120 = ~pi1808 & n34979;
  assign n35121 = ~n35119 & ~n35120;
  assign n35122 = ~pi1636 & n34984;
  assign n35123 = ~pi1859 & n34977;
  assign n35124 = ~n35122 & ~n35123;
  assign n35125 = n35121 & n35124;
  assign n35126 = n34976 & ~n35125;
  assign n35127 = n35062 & n35097;
  assign n35128 = ~pi0578 & n35127;
  assign n35129 = n35033 & n35128;
  assign n35130 = n35059 & n35129;
  assign n35131 = pi0593 & n35130;
  assign n35132 = ~pi0593 & ~n35130;
  assign n35133 = ~n35131 & ~n35132;
  assign n35134 = ~n34976 & n35133;
  assign n35135 = ~n35126 & ~n35134;
  assign n35136 = n34965 & ~n35135;
  assign n35137 = ~n35118 & ~n35136;
  assign n35138 = n35117 & n35137;
  assign n35139 = n35096 & n35138;
  assign n35140 = ~n35081 & n35139;
  assign n35141 = ~n35057 & n35140;
  assign n35142 = ~pi1814 & n34977;
  assign n35143 = ~pi1803 & n34979;
  assign n35144 = ~n35142 & ~n35143;
  assign n35145 = ~pi1659 & n34982;
  assign n35146 = ~pi1652 & n34984;
  assign n35147 = ~n35145 & ~n35146;
  assign n35148 = n35144 & n35147;
  assign n35149 = n34976 & ~n35148;
  assign n35150 = pi0572 & n35099;
  assign n35151 = ~pi0572 & ~n35099;
  assign n35152 = ~n35150 & ~n35151;
  assign n35153 = ~n34976 & n35152;
  assign n35154 = ~n35149 & ~n35153;
  assign n35155 = n34965 & ~n35154;
  assign n35156 = ~n13398 & ~n34965;
  assign n35157 = ~n35155 & ~n35156;
  assign n35158 = n13701 & ~n34965;
  assign n35159 = pi0602 & n35128;
  assign n35160 = ~pi0602 & ~n35128;
  assign n35161 = ~n35159 & ~n35160;
  assign n35162 = ~n34976 & ~n35161;
  assign n35163 = ~pi1651 & n34984;
  assign n35164 = ~pi1801 & n34979;
  assign n35165 = ~n35163 & ~n35164;
  assign n35166 = ~pi1813 & n34977;
  assign n35167 = n35165 & ~n35166;
  assign n35168 = ~pi1658 & n34982;
  assign n35169 = n35167 & ~n35168;
  assign n35170 = n34976 & n35169;
  assign n35171 = ~n35162 & ~n35170;
  assign n35172 = n34965 & ~n35171;
  assign n35173 = ~n35158 & ~n35172;
  assign n35174 = ~pi1633 & n34982;
  assign n35175 = ~pi1639 & n34984;
  assign n35176 = ~n35174 & ~n35175;
  assign n35177 = ~pi1708 & n34977;
  assign n35178 = ~pi1802 & n34979;
  assign n35179 = ~n35177 & ~n35178;
  assign n35180 = n35176 & n35179;
  assign n35181 = n34976 & ~n35180;
  assign n35182 = ~pi0571 & ~n35064;
  assign n35183 = pi0571 & n35064;
  assign n35184 = ~n35182 & ~n35183;
  assign n35185 = ~n34976 & n35184;
  assign n35186 = ~n35181 & ~n35185;
  assign n35187 = n34965 & ~n35186;
  assign n35188 = ~n13121 & ~n34965;
  assign n35189 = ~n35187 & ~n35188;
  assign n35190 = n12726 & ~n34965;
  assign n35191 = ~pi0590 & ~n35040;
  assign n35192 = pi0590 & n35040;
  assign n35193 = ~n35191 & ~n35192;
  assign n35194 = ~n34976 & ~n35193;
  assign n35195 = ~pi1650 & n34984;
  assign n35196 = ~pi1712 & n34979;
  assign n35197 = ~n35195 & ~n35196;
  assign n35198 = ~pi1812 & n34977;
  assign n35199 = n35197 & ~n35198;
  assign n35200 = ~pi1635 & n34982;
  assign n35201 = n35199 & ~n35200;
  assign n35202 = n34976 & n35201;
  assign n35203 = ~n35194 & ~n35202;
  assign n35204 = n34965 & ~n35203;
  assign n35205 = ~n35190 & ~n35204;
  assign n35206 = n35189 & ~n35205;
  assign n35207 = ~n35173 & n35206;
  assign n35208 = n35157 & n35207;
  assign n35209 = n35141 & n35208;
  assign n35210 = n35031 & n35209;
  assign n35211 = n35015 & n35210;
  assign n35212 = n34999 & n35211;
  assign n35213 = ~n13988 & ~n34965;
  assign n35214 = ~pi1709 & n34982;
  assign n35215 = ~pi1811 & n34984;
  assign n35216 = ~n35214 & ~n35215;
  assign n35217 = ~pi1864 & n34977;
  assign n35218 = ~pi1865 & n34979;
  assign n35219 = ~n35217 & ~n35218;
  assign n35220 = n35216 & n35219;
  assign n35221 = n34976 & ~n35220;
  assign n35222 = pi0578 & ~n35036;
  assign n35223 = ~n35037 & ~n35222;
  assign n35224 = ~n34976 & ~n35223;
  assign n35225 = ~n35221 & ~n35224;
  assign n35226 = n34965 & ~n35225;
  assign n35227 = ~n35213 & ~n35226;
  assign n35228 = ~n14816 & ~n34965;
  assign n35229 = pi0603 & ~n35016;
  assign n35230 = ~n35061 & ~n35229;
  assign n35231 = ~n34976 & ~n35230;
  assign n35232 = ~pi1707 & n34977;
  assign n35233 = ~pi1805 & n34979;
  assign n35234 = ~n35232 & ~n35233;
  assign n35235 = ~pi1661 & n34982;
  assign n35236 = ~pi1637 & n34984;
  assign n35237 = ~n35235 & ~n35236;
  assign n35238 = n35234 & n35237;
  assign n35239 = n34976 & ~n35238;
  assign n35240 = ~n35231 & ~n35239;
  assign n35241 = n34965 & ~n35240;
  assign n35242 = ~n35228 & ~n35241;
  assign n35243 = n35227 & n35242;
  assign n35244 = n35212 & n35243;
  assign n35245 = pi0482 & ~n34998;
  assign po0758 = n35244 | n35245;
  assign n35247 = ~n31439 & n31449;
  assign n35248 = ~n31438 & ~n35247;
  assign n35249 = ~n31445 & ~n35248;
  assign n35250 = pi0712 & ~n35249;
  assign n35251 = ~pi0712 & ~n24744;
  assign n35252 = ~n35250 & ~n35251;
  assign n35253 = n32628 & ~n35252;
  assign n35254 = pi0483 & ~n32628;
  assign po0759 = n35253 | n35254;
  assign n35256 = ~pi0712 & ~n24769;
  assign n35257 = ~n35250 & ~n35256;
  assign n35258 = n32628 & ~n35257;
  assign n35259 = pi0484 & ~n32628;
  assign po0760 = n35258 | n35259;
  assign n35261 = ~pi0712 & ~n25699;
  assign n35262 = ~n35250 & ~n35261;
  assign n35263 = n32628 & ~n35262;
  assign n35264 = pi0485 & ~n32628;
  assign po0761 = n35263 | n35264;
  assign n35266 = n32635 & ~n35252;
  assign n35267 = pi0486 & ~n32635;
  assign po0762 = n35266 | n35267;
  assign n35269 = n32635 & ~n35257;
  assign n35270 = pi0487 & ~n32635;
  assign po0763 = n35269 | n35270;
  assign n35272 = n32635 & ~n35262;
  assign n35273 = pi0488 & ~n32635;
  assign po0764 = n35272 | n35273;
  assign n35275 = ~n27714 & n31382;
  assign n35276 = pi0489 & n31381;
  assign n35277 = ~n24289 & n31384;
  assign n35278 = pi0489 & ~n31384;
  assign n35279 = ~n35277 & ~n35278;
  assign n35280 = n31388 & ~n35279;
  assign n35281 = ~n35276 & ~n35280;
  assign n35282 = ~n31391 & n35281;
  assign n35283 = ~n31382 & ~n35282;
  assign po0765 = n35275 | n35283;
  assign n35285 = ~n27714 & n31400;
  assign n35286 = pi0490 & n31399;
  assign n35287 = ~n24289 & n31402;
  assign n35288 = pi0490 & ~n31402;
  assign n35289 = ~n35287 & ~n35288;
  assign n35290 = n31406 & ~n35289;
  assign n35291 = ~n35286 & ~n35290;
  assign n35292 = ~n31409 & n35291;
  assign n35293 = ~n31400 & ~n35292;
  assign po0766 = n35285 | n35293;
  assign n35295 = pi0491 & pi3377;
  assign n35296 = pi1771 & ~pi3377;
  assign n35297 = ~pi0491 & n35296;
  assign n35298 = ~n35295 & ~n35297;
  assign n35299 = ~pi0604 & ~pi3377;
  assign n35300 = pi0491 & n35299;
  assign po0768 = ~n35298 | n35300;
  assign n35302 = pi0729 & pi2765;
  assign n35303 = ~pi0654 & n35302;
  assign n35304 = n34868 & n35303;
  assign n35305 = pi0654 & pi2765;
  assign n35306 = ~pi0729 & n35305;
  assign n35307 = pi0654 & ~pi2765;
  assign n35308 = pi0729 & n35307;
  assign n35309 = ~n35306 & ~n35308;
  assign n35310 = ~n35303 & n35309;
  assign n35311 = ~n35304 & ~n35310;
  assign n35312 = pi0498 & pi0504;
  assign n35313 = pi0497 & n35312;
  assign n35314 = pi0492 & pi0493;
  assign n35315 = n35313 & n35314;
  assign n35316 = n35306 & n35315;
  assign n35317 = pi0552 & pi0553;
  assign n35318 = pi0551 & pi0563;
  assign n35319 = n35317 & n35318;
  assign n35320 = pi0549 & pi0550;
  assign n35321 = pi0548 & n35320;
  assign n35322 = pi0547 & n35321;
  assign n35323 = n35319 & n35322;
  assign n35324 = n35316 & n35323;
  assign po0944 = ~n35311 | n35324;
  assign po3083 = n35316 & ~n35323;
  assign n35327 = ~po0944 & ~po3083;
  assign n35328 = pi0893 & ~n35327;
  assign n35329 = pi0493 & n35313;
  assign n35330 = ~pi0492 & ~n35329;
  assign n35331 = pi0492 & n35329;
  assign n35332 = ~n35330 & ~n35331;
  assign n35333 = n35327 & ~n35332;
  assign n35334 = ~n35328 & ~n35333;
  assign po0771 = pi1697 & ~n35334;
  assign n35336 = ~pi0493 & ~n35313;
  assign n35337 = ~n35329 & ~n35336;
  assign n35338 = n35327 & ~n35337;
  assign n35339 = pi0884 & ~n35327;
  assign n35340 = ~n35338 & ~n35339;
  assign po0772 = ~pi1697 | ~n35340;
  assign n35342 = ~pi0712 & ~n25718;
  assign n35343 = pi0712 & ~n31454;
  assign n35344 = ~n35342 & ~n35343;
  assign n35345 = n32628 & ~n35344;
  assign n35346 = pi0494 & ~n32628;
  assign po0773 = n35345 | n35346;
  assign n35348 = n32635 & ~n35344;
  assign n35349 = pi0495 & ~n32635;
  assign po0774 = n35348 | n35349;
  assign n35351 = pi0496 & ~n31865;
  assign n35352 = n31795 & ~n31803;
  assign n35353 = ~n31804 & ~n35352;
  assign n35354 = pi3641 & ~n35353;
  assign n35355 = pi0496 & ~pi3641;
  assign n35356 = ~n35354 & ~n35355;
  assign n35357 = n31865 & ~n35356;
  assign n35358 = ~n35351 & ~n35357;
  assign n35359 = ~n31777 & ~n35358;
  assign n35360 = pi1706 & n31777;
  assign n35361 = ~n35359 & ~n35360;
  assign n35362 = ~n31779 & ~n35361;
  assign n35363 = ~pi2398 & n31779;
  assign po0775 = n35362 | n35363;
  assign n35365 = ~pi0885 & ~n35327;
  assign n35366 = ~pi0497 & ~n35312;
  assign n35367 = ~n35313 & ~n35366;
  assign n35368 = n35327 & n35367;
  assign n35369 = ~n35365 & ~n35368;
  assign po0776 = ~pi1697 | n35369;
  assign n35371 = ~pi0741 & ~n35327;
  assign n35372 = ~pi0498 & n35327;
  assign n35373 = ~n35371 & ~n35372;
  assign po0777 = ~pi1697 | n35373;
  assign n35375 = pi0959 & pi1746;
  assign n35376 = ~pi0960 & pi3666;
  assign n35377 = pi0960 & ~pi3666;
  assign n35378 = ~n35376 & ~n35377;
  assign n35379 = ~pi0959 & ~n35378;
  assign po0896 = ~n35375 & ~n35379;
  assign n35381 = pi0502 & pi0503;
  assign n35382 = pi0501 & n35381;
  assign n35383 = pi0500 & n35382;
  assign n35384 = ~pi0499 & n35383;
  assign n35385 = pi0499 & ~n35383;
  assign n35386 = ~n35384 & ~n35385;
  assign n35387 = ~pi0899 & ~pi0961;
  assign n35388 = pi3251 & pi3635;
  assign n35389 = ~pi0941 & pi3668;
  assign n35390 = pi0941 & po0032;
  assign n35391 = ~n35389 & ~n35390;
  assign n35392 = pi0954 & ~n35391;
  assign n35393 = ~pi0954 & n35391;
  assign po3571 = ~n35392 & ~n35393;
  assign po2713 = n35388 & po3571;
  assign n35396 = n35387 & po2713;
  assign n35397 = pi0899 & ~pi0961;
  assign n35398 = ~pi2399 & n35397;
  assign n35399 = ~pi0899 & pi0961;
  assign n35400 = pi3549 & n35399;
  assign n35401 = pi3480 & ~n35399;
  assign n35402 = ~n35400 & ~n35401;
  assign n35403 = ~n35397 & ~n35402;
  assign n35404 = ~n35398 & ~n35403;
  assign n35405 = ~n35387 & ~n35404;
  assign n35406 = ~n35396 & ~n35405;
  assign n35407 = ~pi0655 & pi2521;
  assign n35408 = pi0700 & n35407;
  assign n35409 = n35406 & n35408;
  assign n35410 = pi0655 & pi2521;
  assign n35411 = ~pi0700 & n35410;
  assign n35412 = pi0655 & ~pi2521;
  assign n35413 = pi0700 & n35412;
  assign n35414 = ~n35411 & ~n35413;
  assign n35415 = ~n35408 & n35414;
  assign n35416 = ~n35409 & ~n35415;
  assign n35417 = pi0499 & pi0500;
  assign n35418 = n35382 & n35417;
  assign n35419 = n35411 & n35418;
  assign n35420 = pi0561 & pi0564;
  assign n35421 = pi0560 & n35420;
  assign n35422 = pi0559 & n35421;
  assign n35423 = pi0557 & pi0558;
  assign n35424 = pi0556 & n35423;
  assign n35425 = pi0555 & n35424;
  assign n35426 = n35422 & n35425;
  assign n35427 = n35419 & n35426;
  assign po0945 = ~n35416 | n35427;
  assign po2836 = n35419 & ~n35426;
  assign n35430 = ~po0945 & ~po2836;
  assign n35431 = ~n35386 & n35430;
  assign n35432 = ~pi0799 & ~n35430;
  assign n35433 = ~n35431 & ~n35432;
  assign po0780 = pi1696 & n35433;
  assign n35435 = ~pi0500 & ~n35382;
  assign n35436 = ~n35383 & ~n35435;
  assign n35437 = n35430 & n35436;
  assign n35438 = ~pi0957 & ~n35430;
  assign n35439 = ~n35437 & ~n35438;
  assign po0781 = ~pi1696 | n35439;
  assign n35441 = ~pi0501 & ~n35381;
  assign n35442 = ~n35382 & ~n35441;
  assign n35443 = n35430 & n35442;
  assign n35444 = ~pi1009 & ~n35430;
  assign n35445 = ~n35443 & ~n35444;
  assign po0782 = ~pi1696 | n35445;
  assign n35447 = ~pi0502 & ~pi0503;
  assign n35448 = ~n35381 & ~n35447;
  assign n35449 = n35430 & n35448;
  assign n35450 = ~pi0793 & ~n35430;
  assign n35451 = ~n35449 & ~n35450;
  assign po0783 = ~pi1696 | n35451;
  assign n35453 = ~pi0503 & n35430;
  assign n35454 = ~pi0795 & ~n35430;
  assign n35455 = ~n35453 & ~n35454;
  assign po0784 = ~pi1696 | n35455;
  assign n35457 = ~pi0739 & ~n35327;
  assign n35458 = ~pi0498 & ~pi0504;
  assign n35459 = ~n35312 & ~n35458;
  assign n35460 = n35327 & n35459;
  assign n35461 = ~n35457 & ~n35460;
  assign po0785 = ~pi1697 | n35461;
  assign n35463 = ~pi1011 & n9365;
  assign n35464 = pi0408 & n8615;
  assign n35465 = ~pi0427 & ~n8615;
  assign n35466 = ~n35464 & ~n35465;
  assign n35467 = n9424 & ~n35466;
  assign n35468 = pi1734 & n9419;
  assign n35469 = pi1729 & n9420;
  assign n35470 = pi1443 & n9422;
  assign n35471 = ~n35469 & ~n35470;
  assign n35472 = ~n35468 & n35471;
  assign n35473 = pi1438 & n8568;
  assign n35474 = n35472 & ~n35473;
  assign n35475 = ~n9424 & ~n35474;
  assign n35476 = ~n35467 & ~n35475;
  assign n35477 = ~po3855 & ~n35476;
  assign n35478 = ~pi3244 & po3855;
  assign n35479 = ~n35477 & ~n35478;
  assign n35480 = pi0413 & n8615;
  assign n35481 = ~pi0407 & ~n8615;
  assign n35482 = ~n35480 & ~n35481;
  assign n35483 = n9424 & ~n35482;
  assign n35484 = pi1437 & n8568;
  assign n35485 = pi1733 & n9419;
  assign n35486 = ~n35484 & ~n35485;
  assign n35487 = pi1442 & n9422;
  assign n35488 = n35486 & ~n35487;
  assign n35489 = pi1728 & n9420;
  assign n35490 = n35488 & ~n35489;
  assign n35491 = ~n9424 & ~n35490;
  assign n35492 = ~n35483 & ~n35491;
  assign n35493 = ~po3855 & ~n35492;
  assign n35494 = ~pi3292 & po3855;
  assign n35495 = ~n35493 & ~n35494;
  assign n35496 = ~n35479 & n35495;
  assign n35497 = ~n35463 & n35496;
  assign n35498 = pi2232 & n35497;
  assign n35499 = ~pi0983 & n9365;
  assign n35500 = n35479 & ~n35495;
  assign n35501 = ~n35499 & n35500;
  assign n35502 = pi2218 & n35501;
  assign n35503 = n35479 & ~n35499;
  assign n35504 = ~pi1050 & n9365;
  assign n35505 = ~n35479 & ~n35504;
  assign n35506 = ~n35503 & ~n35505;
  assign n35507 = ~n35495 & n35506;
  assign n35508 = ~n13398 & n35507;
  assign n35509 = ~n35502 & ~n35508;
  assign n35510 = ~n35479 & ~n35495;
  assign n35511 = ~n35504 & n35510;
  assign n35512 = pi2204 & n35511;
  assign n35513 = n35509 & ~n35512;
  assign n35514 = ~pi0984 & n9365;
  assign n35515 = n35479 & n35514;
  assign n35516 = n35463 & ~n35479;
  assign n35517 = ~n35515 & ~n35516;
  assign n35518 = n35495 & ~n35517;
  assign n35519 = ~n13398 & n35518;
  assign n35520 = n35513 & ~n35519;
  assign n35521 = n35479 & n35495;
  assign n35522 = ~n35514 & n35521;
  assign n35523 = pi2246 & n35522;
  assign n35524 = n35520 & ~n35523;
  assign n35525 = ~n35498 & n35524;
  assign n35526 = ~n9426 & ~po3855;
  assign n35527 = ~n8615 & ~n8619;
  assign n35528 = ~n8612 & ~n10807;
  assign n35529 = n35527 & n35528;
  assign n35530 = ~pi0405 & ~pi0420;
  assign n35531 = pi0419 & pi0421;
  assign n35532 = n35530 & n35531;
  assign n35533 = n9373 & n35532;
  assign n35534 = pi0408 & n35533;
  assign n35535 = ~n10811 & ~n35534;
  assign n35536 = ~n10808 & n35535;
  assign n35537 = n35529 & n35536;
  assign n35538 = ~n8561 & ~n35537;
  assign n35539 = n35526 & ~n35538;
  assign n35540 = ~n35525 & ~n35539;
  assign n35541 = pi0505 & n35539;
  assign po0787 = n35540 | n35541;
  assign n35543 = pi2233 & n35497;
  assign n35544 = pi2219 & n35501;
  assign n35545 = ~n13988 & n35507;
  assign n35546 = ~n35544 & ~n35545;
  assign n35547 = pi2205 & n35511;
  assign n35548 = n35546 & ~n35547;
  assign n35549 = ~n13988 & n35518;
  assign n35550 = n35548 & ~n35549;
  assign n35551 = pi2247 & n35522;
  assign n35552 = n35550 & ~n35551;
  assign n35553 = ~n35543 & n35552;
  assign n35554 = ~n35539 & ~n35553;
  assign n35555 = pi0506 & n35539;
  assign po0788 = n35554 | n35555;
  assign n35557 = pi2220 & n35501;
  assign n35558 = pi2234 & n35497;
  assign n35559 = ~n12415 & n35518;
  assign n35560 = ~n35558 & ~n35559;
  assign n35561 = pi2248 & n35522;
  assign n35562 = n35560 & ~n35561;
  assign n35563 = ~n12415 & n35507;
  assign n35564 = n35562 & ~n35563;
  assign n35565 = pi2206 & n35511;
  assign n35566 = n35564 & ~n35565;
  assign n35567 = ~n35557 & n35566;
  assign n35568 = ~n35539 & ~n35567;
  assign n35569 = pi0507 & n35539;
  assign po0789 = n35568 | n35569;
  assign n35571 = pi2221 & n35501;
  assign n35572 = pi2235 & n35497;
  assign n35573 = ~n14816 & n35518;
  assign n35574 = ~n35572 & ~n35573;
  assign n35575 = pi2249 & n35522;
  assign n35576 = n35574 & ~n35575;
  assign n35577 = ~n14816 & n35507;
  assign n35578 = n35576 & ~n35577;
  assign n35579 = pi2207 & n35511;
  assign n35580 = n35578 & ~n35579;
  assign n35581 = ~n35571 & n35580;
  assign n35582 = ~n35539 & ~n35581;
  assign n35583 = pi0508 & n35539;
  assign po0790 = n35582 | n35583;
  assign n35585 = pi2222 & n35501;
  assign n35586 = pi2236 & n35497;
  assign n35587 = ~n15115 & n35507;
  assign n35588 = ~n35586 & ~n35587;
  assign n35589 = pi2250 & n35522;
  assign n35590 = n35588 & ~n35589;
  assign n35591 = ~n15115 & n35518;
  assign n35592 = n35590 & ~n35591;
  assign n35593 = pi2208 & n35511;
  assign n35594 = n35592 & ~n35593;
  assign n35595 = ~n35585 & n35594;
  assign n35596 = ~n35539 & ~n35595;
  assign n35597 = pi0509 & n35539;
  assign po0791 = n35596 | n35597;
  assign n35599 = pi2223 & n35501;
  assign n35600 = pi2237 & n35497;
  assign n35601 = ~n12061 & n35507;
  assign n35602 = ~n35600 & ~n35601;
  assign n35603 = pi2251 & n35522;
  assign n35604 = n35602 & ~n35603;
  assign n35605 = ~n12061 & n35518;
  assign n35606 = n35604 & ~n35605;
  assign n35607 = pi2209 & n35511;
  assign n35608 = n35606 & ~n35607;
  assign n35609 = ~n35599 & n35608;
  assign n35610 = ~n35539 & ~n35609;
  assign n35611 = pi0510 & n35539;
  assign po0792 = n35610 | n35611;
  assign n35613 = ~pi0407 & n9424;
  assign n35614 = ~n35491 & ~n35613;
  assign n35615 = ~po3855 & ~n35614;
  assign n35616 = ~pi3330 & po3855;
  assign n35617 = ~n35615 & ~n35616;
  assign n35618 = ~pi0427 & n9424;
  assign n35619 = ~n35475 & ~n35618;
  assign n35620 = ~po3855 & ~n35619;
  assign n35621 = ~pi3394 & po3855;
  assign n35622 = ~n35620 & ~n35621;
  assign n35623 = ~pi0985 & n9365;
  assign n35624 = n35622 & ~n35623;
  assign n35625 = ~pi0986 & n9365;
  assign n35626 = ~n35622 & ~n35625;
  assign n35627 = ~n35624 & ~n35626;
  assign n35628 = ~n35617 & n35627;
  assign n35629 = ~n12726 & n35628;
  assign n35630 = ~pi0945 & n9365;
  assign n35631 = n35617 & n35622;
  assign n35632 = ~n35630 & n35631;
  assign n35633 = pi2314 & n35632;
  assign n35634 = ~n35629 & ~n35633;
  assign n35635 = ~pi0760 & n9365;
  assign n35636 = n35617 & ~n35622;
  assign n35637 = ~n35635 & n35636;
  assign n35638 = pi2303 & n35637;
  assign n35639 = n35634 & ~n35638;
  assign n35640 = n35622 & n35630;
  assign n35641 = ~n35622 & n35635;
  assign n35642 = ~n35640 & ~n35641;
  assign n35643 = n35617 & ~n35642;
  assign n35644 = ~n12726 & n35643;
  assign n35645 = n35639 & ~n35644;
  assign n35646 = ~n35617 & n35622;
  assign n35647 = ~n35623 & n35646;
  assign n35648 = pi2292 & n35647;
  assign n35649 = ~n35617 & ~n35625;
  assign n35650 = ~n35622 & n35649;
  assign n35651 = pi2279 & n35650;
  assign n35652 = ~n35648 & ~n35651;
  assign n35653 = n35645 & n35652;
  assign n35654 = ~n8615 & ~n10794;
  assign n35655 = ~pi0408 & n35533;
  assign n35656 = ~n10791 & ~n35655;
  assign n35657 = ~n10800 & n35656;
  assign n35658 = n35654 & n35657;
  assign n35659 = ~n8561 & ~n35658;
  assign n35660 = n35526 & ~n35659;
  assign n35661 = ~n35653 & ~n35660;
  assign n35662 = pi0511 & n35660;
  assign po0794 = n35661 | n35662;
  assign n35664 = ~n13701 & n35643;
  assign n35665 = pi2315 & n35632;
  assign n35666 = ~n35664 & ~n35665;
  assign n35667 = pi2089 & n35637;
  assign n35668 = n35666 & ~n35667;
  assign n35669 = ~n13701 & n35628;
  assign n35670 = n35668 & ~n35669;
  assign n35671 = pi2067 & n35647;
  assign n35672 = pi2280 & n35650;
  assign n35673 = ~n35671 & ~n35672;
  assign n35674 = n35670 & n35673;
  assign n35675 = ~n35660 & ~n35674;
  assign n35676 = pi0512 & n35660;
  assign po0795 = n35675 | n35676;
  assign n35678 = pi2294 & n35647;
  assign n35679 = pi2317 & n35632;
  assign n35680 = ~n13398 & n35643;
  assign n35681 = ~n35679 & ~n35680;
  assign n35682 = pi2305 & n35637;
  assign n35683 = n35681 & ~n35682;
  assign n35684 = ~n13398 & n35628;
  assign n35685 = n35683 & ~n35684;
  assign n35686 = pi2282 & n35650;
  assign n35687 = n35685 & ~n35686;
  assign n35688 = ~n35678 & n35687;
  assign n35689 = ~n35660 & ~n35688;
  assign n35690 = pi0513 & n35660;
  assign po0796 = n35689 | n35690;
  assign n35692 = pi2295 & n35647;
  assign n35693 = pi2318 & n35632;
  assign n35694 = ~n13988 & n35628;
  assign n35695 = ~n35693 & ~n35694;
  assign n35696 = pi2084 & n35637;
  assign n35697 = n35695 & ~n35696;
  assign n35698 = ~n13988 & n35643;
  assign n35699 = n35697 & ~n35698;
  assign n35700 = pi2283 & n35650;
  assign n35701 = n35699 & ~n35700;
  assign n35702 = ~n35692 & n35701;
  assign n35703 = ~n35660 & ~n35702;
  assign n35704 = pi0514 & n35660;
  assign po0797 = n35703 | n35704;
  assign n35706 = pi2296 & n35647;
  assign n35707 = pi2319 & n35632;
  assign n35708 = ~n12415 & n35643;
  assign n35709 = ~n35707 & ~n35708;
  assign n35710 = pi2087 & n35637;
  assign n35711 = n35709 & ~n35710;
  assign n35712 = ~n12415 & n35628;
  assign n35713 = n35711 & ~n35712;
  assign n35714 = pi2284 & n35650;
  assign n35715 = n35713 & ~n35714;
  assign n35716 = ~n35706 & n35715;
  assign n35717 = ~n35660 & ~n35716;
  assign n35718 = pi0515 & n35660;
  assign po0798 = n35717 | n35718;
  assign n35720 = pi2321 & n35632;
  assign n35721 = pi2298 & n35647;
  assign n35722 = ~n15115 & n35628;
  assign n35723 = ~n35721 & ~n35722;
  assign n35724 = pi2286 & n35650;
  assign n35725 = n35723 & ~n35724;
  assign n35726 = ~n15115 & n35643;
  assign n35727 = n35725 & ~n35726;
  assign n35728 = pi2307 & n35637;
  assign n35729 = n35727 & ~n35728;
  assign n35730 = ~n35720 & n35729;
  assign n35731 = ~n35660 & ~n35730;
  assign n35732 = pi0516 & n35660;
  assign po0799 = n35731 | n35732;
  assign n35734 = pi2322 & n35632;
  assign n35735 = pi2299 & n35647;
  assign n35736 = ~n12061 & n35643;
  assign n35737 = ~n35735 & ~n35736;
  assign n35738 = pi2068 & n35650;
  assign n35739 = n35737 & ~n35738;
  assign n35740 = ~n12061 & n35628;
  assign n35741 = n35739 & ~n35740;
  assign n35742 = pi2308 & n35637;
  assign n35743 = n35741 & ~n35742;
  assign n35744 = ~n35734 & n35743;
  assign n35745 = ~n35660 & ~n35744;
  assign n35746 = pi0517 & n35660;
  assign po0800 = n35745 | n35746;
  assign n35748 = ~n9825 & n35643;
  assign n35749 = pi2300 & n35647;
  assign n35750 = ~n35748 & ~n35749;
  assign n35751 = pi2287 & n35650;
  assign n35752 = n35750 & ~n35751;
  assign n35753 = ~n9825 & n35628;
  assign n35754 = n35752 & ~n35753;
  assign n35755 = pi2323 & n35632;
  assign n35756 = pi2309 & n35637;
  assign n35757 = ~n35755 & ~n35756;
  assign n35758 = n35754 & n35757;
  assign n35759 = ~n35660 & ~n35758;
  assign n35760 = pi0518 & n35660;
  assign po0801 = n35759 | n35760;
  assign n35762 = ~n15426 & n35643;
  assign n35763 = pi2325 & n35632;
  assign n35764 = ~n35762 & ~n35763;
  assign n35765 = pi2311 & n35637;
  assign n35766 = n35764 & ~n35765;
  assign n35767 = ~n15426 & n35628;
  assign n35768 = n35766 & ~n35767;
  assign n35769 = pi2088 & n35647;
  assign n35770 = pi2289 & n35650;
  assign n35771 = ~n35769 & ~n35770;
  assign n35772 = n35768 & n35771;
  assign n35773 = ~n35660 & ~n35772;
  assign n35774 = pi0519 & n35660;
  assign po0802 = n35773 | n35774;
  assign n35776 = ~n14403 & n35643;
  assign n35777 = pi2301 & n35647;
  assign n35778 = ~n35776 & ~n35777;
  assign n35779 = pi2290 & n35650;
  assign n35780 = n35778 & ~n35779;
  assign n35781 = ~n14403 & n35628;
  assign n35782 = n35780 & ~n35781;
  assign n35783 = pi2326 & n35632;
  assign n35784 = pi2312 & n35637;
  assign n35785 = ~n35783 & ~n35784;
  assign n35786 = n35782 & n35785;
  assign n35787 = ~n35660 & ~n35786;
  assign n35788 = pi0520 & n35660;
  assign po0803 = n35787 | n35788;
  assign n35790 = pi2327 & n35632;
  assign n35791 = pi2302 & n35647;
  assign n35792 = ~n11181 & n35628;
  assign n35793 = ~n35791 & ~n35792;
  assign n35794 = pi2291 & n35650;
  assign n35795 = n35793 & ~n35794;
  assign n35796 = ~n11181 & n35643;
  assign n35797 = n35795 & ~n35796;
  assign n35798 = pi2313 & n35637;
  assign n35799 = n35797 & ~n35798;
  assign n35800 = ~n35790 & n35799;
  assign n35801 = ~n35660 & ~n35800;
  assign n35802 = pi0521 & n35660;
  assign po0804 = n35801 | n35802;
  assign n35804 = pi1597 & ~po3627;
  assign n35805 = pi3237 & ~n35804;
  assign n35806 = ~pi0875 & pi1444;
  assign n35807 = ~pi1444 & ~pi3300;
  assign n35808 = pi3141 & n35807;
  assign n35809 = ~n35806 & ~n35808;
  assign n35810 = pi0522 & n35809;
  assign n35811 = pi3372 & n35810;
  assign po0805 = n35805 & ~n35811;
  assign n35813 = pi0419 & n10752;
  assign n35814 = pi0419 & pi0420;
  assign n35815 = pi0421 & n35814;
  assign n35816 = n9373 & n35815;
  assign n35817 = ~pi0405 & n35816;
  assign n35818 = pi0409 & n35817;
  assign n35819 = pi0420 & n10752;
  assign n35820 = pi0410 & n35817;
  assign n35821 = ~n35819 & ~n35820;
  assign n35822 = ~n35818 & n35821;
  assign n35823 = ~n35813 & n35822;
  assign n35824 = ~n10752 & ~n24815;
  assign n35825 = n8607 & n24807;
  assign n35826 = pi0421 & n35825;
  assign n35827 = n9373 & n35826;
  assign n35828 = pi0405 & n35816;
  assign n35829 = ~n35827 & ~n35828;
  assign n35830 = ~n35817 & n35829;
  assign n35831 = n35824 & n35830;
  assign n35832 = pi0408 & n35831;
  assign n35833 = ~pi0427 & ~n35831;
  assign n35834 = ~n35832 & ~n35833;
  assign n35835 = pi0419 & n10749;
  assign n35836 = pi0418 & n10752;
  assign n35837 = ~n35817 & ~n35836;
  assign n35838 = ~n8612 & ~n10759;
  assign n35839 = ~n35827 & n35838;
  assign n35840 = pi0422 & ~n35839;
  assign n35841 = ~n35828 & ~n35840;
  assign n35842 = pi0419 & n8619;
  assign n35843 = n35841 & ~n35842;
  assign n35844 = ~n24815 & n35843;
  assign n35845 = n35837 & n35844;
  assign n35846 = ~n35835 & n35845;
  assign n35847 = ~n35834 & ~n35846;
  assign n35848 = n35823 & n35847;
  assign n35849 = pi0411 & n35831;
  assign n35850 = pi0414 & ~n35831;
  assign n35851 = ~n35849 & ~n35850;
  assign n35852 = pi0413 & n35831;
  assign n35853 = ~pi0407 & ~n35831;
  assign n35854 = ~n35852 & ~n35853;
  assign n35855 = ~pi0412 & n35831;
  assign n35856 = ~pi0415 & ~n35831;
  assign n35857 = ~n35855 & ~n35856;
  assign n35858 = n35854 & n35857;
  assign n35859 = ~n35851 & n35858;
  assign n35860 = n35848 & n35859;
  assign n35861 = ~n35854 & n35857;
  assign n35862 = ~n35846 & n35851;
  assign n35863 = n35823 & n35862;
  assign n35864 = n35834 & n35863;
  assign n35865 = n35861 & n35864;
  assign n35866 = ~n35834 & n35863;
  assign n35867 = n35861 & n35866;
  assign n35868 = n35834 & ~n35846;
  assign n35869 = n35823 & n35868;
  assign n35870 = n35851 & ~n35857;
  assign n35871 = ~n35854 & n35870;
  assign n35872 = n35869 & n35871;
  assign n35873 = n35848 & ~n35854;
  assign n35874 = n35870 & n35873;
  assign n35875 = ~n35872 & ~n35874;
  assign n35876 = ~n35867 & n35875;
  assign n35877 = ~n35865 & n35876;
  assign n35878 = n35847 & ~n35851;
  assign n35879 = ~n35854 & ~n35857;
  assign n35880 = n35823 & n35879;
  assign n35881 = n35878 & n35880;
  assign n35882 = n35877 & ~n35881;
  assign n35883 = n35859 & n35869;
  assign n35884 = n35882 & ~n35883;
  assign n35885 = ~n35860 & n35884;
  assign n35886 = ~n8612 & ~n8619;
  assign n35887 = ~n8561 & ~n35886;
  assign n35888 = ~n35885 & n35887;
  assign n35889 = pi0523 & n8561;
  assign po0807 = n35888 | n35889;
  assign n35891 = ~n8561 & n35886;
  assign n35892 = ~n35885 & n35891;
  assign n35893 = pi0524 & n8561;
  assign po0808 = n35892 | n35893;
  assign n35895 = pi0526 & pi0531;
  assign n35896 = pi0525 & n35895;
  assign n35897 = ~pi0525 & ~n35895;
  assign n35898 = ~n35896 & ~n35897;
  assign n35899 = ~n34848 & n35327;
  assign po0809 = ~n35898 & n35899;
  assign n35901 = ~pi0526 & ~pi0531;
  assign n35902 = ~n35895 & ~n35901;
  assign po0810 = n35899 & ~n35902;
  assign n35904 = ~pi0527 & n35896;
  assign n35905 = pi0527 & ~n35896;
  assign n35906 = ~n35904 & ~n35905;
  assign po0811 = n35899 & n35906;
  assign n35908 = pi0528 & pi0529;
  assign n35909 = ~pi0528 & ~pi0529;
  assign n35910 = ~n35908 & ~n35909;
  assign n35911 = pi0530 & pi0532;
  assign n35912 = pi0529 & pi0542;
  assign n35913 = pi0528 & n35912;
  assign n35914 = n35911 & n35913;
  assign n35915 = n35430 & ~n35914;
  assign po0812 = ~n35910 & n35915;
  assign po0813 = pi0529 & n35915;
  assign n35918 = pi0532 & n35908;
  assign n35919 = ~pi0530 & n35918;
  assign n35920 = pi0530 & ~n35918;
  assign n35921 = ~n35919 & ~n35920;
  assign po0814 = n35915 & n35921;
  assign po0815 = pi0531 & n35899;
  assign n35924 = ~pi0532 & ~n35908;
  assign n35925 = ~n35918 & ~n35924;
  assign po0816 = n35915 & ~n35925;
  assign n35927 = ~n12726 & n35518;
  assign n35928 = pi2215 & n35501;
  assign n35929 = ~n35927 & ~n35928;
  assign n35930 = pi2201 & n35511;
  assign n35931 = n35929 & ~n35930;
  assign n35932 = ~n12726 & n35507;
  assign n35933 = n35931 & ~n35932;
  assign n35934 = pi2229 & n35497;
  assign n35935 = pi2243 & n35522;
  assign n35936 = ~n35934 & ~n35935;
  assign n35937 = n35933 & n35936;
  assign n35938 = ~n35539 & ~n35937;
  assign n35939 = pi0533 & n35539;
  assign po0817 = n35938 | n35939;
  assign n35941 = ~n10608 & n35507;
  assign n35942 = pi2239 & n35497;
  assign n35943 = ~n35941 & ~n35942;
  assign n35944 = pi2253 & n35522;
  assign n35945 = n35943 & ~n35944;
  assign n35946 = ~n10608 & n35518;
  assign n35947 = n35945 & ~n35946;
  assign n35948 = pi2225 & n35501;
  assign n35949 = pi2211 & n35511;
  assign n35950 = ~n35948 & ~n35949;
  assign n35951 = n35947 & n35950;
  assign n35952 = ~n35539 & ~n35951;
  assign n35953 = pi0534 & n35539;
  assign po0818 = n35952 | n35953;
  assign n35955 = ~n15426 & n35518;
  assign n35956 = pi2226 & n35501;
  assign n35957 = ~n35955 & ~n35956;
  assign n35958 = pi2212 & n35511;
  assign n35959 = n35957 & ~n35958;
  assign n35960 = ~n15426 & n35507;
  assign n35961 = n35959 & ~n35960;
  assign n35962 = pi2240 & n35497;
  assign n35963 = pi2254 & n35522;
  assign n35964 = ~n35962 & ~n35963;
  assign n35965 = n35961 & n35964;
  assign n35966 = ~n35539 & ~n35965;
  assign n35967 = pi0535 & n35539;
  assign po0819 = n35966 | n35967;
  assign n35969 = ~n14403 & n35507;
  assign n35970 = pi2227 & n35501;
  assign n35971 = ~n35969 & ~n35970;
  assign n35972 = pi2213 & n35511;
  assign n35973 = n35971 & ~n35972;
  assign n35974 = ~n14403 & n35518;
  assign n35975 = n35973 & ~n35974;
  assign n35976 = pi2241 & n35497;
  assign n35977 = pi2255 & n35522;
  assign n35978 = ~n35976 & ~n35977;
  assign n35979 = n35975 & n35978;
  assign n35980 = ~n35539 & ~n35979;
  assign n35981 = pi0536 & n35539;
  assign po0820 = n35980 | n35981;
  assign n35983 = ~n35851 & n35861;
  assign n35984 = n35869 & n35983;
  assign n35985 = ~n35851 & n35854;
  assign n35986 = ~n35857 & n35985;
  assign n35987 = n35848 & n35986;
  assign n35988 = ~n35984 & ~n35987;
  assign n35989 = n35869 & n35986;
  assign n35990 = pi0420 & ~n35817;
  assign n35991 = ~n35820 & ~n35990;
  assign n35992 = ~n35837 & ~n35991;
  assign n35993 = ~pi0407 & pi0415;
  assign n35994 = ~pi0414 & n35993;
  assign n35995 = pi0419 & ~n35817;
  assign n35996 = ~n35818 & ~n35995;
  assign n35997 = pi0427 & ~n35996;
  assign n35998 = n35994 & n35997;
  assign n35999 = n35992 & n35998;
  assign n36000 = n35848 & n35983;
  assign n36001 = ~n35999 & ~n36000;
  assign n36002 = ~n35989 & n36001;
  assign n36003 = n35988 & n36002;
  assign n36004 = n35887 & ~n36003;
  assign n36005 = pi0537 & n8561;
  assign po0821 = n36004 | n36005;
  assign n36007 = n35891 & ~n36003;
  assign n36008 = pi0538 & n8561;
  assign po0822 = n36007 | n36008;
  assign n36010 = ~n35837 & n35996;
  assign n36011 = n20498 & n36010;
  assign n36012 = ~pi0414 & ~n35991;
  assign n36013 = ~pi0415 & n36012;
  assign n36014 = n36011 & n36013;
  assign n36015 = ~pi0407 & pi0427;
  assign n36016 = n36010 & n36015;
  assign n36017 = n36013 & n36016;
  assign n36018 = ~pi0415 & n36010;
  assign n36019 = pi0414 & ~n35991;
  assign n36020 = n20498 & n36019;
  assign n36021 = n36018 & n36020;
  assign n36022 = n36015 & n36019;
  assign n36023 = n36018 & n36022;
  assign n36024 = pi0415 & n36012;
  assign n36025 = n36016 & n36024;
  assign n36026 = n36011 & n36024;
  assign n36027 = pi0407 & ~pi0427;
  assign n36028 = n36010 & n36027;
  assign n36029 = n36024 & n36028;
  assign n36030 = pi0407 & pi0427;
  assign n36031 = pi0415 & n36030;
  assign n36032 = n36010 & n36012;
  assign n36033 = n36031 & n36032;
  assign n36034 = ~n36029 & ~n36033;
  assign n36035 = ~n36026 & n36034;
  assign n36036 = ~n36025 & n36035;
  assign n36037 = n36018 & n36019;
  assign n36038 = n36027 & n36037;
  assign n36039 = n36036 & ~n36038;
  assign n36040 = n36010 & n36019;
  assign n36041 = ~pi0415 & n36030;
  assign n36042 = n36040 & n36041;
  assign n36043 = n36039 & ~n36042;
  assign n36044 = ~n36023 & n36043;
  assign n36045 = ~n36021 & n36044;
  assign n36046 = ~pi0427 & ~n35996;
  assign n36047 = n35992 & n36046;
  assign n36048 = n35994 & n36047;
  assign n36049 = n36045 & ~n36048;
  assign n36050 = n36013 & n36028;
  assign n36051 = n36032 & n36041;
  assign n36052 = ~n36050 & ~n36051;
  assign n36053 = n36049 & n36052;
  assign n36054 = ~n36017 & n36053;
  assign n36055 = ~n36014 & n36054;
  assign n36056 = ~n8561 & ~n36055;
  assign n36057 = pi0539 & n8561;
  assign po0823 = n36056 | n36057;
  assign n36059 = ~n8561 & po3627;
  assign n36060 = n9345 & n36059;
  assign n36061 = ~pi0412 & n35817;
  assign n36062 = ~pi0415 & ~n35817;
  assign n36063 = ~n36061 & ~n36062;
  assign n36064 = pi0408 & n35817;
  assign n36065 = ~pi0427 & ~n35817;
  assign n36066 = ~n36064 & ~n36065;
  assign n36067 = pi0413 & n35817;
  assign n36068 = ~pi0407 & ~n35817;
  assign n36069 = ~n36067 & ~n36068;
  assign n36070 = ~n36066 & ~n36069;
  assign n36071 = n36063 & n36070;
  assign n36072 = pi0425 & n35817;
  assign n36073 = ~n35995 & ~n36072;
  assign n36074 = pi0419 & n24811;
  assign n36075 = pi0403 & n36074;
  assign n36076 = ~n10753 & ~n36075;
  assign n36077 = ~n35817 & n36076;
  assign n36078 = n36073 & ~n36077;
  assign n36079 = pi0426 & n35817;
  assign n36080 = ~n35990 & ~n36079;
  assign n36081 = pi0411 & n35817;
  assign n36082 = pi0414 & ~n35817;
  assign n36083 = ~n36081 & ~n36082;
  assign n36084 = ~n36080 & ~n36083;
  assign n36085 = n36078 & n36084;
  assign n36086 = n36071 & n36085;
  assign n36087 = ~pi0411 & ~pi0413;
  assign n36088 = ~pi0424 & n36087;
  assign n36089 = n9373 & n35531;
  assign n36090 = pi0405 & n36089;
  assign n36091 = ~pi0420 & n36090;
  assign n36092 = ~n36088 & n36091;
  assign n36093 = ~n36086 & ~n36092;
  assign n36094 = ~n36063 & n36069;
  assign n36095 = ~n36077 & ~n36080;
  assign n36096 = n36066 & ~n36073;
  assign n36097 = n36083 & n36096;
  assign n36098 = n36095 & n36097;
  assign n36099 = n36094 & n36098;
  assign n36100 = ~n36066 & ~n36073;
  assign n36101 = n36095 & n36100;
  assign n36102 = n36063 & ~n36069;
  assign n36103 = n36101 & n36102;
  assign n36104 = ~n36083 & n36103;
  assign n36105 = ~n36063 & ~n36069;
  assign n36106 = n36083 & n36101;
  assign n36107 = n36105 & n36106;
  assign n36108 = n36094 & n36106;
  assign n36109 = ~n36107 & ~n36108;
  assign n36110 = ~n36104 & n36109;
  assign n36111 = pi0419 & n8609;
  assign n36112 = pi0418 & n36111;
  assign n36113 = n35993 & n36047;
  assign n36114 = pi0414 & n36113;
  assign n36115 = pi0405 & n34038;
  assign n36116 = pi0421 & n36115;
  assign n36117 = ~n36114 & ~n36116;
  assign n36118 = ~n36112 & n36117;
  assign n36119 = n36110 & n36118;
  assign n36120 = n36066 & ~n36069;
  assign n36121 = n36063 & n36078;
  assign n36122 = n36084 & n36121;
  assign n36123 = n36120 & n36122;
  assign n36124 = n36119 & ~n36123;
  assign n36125 = ~n36099 & n36124;
  assign n36126 = n36093 & n36125;
  assign n36127 = n36060 & ~n36126;
  assign n36128 = n8561 & po3627;
  assign n36129 = pi0540 & n36128;
  assign po0824 = n36127 | n36129;
  assign n36131 = ~n24863 & n24878;
  assign n36132 = ~n24867 & n36131;
  assign n36133 = ~n24870 & n36132;
  assign n36134 = n19553 & ~n36133;
  assign n36135 = ~pi1666 & n36134;
  assign n36136 = n19553 & n24840;
  assign n36137 = ~pi1667 & n36136;
  assign n36138 = n25516 & n36137;
  assign n36139 = ~n36135 & ~n36138;
  assign n36140 = n25623 & ~n36139;
  assign n36141 = pi0541 & n8561;
  assign n36142 = ~n36140 & ~n36141;
  assign po0825 = po3627 & ~n36142;
  assign n36144 = n35908 & n35911;
  assign n36145 = ~pi0542 & n36144;
  assign n36146 = pi0542 & ~n36144;
  assign n36147 = ~n36145 & ~n36146;
  assign n36148 = ~n35914 & n36147;
  assign po0826 = ~n35430 | n36148;
  assign n36150 = ~n34868 & n35303;
  assign n36151 = n35306 & ~n35315;
  assign n36152 = ~n36150 & ~n36151;
  assign po1022 = n35308 | ~n36152;
  assign n36154 = ~po0944 & po1022;
  assign n36155 = ~n35306 & n36154;
  assign po0827 = ~po3083 & n36155;
  assign n36157 = pi2018 & ~po3627;
  assign n36158 = pi3068 & ~n36157;
  assign n36159 = pi0544 & ~pi3373;
  assign n36160 = n36158 & ~n36159;
  assign n36161 = ~pi1447 & ~pi2820;
  assign n36162 = ~pi0877 & pi1447;
  assign n36163 = ~n36161 & ~n36162;
  assign n36164 = n36158 & ~n36163;
  assign po0828 = n36160 | n36164;
  assign n36166 = pi0545 & pi3186;
  assign n36167 = ~pi0687 & ~pi0724;
  assign n36168 = ~pi0725 & ~pi0726;
  assign n36169 = n36167 & n36168;
  assign n36170 = ~pi0772 & ~pi0786;
  assign n36171 = ~pi0771 & n36170;
  assign n36172 = ~pi0782 & n36171;
  assign n36173 = n36169 & n36172;
  assign n36174 = ~po3616 & n8380;
  assign n36175 = pi3323 & n36174;
  assign n36176 = pi3324 & n8200;
  assign n36177 = n36175 & n36176;
  assign n36178 = pi3294 & n8194;
  assign n36179 = pi3322 & n36174;
  assign n36180 = n36178 & n36179;
  assign n36181 = ~n36177 & ~n36180;
  assign n36182 = pi2986 & n10770;
  assign n36183 = ~n36181 & n36182;
  assign n36184 = pi2048 & ~n36181;
  assign n36185 = ~pi2986 & n10770;
  assign n36186 = n36184 & n36185;
  assign n36187 = ~n36183 & ~n36186;
  assign n36188 = ~n8598 & ~n16213;
  assign n36189 = ~n36181 & ~n36188;
  assign n36190 = n36187 & ~n36189;
  assign n36191 = n36173 & ~n36190;
  assign n36192 = ~pi0723 & ~pi0732;
  assign n36193 = ~pi0769 & ~pi0770;
  assign n36194 = n36192 & n36193;
  assign n36195 = n36191 & n36194;
  assign n36196 = pi0787 & n36195;
  assign n36197 = ~pi0733 & n36196;
  assign n36198 = n8563 & n36197;
  assign n36199 = pi3490 & pi3544;
  assign n36200 = ~n36198 & ~n36199;
  assign n36201 = n36166 & n36200;
  assign n36202 = pi2975 & ~n36201;
  assign n36203 = pi1598 & ~po3627;
  assign po0829 = n36202 & ~n36203;
  assign n36205 = pi1049 & ~po3627;
  assign n36206 = pi2976 & ~n36205;
  assign n36207 = pi1931 & n36206;
  assign n36208 = ~pi0879 & pi1738;
  assign n36209 = ~pi1738 & ~pi3302;
  assign n36210 = ~n36208 & ~n36209;
  assign n36211 = n36207 & ~n36210;
  assign n36212 = pi1931 & ~pi3189;
  assign n36213 = pi0546 & ~n36212;
  assign n36214 = n36206 & ~n36213;
  assign po0830 = n36211 | n36214;
  assign n36216 = pi0550 & pi0563;
  assign n36217 = pi0551 & n35317;
  assign n36218 = n36216 & n36217;
  assign n36219 = pi0548 & n36218;
  assign n36220 = pi0549 & n36219;
  assign n36221 = ~pi0547 & n36220;
  assign n36222 = pi0547 & ~n36220;
  assign n36223 = ~n36221 & ~n36222;
  assign n36224 = po3083 & ~n36223;
  assign n36225 = pi0547 & ~po3083;
  assign n36226 = ~n36224 & ~n36225;
  assign n36227 = ~po0944 & n36226;
  assign n36228 = pi0948 & po0944;
  assign po0831 = n36227 | n36228;
  assign n36230 = n35319 & n35320;
  assign n36231 = pi0548 & n36230;
  assign n36232 = ~pi0548 & ~n36230;
  assign n36233 = ~n36231 & ~n36232;
  assign n36234 = po3083 & ~n36233;
  assign n36235 = ~pi0548 & ~po3083;
  assign n36236 = ~n36234 & ~n36235;
  assign n36237 = ~po0944 & ~n36236;
  assign n36238 = pi0949 & po0944;
  assign po0832 = n36237 | n36238;
  assign n36240 = pi0553 & n36216;
  assign n36241 = pi0551 & n36240;
  assign n36242 = pi0552 & n36241;
  assign n36243 = ~pi0549 & n36242;
  assign n36244 = pi0549 & ~n36242;
  assign n36245 = ~n36243 & ~n36244;
  assign n36246 = po3083 & ~n36245;
  assign n36247 = pi0549 & ~po3083;
  assign n36248 = ~n36246 & ~n36247;
  assign n36249 = ~po0944 & n36248;
  assign n36250 = pi0950 & po0944;
  assign po0833 = n36249 | n36250;
  assign n36252 = pi0563 & n36217;
  assign n36253 = ~pi0550 & ~n36252;
  assign n36254 = pi0550 & n36252;
  assign n36255 = ~n36253 & ~n36254;
  assign n36256 = po3083 & ~n36255;
  assign n36257 = ~pi0550 & ~po3083;
  assign n36258 = ~n36256 & ~n36257;
  assign n36259 = ~po0944 & ~n36258;
  assign n36260 = pi0951 & po0944;
  assign po0834 = n36259 | n36260;
  assign n36262 = ~pi0551 & ~n35317;
  assign n36263 = ~n36217 & ~n36262;
  assign n36264 = po3083 & n36263;
  assign n36265 = pi0551 & ~po3083;
  assign n36266 = ~n36264 & ~n36265;
  assign n36267 = ~po0944 & n36266;
  assign n36268 = pi0892 & po0944;
  assign po0835 = n36267 | n36268;
  assign n36270 = ~pi0552 & ~pi0553;
  assign n36271 = ~n35317 & ~n36270;
  assign n36272 = po3083 & n36271;
  assign n36273 = pi0552 & ~po3083;
  assign n36274 = ~n36272 & ~n36273;
  assign n36275 = ~po0944 & n36274;
  assign n36276 = pi0952 & po0944;
  assign po0836 = n36275 | n36276;
  assign n36278 = ~pi0553 & ~po3083;
  assign n36279 = pi0553 & po3083;
  assign n36280 = ~n36278 & ~n36279;
  assign n36281 = ~po0944 & ~n36280;
  assign n36282 = pi0953 & po0944;
  assign po0837 = n36281 | n36282;
  assign n36284 = n34845 & n35895;
  assign n36285 = pi0554 & ~n36284;
  assign n36286 = ~pi0554 & n36284;
  assign n36287 = ~n36285 & ~n36286;
  assign n36288 = ~n34848 & n36287;
  assign po0838 = ~n35327 | n36288;
  assign n36290 = pi0558 & pi0559;
  assign n36291 = n35421 & n36290;
  assign n36292 = pi0556 & n36291;
  assign n36293 = pi0557 & n36292;
  assign n36294 = ~pi0555 & n36293;
  assign n36295 = pi0555 & ~n36293;
  assign n36296 = ~n36294 & ~n36295;
  assign n36297 = po2836 & ~n36296;
  assign n36298 = pi0555 & ~po2836;
  assign n36299 = ~n36297 & ~n36298;
  assign n36300 = ~po0945 & n36299;
  assign n36301 = pi0963 & po0945;
  assign po0839 = n36300 | n36301;
  assign n36303 = n35422 & n35423;
  assign n36304 = pi0556 & n36303;
  assign n36305 = ~pi0556 & ~n36303;
  assign n36306 = ~n36304 & ~n36305;
  assign n36307 = po2836 & ~n36306;
  assign n36308 = ~pi0556 & ~po2836;
  assign n36309 = ~n36307 & ~n36308;
  assign n36310 = ~po0945 & ~n36309;
  assign n36311 = pi0964 & po0945;
  assign po0840 = n36310 | n36311;
  assign n36313 = pi0561 & n36290;
  assign n36314 = pi0560 & n36313;
  assign n36315 = pi0564 & n36314;
  assign n36316 = ~pi0557 & n36315;
  assign n36317 = pi0557 & ~n36315;
  assign n36318 = ~n36316 & ~n36317;
  assign n36319 = po2836 & ~n36318;
  assign n36320 = pi0557 & ~po2836;
  assign n36321 = ~n36319 & ~n36320;
  assign n36322 = ~po0945 & n36321;
  assign n36323 = pi0965 & po0945;
  assign po0841 = n36322 | n36323;
  assign n36325 = ~pi0558 & ~n35422;
  assign n36326 = pi0558 & n35422;
  assign n36327 = ~n36325 & ~n36326;
  assign n36328 = po2836 & ~n36327;
  assign n36329 = ~pi0558 & ~po2836;
  assign n36330 = ~n36328 & ~n36329;
  assign n36331 = ~po0945 & ~n36330;
  assign n36332 = pi0900 & po0945;
  assign po0842 = n36331 | n36332;
  assign n36334 = ~pi0559 & ~n35421;
  assign n36335 = ~n35422 & ~n36334;
  assign n36336 = po2836 & n36335;
  assign n36337 = pi0559 & ~po2836;
  assign n36338 = ~n36336 & ~n36337;
  assign n36339 = ~po0945 & n36338;
  assign n36340 = pi0797 & po0945;
  assign po0843 = n36339 | n36340;
  assign n36342 = ~pi0560 & ~n35420;
  assign n36343 = ~n35421 & ~n36342;
  assign n36344 = po2836 & n36343;
  assign n36345 = pi0560 & ~po2836;
  assign n36346 = ~n36344 & ~n36345;
  assign n36347 = ~po0945 & n36346;
  assign n36348 = pi0798 & po0945;
  assign po0844 = n36347 | n36348;
  assign n36350 = ~pi0561 & ~po2836;
  assign n36351 = pi0561 & po2836;
  assign n36352 = ~n36350 & ~n36351;
  assign n36353 = ~po0945 & ~n36352;
  assign n36354 = pi0967 & po0945;
  assign po0845 = n36353 | n36354;
  assign n36356 = ~n35406 & n35408;
  assign n36357 = n35411 & ~n35418;
  assign n36358 = ~n36356 & ~n36357;
  assign po0993 = n35413 | ~n36358;
  assign n36360 = ~po0945 & po0993;
  assign n36361 = ~n35411 & n36360;
  assign po0846 = ~po2836 & n36361;
  assign n36363 = ~pi0563 & ~n36217;
  assign n36364 = ~n36252 & ~n36363;
  assign n36365 = po3083 & n36364;
  assign n36366 = pi0563 & ~po3083;
  assign n36367 = ~n36365 & ~n36366;
  assign n36368 = ~po0944 & n36367;
  assign n36369 = pi0891 & po0944;
  assign po0847 = n36368 | n36369;
  assign n36371 = ~pi0561 & ~pi0564;
  assign n36372 = ~n35420 & ~n36371;
  assign n36373 = po2836 & n36372;
  assign n36374 = pi0564 & ~po2836;
  assign n36375 = ~n36373 & ~n36374;
  assign n36376 = ~po0945 & n36375;
  assign n36377 = pi0966 & po0945;
  assign po0848 = n36376 | n36377;
  assign po0849 = pi3479 | pi3682;
  assign po0850 = pi3479 | ~pi3682;
  assign n36381 = pi0422 & n10759;
  assign n36382 = ~n35835 & ~n35836;
  assign n36383 = ~n10793 & n36382;
  assign n36384 = ~n36381 & n36383;
  assign n36385 = n10762 & n36384;
  assign n36386 = pi2978 & ~n36385;
  assign n36387 = ~n9361 & ~n10812;
  assign n36388 = ~n9415 & n10805;
  assign n36389 = n36387 & n36388;
  assign n36390 = pi0830 & ~n10805;
  assign n36391 = n10812 & n36390;
  assign n36392 = ~n36389 & ~n36391;
  assign n36393 = n11200 & n36392;
  assign n36394 = n11682 & ~n36392;
  assign n36395 = ~n36393 & ~n36394;
  assign n36396 = ~n10854 & ~n10873;
  assign n36397 = ~n10805 & n36396;
  assign n36398 = n9415 & n10805;
  assign n36399 = ~n10805 & ~n10812;
  assign n36400 = ~n36398 & ~n36399;
  assign n36401 = ~n10806 & n36400;
  assign n36402 = ~n10813 & n36401;
  assign n36403 = ~n36397 & n36402;
  assign n36404 = ~n36395 & n36403;
  assign n36405 = n9415 & ~n10812;
  assign n36406 = ~n10384 & n36405;
  assign n36407 = pi0421 & n10752;
  assign n36408 = ~n36406 & ~n36407;
  assign n36409 = n36392 & n36408;
  assign n36410 = n10372 & ~n36392;
  assign n36411 = ~n36409 & ~n36410;
  assign n36412 = ~n36403 & ~n36411;
  assign n36413 = ~n36404 & ~n36412;
  assign n36414 = n9361 & ~n10812;
  assign n36415 = n36388 & n36414;
  assign n36416 = ~n10805 & n10812;
  assign n36417 = ~n10854 & n36416;
  assign n36418 = ~n36415 & ~n36417;
  assign n36419 = ~n36413 & n36418;
  assign n36420 = ~n9825 & n36392;
  assign n36421 = ~n11181 & ~n36392;
  assign n36422 = ~n36420 & ~n36421;
  assign n36423 = n36403 & n36422;
  assign n36424 = n11752 & n36392;
  assign n36425 = n11674 & ~n36392;
  assign n36426 = ~n36424 & ~n36425;
  assign n36427 = ~n36403 & ~n36426;
  assign n36428 = ~n36423 & ~n36427;
  assign n36429 = ~n36418 & ~n36428;
  assign n36430 = ~n36419 & ~n36429;
  assign n36431 = n36386 & ~n36430;
  assign n36432 = pi0422 & n8612;
  assign n36433 = ~n35842 & ~n36432;
  assign n36434 = n8621 & n36433;
  assign n36435 = pi2409 & ~n36434;
  assign n36436 = n9415 & ~n10384;
  assign n36437 = ~n9415 & ~n9825;
  assign n36438 = ~n36436 & ~n36437;
  assign n36439 = n9361 & n36438;
  assign n36440 = ~n9415 & ~n10372;
  assign n36441 = ~n36436 & ~n36440;
  assign n36442 = ~n9361 & n36441;
  assign n36443 = ~n36439 & ~n36442;
  assign n36444 = n9415 & ~n10661;
  assign n36445 = ~n9415 & ~n10608;
  assign n36446 = ~n36444 & ~n36445;
  assign n36447 = n9361 & n36446;
  assign n36448 = ~n9415 & ~n10653;
  assign n36449 = ~n36444 & ~n36448;
  assign n36450 = ~n9361 & n36449;
  assign n36451 = ~n36447 & ~n36450;
  assign n36452 = ~pi3680 & n36451;
  assign n36453 = ~pi3680 & ~n36452;
  assign n36454 = n36443 & ~n36453;
  assign n36455 = n36435 & n36454;
  assign n36456 = ~n36431 & ~n36455;
  assign n36457 = ~n35827 & n36456;
  assign n36458 = n9345 & ~n36457;
  assign n36459 = ~pi3682 & ~n36458;
  assign n36460 = ~n8561 & ~n36459;
  assign n36461 = pi0565 & n8561;
  assign po0851 = n36460 | n36461;
  assign n36463 = pi2216 & n35501;
  assign n36464 = pi2202 & n35511;
  assign n36465 = ~n36463 & ~n36464;
  assign n36466 = pi2230 & n35497;
  assign n36467 = pi2244 & n35522;
  assign n36468 = ~n36466 & ~n36467;
  assign n36469 = n36465 & n36468;
  assign n36470 = ~n35507 & ~n35518;
  assign n36471 = ~n13701 & ~n36470;
  assign n36472 = n36469 & ~n36471;
  assign n36473 = ~n35539 & ~n36472;
  assign n36474 = pi0566 & n35539;
  assign po0852 = n36473 | n36474;
  assign n36476 = pi2231 & n35497;
  assign n36477 = pi2245 & n35522;
  assign n36478 = ~n36476 & ~n36477;
  assign n36479 = pi2217 & n35501;
  assign n36480 = pi2203 & n35511;
  assign n36481 = ~n36479 & ~n36480;
  assign n36482 = n36478 & n36481;
  assign n36483 = ~n13121 & ~n36470;
  assign n36484 = n36482 & ~n36483;
  assign n36485 = ~n35539 & ~n36484;
  assign n36486 = pi0567 & n35539;
  assign po0853 = n36485 | n36486;
  assign n36488 = ~n9825 & ~n36470;
  assign n36489 = pi2238 & n35497;
  assign n36490 = pi2252 & n35522;
  assign n36491 = ~n36489 & ~n36490;
  assign n36492 = pi2224 & n35501;
  assign n36493 = pi2210 & n35511;
  assign n36494 = ~n36492 & ~n36493;
  assign n36495 = n36491 & n36494;
  assign n36496 = ~n36488 & n36495;
  assign n36497 = ~n35539 & ~n36496;
  assign n36498 = pi0568 & n35539;
  assign po0854 = n36497 | n36498;
  assign n36500 = pi2242 & n35497;
  assign n36501 = pi2256 & n35522;
  assign n36502 = ~n36500 & ~n36501;
  assign n36503 = pi2228 & n35501;
  assign n36504 = pi2214 & n35511;
  assign n36505 = ~n36503 & ~n36504;
  assign n36506 = n36502 & n36505;
  assign n36507 = ~n11181 & ~n36470;
  assign n36508 = n36506 & ~n36507;
  assign n36509 = ~n35539 & ~n36508;
  assign n36510 = pi0569 & n35539;
  assign po0855 = n36509 | n36510;
  assign n36512 = pi1048 & ~po3627;
  assign n36513 = pi3239 & ~n36512;
  assign n36514 = pi1931 & ~pi3226;
  assign n36515 = pi0570 & ~n36514;
  assign n36516 = pi1931 & ~pi3144;
  assign n36517 = ~pi1735 & ~pi3303;
  assign n36518 = n36516 & n36517;
  assign n36519 = pi1735 & pi1931;
  assign n36520 = pi0878 & n36519;
  assign n36521 = ~n36518 & ~n36520;
  assign n36522 = n36515 & n36521;
  assign po0856 = n36513 & ~n36522;
  assign n36524 = ~pi3291 & ~n34969;
  assign n36525 = n34994 & n36524;
  assign n36526 = n34998 & ~n36525;
  assign n36527 = ~n35189 & n36526;
  assign n36528 = pi0571 & ~n36526;
  assign po0857 = n36527 | n36528;
  assign n36530 = ~n35157 & n36526;
  assign n36531 = pi0572 & ~n36526;
  assign po0858 = n36530 | n36531;
  assign n36533 = n35057 & n36526;
  assign n36534 = pi0573 & ~n36526;
  assign po0859 = n36533 | n36534;
  assign n36536 = n35858 & n35866;
  assign n36537 = ~pi0414 & n35992;
  assign n36538 = n20417 & n35997;
  assign n36539 = n36537 & n36538;
  assign n36540 = ~n35851 & n35868;
  assign n36541 = n35880 & n36540;
  assign n36542 = ~n35846 & ~n35857;
  assign n36543 = n35851 & n35854;
  assign n36544 = n35823 & n36543;
  assign n36545 = n35834 & n36544;
  assign n36546 = n36542 & n36545;
  assign n36547 = ~n35834 & n36544;
  assign n36548 = n36542 & n36547;
  assign n36549 = ~n36546 & ~n36548;
  assign n36550 = ~n36541 & n36549;
  assign n36551 = n35858 & n35864;
  assign n36552 = n36550 & ~n36551;
  assign n36553 = ~n36539 & n36552;
  assign n36554 = ~n36536 & n36553;
  assign n36555 = n35887 & ~n36554;
  assign n36556 = pi0574 & n8561;
  assign po0860 = n36555 | n36556;
  assign n36558 = ~n8561 & n8615;
  assign n36559 = n8607 & n36558;
  assign n36560 = ~pi0403 & ~pi0416;
  assign n36561 = pi0417 & n36560;
  assign n36562 = pi0418 & n36561;
  assign n36563 = ~n35827 & ~n36562;
  assign n36564 = ~n10752 & n36563;
  assign n36565 = ~n36075 & n36564;
  assign n36566 = ~pi0412 & n36565;
  assign n36567 = ~pi0415 & ~n36565;
  assign n36568 = ~n36566 & ~n36567;
  assign n36569 = ~n8620 & ~n10750;
  assign n36570 = ~pi0422 & ~n35839;
  assign n36571 = ~n35817 & ~n36570;
  assign n36572 = ~n35828 & n36571;
  assign n36573 = n36569 & n36572;
  assign n36574 = ~n36562 & n36573;
  assign n36575 = n36076 & n36574;
  assign n36576 = ~n24815 & n36575;
  assign n36577 = ~n36568 & ~n36576;
  assign n36578 = ~n8561 & n36577;
  assign n36579 = pi0411 & n36565;
  assign n36580 = pi0414 & ~n36565;
  assign n36581 = ~n36579 & ~n36580;
  assign n36582 = pi0420 & n36075;
  assign n36583 = ~n35819 & ~n36582;
  assign n36584 = ~n36079 & n36583;
  assign n36585 = n36581 & n36584;
  assign n36586 = pi0408 & n36565;
  assign n36587 = ~pi0427 & ~n36565;
  assign n36588 = ~n36586 & ~n36587;
  assign n36589 = pi0413 & n36565;
  assign n36590 = ~pi0407 & ~n36565;
  assign n36591 = ~n36589 & ~n36590;
  assign n36592 = pi0419 & n36075;
  assign n36593 = ~n35813 & ~n36592;
  assign n36594 = ~n36072 & n36593;
  assign n36595 = n36591 & n36594;
  assign n36596 = n36588 & n36595;
  assign n36597 = n36585 & n36596;
  assign n36598 = n36578 & n36597;
  assign n36599 = ~n36559 & ~n36598;
  assign n36600 = po3627 & ~n36599;
  assign n36601 = ~pi0575 & n36128;
  assign po0861 = n36600 | n36601;
  assign n36603 = n35891 & ~n36554;
  assign n36604 = pi0576 & n8561;
  assign po0862 = n36603 | n36604;
  assign n36606 = n31797 & ~n31802;
  assign n36607 = ~n31803 & ~n36606;
  assign n36608 = n31865 & ~n36607;
  assign n36609 = pi3641 & n36608;
  assign n36610 = pi0577 & ~n32073;
  assign n36611 = ~n36609 & ~n36610;
  assign n36612 = ~n31777 & ~n36611;
  assign n36613 = pi1716 & n31777;
  assign n36614 = ~n36612 & ~n36613;
  assign n36615 = ~n31779 & ~n36614;
  assign n36616 = ~pi2092 & n31779;
  assign po0863 = n36615 | n36616;
  assign n36618 = ~n35227 & n36526;
  assign n36619 = pi0578 & ~n36526;
  assign po0864 = n36618 | n36619;
  assign n36621 = ~n36576 & n36588;
  assign n36622 = n36584 & n36594;
  assign n36623 = n36621 & n36622;
  assign n36624 = n36581 & ~n36591;
  assign n36625 = ~n36568 & n36624;
  assign n36626 = n36623 & n36625;
  assign n36627 = pi0419 & ~pi0420;
  assign n36628 = n8615 & n36627;
  assign n36629 = ~n36626 & ~n36628;
  assign n36630 = ~n8561 & ~n36629;
  assign n36631 = ~pi0579 & n8561;
  assign n36632 = ~n36630 & ~n36631;
  assign po0865 = po3627 & ~n36632;
  assign n36634 = pi0580 & n8561;
  assign n36635 = pi0403 & ~pi0418;
  assign n36636 = n8615 & n36635;
  assign n36637 = n36568 & ~n36591;
  assign n36638 = ~n36576 & n36581;
  assign n36639 = n36622 & n36638;
  assign n36640 = n36588 & n36639;
  assign n36641 = n36637 & n36640;
  assign n36642 = ~n36636 & ~n36641;
  assign n36643 = ~n8561 & n36642;
  assign n36644 = ~n36634 & ~n36643;
  assign po0866 = po3627 & n36644;
  assign n36646 = ~n27717 & n31382;
  assign n36647 = pi0583 & n31381;
  assign n36648 = ~n24446 & n31384;
  assign n36649 = pi0583 & ~n31384;
  assign n36650 = ~n36648 & ~n36649;
  assign n36651 = n31388 & ~n36650;
  assign n36652 = ~n36647 & ~n36651;
  assign n36653 = ~n31391 & n36652;
  assign n36654 = ~n31382 & ~n36653;
  assign po0869 = n36646 | n36654;
  assign n36656 = ~n27717 & n31400;
  assign n36657 = pi0584 & n31399;
  assign n36658 = ~n24446 & n31402;
  assign n36659 = pi0584 & ~n31402;
  assign n36660 = ~n36658 & ~n36659;
  assign n36661 = n31406 & ~n36660;
  assign n36662 = ~n36657 & ~n36661;
  assign n36663 = ~n31409 & n36662;
  assign n36664 = ~n31400 & ~n36663;
  assign po0870 = n36656 | n36664;
  assign n36666 = ~n34993 & n36526;
  assign n36667 = pi0585 & ~n36526;
  assign po0871 = n36666 | n36667;
  assign n36669 = n19553 & n32625;
  assign n36670 = ~n9352 & n36669;
  assign n36671 = ~n19551 & ~n36670;
  assign n36672 = ~n19543 & n36671;
  assign n36673 = pi0586 & ~po3897;
  assign n36674 = n36672 & n36673;
  assign n36675 = n25053 & n31437;
  assign n36676 = ~n25053 & ~n31437;
  assign n36677 = ~n36675 & ~n36676;
  assign n36678 = n36669 & ~n36677;
  assign n36679 = ~pi0835 & ~n13121;
  assign n36680 = ~n36678 & ~n36679;
  assign n36681 = ~pi1513 & n20345;
  assign n36682 = ~pi1532 & n20347;
  assign n36683 = ~n36681 & ~n36682;
  assign n36684 = ~pi1614 & n20350;
  assign n36685 = ~pi1566 & n20353;
  assign n36686 = ~pi1410 & n20356;
  assign n36687 = ~n36685 & ~n36686;
  assign n36688 = ~pi1495 & n20360;
  assign n36689 = ~pi1402 & n20363;
  assign n36690 = ~n36688 & ~n36689;
  assign n36691 = n36687 & n36690;
  assign n36692 = ~n36684 & n36691;
  assign n36693 = n36683 & n36692;
  assign n36694 = n19550 & ~n36693;
  assign n36695 = n36680 & ~n36694;
  assign n36696 = ~n36672 & ~n36695;
  assign n36697 = ~po3897 & n36696;
  assign po0872 = n36674 | n36697;
  assign n36699 = pi2316 & n35632;
  assign n36700 = pi2304 & n35637;
  assign n36701 = ~n36699 & ~n36700;
  assign n36702 = pi2293 & n35647;
  assign n36703 = pi2281 & n35650;
  assign n36704 = ~n36702 & ~n36703;
  assign n36705 = n36701 & n36704;
  assign n36706 = ~n35628 & ~n35643;
  assign n36707 = ~n13121 & ~n36706;
  assign n36708 = n36705 & ~n36707;
  assign n36709 = ~n35660 & ~n36708;
  assign n36710 = pi0587 & n35660;
  assign po0873 = n36709 | n36710;
  assign n36712 = pi2297 & n35647;
  assign n36713 = pi2285 & n35650;
  assign n36714 = ~n36712 & ~n36713;
  assign n36715 = pi2320 & n35632;
  assign n36716 = pi2306 & n35637;
  assign n36717 = ~n36715 & ~n36716;
  assign n36718 = n36714 & n36717;
  assign n36719 = ~n14816 & ~n36706;
  assign n36720 = n36718 & ~n36719;
  assign n36721 = ~n35660 & ~n36720;
  assign n36722 = pi0588 & n35660;
  assign po0874 = n36721 | n36722;
  assign n36724 = pi2324 & n35632;
  assign n36725 = pi2310 & n35637;
  assign n36726 = ~n36724 & ~n36725;
  assign n36727 = pi2122 & n35647;
  assign n36728 = pi2288 & n35650;
  assign n36729 = ~n36727 & ~n36728;
  assign n36730 = n36726 & n36729;
  assign n36731 = ~n10608 & ~n36706;
  assign n36732 = n36730 & ~n36731;
  assign n36733 = ~n35660 & ~n36732;
  assign n36734 = pi0589 & n35660;
  assign po0875 = n36733 | n36734;
  assign n36736 = n35205 & n36526;
  assign n36737 = pi0590 & ~n36526;
  assign po0876 = n36736 | n36737;
  assign n36739 = ~n35096 & n36526;
  assign n36740 = pi0591 & ~n36526;
  assign po0877 = n36739 | n36740;
  assign n36742 = ~n35031 & n36526;
  assign n36743 = pi0592 & ~n36526;
  assign po0878 = n36742 | n36743;
  assign n36745 = ~n35137 & n36526;
  assign n36746 = pi0593 & ~n36526;
  assign po0879 = n36745 | n36746;
  assign n36748 = ~n35117 & n36526;
  assign n36749 = pi0594 & ~n36526;
  assign po0880 = n36748 | n36749;
  assign n36751 = n35081 & n36526;
  assign n36752 = pi0595 & ~n36526;
  assign po0881 = n36751 | n36752;
  assign n36754 = pi0596 & n8561;
  assign n36755 = pi0403 & pi0418;
  assign n36756 = n8615 & n36755;
  assign n36757 = ~n36588 & n36639;
  assign n36758 = n36637 & n36757;
  assign n36759 = ~n36756 & ~n36758;
  assign n36760 = ~n8561 & n36759;
  assign n36761 = ~n36754 & ~n36760;
  assign po0882 = po3627 & n36761;
  assign n36763 = ~n36576 & ~n36588;
  assign n36764 = n36622 & n36763;
  assign n36765 = n36625 & n36764;
  assign n36766 = n8615 & n35814;
  assign n36767 = ~n36765 & ~n36766;
  assign n36768 = ~n8561 & ~n36767;
  assign n36769 = ~pi0597 & n8561;
  assign n36770 = ~n36768 & ~n36769;
  assign po0883 = po3627 & ~n36770;
  assign n36772 = pi0598 & n8561;
  assign n36773 = ~pi0403 & pi0418;
  assign n36774 = n8615 & n36773;
  assign n36775 = n36568 & n36591;
  assign n36776 = n36757 & n36775;
  assign n36777 = ~n36774 & ~n36776;
  assign n36778 = ~n8561 & n36777;
  assign n36779 = ~n36772 & ~n36778;
  assign po0884 = po3627 & n36779;
  assign n36781 = pi0599 & n8561;
  assign n36782 = ~pi0403 & ~pi0418;
  assign n36783 = n8615 & n36782;
  assign n36784 = n36640 & n36775;
  assign n36785 = ~n36783 & ~n36784;
  assign n36786 = ~n8561 & n36785;
  assign n36787 = ~n36781 & ~n36786;
  assign po0885 = po3627 & n36787;
  assign n36789 = pi0600 & ~pi3647;
  assign n36790 = ~pi0931 & ~pi1067;
  assign n36791 = ~pi1088 & n36790;
  assign n36792 = ~pi1069 & n36791;
  assign n36793 = ~pi1068 & n36792;
  assign n36794 = ~pi0932 & ~pi1083;
  assign n36795 = n36793 & n36794;
  assign n36796 = ~pi0847 & n36795;
  assign n36797 = ~pi1085 & n36796;
  assign n36798 = ~pi0940 & n36797;
  assign n36799 = ~pi0689 & n36798;
  assign n36800 = ~pi0651 & ~pi0727;
  assign n36801 = n36799 & n36800;
  assign n36802 = ~pi0617 & n36801;
  assign n36803 = ~pi1087 & n36802;
  assign n36804 = ~pi0600 & n36803;
  assign n36805 = pi0600 & ~n36803;
  assign n36806 = ~n36804 & ~n36805;
  assign n36807 = pi3647 & ~n36806;
  assign n36808 = ~n36789 & ~n36807;
  assign n36809 = pi0742 & pi0940;
  assign n36810 = ~pi0742 & ~pi0940;
  assign n36811 = ~n36809 & ~n36810;
  assign n36812 = pi0743 & pi0932;
  assign n36813 = ~pi0743 & ~pi0932;
  assign n36814 = ~n36812 & ~n36813;
  assign n36815 = n36811 & n36814;
  assign n36816 = pi0744 & pi1083;
  assign n36817 = ~pi0744 & ~pi1083;
  assign n36818 = ~n36816 & ~n36817;
  assign n36819 = pi0745 & pi1068;
  assign n36820 = ~pi0745 & ~pi1068;
  assign n36821 = ~n36819 & ~n36820;
  assign n36822 = n36818 & n36821;
  assign n36823 = pi0746 & pi1069;
  assign n36824 = ~pi0746 & ~pi1069;
  assign n36825 = ~n36823 & ~n36824;
  assign n36826 = pi0737 & pi1088;
  assign n36827 = ~pi0737 & ~pi1088;
  assign n36828 = ~n36826 & ~n36827;
  assign n36829 = n36825 & n36828;
  assign n36830 = pi0747 & pi1067;
  assign n36831 = ~pi0747 & ~pi1067;
  assign n36832 = ~n36830 & ~n36831;
  assign n36833 = pi0748 & pi0931;
  assign n36834 = ~pi0748 & ~pi0931;
  assign n36835 = ~n36833 & ~n36834;
  assign n36836 = n36832 & n36835;
  assign n36837 = n36829 & n36836;
  assign n36838 = n36822 & n36837;
  assign n36839 = n36815 & n36838;
  assign n36840 = pi0600 & pi0895;
  assign n36841 = ~pi0600 & ~pi0895;
  assign n36842 = ~n36840 & ~n36841;
  assign n36843 = pi0617 & pi0896;
  assign n36844 = ~pi0617 & ~pi0896;
  assign n36845 = ~n36843 & ~n36844;
  assign n36846 = n36842 & n36845;
  assign n36847 = pi0870 & pi1087;
  assign n36848 = ~pi0870 & ~pi1087;
  assign n36849 = ~n36847 & ~n36848;
  assign n36850 = pi0727 & pi0897;
  assign n36851 = ~pi0727 & ~pi0897;
  assign n36852 = ~n36850 & ~n36851;
  assign n36853 = n36849 & n36852;
  assign n36854 = pi0651 & pi0872;
  assign n36855 = ~pi0651 & ~pi0872;
  assign n36856 = ~n36854 & ~n36855;
  assign n36857 = pi0689 & pi0871;
  assign n36858 = ~pi0689 & ~pi0871;
  assign n36859 = ~n36857 & ~n36858;
  assign n36860 = n36856 & n36859;
  assign n36861 = pi0869 & pi1085;
  assign n36862 = ~pi0869 & ~pi1085;
  assign n36863 = ~n36861 & ~n36862;
  assign n36864 = pi0847 & pi0894;
  assign n36865 = ~pi0847 & ~pi0894;
  assign n36866 = ~n36864 & ~n36865;
  assign n36867 = n36863 & n36866;
  assign n36868 = n36860 & n36867;
  assign n36869 = n36853 & n36868;
  assign n36870 = n36846 & n36869;
  assign n36871 = n36839 & n36870;
  assign n36872 = ~pi0738 & ~pi0790;
  assign n36873 = ~n36871 & ~n36872;
  assign n36874 = pi1931 & ~n36873;
  assign n36875 = pi3647 & n36874;
  assign n36876 = pi3575 & pi3647;
  assign n36877 = ~n36875 & ~n36876;
  assign n36878 = n36808 & n36877;
  assign n36879 = pi0895 & n36876;
  assign po0887 = n36878 | n36879;
  assign n36881 = pi0601 & ~pi3635;
  assign n36882 = ~pi0934 & ~pi1026;
  assign n36883 = ~pi0933 & ~pi1071;
  assign n36884 = ~pi1040 & n36883;
  assign n36885 = ~pi1072 & n36884;
  assign n36886 = n36882 & n36885;
  assign n36887 = ~pi1027 & n36886;
  assign n36888 = ~pi0848 & n36887;
  assign n36889 = ~pi1091 & n36888;
  assign n36890 = ~pi0935 & n36889;
  assign n36891 = ~pi0690 & n36890;
  assign n36892 = ~pi0652 & ~pi0698;
  assign n36893 = n36891 & n36892;
  assign n36894 = ~pi0618 & n36893;
  assign n36895 = ~pi1070 & n36894;
  assign n36896 = ~pi0601 & n36895;
  assign n36897 = pi0601 & ~n36895;
  assign n36898 = ~n36896 & ~n36897;
  assign n36899 = pi3635 & ~n36898;
  assign n36900 = ~n36881 & ~n36899;
  assign n36901 = pi0800 & pi0935;
  assign n36902 = ~pi0800 & ~pi0935;
  assign n36903 = ~n36901 & ~n36902;
  assign n36904 = pi0801 & pi0934;
  assign n36905 = ~pi0801 & ~pi0934;
  assign n36906 = ~n36904 & ~n36905;
  assign n36907 = n36903 & n36906;
  assign n36908 = pi0802 & pi1026;
  assign n36909 = ~pi0802 & ~pi1026;
  assign n36910 = ~n36908 & ~n36909;
  assign n36911 = pi0850 & pi1027;
  assign n36912 = ~pi0850 & ~pi1027;
  assign n36913 = ~n36911 & ~n36912;
  assign n36914 = n36910 & n36913;
  assign n36915 = pi0805 & pi0933;
  assign n36916 = ~pi0805 & ~pi0933;
  assign n36917 = ~n36915 & ~n36916;
  assign n36918 = pi0803 & pi1072;
  assign n36919 = ~pi0803 & ~pi1072;
  assign n36920 = ~n36918 & ~n36919;
  assign n36921 = n36917 & n36920;
  assign n36922 = pi0846 & pi1040;
  assign n36923 = ~pi0846 & ~pi1040;
  assign n36924 = ~n36922 & ~n36923;
  assign n36925 = pi0804 & pi1071;
  assign n36926 = ~pi0804 & ~pi1071;
  assign n36927 = ~n36925 & ~n36926;
  assign n36928 = n36924 & n36927;
  assign n36929 = n36921 & n36928;
  assign n36930 = n36914 & n36929;
  assign n36931 = n36907 & n36930;
  assign n36932 = pi0601 & pi0969;
  assign n36933 = ~pi0601 & ~pi0969;
  assign n36934 = ~n36932 & ~n36933;
  assign n36935 = pi0618 & pi0970;
  assign n36936 = ~pi0618 & ~pi0970;
  assign n36937 = ~n36935 & ~n36936;
  assign n36938 = n36934 & n36937;
  assign n36939 = pi0981 & pi1070;
  assign n36940 = ~pi0981 & ~pi1070;
  assign n36941 = ~n36939 & ~n36940;
  assign n36942 = pi0698 & pi0972;
  assign n36943 = ~pi0698 & ~pi0972;
  assign n36944 = ~n36942 & ~n36943;
  assign n36945 = n36941 & n36944;
  assign n36946 = pi0652 & pi0971;
  assign n36947 = ~pi0652 & ~pi0971;
  assign n36948 = ~n36946 & ~n36947;
  assign n36949 = pi0690 & pi0978;
  assign n36950 = ~pi0690 & ~pi0978;
  assign n36951 = ~n36949 & ~n36950;
  assign n36952 = n36948 & n36951;
  assign n36953 = pi0977 & pi1091;
  assign n36954 = ~pi0977 & ~pi1091;
  assign n36955 = ~n36953 & ~n36954;
  assign n36956 = pi0848 & pi0968;
  assign n36957 = ~pi0848 & ~pi0968;
  assign n36958 = ~n36956 & ~n36957;
  assign n36959 = n36955 & n36958;
  assign n36960 = n36952 & n36959;
  assign n36961 = n36945 & n36960;
  assign n36962 = n36938 & n36961;
  assign n36963 = n36931 & n36962;
  assign n36964 = ~pi0792 & ~pi0941;
  assign n36965 = ~n36963 & ~n36964;
  assign n36966 = pi2111 & ~n36965;
  assign n36967 = pi3635 & n36966;
  assign n36968 = pi3576 & pi3635;
  assign n36969 = ~n36967 & ~n36968;
  assign n36970 = n36900 & n36969;
  assign n36971 = pi0969 & n36968;
  assign po0889 = n36970 | n36971;
  assign n36973 = n35173 & n36526;
  assign n36974 = pi0602 & ~n36526;
  assign po0890 = n36973 | n36974;
  assign n36976 = ~n35242 & n36526;
  assign n36977 = pi0603 & ~n36526;
  assign po0891 = n36976 | n36977;
  assign po1085 = pi3100 & n36197;
  assign n36980 = pi0789 & pi3540;
  assign po0892 = po1085 | ~n36980;
  assign n36982 = ~pi0625 & n31013;
  assign n36983 = ~n31016 & ~n36982;
  assign n36984 = ~pi0605 & n31016;
  assign n36985 = ~n36983 & ~n36984;
  assign n36986 = pi0248 & pi0479;
  assign n36987 = ~n31038 & ~n31069;
  assign n36988 = ~n31026 & n36987;
  assign n36989 = n36986 & n36988;
  assign n36990 = pi0350 & n36989;
  assign n36991 = ~pi0247 & pi0329;
  assign n36992 = n36990 & n36991;
  assign n36993 = pi0955 & ~n36992;
  assign n36994 = ~pi0247 & ~pi1017;
  assign n36995 = n36993 & n36994;
  assign n36996 = ~n31347 & ~n36995;
  assign n36997 = ~pi2599 & ~n36996;
  assign n36998 = pi0605 & n31889;
  assign n36999 = ~n36997 & ~n36998;
  assign n37000 = ~n31013 & ~n36999;
  assign n37001 = ~n17368 & n31350;
  assign n37002 = ~n37000 & ~n37001;
  assign n37003 = ~n31016 & ~n37002;
  assign po0893 = n36985 | n37003;
  assign n37005 = ~pi0623 & n31013;
  assign n37006 = ~n31016 & ~n37005;
  assign n37007 = ~pi0606 & n31016;
  assign n37008 = ~n37006 & ~n37007;
  assign n37009 = pi0606 & n31889;
  assign n37010 = ~n36997 & ~n37009;
  assign n37011 = ~n31013 & ~n37010;
  assign n37012 = ~n9825 & n31350;
  assign n37013 = ~n37011 & ~n37012;
  assign n37014 = ~n31016 & ~n37013;
  assign po0894 = n37008 | n37014;
  assign n37016 = ~pi0624 & n31013;
  assign n37017 = ~n31016 & ~n37016;
  assign n37018 = ~pi0607 & n31016;
  assign n37019 = ~n37017 & ~n37018;
  assign n37020 = pi0607 & n31889;
  assign n37021 = ~n36997 & ~n37020;
  assign n37022 = ~n31013 & ~n37021;
  assign n37023 = ~n17199 & n31350;
  assign n37024 = ~n37022 & ~n37023;
  assign n37025 = ~n31016 & ~n37024;
  assign po0895 = n37019 | n37025;
  assign n37027 = ~pi0655 & n35406;
  assign n37028 = ~n35914 & ~n37027;
  assign n37029 = pi0562 & n37028;
  assign n37030 = ~pi0631 & n37029;
  assign n37031 = ~pi0955 & ~pi1017;
  assign n37032 = ~pi0562 & ~pi0693;
  assign n37033 = n37028 & n37032;
  assign n37034 = ~n37031 & n37033;
  assign n37035 = ~pi0608 & ~n37028;
  assign n37036 = ~n37034 & ~n37035;
  assign po0897 = n37030 | ~n37036;
  assign n37038 = n14475 & n36392;
  assign n37039 = n14545 & ~n36392;
  assign n37040 = ~n37038 & ~n37039;
  assign n37041 = n36403 & ~n37040;
  assign n37042 = ~n14502 & n36405;
  assign n37043 = pi0423 & n10752;
  assign n37044 = ~n37042 & ~n37043;
  assign n37045 = n36392 & n37044;
  assign n37046 = n14458 & ~n36392;
  assign n37047 = ~n37045 & ~n37046;
  assign n37048 = ~n36403 & ~n37047;
  assign n37049 = ~n37041 & ~n37048;
  assign n37050 = n36418 & ~n37049;
  assign n37051 = ~n14403 & n36392;
  assign n37052 = ~n14816 & ~n36392;
  assign n37053 = ~n37051 & ~n37052;
  assign n37054 = n36403 & n37053;
  assign n37055 = n14430 & n36392;
  assign n37056 = n14537 & ~n36392;
  assign n37057 = ~n37055 & ~n37056;
  assign n37058 = ~n36403 & ~n37057;
  assign n37059 = ~n37054 & ~n37058;
  assign n37060 = ~n36418 & ~n37059;
  assign n37061 = ~n37050 & ~n37060;
  assign n37062 = n11795 & n36392;
  assign n37063 = n12114 & ~n36392;
  assign n37064 = ~n37062 & ~n37063;
  assign n37065 = n36403 & ~n37064;
  assign n37066 = ~n10661 & n36405;
  assign n37067 = pi0405 & n10752;
  assign n37068 = ~n37066 & ~n37067;
  assign n37069 = n36392 & n37068;
  assign n37070 = n10653 & ~n36392;
  assign n37071 = ~n37069 & ~n37070;
  assign n37072 = ~n36403 & ~n37071;
  assign n37073 = ~n37065 & ~n37072;
  assign n37074 = n36418 & ~n37073;
  assign n37075 = ~n10608 & n36392;
  assign n37076 = ~n12061 & ~n36392;
  assign n37077 = ~n37075 & ~n37076;
  assign n37078 = n36403 & n37077;
  assign n37079 = n11781 & n36392;
  assign n37080 = n12106 & ~n36392;
  assign n37081 = ~n37079 & ~n37080;
  assign n37082 = ~n36403 & ~n37081;
  assign n37083 = ~n37078 & ~n37082;
  assign n37084 = ~n36418 & ~n37083;
  assign n37085 = ~n37074 & ~n37084;
  assign n37086 = n37061 & n37085;
  assign n37087 = n12138 & n36392;
  assign n37088 = n12493 & ~n36392;
  assign n37089 = ~n37087 & ~n37088;
  assign n37090 = n36403 & ~n37089;
  assign n37091 = ~n12163 & n36405;
  assign n37092 = pi0424 & n10752;
  assign n37093 = ~n37091 & ~n37092;
  assign n37094 = n36392 & n37093;
  assign n37095 = n12445 & ~n36392;
  assign n37096 = ~n37094 & ~n37095;
  assign n37097 = ~n36403 & ~n37096;
  assign n37098 = ~n37090 & ~n37097;
  assign n37099 = n36418 & ~n37098;
  assign n37100 = ~n12726 & n36392;
  assign n37101 = ~n12415 & ~n36392;
  assign n37102 = ~n37100 & ~n37101;
  assign n37103 = n36403 & n37102;
  assign n37104 = n12751 & n36392;
  assign n37105 = n12485 & ~n36392;
  assign n37106 = ~n37104 & ~n37105;
  assign n37107 = ~n36403 & ~n37106;
  assign n37108 = ~n37103 & ~n37107;
  assign n37109 = ~n36418 & ~n37108;
  assign n37110 = ~n37099 & ~n37109;
  assign n37111 = n12819 & n36392;
  assign n37112 = n12870 & ~n36392;
  assign n37113 = ~n37111 & ~n37112;
  assign n37114 = n36403 & ~n37113;
  assign n37115 = ~n12801 & n36405;
  assign n37116 = pi0425 & n10752;
  assign n37117 = ~n37115 & ~n37116;
  assign n37118 = n36392 & n37117;
  assign n37119 = n12785 & ~n36392;
  assign n37120 = ~n37118 & ~n37119;
  assign n37121 = ~n36403 & ~n37120;
  assign n37122 = ~n37114 & ~n37121;
  assign n37123 = n36418 & ~n37122;
  assign n37124 = n13121 & n36392;
  assign n37125 = n13398 & ~n36392;
  assign n37126 = ~n37124 & ~n37125;
  assign n37127 = n36403 & ~n37126;
  assign n37128 = n13149 & n36392;
  assign n37129 = n12862 & ~n36392;
  assign n37130 = ~n37128 & ~n37129;
  assign n37131 = ~n36403 & ~n37130;
  assign n37132 = ~n37127 & ~n37131;
  assign n37133 = ~n36418 & ~n37132;
  assign n37134 = ~n37123 & ~n37133;
  assign n37135 = n13710 & n36392;
  assign n37136 = n14095 & ~n36392;
  assign n37137 = ~n37135 & ~n37136;
  assign n37138 = n36403 & ~n37137;
  assign n37139 = ~n13735 & n36405;
  assign n37140 = pi0409 & n10752;
  assign n37141 = ~n37139 & ~n37140;
  assign n37142 = n36392 & n37141;
  assign n37143 = n14046 & ~n36392;
  assign n37144 = ~n37142 & ~n37143;
  assign n37145 = ~n36403 & ~n37144;
  assign n37146 = ~n37138 & ~n37145;
  assign n37147 = n36418 & ~n37146;
  assign n37148 = n13988 & n36392;
  assign n37149 = n13701 & ~n36392;
  assign n37150 = ~n37148 & ~n37149;
  assign n37151 = n36403 & ~n37150;
  assign n37152 = n14016 & n36392;
  assign n37153 = n14087 & ~n36392;
  assign n37154 = ~n37152 & ~n37153;
  assign n37155 = ~n36403 & ~n37154;
  assign n37156 = ~n37151 & ~n37155;
  assign n37157 = ~n36418 & ~n37156;
  assign n37158 = ~n37147 & ~n37157;
  assign n37159 = n37134 & n37158;
  assign n37160 = n14095 & n36392;
  assign n37161 = n13710 & ~n36392;
  assign n37162 = ~n37160 & ~n37161;
  assign n37163 = n36403 & ~n37162;
  assign n37164 = ~n14152 & n36405;
  assign n37165 = pi0406 & n10752;
  assign n37166 = ~n37164 & ~n37165;
  assign n37167 = n36392 & n37166;
  assign n37168 = n14134 & ~n36392;
  assign n37169 = ~n37167 & ~n37168;
  assign n37170 = ~n36403 & ~n37169;
  assign n37171 = ~n37163 & ~n37170;
  assign n37172 = n36418 & ~n37171;
  assign n37173 = ~n13701 & n36392;
  assign n37174 = ~n13988 & ~n36392;
  assign n37175 = ~n37173 & ~n37174;
  assign n37176 = n36403 & n37175;
  assign n37177 = n14087 & n36392;
  assign n37178 = n14016 & ~n36392;
  assign n37179 = ~n37177 & ~n37178;
  assign n37180 = ~n36403 & ~n37179;
  assign n37181 = ~n37176 & ~n37180;
  assign n37182 = ~n36418 & ~n37181;
  assign n37183 = ~n37172 & ~n37182;
  assign n37184 = n12870 & n36392;
  assign n37185 = n12819 & ~n36392;
  assign n37186 = ~n37184 & ~n37185;
  assign n37187 = n36403 & ~n37186;
  assign n37188 = ~n13424 & n36405;
  assign n37189 = pi0426 & n10752;
  assign n37190 = ~n37188 & ~n37189;
  assign n37191 = n36392 & n37190;
  assign n37192 = n13451 & ~n36392;
  assign n37193 = ~n37191 & ~n37192;
  assign n37194 = ~n36403 & ~n37193;
  assign n37195 = ~n37187 & ~n37194;
  assign n37196 = n36418 & ~n37195;
  assign n37197 = n13398 & n36392;
  assign n37198 = n13121 & ~n36392;
  assign n37199 = ~n37197 & ~n37198;
  assign n37200 = n36403 & ~n37199;
  assign n37201 = n12862 & n36392;
  assign n37202 = n13149 & ~n36392;
  assign n37203 = ~n37201 & ~n37202;
  assign n37204 = ~n36403 & ~n37203;
  assign n37205 = ~n37200 & ~n37204;
  assign n37206 = ~n36418 & ~n37205;
  assign n37207 = ~n37196 & ~n37206;
  assign n37208 = n36430 & n37207;
  assign n37209 = ~n36384 & n37208;
  assign n37210 = n37183 & n37209;
  assign n37211 = n37159 & n37210;
  assign n37212 = n14832 & n36392;
  assign n37213 = n15195 & ~n36392;
  assign n37214 = ~n37212 & ~n37213;
  assign n37215 = n36403 & ~n37214;
  assign n37216 = ~n14857 & n36405;
  assign n37217 = pi0422 & n10752;
  assign n37218 = ~n37216 & ~n37217;
  assign n37219 = n36392 & n37218;
  assign n37220 = n15146 & ~n36392;
  assign n37221 = ~n37219 & ~n37220;
  assign n37222 = ~n36403 & ~n37221;
  assign n37223 = ~n37215 & ~n37222;
  assign n37224 = n36418 & ~n37223;
  assign n37225 = ~n15426 & n36392;
  assign n37226 = ~n15115 & ~n36392;
  assign n37227 = ~n37225 & ~n37226;
  assign n37228 = n36403 & n37227;
  assign n37229 = n15454 & n36392;
  assign n37230 = n15187 & ~n36392;
  assign n37231 = ~n37229 & ~n37230;
  assign n37232 = ~n36403 & ~n37231;
  assign n37233 = ~n37228 & ~n37232;
  assign n37234 = ~n36418 & ~n37233;
  assign n37235 = ~n37224 & ~n37234;
  assign n37236 = n37211 & n37235;
  assign n37237 = n37110 & n37236;
  assign n37238 = n37086 & n37237;
  assign n37239 = ~n8561 & ~n37238;
  assign n37240 = ~pi0609 & n8561;
  assign po0899 = n37239 | n37240;
  assign n37242 = ~pi0622 & n37028;
  assign n37243 = pi0562 & n37242;
  assign n37244 = ~pi0610 & ~n37028;
  assign n37245 = ~n37034 & ~n37244;
  assign po0900 = n37243 | ~n37245;
  assign n37247 = ~pi0628 & n37028;
  assign n37248 = pi0562 & n37247;
  assign n37249 = ~pi0611 & ~n37028;
  assign n37250 = ~n37034 & ~n37249;
  assign po0901 = n37248 | ~n37250;
  assign n37252 = ~pi0989 & n9365;
  assign n37253 = ~n9384 & n9424;
  assign n37254 = ~n9424 & ~n9440;
  assign n37255 = ~n37253 & ~n37254;
  assign n37256 = ~po3855 & n37255;
  assign n37257 = ~pi3391 & po3855;
  assign n37258 = ~n37256 & ~n37257;
  assign n37259 = n9381 & n9424;
  assign n37260 = ~n9424 & ~n9433;
  assign n37261 = ~n37259 & ~n37260;
  assign n37262 = ~po3855 & n37261;
  assign n37263 = ~pi3367 & po3855;
  assign n37264 = ~n37262 & ~n37263;
  assign n37265 = ~n37258 & n37264;
  assign n37266 = n37252 & n37265;
  assign n37267 = ~pi1010 & n9365;
  assign n37268 = ~n37258 & ~n37264;
  assign n37269 = n37267 & n37268;
  assign n37270 = ~n37266 & ~n37269;
  assign n37271 = ~n12726 & ~n37270;
  assign n37272 = ~pi0988 & n9365;
  assign n37273 = n37258 & ~n37264;
  assign n37274 = ~n37272 & n37273;
  assign n37275 = pi2661 & n37274;
  assign n37276 = ~n37271 & ~n37275;
  assign n37277 = ~pi0987 & n9365;
  assign n37278 = n37258 & n37264;
  assign n37279 = ~n37277 & n37278;
  assign n37280 = pi2550 & n37279;
  assign n37281 = n37276 & ~n37280;
  assign n37282 = n37277 & n37278;
  assign n37283 = n37272 & n37273;
  assign n37284 = ~n37282 & ~n37283;
  assign n37285 = ~n12726 & ~n37284;
  assign n37286 = n37281 & ~n37285;
  assign n37287 = ~n37267 & n37268;
  assign n37288 = pi2602 & n37287;
  assign n37289 = ~n37252 & n37265;
  assign n37290 = pi2675 & n37289;
  assign n37291 = ~n37288 & ~n37290;
  assign n37292 = n37286 & n37291;
  assign n37293 = ~n35539 & ~n37292;
  assign n37294 = pi0612 & n35539;
  assign po0902 = n37293 | n37294;
  assign n37296 = ~n10608 & ~n37270;
  assign n37297 = pi2671 & n37274;
  assign n37298 = ~n37296 & ~n37297;
  assign n37299 = pi2657 & n37279;
  assign n37300 = n37298 & ~n37299;
  assign n37301 = ~n10608 & ~n37284;
  assign n37302 = n37300 & ~n37301;
  assign n37303 = pi2695 & n37287;
  assign n37304 = pi2685 & n37289;
  assign n37305 = ~n37303 & ~n37304;
  assign n37306 = n37302 & n37305;
  assign n37307 = ~n35539 & ~n37306;
  assign n37308 = pi0613 & n35539;
  assign po0903 = n37307 | n37308;
  assign n37310 = ~n15426 & ~n37270;
  assign n37311 = pi2672 & n37274;
  assign n37312 = ~n37310 & ~n37311;
  assign n37313 = pi2658 & n37279;
  assign n37314 = n37312 & ~n37313;
  assign n37315 = ~n15426 & ~n37284;
  assign n37316 = n37314 & ~n37315;
  assign n37317 = pi2696 & n37287;
  assign n37318 = pi2615 & n37289;
  assign n37319 = ~n37317 & ~n37318;
  assign n37320 = n37316 & n37319;
  assign n37321 = ~n35539 & ~n37320;
  assign n37322 = pi0614 & n35539;
  assign po0904 = n37321 | n37322;
  assign n37324 = ~pi0686 & ~pi0921;
  assign n37325 = pi0615 & n34979;
  assign n37326 = ~pi3291 & ~n34974;
  assign n37327 = ~n34969 & n37326;
  assign n37328 = ~n37324 & n37327;
  assign n37329 = ~n37325 & ~n37328;
  assign n37330 = ~n9352 & n37329;
  assign n37331 = n37324 & n37330;
  assign n37332 = ~n9352 & ~n34975;
  assign n37333 = pi0615 & n37332;
  assign n37334 = ~n37328 & n37333;
  assign n37335 = ~n37331 & ~n37334;
  assign n37336 = ~pi0615 & n37335;
  assign n37337 = ~pi0615 & n34977;
  assign n37338 = pi0615 & ~n34977;
  assign n37339 = ~n37337 & ~n37338;
  assign n37340 = ~n9352 & n37324;
  assign n37341 = ~n37325 & n37340;
  assign n37342 = ~n37339 & ~n37341;
  assign n37343 = ~pi0615 & ~n34979;
  assign n37344 = ~n37325 & ~n37343;
  assign n37345 = n37341 & n37344;
  assign n37346 = ~n37342 & ~n37345;
  assign n37347 = ~n37335 & n37346;
  assign po0905 = n37336 | n37347;
  assign n37349 = ~pi0616 & n37335;
  assign n37350 = pi0616 & ~n37335;
  assign po0906 = n37349 | n37350;
  assign n37352 = pi0617 & ~pi3647;
  assign n37353 = ~pi0932 & ~pi0940;
  assign n37354 = ~pi1083 & n36793;
  assign n37355 = ~pi0847 & ~pi1085;
  assign n37356 = n37354 & n37355;
  assign n37357 = n37353 & n37356;
  assign n37358 = ~pi0651 & ~pi0689;
  assign n37359 = n37357 & n37358;
  assign n37360 = ~pi1087 & n37359;
  assign n37361 = ~pi0727 & n37360;
  assign n37362 = ~pi0617 & n37361;
  assign n37363 = pi0617 & ~n37361;
  assign n37364 = ~n37362 & ~n37363;
  assign n37365 = pi3647 & ~n37364;
  assign n37366 = ~n37352 & ~n37365;
  assign n37367 = n36877 & n37366;
  assign n37368 = pi0896 & n36876;
  assign po0907 = n37367 | n37368;
  assign n37370 = pi0618 & ~pi3635;
  assign n37371 = ~pi0934 & ~pi0935;
  assign n37372 = ~pi1027 & n36885;
  assign n37373 = ~pi1026 & n37372;
  assign n37374 = ~pi0848 & ~pi1091;
  assign n37375 = n37373 & n37374;
  assign n37376 = n37371 & n37375;
  assign n37377 = ~pi0652 & ~pi0690;
  assign n37378 = n37376 & n37377;
  assign n37379 = ~pi1070 & n37378;
  assign n37380 = ~pi0698 & n37379;
  assign n37381 = ~pi0618 & n37380;
  assign n37382 = pi0618 & ~n37380;
  assign n37383 = ~n37381 & ~n37382;
  assign n37384 = pi3635 & ~n37383;
  assign n37385 = ~n37370 & ~n37384;
  assign n37386 = n36969 & n37385;
  assign n37387 = pi0970 & n36968;
  assign po0908 = n37386 | n37387;
  assign n37389 = ~pi3681 & n31863;
  assign n37390 = ~n31856 & ~n37389;
  assign n37391 = pi3439 & ~pi3469;
  assign n37392 = ~pi3681 & n37391;
  assign n37393 = n37390 & ~n37392;
  assign n37394 = pi1428 & ~n37393;
  assign n37395 = ~pi3681 & ~n31860;
  assign n37396 = ~pi1370 & n37395;
  assign n37397 = ~pi0691 & n37396;
  assign n37398 = ~pi0619 & n37397;
  assign n37399 = pi0619 & ~n37397;
  assign n37400 = ~n37398 & ~n37399;
  assign n37401 = pi0691 & ~n37396;
  assign n37402 = ~n37397 & ~n37401;
  assign n37403 = pi1370 & ~n37395;
  assign n37404 = ~n37396 & ~n37403;
  assign n37405 = ~n37402 & ~n37404;
  assign n37406 = ~n37400 & n37405;
  assign n37407 = n37400 & ~n37405;
  assign n37408 = ~n37406 & ~n37407;
  assign n37409 = pi3641 & ~n37408;
  assign n37410 = ~pi0619 & ~pi3641;
  assign n37411 = ~n37409 & ~n37410;
  assign n37412 = n37390 & ~n37411;
  assign n37413 = ~n37392 & n37412;
  assign po0909 = n37394 | n37413;
  assign n37415 = ~pi0620 & ~pi3641;
  assign n37416 = pi0620 & ~n37398;
  assign n37417 = ~pi0620 & n37398;
  assign n37418 = ~n37416 & ~n37417;
  assign n37419 = n37406 & ~n37418;
  assign n37420 = ~n37406 & n37418;
  assign n37421 = ~n37419 & ~n37420;
  assign n37422 = pi3641 & ~n37421;
  assign n37423 = ~n37415 & ~n37422;
  assign n37424 = n37393 & ~n37423;
  assign n37425 = pi1427 & ~n37393;
  assign po0910 = n37424 | n37425;
  assign n37427 = ~pi0608 & n37029;
  assign n37428 = ~pi0621 & ~n37028;
  assign n37429 = ~n37034 & ~n37428;
  assign po0911 = n37427 | ~n37429;
  assign n37431 = ~pi0621 & n37028;
  assign n37432 = pi0562 & n37431;
  assign n37433 = ~pi0622 & ~n37028;
  assign n37434 = ~n37034 & ~n37433;
  assign po0912 = n37432 | ~n37434;
  assign n37436 = ~pi0610 & n37028;
  assign n37437 = pi0562 & n37436;
  assign n37438 = ~pi0623 & ~n37028;
  assign n37439 = ~n37034 & ~n37438;
  assign po0913 = n37437 | ~n37439;
  assign n37441 = ~pi0623 & n37028;
  assign n37442 = pi0562 & n37441;
  assign n37443 = ~pi0624 & ~n37028;
  assign n37444 = ~n37034 & ~n37443;
  assign po0914 = n37442 | ~n37444;
  assign n37446 = ~pi0624 & n37028;
  assign n37447 = pi0562 & n37446;
  assign n37448 = ~pi0625 & ~n37028;
  assign n37449 = ~n37034 & ~n37448;
  assign po0915 = n37447 | ~n37449;
  assign n37451 = ~pi0694 & n37028;
  assign n37452 = pi0562 & n37451;
  assign n37453 = ~pi0626 & ~n37028;
  assign n37454 = ~n37034 & ~n37453;
  assign po0916 = n37452 | ~n37454;
  assign n37456 = ~pi0626 & n37028;
  assign n37457 = pi0562 & n37456;
  assign n37458 = ~pi0627 & ~n37028;
  assign n37459 = ~n37034 & ~n37458;
  assign po0917 = n37457 | ~n37459;
  assign n37461 = ~pi0627 & n37028;
  assign n37462 = pi0562 & n37461;
  assign n37463 = ~pi0628 & ~n37028;
  assign n37464 = ~n37034 & ~n37463;
  assign po0918 = n37462 | ~n37464;
  assign n37466 = ~pi0611 & n37028;
  assign n37467 = pi0562 & n37466;
  assign n37468 = ~pi0629 & ~n37028;
  assign n37469 = ~n37034 & ~n37468;
  assign po0919 = n37467 | ~n37469;
  assign n37471 = ~pi0629 & n37028;
  assign n37472 = pi0562 & n37471;
  assign n37473 = ~pi0630 & ~n37028;
  assign n37474 = ~n37034 & ~n37473;
  assign po0920 = n37472 | ~n37474;
  assign n37476 = ~pi0630 & n37028;
  assign n37477 = pi0562 & n37476;
  assign n37478 = ~pi0631 & ~n37028;
  assign n37479 = ~n37034 & ~n37478;
  assign po0921 = n37477 | ~n37479;
  assign n37481 = ~n35015 & n36526;
  assign n37482 = pi0632 & ~n36526;
  assign po0922 = n37481 | n37482;
  assign po0923 = ~pi0700 & ~po0993;
  assign n37485 = pi2653 & n37279;
  assign n37486 = ~n14816 & ~n37284;
  assign n37487 = pi2667 & n37274;
  assign n37488 = ~n14816 & ~n37270;
  assign n37489 = ~n37487 & ~n37488;
  assign n37490 = ~n37486 & n37489;
  assign n37491 = ~n37485 & n37490;
  assign n37492 = pi2691 & n37287;
  assign n37493 = pi2681 & n37289;
  assign n37494 = ~n37492 & ~n37493;
  assign n37495 = n37491 & n37494;
  assign n37496 = ~n35539 & ~n37495;
  assign n37497 = pi0634 & n35539;
  assign po0924 = n37496 | n37497;
  assign po0925 = ~pi0729 & ~po1022;
  assign n37500 = pi2649 & n37279;
  assign n37501 = ~n13121 & ~n37284;
  assign n37502 = pi2663 & n37274;
  assign n37503 = ~n13121 & ~n37270;
  assign n37504 = ~n37502 & ~n37503;
  assign n37505 = ~n37501 & n37504;
  assign n37506 = ~n37500 & n37505;
  assign n37507 = pi2688 & n37287;
  assign n37508 = pi2677 & n37289;
  assign n37509 = ~n37507 & ~n37508;
  assign n37510 = n37506 & n37509;
  assign n37511 = ~n35539 & ~n37510;
  assign n37512 = pi0636 & n35539;
  assign po0926 = n37511 | n37512;
  assign n37514 = pi2650 & n37279;
  assign n37515 = ~n13398 & ~n37284;
  assign n37516 = pi2664 & n37274;
  assign n37517 = ~n13398 & ~n37270;
  assign n37518 = ~n37516 & ~n37517;
  assign n37519 = ~n37515 & n37518;
  assign n37520 = ~n37514 & n37519;
  assign n37521 = pi2563 & n37287;
  assign n37522 = pi2678 & n37289;
  assign n37523 = ~n37521 & ~n37522;
  assign n37524 = n37520 & n37523;
  assign n37525 = ~n35539 & ~n37524;
  assign n37526 = pi0637 & n35539;
  assign po0927 = n37525 | n37526;
  assign n37528 = pi2680 & n37289;
  assign n37529 = ~n12415 & ~n37284;
  assign n37530 = pi2690 & n37287;
  assign n37531 = ~n12415 & ~n37270;
  assign n37532 = ~n37530 & ~n37531;
  assign n37533 = ~n37529 & n37532;
  assign n37534 = ~n37528 & n37533;
  assign n37535 = pi2666 & n37274;
  assign n37536 = pi2652 & n37279;
  assign n37537 = ~n37535 & ~n37536;
  assign n37538 = n37534 & n37537;
  assign n37539 = ~n35539 & ~n37538;
  assign n37540 = pi0638 & n35539;
  assign po0928 = n37539 | n37540;
  assign n37542 = pi2654 & n37279;
  assign n37543 = ~n15115 & ~n37284;
  assign n37544 = pi2668 & n37274;
  assign n37545 = ~n15115 & ~n37270;
  assign n37546 = ~n37544 & ~n37545;
  assign n37547 = ~n37543 & n37546;
  assign n37548 = ~n37542 & n37547;
  assign n37549 = pi2692 & n37287;
  assign n37550 = pi2682 & n37289;
  assign n37551 = ~n37549 & ~n37550;
  assign n37552 = n37548 & n37551;
  assign n37553 = ~n35539 & ~n37552;
  assign n37554 = pi0639 & n35539;
  assign po0929 = n37553 | n37554;
  assign n37556 = pi2683 & n37289;
  assign n37557 = ~n12061 & ~n37284;
  assign n37558 = pi2693 & n37287;
  assign n37559 = ~n12061 & ~n37270;
  assign n37560 = ~n37558 & ~n37559;
  assign n37561 = ~n37557 & n37560;
  assign n37562 = ~n37556 & n37561;
  assign n37563 = pi2669 & n37274;
  assign n37564 = pi2655 & n37279;
  assign n37565 = ~n37563 & ~n37564;
  assign n37566 = n37562 & n37565;
  assign n37567 = ~n35539 & ~n37566;
  assign n37568 = pi0640 & n35539;
  assign po0930 = n37567 | n37568;
  assign n37570 = pi2660 & n37279;
  assign n37571 = ~n11181 & ~n37284;
  assign n37572 = pi2674 & n37274;
  assign n37573 = ~n11181 & ~n37270;
  assign n37574 = ~n37572 & ~n37573;
  assign n37575 = ~n37571 & n37574;
  assign n37576 = ~n37570 & n37575;
  assign n37577 = pi2562 & n37287;
  assign n37578 = pi2603 & n37289;
  assign n37579 = ~n37577 & ~n37578;
  assign n37580 = n37576 & n37579;
  assign n37581 = ~n35539 & ~n37580;
  assign n37582 = pi0641 & n35539;
  assign po0931 = n37581 | n37582;
  assign n37584 = ~n9361 & ~n13451;
  assign n37585 = n9361 & ~n13398;
  assign n37586 = ~n37584 & ~n37585;
  assign n37587 = ~n9372 & n37265;
  assign n37588 = ~n9404 & n37268;
  assign n37589 = ~n37587 & ~n37588;
  assign n37590 = ~n37586 & ~n37589;
  assign n37591 = n9404 & n37268;
  assign n37592 = pi1977 & n37591;
  assign n37593 = ~n37590 & ~n37592;
  assign n37594 = n9372 & n37265;
  assign n37595 = pi2272 & n37594;
  assign n37596 = n37593 & ~n37595;
  assign n37597 = ~n9411 & n37273;
  assign n37598 = ~n9394 & n37278;
  assign n37599 = ~n37597 & ~n37598;
  assign n37600 = ~n37586 & ~n37599;
  assign n37601 = n37596 & ~n37600;
  assign n37602 = n9394 & n37278;
  assign n37603 = pi2258 & n37602;
  assign n37604 = n9411 & n37273;
  assign n37605 = pi2262 & n37604;
  assign n37606 = ~n37603 & ~n37605;
  assign n37607 = n37601 & n37606;
  assign n37608 = ~n35539 & ~n37607;
  assign n37609 = pi0642 & n35539;
  assign po0932 = n37608 | n37609;
  assign n37611 = n9361 & ~n10608;
  assign n37612 = ~n9361 & ~n10653;
  assign n37613 = ~n37611 & ~n37612;
  assign n37614 = ~n37589 & ~n37613;
  assign n37615 = pi1984 & n37591;
  assign n37616 = ~n37614 & ~n37615;
  assign n37617 = pi2446 & n37594;
  assign n37618 = n37616 & ~n37617;
  assign n37619 = ~n37599 & ~n37613;
  assign n37620 = n37618 & ~n37619;
  assign n37621 = pi2436 & n37602;
  assign n37622 = pi2269 & n37604;
  assign n37623 = ~n37621 & ~n37622;
  assign n37624 = n37620 & n37623;
  assign n37625 = ~n35539 & ~n37624;
  assign n37626 = pi0643 & n35539;
  assign po0933 = n37625 | n37626;
  assign n37628 = ~pi0920 & n9365;
  assign n37629 = pi0414 & n9424;
  assign n37630 = ~n37254 & ~n37629;
  assign n37631 = ~po3855 & n37630;
  assign n37632 = ~pi3398 & po3855;
  assign n37633 = ~n37631 & ~n37632;
  assign n37634 = pi0415 & n9424;
  assign n37635 = ~n37260 & ~n37634;
  assign n37636 = ~po3855 & n37635;
  assign n37637 = ~pi3392 & po3855;
  assign n37638 = ~n37636 & ~n37637;
  assign n37639 = ~n37633 & n37638;
  assign n37640 = n37628 & n37639;
  assign n37641 = ~pi0991 & n9365;
  assign n37642 = ~n37633 & ~n37638;
  assign n37643 = n37641 & n37642;
  assign n37644 = ~n37640 & ~n37643;
  assign n37645 = ~n13701 & ~n37644;
  assign n37646 = ~pi0990 & n9365;
  assign n37647 = n37633 & ~n37638;
  assign n37648 = ~n37646 & n37647;
  assign n37649 = pi2720 & n37648;
  assign n37650 = ~n37645 & ~n37649;
  assign n37651 = ~pi1051 & n9365;
  assign n37652 = n37633 & n37638;
  assign n37653 = ~n37651 & n37652;
  assign n37654 = pi2709 & n37653;
  assign n37655 = n37650 & ~n37654;
  assign n37656 = n37651 & n37652;
  assign n37657 = n37646 & n37647;
  assign n37658 = ~n37656 & ~n37657;
  assign n37659 = ~n13701 & ~n37658;
  assign n37660 = n37655 & ~n37659;
  assign n37661 = ~n37641 & n37642;
  assign n37662 = pi2739 & n37661;
  assign n37663 = ~n37628 & n37639;
  assign n37664 = pi2566 & n37663;
  assign n37665 = ~n37662 & ~n37664;
  assign n37666 = n37660 & n37665;
  assign n37667 = ~n35660 & ~n37666;
  assign n37668 = pi0644 & n35660;
  assign po0934 = n37667 | n37668;
  assign n37670 = ~n9825 & ~n37644;
  assign n37671 = pi2774 & n37648;
  assign n37672 = ~n37670 & ~n37671;
  assign n37673 = pi2716 & n37653;
  assign n37674 = n37672 & ~n37673;
  assign n37675 = ~n9825 & ~n37658;
  assign n37676 = n37674 & ~n37675;
  assign n37677 = pi2744 & n37661;
  assign n37678 = pi2561 & n37663;
  assign n37679 = ~n37677 & ~n37678;
  assign n37680 = n37676 & n37679;
  assign n37681 = ~n35660 & ~n37680;
  assign n37682 = pi0645 & n35660;
  assign po0935 = n37681 | n37682;
  assign n37684 = ~n10608 & ~n37644;
  assign n37685 = pi2725 & n37648;
  assign n37686 = ~n37684 & ~n37685;
  assign n37687 = pi2717 & n37653;
  assign n37688 = n37686 & ~n37687;
  assign n37689 = ~n10608 & ~n37658;
  assign n37690 = n37688 & ~n37689;
  assign n37691 = pi2543 & n37661;
  assign n37692 = pi2735 & n37663;
  assign n37693 = ~n37691 & ~n37692;
  assign n37694 = n37690 & n37693;
  assign n37695 = ~n35660 & ~n37694;
  assign n37696 = pi0646 & n35660;
  assign po0936 = n37695 | n37696;
  assign n37698 = ~n34977 & ~n34979;
  assign n37699 = ~n37341 & n37698;
  assign n37700 = ~n34982 & ~n34984;
  assign n37701 = n37341 & n37700;
  assign n37702 = ~n37699 & ~n37701;
  assign n37703 = ~n37335 & n37702;
  assign n37704 = ~pi0647 & n37335;
  assign po0937 = n37703 | n37704;
  assign n37706 = pi1330 & ~po3627;
  assign n37707 = pi3227 & ~n37706;
  assign n37708 = ~pi1641 & ~pi3681;
  assign n37709 = pi1096 & n37708;
  assign n37710 = pi3238 & ~n37709;
  assign n37711 = pi0648 & n37710;
  assign po0938 = n37707 & ~n37711;
  assign n37713 = ~pi0419 & pi0420;
  assign n37714 = n8615 & n37713;
  assign n37715 = ~n36588 & n36595;
  assign n37716 = n36577 & n36585;
  assign n37717 = n37715 & n37716;
  assign n37718 = ~n37714 & ~n37717;
  assign n37719 = ~n8561 & ~n37718;
  assign n37720 = ~pi0649 & n8561;
  assign n37721 = ~n37719 & ~n37720;
  assign po0939 = po3627 & ~n37721;
  assign n37723 = pi0650 & n8561;
  assign n37724 = pi0415 & n36010;
  assign n37725 = n36022 & n37724;
  assign n37726 = n36020 & n37724;
  assign n37727 = pi0407 & pi0415;
  assign n37728 = ~pi0414 & n36046;
  assign n37729 = n37727 & n37728;
  assign n37730 = n35992 & n37729;
  assign n37731 = ~n36114 & ~n37730;
  assign n37732 = ~n37726 & n37731;
  assign n37733 = ~n37725 & n37732;
  assign n37734 = ~n8561 & ~n37733;
  assign n37735 = ~n37723 & ~n37734;
  assign n37736 = n36031 & n36040;
  assign n37737 = ~n10793 & ~n36562;
  assign n37738 = ~n36075 & n37737;
  assign n37739 = ~n37736 & n37738;
  assign n37740 = ~n8561 & ~n37739;
  assign n37741 = n20417 & n35992;
  assign n37742 = n37728 & n37741;
  assign n37743 = n20460 & n35992;
  assign n37744 = n37728 & n37743;
  assign n37745 = n36537 & n37727;
  assign n37746 = n35997 & n37745;
  assign n37747 = n20460 & n35997;
  assign n37748 = n36537 & n37747;
  assign n37749 = ~n37746 & ~n37748;
  assign n37750 = ~n37744 & n37749;
  assign n37751 = ~n37742 & n37750;
  assign n37752 = ~n8561 & ~n37751;
  assign n37753 = ~n37740 & ~n37752;
  assign po0940 = ~n37735 | ~n37753;
  assign n37755 = pi0651 & ~pi3647;
  assign n37756 = pi0651 & n36799;
  assign n37757 = ~pi0651 & ~n36799;
  assign n37758 = ~n37756 & ~n37757;
  assign n37759 = pi3647 & n37758;
  assign n37760 = ~n37755 & ~n37759;
  assign n37761 = n36877 & n37760;
  assign n37762 = pi0872 & n36876;
  assign po0941 = n37761 | n37762;
  assign n37764 = pi0652 & ~pi3635;
  assign n37765 = pi0652 & n36891;
  assign n37766 = ~pi0652 & ~n36891;
  assign n37767 = ~n37765 & ~n37766;
  assign n37768 = pi3635 & n37767;
  assign n37769 = ~n37764 & ~n37768;
  assign n37770 = n36969 & n37769;
  assign n37771 = pi0971 & n36968;
  assign po0942 = n37770 | n37771;
  assign n37773 = n31799 & n31801;
  assign n37774 = ~n31802 & ~n37773;
  assign n37775 = n31865 & ~n37774;
  assign n37776 = pi3641 & n37775;
  assign n37777 = pi0653 & ~n32073;
  assign n37778 = ~n37776 & ~n37777;
  assign n37779 = ~n31777 & ~n37778;
  assign n37780 = pi1717 & n31777;
  assign n37781 = ~n37779 & ~n37780;
  assign n37782 = ~n31779 & ~n37781;
  assign n37783 = ~pi2393 & n31779;
  assign po0943 = n37782 | n37783;
  assign n37785 = pi2552 & n37663;
  assign n37786 = ~n11181 & ~n37644;
  assign n37787 = pi2542 & n37661;
  assign n37788 = ~n11181 & ~n37658;
  assign n37789 = ~n37787 & ~n37788;
  assign n37790 = ~n37786 & n37789;
  assign n37791 = ~n37785 & n37790;
  assign n37792 = pi2727 & n37648;
  assign n37793 = pi2532 & n37653;
  assign n37794 = ~n37792 & ~n37793;
  assign n37795 = n37791 & n37794;
  assign n37796 = ~n35660 & ~n37795;
  assign n37797 = pi0656 & n35660;
  assign po0946 = n37796 | n37797;
  assign n37799 = pi2733 & n37663;
  assign n37800 = ~n14816 & ~n37644;
  assign n37801 = pi2742 & n37661;
  assign n37802 = ~n14816 & ~n37658;
  assign n37803 = ~n37801 & ~n37802;
  assign n37804 = ~n37800 & n37803;
  assign n37805 = ~n37799 & n37804;
  assign n37806 = pi2723 & n37648;
  assign n37807 = pi2713 & n37653;
  assign n37808 = ~n37806 & ~n37807;
  assign n37809 = n37805 & n37808;
  assign n37810 = ~n35660 & ~n37809;
  assign n37811 = pi0657 & n35660;
  assign po0947 = n37810 | n37811;
  assign n37813 = ~n13701 & ~n37284;
  assign n37814 = pi2662 & n37274;
  assign n37815 = ~n37813 & ~n37814;
  assign n37816 = pi2648 & n37279;
  assign n37817 = n37815 & ~n37816;
  assign n37818 = ~n13701 & ~n37270;
  assign n37819 = n37817 & ~n37818;
  assign n37820 = pi2687 & n37287;
  assign n37821 = pi2676 & n37289;
  assign n37822 = ~n37820 & ~n37821;
  assign n37823 = n37819 & n37822;
  assign n37824 = ~n35539 & ~n37823;
  assign n37825 = pi0658 & n35539;
  assign po0948 = n37824 | n37825;
  assign n37827 = ~pi0659 & n20459;
  assign n37828 = ~n20459 & n20479;
  assign n37829 = ~n37827 & ~n37828;
  assign po0949 = ~po3897 & n37829;
  assign n37831 = n9361 & ~n12726;
  assign n37832 = ~n9361 & ~n12445;
  assign n37833 = ~n37831 & ~n37832;
  assign n37834 = ~n37599 & ~n37833;
  assign n37835 = pi1976 & n37591;
  assign n37836 = ~n37834 & ~n37835;
  assign n37837 = pi2271 & n37594;
  assign n37838 = n37836 & ~n37837;
  assign n37839 = ~n37589 & ~n37833;
  assign n37840 = n37838 & ~n37839;
  assign n37841 = pi2257 & n37602;
  assign n37842 = pi2261 & n37604;
  assign n37843 = ~n37841 & ~n37842;
  assign n37844 = n37840 & n37843;
  assign n37845 = ~n35539 & ~n37844;
  assign n37846 = pi0660 & n35539;
  assign po0950 = n37845 | n37846;
  assign n37848 = ~n9361 & ~n14046;
  assign n37849 = n9361 & ~n13988;
  assign n37850 = ~n37848 & ~n37849;
  assign n37851 = ~n37599 & ~n37850;
  assign n37852 = pi1978 & n37591;
  assign n37853 = ~n37851 & ~n37852;
  assign n37854 = pi2442 & n37594;
  assign n37855 = n37853 & ~n37854;
  assign n37856 = ~n37589 & ~n37850;
  assign n37857 = n37855 & ~n37856;
  assign n37858 = pi2432 & n37602;
  assign n37859 = pi2263 & n37604;
  assign n37860 = ~n37858 & ~n37859;
  assign n37861 = n37857 & n37860;
  assign n37862 = ~n35539 & ~n37861;
  assign n37863 = pi0661 & n35539;
  assign po0951 = n37862 | n37863;
  assign n37865 = ~n9361 & ~n17983;
  assign n37866 = n9361 & ~n12415;
  assign n37867 = ~n37865 & ~n37866;
  assign n37868 = ~n37599 & ~n37867;
  assign n37869 = pi1979 & n37591;
  assign n37870 = ~n37868 & ~n37869;
  assign n37871 = pi2273 & n37594;
  assign n37872 = n37870 & ~n37871;
  assign n37873 = ~n37589 & ~n37867;
  assign n37874 = n37872 & ~n37873;
  assign n37875 = pi2259 & n37602;
  assign n37876 = pi2264 & n37604;
  assign n37877 = ~n37875 & ~n37876;
  assign n37878 = n37874 & n37877;
  assign n37879 = ~n35539 & ~n37878;
  assign n37880 = pi0662 & n35539;
  assign po0952 = n37879 | n37880;
  assign n37882 = ~n9361 & ~n17927;
  assign n37883 = n9361 & ~n14816;
  assign n37884 = ~n37882 & ~n37883;
  assign n37885 = ~n37599 & ~n37884;
  assign n37886 = pi2265 & n37604;
  assign n37887 = ~n37885 & ~n37886;
  assign n37888 = pi2260 & n37602;
  assign n37889 = n37887 & ~n37888;
  assign n37890 = ~n37589 & ~n37884;
  assign n37891 = n37889 & ~n37890;
  assign n37892 = pi2443 & n37594;
  assign n37893 = pi1980 & n37591;
  assign n37894 = ~n37892 & ~n37893;
  assign n37895 = n37891 & n37894;
  assign n37896 = ~n35539 & ~n37895;
  assign n37897 = pi0663 & n35539;
  assign po0953 = n37896 | n37897;
  assign n37899 = ~n9361 & ~n17866;
  assign n37900 = n9361 & ~n15115;
  assign n37901 = ~n37899 & ~n37900;
  assign n37902 = ~n37599 & ~n37901;
  assign n37903 = pi1981 & n37591;
  assign n37904 = ~n37902 & ~n37903;
  assign n37905 = pi2274 & n37594;
  assign n37906 = n37904 & ~n37905;
  assign n37907 = ~n37589 & ~n37901;
  assign n37908 = n37906 & ~n37907;
  assign n37909 = pi2433 & n37602;
  assign n37910 = pi2266 & n37604;
  assign n37911 = ~n37909 & ~n37910;
  assign n37912 = n37908 & n37911;
  assign n37913 = ~n35539 & ~n37912;
  assign n37914 = pi0664 & n35539;
  assign po0954 = n37913 | n37914;
  assign n37916 = ~n9361 & ~n17809;
  assign n37917 = n9361 & ~n12061;
  assign n37918 = ~n37916 & ~n37917;
  assign n37919 = ~n37599 & ~n37918;
  assign n37920 = pi2267 & n37604;
  assign n37921 = ~n37919 & ~n37920;
  assign n37922 = pi2434 & n37602;
  assign n37923 = n37921 & ~n37922;
  assign n37924 = ~n37589 & ~n37918;
  assign n37925 = n37923 & ~n37924;
  assign n37926 = pi2444 & n37594;
  assign n37927 = pi1982 & n37591;
  assign n37928 = ~n37926 & ~n37927;
  assign n37929 = n37925 & n37928;
  assign n37930 = ~n35539 & ~n37929;
  assign n37931 = pi0665 & n35539;
  assign po0955 = n37930 | n37931;
  assign n37933 = n9361 & ~n9825;
  assign n37934 = ~n9361 & ~n10372;
  assign n37935 = ~n37933 & ~n37934;
  assign n37936 = ~n37599 & ~n37935;
  assign n37937 = pi2268 & n37604;
  assign n37938 = ~n37936 & ~n37937;
  assign n37939 = pi2435 & n37602;
  assign n37940 = n37938 & ~n37939;
  assign n37941 = ~n37589 & ~n37935;
  assign n37942 = n37940 & ~n37941;
  assign n37943 = pi2445 & n37594;
  assign n37944 = pi1983 & n37591;
  assign n37945 = ~n37943 & ~n37944;
  assign n37946 = n37942 & n37945;
  assign n37947 = ~n35539 & ~n37946;
  assign n37948 = pi0666 & n35539;
  assign po0956 = n37947 | n37948;
  assign n37950 = ~n9361 & ~n17751;
  assign n37951 = n9361 & ~n11181;
  assign n37952 = ~n37950 & ~n37951;
  assign n37953 = ~n37599 & ~n37952;
  assign n37954 = pi1985 & n37591;
  assign n37955 = ~n37953 & ~n37954;
  assign n37956 = pi2447 & n37594;
  assign n37957 = n37955 & ~n37956;
  assign n37958 = ~n37589 & ~n37952;
  assign n37959 = n37957 & ~n37958;
  assign n37960 = pi2437 & n37602;
  assign n37961 = pi2270 & n37604;
  assign n37962 = ~n37960 & ~n37961;
  assign n37963 = n37959 & n37962;
  assign n37964 = ~n35539 & ~n37963;
  assign n37965 = pi0667 & n35539;
  assign po0957 = n37964 | n37965;
  assign n37967 = ~n12726 & ~n37658;
  assign n37968 = pi2738 & n37661;
  assign n37969 = ~n37967 & ~n37968;
  assign n37970 = pi2728 & n37663;
  assign n37971 = n37969 & ~n37970;
  assign n37972 = ~n12726 & ~n37644;
  assign n37973 = n37971 & ~n37972;
  assign n37974 = pi2719 & n37648;
  assign n37975 = pi2708 & n37653;
  assign n37976 = ~n37974 & ~n37975;
  assign n37977 = n37973 & n37976;
  assign n37978 = ~n35660 & ~n37977;
  assign n37979 = pi0668 & n35660;
  assign po0958 = n37978 | n37979;
  assign n37981 = pi2710 & n37653;
  assign n37982 = ~n13121 & ~n37644;
  assign n37983 = pi2531 & n37648;
  assign n37984 = ~n13121 & ~n37658;
  assign n37985 = ~n37983 & ~n37984;
  assign n37986 = ~n37982 & n37985;
  assign n37987 = ~n37981 & n37986;
  assign n37988 = pi2548 & n37661;
  assign n37989 = pi2729 & n37663;
  assign n37990 = ~n37988 & ~n37989;
  assign n37991 = n37987 & n37990;
  assign n37992 = ~n35660 & ~n37991;
  assign n37993 = pi0669 & n35660;
  assign po0959 = n37992 | n37993;
  assign n37995 = pi2730 & n37663;
  assign n37996 = ~n13398 & ~n37644;
  assign n37997 = pi2740 & n37661;
  assign n37998 = ~n13398 & ~n37658;
  assign n37999 = ~n37997 & ~n37998;
  assign n38000 = ~n37996 & n37999;
  assign n38001 = ~n37995 & n38000;
  assign n38002 = pi2528 & n37648;
  assign n38003 = pi2711 & n37653;
  assign n38004 = ~n38002 & ~n38003;
  assign n38005 = n38001 & n38004;
  assign n38006 = ~n35660 & ~n38005;
  assign n38007 = pi0670 & n35660;
  assign po0960 = n38006 | n38007;
  assign n38009 = pi2731 & n37663;
  assign n38010 = ~n13988 & ~n37658;
  assign n38011 = pi2741 & n37661;
  assign n38012 = ~n13988 & ~n37644;
  assign n38013 = ~n38011 & ~n38012;
  assign n38014 = ~n38010 & n38013;
  assign n38015 = ~n38009 & n38014;
  assign n38016 = pi2721 & n37648;
  assign n38017 = pi2536 & n37653;
  assign n38018 = ~n38016 & ~n38017;
  assign n38019 = n38015 & n38018;
  assign n38020 = ~n35660 & ~n38019;
  assign n38021 = pi0671 & n35660;
  assign po0961 = n38020 | n38021;
  assign n38023 = pi2732 & n37663;
  assign n38024 = ~n12415 & ~n37658;
  assign n38025 = pi2546 & n37661;
  assign n38026 = ~n12415 & ~n37644;
  assign n38027 = ~n38025 & ~n38026;
  assign n38028 = ~n38024 & n38027;
  assign n38029 = ~n38023 & n38028;
  assign n38030 = pi2722 & n37648;
  assign n38031 = pi2712 & n37653;
  assign n38032 = ~n38030 & ~n38031;
  assign n38033 = n38029 & n38032;
  assign n38034 = ~n35660 & ~n38033;
  assign n38035 = pi0672 & n35660;
  assign po0962 = n38034 | n38035;
  assign n38037 = pi2715 & n37653;
  assign n38038 = ~n12061 & ~n37644;
  assign n38039 = pi2773 & n37648;
  assign n38040 = ~n12061 & ~n37658;
  assign n38041 = ~n38039 & ~n38040;
  assign n38042 = ~n38038 & n38041;
  assign n38043 = ~n38037 & n38042;
  assign n38044 = pi2743 & n37661;
  assign n38045 = pi2734 & n37663;
  assign n38046 = ~n38044 & ~n38045;
  assign n38047 = n38043 & n38046;
  assign n38048 = ~n35660 & ~n38047;
  assign n38049 = pi0673 & n35660;
  assign po0963 = n38048 | n38049;
  assign n38051 = pi2560 & n37663;
  assign n38052 = ~n15115 & ~n37644;
  assign n38053 = pi2547 & n37661;
  assign n38054 = ~n15115 & ~n37658;
  assign n38055 = ~n38053 & ~n38054;
  assign n38056 = ~n38052 & n38055;
  assign n38057 = ~n38051 & n38056;
  assign n38058 = pi2724 & n37648;
  assign n38059 = pi2714 & n37653;
  assign n38060 = ~n38058 & ~n38059;
  assign n38061 = n38057 & n38060;
  assign n38062 = ~n35660 & ~n38061;
  assign n38063 = pi0674 & n35660;
  assign po0964 = n38062 | n38063;
  assign n38065 = ~n15426 & ~n37658;
  assign n38066 = pi2545 & n37661;
  assign n38067 = ~n38065 & ~n38066;
  assign n38068 = pi2736 & n37663;
  assign n38069 = n38067 & ~n38068;
  assign n38070 = ~n15426 & ~n37644;
  assign n38071 = n38069 & ~n38070;
  assign n38072 = pi2565 & n37648;
  assign n38073 = pi2534 & n37653;
  assign n38074 = ~n38072 & ~n38073;
  assign n38075 = n38071 & n38074;
  assign n38076 = ~n35660 & ~n38075;
  assign n38077 = pi0675 & n35660;
  assign po0965 = n38076 | n38077;
  assign n38079 = ~n14403 & ~n37658;
  assign n38080 = pi2745 & n37661;
  assign n38081 = ~n38079 & ~n38080;
  assign n38082 = pi2737 & n37663;
  assign n38083 = n38081 & ~n38082;
  assign n38084 = ~n14403 & ~n37644;
  assign n38085 = n38083 & ~n38084;
  assign n38086 = pi2726 & n37648;
  assign n38087 = pi2718 & n37653;
  assign n38088 = ~n38086 & ~n38087;
  assign n38089 = n38085 & n38088;
  assign n38090 = ~n35660 & ~n38089;
  assign n38091 = pi0676 & n35660;
  assign po0966 = n38090 | n38091;
  assign n38093 = n10873 & n13701;
  assign n38094 = ~n10873 & n14087;
  assign n38095 = ~n38093 & ~n38094;
  assign n38096 = ~n10843 & n37639;
  assign n38097 = ~n10835 & n37642;
  assign n38098 = ~n38096 & ~n38097;
  assign n38099 = n38095 & ~n38098;
  assign n38100 = n10850 & n37647;
  assign n38101 = pi2520 & n38100;
  assign n38102 = ~n38099 & ~n38101;
  assign n38103 = n10825 & n37652;
  assign n38104 = pi2535 & n38103;
  assign n38105 = n38102 & ~n38104;
  assign n38106 = ~n10850 & n37647;
  assign n38107 = ~n10825 & n37652;
  assign n38108 = ~n38106 & ~n38107;
  assign n38109 = n38095 & ~n38108;
  assign n38110 = n38105 & ~n38109;
  assign n38111 = n10843 & n37639;
  assign n38112 = pi2752 & n38111;
  assign n38113 = n10835 & n37642;
  assign n38114 = pi2412 & n38113;
  assign n38115 = ~n38112 & ~n38114;
  assign n38116 = n38110 & n38115;
  assign n38117 = ~n35660 & ~n38116;
  assign n38118 = pi0677 & n35660;
  assign po0967 = n38117 | n38118;
  assign n38120 = n10873 & n13988;
  assign n38121 = ~n10873 & n14016;
  assign n38122 = ~n38120 & ~n38121;
  assign n38123 = ~n38108 & n38122;
  assign n38124 = pi2527 & n38100;
  assign n38125 = ~n38123 & ~n38124;
  assign n38126 = pi2746 & n38103;
  assign n38127 = n38125 & ~n38126;
  assign n38128 = ~n38098 & n38122;
  assign n38129 = n38127 & ~n38128;
  assign n38130 = pi2753 & n38111;
  assign n38131 = pi2463 & n38113;
  assign n38132 = ~n38130 & ~n38131;
  assign n38133 = n38129 & n38132;
  assign n38134 = ~n35660 & ~n38133;
  assign n38135 = pi0678 & n35660;
  assign po0968 = n38134 | n38135;
  assign n38137 = n10873 & n12061;
  assign n38138 = ~n10873 & n12106;
  assign n38139 = ~n38137 & ~n38138;
  assign n38140 = ~n38098 & n38139;
  assign n38141 = pi2466 & n38113;
  assign n38142 = ~n38140 & ~n38141;
  assign n38143 = pi2754 & n38111;
  assign n38144 = n38142 & ~n38143;
  assign n38145 = ~n38108 & n38139;
  assign n38146 = n38144 & ~n38145;
  assign n38147 = pi2747 & n38103;
  assign n38148 = pi2457 & n38100;
  assign n38149 = ~n38147 & ~n38148;
  assign n38150 = n38146 & n38149;
  assign n38151 = ~n35660 & ~n38150;
  assign n38152 = pi0679 & n35660;
  assign po0969 = n38151 | n38152;
  assign n38154 = n9825 & n10873;
  assign n38155 = ~n10873 & n11752;
  assign n38156 = ~n38154 & ~n38155;
  assign n38157 = ~n38098 & n38156;
  assign n38158 = pi2410 & n38113;
  assign n38159 = ~n38157 & ~n38158;
  assign n38160 = pi2530 & n38111;
  assign n38161 = n38159 & ~n38160;
  assign n38162 = ~n38108 & n38156;
  assign n38163 = n38161 & ~n38162;
  assign n38164 = pi2748 & n38103;
  assign n38165 = pi2458 & n38100;
  assign n38166 = ~n38164 & ~n38165;
  assign n38167 = n38163 & n38166;
  assign n38168 = ~n35660 & ~n38167;
  assign n38169 = pi0680 & n35660;
  assign po0970 = n38168 | n38169;
  assign n38171 = n10608 & n10873;
  assign n38172 = ~n10873 & n11781;
  assign n38173 = ~n38171 & ~n38172;
  assign n38174 = ~n38108 & n38173;
  assign n38175 = pi2525 & n38100;
  assign n38176 = ~n38174 & ~n38175;
  assign n38177 = pi2533 & n38103;
  assign n38178 = n38176 & ~n38177;
  assign n38179 = ~n38098 & n38173;
  assign n38180 = n38178 & ~n38179;
  assign n38181 = pi2755 & n38111;
  assign n38182 = pi2467 & n38113;
  assign n38183 = ~n38181 & ~n38182;
  assign n38184 = n38180 & n38183;
  assign n38185 = ~n35660 & ~n38184;
  assign n38186 = pi0681 & n35660;
  assign po0971 = n38185 | n38186;
  assign n38188 = n10873 & n15426;
  assign n38189 = ~n10873 & n15454;
  assign n38190 = ~n38188 & ~n38189;
  assign n38191 = ~n38108 & n38190;
  assign n38192 = pi2459 & n38100;
  assign n38193 = ~n38191 & ~n38192;
  assign n38194 = pi2749 & n38103;
  assign n38195 = n38193 & ~n38194;
  assign n38196 = ~n38098 & n38190;
  assign n38197 = n38195 & ~n38196;
  assign n38198 = pi2544 & n38111;
  assign n38199 = pi2468 & n38113;
  assign n38200 = ~n38198 & ~n38199;
  assign n38201 = n38197 & n38200;
  assign n38202 = ~n35660 & ~n38201;
  assign n38203 = pi0682 & n35660;
  assign po0972 = n38202 | n38203;
  assign n38205 = n10873 & n14403;
  assign n38206 = ~n10873 & n14430;
  assign n38207 = ~n38205 & ~n38206;
  assign n38208 = ~n38098 & n38207;
  assign n38209 = pi2460 & n38100;
  assign n38210 = ~n38208 & ~n38209;
  assign n38211 = pi2750 & n38103;
  assign n38212 = n38210 & ~n38211;
  assign n38213 = ~n38108 & n38207;
  assign n38214 = n38212 & ~n38213;
  assign n38215 = pi2756 & n38111;
  assign n38216 = pi2469 & n38113;
  assign n38217 = ~n38215 & ~n38216;
  assign n38218 = n38214 & n38217;
  assign n38219 = ~n35660 & ~n38218;
  assign n38220 = pi0683 & n35660;
  assign po0973 = n38219 | n38220;
  assign n38222 = pi1046 & pi3481;
  assign n38223 = ~pi1931 & ~pi2403;
  assign n38224 = ~pi0570 & pi1931;
  assign n38225 = ~n38223 & ~n38224;
  assign n38226 = pi0918 & ~n38225;
  assign n38227 = pi3641 & n38226;
  assign n38228 = pi0980 & pi3641;
  assign n38229 = ~pi0545 & n38228;
  assign n38230 = ~n38227 & ~n38229;
  assign n38231 = ~pi1931 & ~pi2401;
  assign n38232 = ~pi0546 & pi1931;
  assign n38233 = ~n38231 & ~n38232;
  assign n38234 = pi0919 & ~n38233;
  assign n38235 = pi3641 & n38234;
  assign n38236 = n38230 & ~n38235;
  assign n38237 = ~pi0544 & pi0917;
  assign n38238 = pi3641 & n38237;
  assign n38239 = pi3539 & pi3641;
  assign n38240 = pi0915 & n38239;
  assign n38241 = pi0916 & ~pi1822;
  assign n38242 = pi3641 & n38241;
  assign n38243 = ~n38240 & ~n38242;
  assign n38244 = ~n38238 & n38243;
  assign n38245 = ~pi0648 & pi0708;
  assign n38246 = pi3641 & n38245;
  assign n38247 = ~pi0522 & pi0914;
  assign n38248 = pi3641 & n38247;
  assign n38249 = pi0913 & ~pi2381;
  assign n38250 = pi3641 & n38249;
  assign n38251 = pi0912 & pi3538;
  assign n38252 = pi3641 & n38251;
  assign n38253 = ~pi2402 & pi3641;
  assign n38254 = ~n38252 & ~n38253;
  assign n38255 = ~n38250 & n38254;
  assign n38256 = ~n38248 & n38255;
  assign n38257 = ~n38246 & n38256;
  assign n38258 = n38244 & n38257;
  assign n38259 = n38236 & n38258;
  assign n38260 = ~pi3481 & ~n38259;
  assign n38261 = ~n38222 & ~n38260;
  assign n38262 = ~pi3203 & po3831;
  assign n38263 = ~n38261 & n38262;
  assign n38264 = n9345 & n38263;
  assign n38265 = pi0684 & ~n38262;
  assign po0975 = n38264 | n38265;
  assign n38267 = ~n37332 & ~n37340;
  assign n38268 = ~n37338 & ~n38267;
  assign n38269 = n37332 & n38268;
  assign n38270 = pi0685 & n38267;
  assign po0976 = n38269 | n38270;
  assign n38272 = ~pi0615 & n37332;
  assign n38273 = ~pi0686 & ~n38272;
  assign n38274 = ~n9352 & ~n34965;
  assign po0977 = n38273 | n38274;
  assign n38276 = pi2789 & ~n9352;
  assign n38277 = ~pi3426 & n38276;
  assign n38278 = n9653 & n38277;
  assign n38279 = ~pi0723 & ~pi0724;
  assign n38280 = ~pi0772 & ~pi0782;
  assign n38281 = ~pi0733 & ~pi0787;
  assign n38282 = ~pi0786 & n38281;
  assign n38283 = n38280 & n38282;
  assign n38284 = ~pi0771 & n38283;
  assign n38285 = ~pi0770 & n38284;
  assign n38286 = ~pi0732 & ~pi0769;
  assign n38287 = n38285 & n38286;
  assign n38288 = n38279 & n38287;
  assign n38289 = n36168 & n38288;
  assign n38290 = pi0687 & n38289;
  assign n38291 = ~pi0687 & ~n38289;
  assign n38292 = ~n38290 & ~n38291;
  assign n38293 = ~n36190 & n38292;
  assign n38294 = pi0687 & n36190;
  assign n38295 = ~n38293 & ~n38294;
  assign n38296 = ~n38278 & ~n38295;
  assign n38297 = ~n9825 & n38278;
  assign po0979 = n38296 | n38297;
  assign n38299 = pi0688 & n36181;
  assign n38300 = pi1467 & pi1603;
  assign n38301 = pi2061 & n8598;
  assign n38302 = pi2059 & ~n8598;
  assign n38303 = ~pi2061 & ~n8598;
  assign n38304 = n38302 & ~n38303;
  assign n38305 = ~n38301 & ~n38304;
  assign n38306 = pi2058 & ~n38305;
  assign n38307 = pi1841 & n38306;
  assign n38308 = pi1474 & pi1602;
  assign n38309 = n38307 & n38308;
  assign n38310 = n38300 & n38309;
  assign n38311 = pi0928 & pi1066;
  assign n38312 = n38310 & n38311;
  assign n38313 = pi1090 & n38312;
  assign n38314 = pi0930 & n38313;
  assign n38315 = pi0688 & n38314;
  assign n38316 = ~pi0688 & ~n38314;
  assign n38317 = ~n38315 & ~n38316;
  assign n38318 = ~n36181 & n38317;
  assign n38319 = ~n38299 & ~n38318;
  assign n38320 = n9675 & n38277;
  assign n38321 = ~n38319 & ~n38320;
  assign n38322 = ~n10608 & n38320;
  assign po0981 = n38321 | n38322;
  assign n38324 = pi0689 & ~pi3647;
  assign n38325 = ~pi0689 & n37357;
  assign n38326 = pi0689 & ~n37357;
  assign n38327 = ~n38325 & ~n38326;
  assign n38328 = pi3647 & ~n38327;
  assign n38329 = ~n38324 & ~n38328;
  assign n38330 = n36877 & n38329;
  assign n38331 = pi0871 & n36876;
  assign po0982 = n38330 | n38331;
  assign n38333 = pi0690 & ~pi3635;
  assign n38334 = ~pi0690 & n37376;
  assign n38335 = pi0690 & ~n37376;
  assign n38336 = ~n38334 & ~n38335;
  assign n38337 = pi3635 & ~n38336;
  assign n38338 = ~n38333 & ~n38337;
  assign n38339 = n36969 & n38338;
  assign n38340 = pi0978 & n36968;
  assign po0983 = n38339 | n38340;
  assign n38342 = pi1429 & ~n37393;
  assign n38343 = n37402 & n37404;
  assign n38344 = ~n37405 & ~n38343;
  assign n38345 = pi3641 & ~n38344;
  assign n38346 = ~pi0691 & ~pi3641;
  assign n38347 = ~n38345 & ~n38346;
  assign n38348 = n37390 & ~n38347;
  assign n38349 = ~n37392 & n38348;
  assign po0984 = n38342 | n38349;
  assign n38351 = ~n8561 & ~n36457;
  assign n38352 = pi0692 & n8561;
  assign po0985 = n38351 | n38352;
  assign n38354 = ~pi0693 & ~n37028;
  assign n38355 = pi0958 & ~n8454;
  assign n38356 = ~pi0958 & pi3664;
  assign n38357 = ~n38355 & ~n38356;
  assign n38358 = n37028 & ~n38357;
  assign po0986 = n38354 | n38358;
  assign n38360 = ~pi0694 & ~n37028;
  assign n38361 = ~pi0693 & n37028;
  assign po0987 = n38360 | n38361;
  assign n38363 = ~n36568 & ~n36591;
  assign n38364 = ~n8561 & n38363;
  assign n38365 = ~n36581 & n38364;
  assign n38366 = n36764 & n38365;
  assign n38367 = ~pi0695 & n8561;
  assign n38368 = ~n38366 & ~n38367;
  assign po0988 = po3627 & ~n38368;
  assign n38370 = ~pi0696 & ~n34870;
  assign n38371 = pi0886 & ~n8503;
  assign n38372 = ~pi0886 & pi3665;
  assign n38373 = ~n38371 & ~n38372;
  assign n38374 = n34870 & ~n38373;
  assign po0989 = n38370 | n38374;
  assign n38376 = ~pi0697 & ~n34870;
  assign n38377 = ~pi0696 & n34870;
  assign po0990 = n38376 | n38377;
  assign n38379 = pi0698 & ~pi3635;
  assign n38380 = n37371 & n37373;
  assign n38381 = n37374 & n38380;
  assign n38382 = n37377 & n38381;
  assign n38383 = ~pi0698 & n38382;
  assign n38384 = pi0698 & ~n38382;
  assign n38385 = ~n38383 & ~n38384;
  assign n38386 = pi3635 & ~n38385;
  assign n38387 = ~n38379 & ~n38386;
  assign n38388 = n36969 & n38387;
  assign n38389 = pi0972 & n36968;
  assign po0991 = n38388 | n38389;
  assign n38391 = pi0699 & pi0849;
  assign n38392 = ~n31785 & ~n38391;
  assign n38393 = n31865 & ~n38392;
  assign n38394 = pi3641 & n38393;
  assign n38395 = pi0699 & ~n32073;
  assign n38396 = ~n38394 & ~n38395;
  assign n38397 = ~n31777 & ~n38396;
  assign n38398 = pi1721 & n31777;
  assign n38399 = ~n38397 & ~n38398;
  assign n38400 = ~n31779 & ~n38399;
  assign n38401 = ~pi2396 & n31779;
  assign po0992 = n38400 | n38401;
  assign n38403 = pi2960 & n38103;
  assign n38404 = pi2452 & n38100;
  assign n38405 = ~n38403 & ~n38404;
  assign n38406 = pi2965 & n38111;
  assign n38407 = pi2413 & n38113;
  assign n38408 = ~n38406 & ~n38407;
  assign n38409 = n38405 & n38408;
  assign n38410 = n38098 & n38108;
  assign n38411 = n10873 & ~n12726;
  assign n38412 = ~n10873 & ~n12751;
  assign n38413 = ~n38411 & ~n38412;
  assign n38414 = ~n38410 & ~n38413;
  assign n38415 = n38409 & ~n38414;
  assign n38416 = ~n35660 & ~n38415;
  assign n38417 = pi0701 & n35660;
  assign po0994 = n38416 | n38417;
  assign n38419 = pi2961 & n38103;
  assign n38420 = pi2453 & n38100;
  assign n38421 = ~n38419 & ~n38420;
  assign n38422 = pi3096 & n38111;
  assign n38423 = pi2461 & n38113;
  assign n38424 = ~n38422 & ~n38423;
  assign n38425 = n38421 & n38424;
  assign n38426 = n10873 & ~n13121;
  assign n38427 = ~n10873 & ~n13149;
  assign n38428 = ~n38426 & ~n38427;
  assign n38429 = ~n38410 & ~n38428;
  assign n38430 = n38425 & ~n38429;
  assign n38431 = ~n35660 & ~n38430;
  assign n38432 = pi0702 & n35660;
  assign po0995 = n38431 | n38432;
  assign n38434 = pi2962 & n38103;
  assign n38435 = pi2454 & n38100;
  assign n38436 = ~n38434 & ~n38435;
  assign n38437 = pi3093 & n38111;
  assign n38438 = pi2462 & n38113;
  assign n38439 = ~n38437 & ~n38438;
  assign n38440 = n38436 & n38439;
  assign n38441 = n10873 & ~n13398;
  assign n38442 = ~n10873 & ~n12862;
  assign n38443 = ~n38441 & ~n38442;
  assign n38444 = ~n38410 & ~n38443;
  assign n38445 = n38440 & ~n38444;
  assign n38446 = ~n35660 & ~n38445;
  assign n38447 = pi0703 & n35660;
  assign po0996 = n38446 | n38447;
  assign n38449 = pi2963 & n38103;
  assign n38450 = pi2455 & n38100;
  assign n38451 = ~n38449 & ~n38450;
  assign n38452 = pi2966 & n38111;
  assign n38453 = pi2464 & n38113;
  assign n38454 = ~n38452 & ~n38453;
  assign n38455 = n38451 & n38454;
  assign n38456 = n10873 & ~n12415;
  assign n38457 = ~n10873 & ~n12485;
  assign n38458 = ~n38456 & ~n38457;
  assign n38459 = ~n38410 & ~n38458;
  assign n38460 = n38455 & ~n38459;
  assign n38461 = ~n35660 & ~n38460;
  assign n38462 = pi0704 & n35660;
  assign po0997 = n38461 | n38462;
  assign n38464 = pi2780 & n38103;
  assign n38465 = pi2456 & n38100;
  assign n38466 = ~n38464 & ~n38465;
  assign n38467 = pi2810 & n38111;
  assign n38468 = pi2465 & n38113;
  assign n38469 = ~n38467 & ~n38468;
  assign n38470 = n38466 & n38469;
  assign n38471 = n10873 & ~n14816;
  assign n38472 = ~n10873 & ~n14537;
  assign n38473 = ~n38471 & ~n38472;
  assign n38474 = ~n38410 & ~n38473;
  assign n38475 = n38470 & ~n38474;
  assign n38476 = ~n35660 & ~n38475;
  assign n38477 = pi0705 & n35660;
  assign po0998 = n38476 | n38477;
  assign n38479 = pi2776 & n38103;
  assign n38480 = pi2526 & n38100;
  assign n38481 = ~n38479 & ~n38480;
  assign n38482 = pi2967 & n38111;
  assign n38483 = pi2411 & n38113;
  assign n38484 = ~n38482 & ~n38483;
  assign n38485 = n38481 & n38484;
  assign n38486 = n10873 & ~n15115;
  assign n38487 = ~n10873 & ~n15187;
  assign n38488 = ~n38486 & ~n38487;
  assign n38489 = ~n38410 & ~n38488;
  assign n38490 = n38485 & ~n38489;
  assign n38491 = ~n35660 & ~n38490;
  assign n38492 = pi0706 & n35660;
  assign po0999 = n38491 | n38492;
  assign n38494 = pi2968 & n38111;
  assign n38495 = pi2470 & n38113;
  assign n38496 = ~n38494 & ~n38495;
  assign n38497 = pi2964 & n38103;
  assign n38498 = pi2524 & n38100;
  assign n38499 = ~n38497 & ~n38498;
  assign n38500 = n38496 & n38499;
  assign n38501 = n10873 & ~n11181;
  assign n38502 = ~n10873 & ~n11674;
  assign n38503 = ~n38501 & ~n38502;
  assign n38504 = ~n38410 & ~n38503;
  assign n38505 = n38500 & ~n38504;
  assign n38506 = ~n35660 & ~n38505;
  assign n38507 = pi0707 & n35660;
  assign po1000 = n38506 | n38507;
  assign n38509 = pi3641 & po3948;
  assign n38510 = ~pi1523 & n20345;
  assign n38511 = ~pi1415 & n20347;
  assign n38512 = ~n38510 & ~n38511;
  assign n38513 = ~pi1590 & n20350;
  assign n38514 = ~pi1619 & n20353;
  assign n38515 = ~pi1558 & n20356;
  assign n38516 = ~n38514 & ~n38515;
  assign n38517 = ~pi1624 & n20360;
  assign n38518 = ~pi1486 & n20363;
  assign n38519 = ~n38517 & ~n38518;
  assign n38520 = n38516 & n38519;
  assign n38521 = ~n38513 & n38520;
  assign n38522 = n38512 & n38521;
  assign n38523 = ~pi1007 & ~n38522;
  assign n38524 = pi1007 & ~n14816;
  assign n38525 = ~n38523 & ~n38524;
  assign n38526 = pi1007 & ~n9352;
  assign n38527 = ~n19551 & ~n38526;
  assign n38528 = n38525 & ~n38527;
  assign n38529 = ~pi0708 & n38527;
  assign n38530 = ~n38528 & ~n38529;
  assign n38531 = ~n38509 & n38530;
  assign n38532 = pi0708 & n38509;
  assign n38533 = pi1048 & pi3293;
  assign n38534 = n38532 & n38533;
  assign n38535 = ~n38531 & ~n38534;
  assign n38536 = pi1049 & pi3293;
  assign n38537 = pi1330 & pi3293;
  assign n38538 = ~n38536 & ~n38537;
  assign n38539 = n38532 & ~n38538;
  assign po1001 = ~n38535 | n38539;
  assign n38541 = ~n8561 & n36622;
  assign n38542 = n36763 & n38541;
  assign n38543 = ~n36581 & n36637;
  assign n38544 = n38542 & n38543;
  assign n38545 = pi0709 & n8561;
  assign n38546 = ~n38544 & ~n38545;
  assign po1002 = po3627 & ~n38546;
  assign n38548 = n36621 & n38541;
  assign n38549 = n38543 & n38548;
  assign n38550 = pi0710 & n8561;
  assign n38551 = ~n38549 & ~n38550;
  assign po1003 = po3627 & ~n38551;
  assign n38553 = ~n36568 & n36591;
  assign n38554 = ~n36581 & n38553;
  assign n38555 = n38548 & n38554;
  assign n38556 = ~pi0711 & n8561;
  assign n38557 = ~n38555 & ~n38556;
  assign po1004 = po3627 & ~n38557;
  assign n38559 = n38542 & n38554;
  assign n38560 = ~pi0712 & n8561;
  assign n38561 = ~n38559 & ~n38560;
  assign po1005 = po3627 & ~n38561;
  assign n38563 = ~n36581 & n36775;
  assign n38564 = n38542 & n38563;
  assign n38565 = ~pi0713 & n8561;
  assign n38566 = ~n38564 & ~n38565;
  assign po1006 = po3627 & ~n38566;
  assign n38568 = n38548 & n38563;
  assign n38569 = ~pi0714 & n8561;
  assign n38570 = ~n38568 & ~n38569;
  assign po1007 = po3627 & ~n38570;
  assign n38572 = n36623 & n38365;
  assign n38573 = pi0715 & n8561;
  assign n38574 = ~n38572 & ~n38573;
  assign po1008 = po3627 & ~n38574;
  assign n38576 = pi0716 & n8561;
  assign n38577 = ~n8561 & n36000;
  assign po1009 = n38576 | n38577;
  assign n38579 = pi0717 & n8561;
  assign n38580 = ~n8561 & n35989;
  assign po1010 = n38579 | n38580;
  assign n38582 = ~n8561 & n35987;
  assign n38583 = pi0718 & n8561;
  assign po1011 = n38582 | n38583;
  assign n38585 = pi0719 & n8561;
  assign n38586 = ~n8561 & n35860;
  assign po1012 = n38585 | n38586;
  assign n38588 = pi0720 & n8561;
  assign n38589 = ~n8561 & n35883;
  assign po1013 = n38588 | n38589;
  assign n38591 = ~n8561 & n35881;
  assign n38592 = pi0721 & n8561;
  assign po1014 = n38591 | n38592;
  assign n38594 = pi0722 & n8561;
  assign n38595 = ~pi0414 & n35997;
  assign n38596 = ~n35837 & n35991;
  assign n38597 = n37727 & n38596;
  assign n38598 = n38595 & n38597;
  assign n38599 = n35997 & n38596;
  assign n38600 = n35994 & n38599;
  assign n38601 = n35994 & n38596;
  assign n38602 = n36046 & n38601;
  assign n38603 = n37728 & n38597;
  assign n38604 = ~n38602 & ~n38603;
  assign n38605 = ~n38600 & n38604;
  assign n38606 = ~n38598 & n38605;
  assign n38607 = ~n8561 & ~n38606;
  assign n38608 = ~n38594 & ~n38607;
  assign n38609 = n20460 & n38596;
  assign n38610 = n37728 & n38609;
  assign n38611 = n38595 & n38609;
  assign n38612 = n20417 & n38599;
  assign n38613 = ~pi0414 & n38612;
  assign n38614 = n20417 & n38596;
  assign n38615 = n37728 & n38614;
  assign n38616 = ~n38613 & ~n38615;
  assign n38617 = ~n38611 & n38616;
  assign n38618 = ~n38610 & n38617;
  assign n38619 = pi0414 & n36046;
  assign n38620 = n38614 & n38619;
  assign n38621 = n38609 & n38619;
  assign n38622 = n35997 & n38609;
  assign n38623 = pi0414 & n38622;
  assign n38624 = pi0414 & n38612;
  assign n38625 = ~n38623 & ~n38624;
  assign n38626 = ~n38621 & n38625;
  assign n38627 = ~n38620 & n38626;
  assign n38628 = n38618 & n38627;
  assign n38629 = ~n8561 & ~n38628;
  assign po1015 = ~n38608 | n38629;
  assign n38631 = ~pi0723 & ~n38287;
  assign n38632 = pi0723 & n38287;
  assign n38633 = ~n38631 & ~n38632;
  assign n38634 = ~n36190 & n38633;
  assign n38635 = pi0723 & n36190;
  assign n38636 = ~n38634 & ~n38635;
  assign n38637 = ~n38278 & ~n38636;
  assign n38638 = ~n12726 & n38278;
  assign po1016 = n38637 | n38638;
  assign n38640 = ~pi0772 & n38282;
  assign n38641 = ~pi0782 & n38640;
  assign n38642 = n36193 & n38641;
  assign n38643 = ~pi0771 & n38642;
  assign n38644 = n36192 & n38643;
  assign n38645 = n36168 & n38644;
  assign n38646 = pi0724 & n38645;
  assign n38647 = ~pi0724 & ~n38645;
  assign n38648 = ~n38646 & ~n38647;
  assign n38649 = ~n36190 & n38648;
  assign n38650 = pi0724 & n36190;
  assign n38651 = ~n38649 & ~n38650;
  assign n38652 = ~n38278 & ~n38651;
  assign n38653 = ~n10608 & n38278;
  assign po1017 = n38652 | n38653;
  assign n38655 = ~pi0726 & ~pi0769;
  assign n38656 = ~pi0770 & ~pi0771;
  assign n38657 = n38641 & n38656;
  assign n38658 = n38655 & n38657;
  assign n38659 = n36192 & n38658;
  assign n38660 = pi0725 & n38659;
  assign n38661 = ~pi0725 & ~n38659;
  assign n38662 = ~n38660 & ~n38661;
  assign n38663 = ~n36190 & n38662;
  assign n38664 = pi0725 & n36190;
  assign n38665 = ~n38663 & ~n38664;
  assign n38666 = ~n38278 & ~n38665;
  assign n38667 = ~n15426 & n38278;
  assign po1018 = n38666 | n38667;
  assign n38669 = n36172 & n38281;
  assign n38670 = n36194 & n38669;
  assign n38671 = pi0726 & n38670;
  assign n38672 = ~pi0726 & ~n38670;
  assign n38673 = ~n38671 & ~n38672;
  assign n38674 = ~n36190 & n38673;
  assign n38675 = pi0726 & n36190;
  assign n38676 = ~n38674 & ~n38675;
  assign n38677 = ~n38278 & ~n38676;
  assign n38678 = ~n14403 & n38278;
  assign po1019 = n38677 | n38678;
  assign n38680 = pi0727 & ~pi3647;
  assign n38681 = n37353 & n37354;
  assign n38682 = n37355 & n38681;
  assign n38683 = n37358 & n38682;
  assign n38684 = ~pi0727 & n38683;
  assign n38685 = pi0727 & ~n38683;
  assign n38686 = ~n38684 & ~n38685;
  assign n38687 = pi3647 & ~n38686;
  assign n38688 = ~n38680 & ~n38687;
  assign n38689 = n36877 & n38688;
  assign n38690 = pi0897 & n36876;
  assign po1020 = n38689 | n38690;
  assign n38692 = ~pi0728 & n31785;
  assign n38693 = pi0728 & ~n31785;
  assign n38694 = ~n38692 & ~n38693;
  assign n38695 = n31865 & ~n38694;
  assign n38696 = pi3641 & n38695;
  assign n38697 = pi0728 & ~n32073;
  assign n38698 = ~n38696 & ~n38697;
  assign n38699 = ~n31777 & ~n38698;
  assign n38700 = pi1720 & n31777;
  assign n38701 = ~n38699 & ~n38700;
  assign n38702 = ~n31779 & ~n38701;
  assign n38703 = ~pi2094 & n31779;
  assign po1021 = n38702 | n38703;
  assign n38705 = pi3502 & pi3506;
  assign n38706 = pi3425 & n38705;
  assign n38707 = pi3425 & ~pi3506;
  assign n38708 = pi3502 & ~pi3677;
  assign n38709 = n38707 & n38708;
  assign n38710 = ~n38706 & ~n38709;
  assign n38711 = ~pi3502 & pi3506;
  assign n38712 = ~pi3425 & n38711;
  assign n38713 = ~pi3425 & ~pi3506;
  assign n38714 = pi3502 & n38713;
  assign n38715 = ~n38712 & ~n38714;
  assign n38716 = pi3677 & ~n38715;
  assign n38717 = n38710 & ~n38716;
  assign n38718 = pi3425 & n38711;
  assign n38719 = ~pi3677 & n38718;
  assign n38720 = ~pi3502 & ~pi3677;
  assign n38721 = n38707 & n38720;
  assign n38722 = ~n38719 & ~n38721;
  assign n38723 = n38717 & n38722;
  assign n38724 = ~n38706 & ~n38714;
  assign n38725 = ~pi3425 & pi3506;
  assign n38726 = ~n38707 & ~n38725;
  assign n38727 = n38708 & ~n38726;
  assign n38728 = ~pi3677 & ~n38712;
  assign n38729 = pi3677 & ~n38718;
  assign n38730 = ~n38728 & ~n38729;
  assign n38731 = ~n38727 & ~n38730;
  assign n38732 = n38724 & n38731;
  assign n38733 = ~n38723 & ~n38732;
  assign n38734 = ~pi3677 & n38706;
  assign n38735 = n38713 & n38720;
  assign n38736 = ~n38734 & ~n38735;
  assign n38737 = n38708 & n38725;
  assign n38738 = n38722 & ~n38737;
  assign n38739 = ~pi3677 & n38714;
  assign n38740 = ~n38709 & ~n38739;
  assign n38741 = n38738 & n38740;
  assign n38742 = n38736 & n38741;
  assign n38743 = n38723 & ~n38742;
  assign n38744 = ~n38732 & n38743;
  assign n38745 = ~n38733 & ~n38744;
  assign n38746 = pi0730 & n38745;
  assign n38747 = pi3266 & pi3271;
  assign n38748 = ~pi3246 & pi3255;
  assign n38749 = n38747 & n38748;
  assign n38750 = ~pi2881 & n38749;
  assign n38751 = ~pi3266 & pi3271;
  assign n38752 = n38748 & n38751;
  assign n38753 = ~pi3049 & n38752;
  assign n38754 = ~n38750 & ~n38753;
  assign n38755 = pi3246 & pi3255;
  assign n38756 = pi3266 & ~pi3271;
  assign n38757 = n38755 & n38756;
  assign n38758 = ~pi2995 & n38757;
  assign n38759 = ~pi3266 & ~pi3271;
  assign n38760 = n38748 & n38759;
  assign n38761 = ~pi3018 & n38760;
  assign n38762 = ~n38758 & ~n38761;
  assign n38763 = ~pi3246 & ~pi3255;
  assign n38764 = n38751 & n38763;
  assign n38765 = ~pi2761 & n38764;
  assign n38766 = n38755 & n38759;
  assign n38767 = ~pi3011 & n38766;
  assign n38768 = ~n38765 & ~n38767;
  assign n38769 = n38759 & n38763;
  assign n38770 = n38751 & n38755;
  assign n38771 = ~pi2898 & n38770;
  assign n38772 = n38748 & n38756;
  assign n38773 = ~pi3004 & n38772;
  assign n38774 = ~n38771 & ~n38773;
  assign n38775 = n38747 & n38755;
  assign n38776 = ~pi3090 & n38775;
  assign n38777 = n38774 & ~n38776;
  assign n38778 = pi3246 & ~pi3255;
  assign n38779 = n38747 & n38778;
  assign n38780 = ~pi1386 & n38779;
  assign n38781 = n38747 & n38763;
  assign n38782 = ~pi1361 & n38781;
  assign n38783 = ~n38780 & ~n38782;
  assign n38784 = n38777 & n38783;
  assign n38785 = ~n38769 & n38784;
  assign n38786 = n38768 & n38785;
  assign n38787 = n38751 & n38778;
  assign n38788 = pi0812 & n38787;
  assign n38789 = n38756 & n38778;
  assign n38790 = pi0406 & n38789;
  assign n38791 = ~n38788 & ~n38790;
  assign n38792 = n38756 & n38763;
  assign n38793 = pi0381 & n38792;
  assign n38794 = n38791 & ~n38793;
  assign n38795 = n38786 & n38794;
  assign n38796 = n38762 & n38795;
  assign n38797 = n38754 & n38796;
  assign n38798 = n38733 & n38742;
  assign n38799 = ~n38797 & n38798;
  assign n38800 = n38733 & ~n38742;
  assign n38801 = pi0731 & n38800;
  assign n38802 = pi0859 & ~n38800;
  assign n38803 = ~n38801 & ~n38802;
  assign n38804 = ~n38798 & ~n38803;
  assign n38805 = ~n38799 & ~n38804;
  assign n38806 = ~n38745 & ~n38805;
  assign po1024 = n38746 | n38806;
  assign n38808 = pi0731 & n38745;
  assign n38809 = ~pi3035 & n38749;
  assign n38810 = ~pi3050 & n38752;
  assign n38811 = ~n38809 & ~n38810;
  assign n38812 = ~pi2900 & n38757;
  assign n38813 = ~pi2956 & n38760;
  assign n38814 = ~n38812 & ~n38813;
  assign n38815 = ~pi2884 & n38772;
  assign n38816 = ~pi3092 & n38770;
  assign n38817 = ~n38815 & ~n38816;
  assign n38818 = ~pi3027 & n38775;
  assign n38819 = n38817 & ~n38818;
  assign n38820 = ~pi2643 & n38764;
  assign n38821 = ~pi3056 & n38766;
  assign n38822 = ~n38820 & ~n38821;
  assign n38823 = ~pi1363 & n38779;
  assign n38824 = ~pi1701 & n38781;
  assign n38825 = ~n38823 & ~n38824;
  assign n38826 = n38822 & n38825;
  assign n38827 = ~n38769 & n38826;
  assign n38828 = n38819 & n38827;
  assign n38829 = pi0813 & n38787;
  assign n38830 = pi0425 & n38789;
  assign n38831 = ~n38829 & ~n38830;
  assign n38832 = pi0391 & n38792;
  assign n38833 = n38831 & ~n38832;
  assign n38834 = n38828 & n38833;
  assign n38835 = n38814 & n38834;
  assign n38836 = n38811 & n38835;
  assign n38837 = n38798 & ~n38836;
  assign n38838 = pi0938 & n38800;
  assign n38839 = pi0730 & ~n38800;
  assign n38840 = ~n38838 & ~n38839;
  assign n38841 = ~n38798 & ~n38840;
  assign n38842 = ~n38837 & ~n38841;
  assign n38843 = ~n38745 & ~n38842;
  assign po1025 = n38808 | n38843;
  assign n38845 = pi0732 & n38643;
  assign n38846 = ~pi0732 & ~n38643;
  assign n38847 = ~n38845 & ~n38846;
  assign n38848 = ~n36190 & n38847;
  assign n38849 = pi0732 & n36190;
  assign n38850 = ~n38848 & ~n38849;
  assign n38851 = ~n38278 & ~n38850;
  assign n38852 = ~n13701 & n38278;
  assign po1026 = n38851 | n38852;
  assign n38854 = pi0733 & ~n38278;
  assign n38855 = n36190 & n38854;
  assign n38856 = ~n12061 & n38278;
  assign n38857 = ~n38855 & ~n38856;
  assign n38858 = pi0733 & pi0787;
  assign n38859 = ~n38281 & ~n38858;
  assign n38860 = ~n36190 & ~n38859;
  assign n38861 = ~n38278 & n38860;
  assign po1027 = ~n38857 | n38861;
  assign n38863 = ~n8561 & n36100;
  assign n38864 = n36095 & n38863;
  assign n38865 = n36094 & n38864;
  assign n38866 = ~n36083 & n38865;
  assign n38867 = ~pi0734 & n8561;
  assign n38868 = ~n38866 & ~n38867;
  assign po1028 = po3627 & ~n38868;
  assign n38870 = pi2697 & n37287;
  assign n38871 = pi2686 & n37289;
  assign n38872 = ~n38870 & ~n38871;
  assign n38873 = pi2673 & n37274;
  assign n38874 = pi2659 & n37279;
  assign n38875 = ~n38873 & ~n38874;
  assign n38876 = n38872 & n38875;
  assign n38877 = n37270 & n37284;
  assign n38878 = ~n14403 & ~n38877;
  assign n38879 = n38876 & ~n38878;
  assign n38880 = ~n35539 & ~n38879;
  assign n38881 = pi0735 & n35539;
  assign po1029 = n38880 | n38881;
  assign n38883 = pi2665 & n37274;
  assign n38884 = pi2651 & n37279;
  assign n38885 = ~n38883 & ~n38884;
  assign n38886 = pi2689 & n37287;
  assign n38887 = pi2679 & n37289;
  assign n38888 = ~n38886 & ~n38887;
  assign n38889 = n38885 & n38888;
  assign n38890 = ~n13988 & ~n38877;
  assign n38891 = n38889 & ~n38890;
  assign n38892 = ~n35539 & ~n38891;
  assign n38893 = pi0736 & n35539;
  assign po1030 = n38892 | n38893;
  assign n38895 = pi1013 & pi1032;
  assign n38896 = pi1030 & n38895;
  assign n38897 = pi1031 & n38896;
  assign n38898 = n9641 & n38897;
  assign n38899 = pi1033 & n9700;
  assign n38900 = ~pi1039 & n38899;
  assign n38901 = n38898 & n38900;
  assign n38902 = ~n17199 & n38277;
  assign n38903 = n38901 & n38902;
  assign n38904 = pi0609 & n38903;
  assign n38905 = pi0609 & n38277;
  assign n38906 = n38898 & n38905;
  assign n38907 = n9649 & n9666;
  assign n38908 = n38906 & n38907;
  assign n38909 = ~n38904 & ~n38908;
  assign n38910 = pi0737 & n38909;
  assign n38911 = ~n15115 & ~n38909;
  assign n38912 = ~n38910 & ~n38911;
  assign n38913 = n38903 & ~n38909;
  assign po1031 = ~n38912 | n38913;
  assign n38915 = n9673 & n38906;
  assign n38916 = ~n38904 & ~n38915;
  assign n38917 = pi0738 & n38916;
  assign n38918 = ~n12726 & ~n38916;
  assign n38919 = ~n38917 & ~n38918;
  assign n38920 = n38903 & ~n38916;
  assign po1032 = ~n38919 | n38920;
  assign n38922 = pi0739 & n38916;
  assign n38923 = ~n12061 & ~n38916;
  assign n38924 = ~n38922 & ~n38923;
  assign po1033 = n38920 | ~n38924;
  assign n38926 = pi0740 & n38916;
  assign n38927 = ~n14403 & ~n38916;
  assign n38928 = ~n38926 & ~n38927;
  assign po1034 = n38920 | ~n38928;
  assign n38930 = pi0741 & n38916;
  assign n38931 = ~n11181 & ~n38916;
  assign n38932 = ~n38930 & ~n38931;
  assign po1035 = n38920 | ~n38932;
  assign n38934 = pi0742 & n38909;
  assign n38935 = ~n13121 & ~n38909;
  assign n38936 = ~n38934 & ~n38935;
  assign po1036 = n38913 | ~n38936;
  assign n38938 = pi0743 & n38909;
  assign n38939 = ~n13398 & ~n38909;
  assign n38940 = ~n38938 & ~n38939;
  assign po1037 = n38913 | ~n38940;
  assign n38942 = pi0744 & n38909;
  assign n38943 = ~n13988 & ~n38909;
  assign n38944 = ~n38942 & ~n38943;
  assign po1038 = n38913 | ~n38944;
  assign n38946 = pi0745 & n38909;
  assign n38947 = ~n12415 & ~n38909;
  assign n38948 = ~n38946 & ~n38947;
  assign po1039 = n38913 | ~n38948;
  assign n38950 = pi0746 & n38909;
  assign n38951 = ~n14816 & ~n38909;
  assign n38952 = ~n38950 & ~n38951;
  assign po1040 = n38913 | ~n38952;
  assign n38954 = pi0747 & n38909;
  assign n38955 = ~n12061 & ~n38909;
  assign n38956 = ~n38954 & ~n38955;
  assign po1041 = n38913 | ~n38956;
  assign n38958 = pi0748 & n38909;
  assign n38959 = ~n11181 & ~n38909;
  assign n38960 = ~n38958 & ~n38959;
  assign po1042 = n38913 | ~n38960;
  assign n38962 = n9669 & n38277;
  assign n38963 = ~n11181 & n38962;
  assign n38964 = pi0749 & ~n36190;
  assign n38965 = ~pi0749 & n36190;
  assign n38966 = ~n38964 & ~n38965;
  assign n38967 = ~n38962 & n38966;
  assign po1043 = n38963 | n38967;
  assign n38969 = ~n27705 & n31382;
  assign n38970 = pi0750 & n31381;
  assign n38971 = ~n24488 & n31384;
  assign n38972 = pi0750 & ~n31384;
  assign n38973 = ~n38971 & ~n38972;
  assign n38974 = n31388 & ~n38973;
  assign n38975 = ~n38970 & ~n38974;
  assign n38976 = ~n31391 & n38975;
  assign n38977 = ~n31382 & ~n38976;
  assign po1044 = n38969 | n38977;
  assign n38979 = ~n27705 & n31400;
  assign n38980 = pi0751 & n31399;
  assign n38981 = ~n24488 & n31402;
  assign n38982 = pi0751 & ~n31402;
  assign n38983 = ~n38981 & ~n38982;
  assign n38984 = n31406 & ~n38983;
  assign n38985 = ~n38980 & ~n38984;
  assign n38986 = ~n31409 & n38985;
  assign n38987 = ~n31400 & ~n38986;
  assign po1045 = n38979 | n38987;
  assign n38989 = pi0752 & n36190;
  assign n38990 = pi0777 & pi0778;
  assign n38991 = pi0775 & n38990;
  assign n38992 = pi0776 & n38991;
  assign n38993 = pi0749 & n38992;
  assign n38994 = pi0781 & n38993;
  assign n38995 = pi0773 & pi0774;
  assign n38996 = pi0861 & n38995;
  assign n38997 = pi0862 & n38996;
  assign n38998 = n38994 & n38997;
  assign n38999 = pi0780 & n38998;
  assign n39000 = pi0845 & n38999;
  assign n39001 = pi0779 & n39000;
  assign n39002 = pi0752 & n39001;
  assign n39003 = ~pi0752 & ~n39001;
  assign n39004 = ~n39002 & ~n39003;
  assign n39005 = ~n36190 & n39004;
  assign n39006 = ~n38989 & ~n39005;
  assign n39007 = ~n38962 & ~n39006;
  assign n39008 = ~n9825 & n38962;
  assign po1046 = n39007 | n39008;
  assign n39010 = pi2694 & n37287;
  assign n39011 = pi2684 & n37289;
  assign n39012 = ~n39010 & ~n39011;
  assign n39013 = pi2670 & n37274;
  assign n39014 = pi2656 & n37279;
  assign n39015 = ~n39013 & ~n39014;
  assign n39016 = n39012 & n39015;
  assign n39017 = ~n9825 & ~n38877;
  assign n39018 = n39016 & ~n39017;
  assign n39019 = ~n35539 & ~n39018;
  assign n39020 = pi0753 & n35539;
  assign po1047 = n39019 | n39020;
  assign n39022 = pi2701 & n37594;
  assign n39023 = pi2275 & n37591;
  assign n39024 = ~n39022 & ~n39023;
  assign n39025 = pi2698 & n37602;
  assign n39026 = pi2438 & n37604;
  assign n39027 = ~n39025 & ~n39026;
  assign n39028 = n39024 & n39027;
  assign n39029 = n37589 & n37599;
  assign n39030 = n9361 & ~n13701;
  assign n39031 = ~n9361 & ~n14134;
  assign n39032 = ~n39030 & ~n39031;
  assign n39033 = ~n39029 & ~n39032;
  assign n39034 = n39028 & ~n39033;
  assign n39035 = ~n35539 & ~n39034;
  assign n39036 = pi0754 & n35539;
  assign po1048 = n39035 | n39036;
  assign n39038 = pi2699 & n37602;
  assign n39039 = pi2439 & n37604;
  assign n39040 = ~n39038 & ~n39039;
  assign n39041 = pi2702 & n37594;
  assign n39042 = pi2276 & n37591;
  assign n39043 = ~n39041 & ~n39042;
  assign n39044 = n39040 & n39043;
  assign n39045 = ~n9361 & ~n12785;
  assign n39046 = n9361 & ~n13121;
  assign n39047 = ~n39045 & ~n39046;
  assign n39048 = ~n39029 & ~n39047;
  assign n39049 = n39044 & ~n39048;
  assign n39050 = ~n35539 & ~n39049;
  assign n39051 = pi0755 & n35539;
  assign po1049 = n39050 | n39051;
  assign n39053 = pi2703 & n37594;
  assign n39054 = pi2277 & n37591;
  assign n39055 = ~n39053 & ~n39054;
  assign n39056 = pi2539 & n37602;
  assign n39057 = pi2440 & n37604;
  assign n39058 = ~n39056 & ~n39057;
  assign n39059 = n39055 & n39058;
  assign n39060 = n9361 & ~n15426;
  assign n39061 = ~n9361 & ~n15146;
  assign n39062 = ~n39060 & ~n39061;
  assign n39063 = ~n39029 & ~n39062;
  assign n39064 = n39059 & ~n39063;
  assign n39065 = ~n35539 & ~n39064;
  assign n39066 = pi0756 & n35539;
  assign po1050 = n39065 | n39066;
  assign n39068 = pi2751 & n37594;
  assign n39069 = pi2278 & n37591;
  assign n39070 = ~n39068 & ~n39069;
  assign n39071 = pi2700 & n37602;
  assign n39072 = pi2441 & n37604;
  assign n39073 = ~n39071 & ~n39072;
  assign n39074 = n39070 & n39073;
  assign n39075 = n9361 & ~n14403;
  assign n39076 = ~n9361 & ~n14458;
  assign n39077 = ~n39075 & ~n39076;
  assign n39078 = ~n39029 & ~n39077;
  assign n39079 = n39074 & ~n39078;
  assign n39080 = ~n35539 & ~n39079;
  assign n39081 = pi0757 & n35539;
  assign po1051 = n39080 | n39081;
  assign n39083 = ~n8561 & n36105;
  assign n39084 = n36100 & n39083;
  assign n39085 = n36095 & n39084;
  assign n39086 = ~n36083 & n39085;
  assign n39087 = ~pi0758 & n8561;
  assign n39088 = ~n39086 & ~n39087;
  assign po1052 = po3627 & ~n39088;
  assign n39090 = n36060 & n36104;
  assign n39091 = pi0759 & n36128;
  assign po1053 = n39090 | n39091;
  assign n39093 = ~n36080 & n36083;
  assign n39094 = ~n8561 & n36078;
  assign n39095 = n39093 & n39094;
  assign n39096 = ~n36066 & n36069;
  assign n39097 = n39095 & n39096;
  assign n39098 = n36063 & n39097;
  assign n39099 = ~pi0760 & n8561;
  assign n39100 = ~n39098 & ~n39099;
  assign po1054 = po3627 & ~n39100;
  assign n39102 = pi0761 & n8561;
  assign n39103 = ~n8561 & n35984;
  assign po1055 = n39102 | n39103;
  assign n39105 = pi0414 & n35992;
  assign n39106 = n37747 & n39105;
  assign n39107 = n36538 & n39105;
  assign n39108 = n37743 & n38619;
  assign n39109 = n37741 & n38619;
  assign n39110 = ~n39108 & ~n39109;
  assign n39111 = ~n39107 & n39110;
  assign n39112 = ~n39106 & n39111;
  assign n39113 = ~n8561 & ~n39112;
  assign n39114 = pi0762 & n8561;
  assign po1056 = n39113 | n39114;
  assign n39116 = pi0763 & n8561;
  assign n39117 = ~n8561 & n35867;
  assign po1057 = n39116 | n39117;
  assign n39119 = pi0764 & n8561;
  assign n39120 = ~n8561 & n35865;
  assign po1058 = n39119 | n39120;
  assign n39122 = ~n8561 & n35874;
  assign n39123 = pi0765 & n8561;
  assign po1059 = n39122 | n39123;
  assign n39125 = ~n8561 & n35872;
  assign n39126 = pi0766 & n8561;
  assign po1060 = n39125 | n39126;
  assign n39128 = pi0767 & n8561;
  assign n39129 = ~n8561 & n36536;
  assign po1061 = n39128 | n39129;
  assign n39131 = pi0768 & n8561;
  assign n39132 = ~n8561 & n36551;
  assign po1062 = n39131 | n39132;
  assign n39134 = ~n13121 & n38278;
  assign n39135 = pi0769 & n36190;
  assign n39136 = ~pi0769 & ~n38657;
  assign n39137 = pi0769 & n38657;
  assign n39138 = ~n39136 & ~n39137;
  assign n39139 = ~n36190 & n39138;
  assign n39140 = ~n39135 & ~n39139;
  assign n39141 = ~n38278 & ~n39140;
  assign po1063 = n39134 | n39141;
  assign n39143 = ~n13398 & n38278;
  assign n39144 = pi0770 & n36190;
  assign n39145 = ~pi0770 & ~n38669;
  assign n39146 = pi0770 & n38669;
  assign n39147 = ~n39145 & ~n39146;
  assign n39148 = ~n36190 & n39147;
  assign n39149 = ~n39144 & ~n39148;
  assign n39150 = ~n38278 & ~n39149;
  assign po1064 = n39143 | n39150;
  assign n39152 = ~pi3651 & ~pi3652;
  assign po1065 = pi3525 | n39152;
  assign n39154 = ~pi3525 & ~pi3651;
  assign po1066 = pi3652 | ~n39154;
  assign n39156 = ~n13988 & n38278;
  assign n39157 = pi0771 & n36190;
  assign n39158 = pi0771 & ~n38283;
  assign n39159 = ~n38284 & ~n39158;
  assign n39160 = ~n36190 & ~n39159;
  assign n39161 = ~n39157 & ~n39160;
  assign n39162 = ~n38278 & ~n39161;
  assign po1067 = n39156 | n39162;
  assign n39164 = ~n14816 & n38278;
  assign n39165 = pi0772 & n36190;
  assign n39166 = pi0772 & ~n38282;
  assign n39167 = ~n38640 & ~n39166;
  assign n39168 = ~n36190 & ~n39167;
  assign n39169 = ~n39165 & ~n39168;
  assign n39170 = ~n38278 & ~n39169;
  assign po1068 = n39164 | n39170;
  assign n39172 = ~n13398 & n38962;
  assign n39173 = pi0749 & pi0778;
  assign n39174 = pi0777 & n39173;
  assign n39175 = pi0776 & n39174;
  assign n39176 = pi0775 & n39175;
  assign n39177 = pi0774 & n39176;
  assign n39178 = pi0773 & n39177;
  assign n39179 = ~pi0773 & ~n39177;
  assign n39180 = ~n39178 & ~n39179;
  assign n39181 = ~n36190 & ~n39180;
  assign n39182 = ~pi0773 & n36190;
  assign n39183 = ~n39181 & ~n39182;
  assign n39184 = ~n38962 & n39183;
  assign po1069 = n39172 | n39184;
  assign n39186 = ~n13988 & n38962;
  assign n39187 = ~pi0774 & ~n38993;
  assign n39188 = pi0774 & n38993;
  assign n39189 = ~n39187 & ~n39188;
  assign n39190 = ~n36190 & ~n39189;
  assign n39191 = ~pi0774 & n36190;
  assign n39192 = ~n39190 & ~n39191;
  assign n39193 = ~n38962 & n39192;
  assign po1070 = n39186 | n39193;
  assign n39195 = ~n12415 & n38962;
  assign n39196 = ~pi0775 & ~n39175;
  assign n39197 = ~n39176 & ~n39196;
  assign n39198 = ~n36190 & ~n39197;
  assign n39199 = ~pi0775 & n36190;
  assign n39200 = ~n39198 & ~n39199;
  assign n39201 = ~n38962 & n39200;
  assign po1071 = n39195 | n39201;
  assign n39203 = ~n14816 & n38962;
  assign n39204 = ~pi0776 & ~n39174;
  assign n39205 = ~n39175 & ~n39204;
  assign n39206 = ~n36190 & ~n39205;
  assign n39207 = ~pi0776 & n36190;
  assign n39208 = ~n39206 & ~n39207;
  assign n39209 = ~n38962 & n39208;
  assign po1072 = n39203 | n39209;
  assign n39211 = ~n15115 & n38962;
  assign n39212 = ~pi0777 & ~n39173;
  assign n39213 = ~n39174 & ~n39212;
  assign n39214 = ~n36190 & ~n39213;
  assign n39215 = ~pi0777 & n36190;
  assign n39216 = ~n39214 & ~n39215;
  assign n39217 = ~n38962 & n39216;
  assign po1073 = n39211 | n39217;
  assign n39219 = ~n12061 & n38962;
  assign n39220 = pi0749 & ~pi0778;
  assign n39221 = ~pi0749 & pi0778;
  assign n39222 = ~n39220 & ~n39221;
  assign n39223 = ~n36190 & n39222;
  assign n39224 = ~pi0778 & n36190;
  assign n39225 = ~n39223 & ~n39224;
  assign n39226 = ~n38962 & n39225;
  assign po1074 = n39219 | n39226;
  assign n39228 = pi0779 & n36190;
  assign n39229 = pi0773 & pi0861;
  assign n39230 = n39177 & n39229;
  assign n39231 = pi0845 & pi0862;
  assign n39232 = n39230 & n39231;
  assign n39233 = pi0780 & n39232;
  assign n39234 = pi0781 & n39233;
  assign n39235 = pi0779 & n39234;
  assign n39236 = ~pi0779 & ~n39234;
  assign n39237 = ~n39235 & ~n39236;
  assign n39238 = ~n36190 & n39237;
  assign n39239 = ~n39228 & ~n39238;
  assign n39240 = ~n38962 & ~n39239;
  assign n39241 = ~n10608 & n38962;
  assign po1075 = n39240 | n39241;
  assign n39243 = ~n15426 & n38962;
  assign n39244 = n38995 & n39176;
  assign n39245 = n39231 & n39244;
  assign n39246 = pi0861 & n39245;
  assign n39247 = pi0781 & n39246;
  assign n39248 = pi0780 & n39247;
  assign n39249 = ~pi0780 & ~n39247;
  assign n39250 = ~n39248 & ~n39249;
  assign n39251 = ~n36190 & ~n39250;
  assign n39252 = ~pi0780 & n36190;
  assign n39253 = ~n39251 & ~n39252;
  assign n39254 = ~n38962 & n39253;
  assign po1076 = n39243 | n39254;
  assign n39256 = ~n14403 & n38962;
  assign n39257 = n39229 & n39231;
  assign n39258 = n39177 & n39257;
  assign n39259 = pi0781 & n39258;
  assign n39260 = ~pi0781 & ~n39258;
  assign n39261 = ~n39259 & ~n39260;
  assign n39262 = ~n36190 & ~n39261;
  assign n39263 = ~pi0781 & n36190;
  assign n39264 = ~n39262 & ~n39263;
  assign n39265 = ~n38962 & n39264;
  assign po1077 = n39256 | n39265;
  assign n39267 = ~n12415 & n38278;
  assign n39268 = pi0782 & n36190;
  assign n39269 = pi0782 & ~n38640;
  assign n39270 = ~n38641 & ~n39269;
  assign n39271 = ~n36190 & ~n39270;
  assign n39272 = ~n39268 & ~n39271;
  assign n39273 = ~n38278 & ~n39272;
  assign po1078 = n39267 | n39273;
  assign n39275 = n36194 & n38281;
  assign n39276 = n36173 & n39275;
  assign po1079 = ~n36197 & ~n39276;
  assign po1080 = pi0784 & ~n36197;
  assign n39279 = pi0785 & n38745;
  assign n39280 = ~pi3006 & n38772;
  assign n39281 = ~pi2806 & n38770;
  assign n39282 = ~n39280 & ~n39281;
  assign n39283 = ~pi3057 & n38775;
  assign n39284 = ~n38764 & ~n39283;
  assign n39285 = n39282 & n39284;
  assign n39286 = ~pi1674 & n38781;
  assign n39287 = n39285 & ~n39286;
  assign n39288 = ~pi1086 & n38779;
  assign n39289 = ~pi3014 & n38766;
  assign n39290 = ~n39288 & ~n39289;
  assign n39291 = ~pi2997 & n38757;
  assign n39292 = ~pi2837 & n38760;
  assign n39293 = ~n39291 & ~n39292;
  assign n39294 = pi0816 & n38787;
  assign n39295 = pi0369 & n38792;
  assign n39296 = ~n39294 & ~n39295;
  assign n39297 = ~pi3089 & n38749;
  assign n39298 = ~pi3053 & n38752;
  assign n39299 = ~n39297 & ~n39298;
  assign n39300 = n39296 & n39299;
  assign n39301 = n39293 & n39300;
  assign n39302 = pi0403 & n38789;
  assign n39303 = n38759 & n38778;
  assign n39304 = ~pi3205 & n39303;
  assign n39305 = ~n39302 & ~n39304;
  assign n39306 = n39301 & n39305;
  assign n39307 = n39290 & n39306;
  assign n39308 = n39287 & n39307;
  assign n39309 = n38798 & ~n39308;
  assign n39310 = pi0825 & n38800;
  assign n39311 = pi0854 & ~n38800;
  assign n39312 = ~n39310 & ~n39311;
  assign n39313 = ~n38798 & ~n39312;
  assign n39314 = ~n39309 & ~n39313;
  assign n39315 = ~n38745 & ~n39314;
  assign po1081 = n39279 | n39315;
  assign n39317 = ~n15115 & n38278;
  assign n39318 = pi0786 & n36190;
  assign n39319 = pi0786 & n38281;
  assign n39320 = ~pi0786 & ~n38281;
  assign n39321 = ~n39319 & ~n39320;
  assign n39322 = ~n36190 & n39321;
  assign n39323 = ~n39318 & ~n39322;
  assign n39324 = ~n38278 & ~n39323;
  assign po1082 = n39317 | n39324;
  assign n39326 = ~n11181 & n38278;
  assign n39327 = pi0787 & n36190;
  assign n39328 = ~pi0787 & ~n36190;
  assign n39329 = ~n39327 & ~n39328;
  assign n39330 = ~n38278 & ~n39329;
  assign po1083 = n39326 | n39330;
  assign n39332 = n33317 & n38787;
  assign n39333 = ~po3946 & ~n39332;
  assign n39334 = pi0788 & n39333;
  assign n39335 = pi3420 & po3946;
  assign n39336 = pi0855 & ~po3946;
  assign n39337 = ~n39335 & ~n39336;
  assign n39338 = ~n39333 & ~n39337;
  assign po1084 = n39334 | n39338;
  assign n39340 = ~pi0790 & n38916;
  assign n39341 = n13701 & ~n38916;
  assign n39342 = ~n39340 & ~n39341;
  assign po1086 = n38920 | n39342;
  assign n39344 = ~pi0791 & n38916;
  assign n39345 = n15426 & ~n38916;
  assign n39346 = ~n39344 & ~n39345;
  assign po1087 = n38920 | n39346;
  assign n39348 = ~pi1033 & n9604;
  assign n39349 = pi1039 & n39348;
  assign n39350 = n38898 & n39349;
  assign n39351 = n38902 & n39350;
  assign n39352 = pi0609 & n39351;
  assign n39353 = ~pi1039 & n39348;
  assign n39354 = n38906 & n39353;
  assign n39355 = ~n39352 & ~n39354;
  assign n39356 = pi0792 & n39355;
  assign n39357 = ~n12726 & ~n39355;
  assign n39358 = ~n39356 & ~n39357;
  assign n39359 = n39351 & ~n39355;
  assign po1088 = ~n39358 | n39359;
  assign n39361 = pi0793 & n39355;
  assign n39362 = ~n12061 & ~n39355;
  assign n39363 = ~n39361 & ~n39362;
  assign po1089 = n39359 | ~n39363;
  assign n39365 = pi0794 & n39355;
  assign n39366 = ~n14403 & ~n39355;
  assign n39367 = ~n39365 & ~n39366;
  assign po1090 = n39359 | ~n39367;
  assign n39369 = pi0795 & n39355;
  assign n39370 = ~n11181 & ~n39355;
  assign n39371 = ~n39369 & ~n39370;
  assign po1091 = n39359 | ~n39371;
  assign n39373 = n38905 & n39350;
  assign n39374 = ~n39352 & ~n39373;
  assign n39375 = ~n17199 & ~n39374;
  assign n39376 = pi0796 & n39374;
  assign n39377 = ~n39375 & ~n39376;
  assign n39378 = n39351 & ~n39374;
  assign po1092 = ~n39377 | n39378;
  assign n39380 = ~n14816 & ~n39374;
  assign n39381 = pi0797 & n39374;
  assign n39382 = ~n39380 & ~n39381;
  assign po1093 = n39378 | ~n39382;
  assign n39384 = ~n15115 & ~n39374;
  assign n39385 = pi0798 & n39374;
  assign n39386 = ~n39384 & ~n39385;
  assign po1094 = n39378 | ~n39386;
  assign n39388 = ~n17368 & ~n39374;
  assign n39389 = pi0799 & n39374;
  assign n39390 = ~n39388 & ~n39389;
  assign po1095 = n39378 | ~n39390;
  assign n39392 = n9651 & n38906;
  assign n39393 = ~n39352 & ~n39392;
  assign n39394 = pi0800 & n39393;
  assign n39395 = ~n13121 & ~n39393;
  assign n39396 = ~n39394 & ~n39395;
  assign n39397 = n39351 & ~n39393;
  assign po1096 = ~n39396 | n39397;
  assign n39399 = pi0801 & n39393;
  assign n39400 = ~n13398 & ~n39393;
  assign n39401 = ~n39399 & ~n39400;
  assign po1097 = n39397 | ~n39401;
  assign n39403 = pi0802 & n39393;
  assign n39404 = ~n13988 & ~n39393;
  assign n39405 = ~n39403 & ~n39404;
  assign po1098 = n39397 | ~n39405;
  assign n39407 = pi0803 & n39393;
  assign n39408 = ~n14816 & ~n39393;
  assign n39409 = ~n39407 & ~n39408;
  assign po1099 = n39397 | ~n39409;
  assign n39411 = pi0804 & n39393;
  assign n39412 = ~n12061 & ~n39393;
  assign n39413 = ~n39411 & ~n39412;
  assign po1100 = n39397 | ~n39413;
  assign n39415 = pi0805 & n39393;
  assign n39416 = ~n11181 & ~n39393;
  assign n39417 = ~n39415 & ~n39416;
  assign po1101 = n39397 | ~n39417;
  assign n39419 = pi0806 & n39333;
  assign n39420 = pi3411 & po3946;
  assign n39421 = pi0856 & ~po3946;
  assign n39422 = ~n39420 & ~n39421;
  assign n39423 = ~n39333 & ~n39422;
  assign po1102 = n39419 | n39423;
  assign n39425 = pi0807 & n39333;
  assign n39426 = pi3406 & po3946;
  assign n39427 = pi0857 & ~po3946;
  assign n39428 = ~n39426 & ~n39427;
  assign n39429 = ~n39333 & ~n39428;
  assign po1103 = n39425 | n39429;
  assign n39431 = pi0808 & n39333;
  assign n39432 = pi3413 & po3946;
  assign n39433 = pi0858 & ~po3946;
  assign n39434 = ~n39432 & ~n39433;
  assign n39435 = ~n39333 & ~n39434;
  assign po1104 = n39431 | n39435;
  assign n39437 = pi0809 & n39333;
  assign n39438 = pi3405 & po3946;
  assign n39439 = pi0824 & ~po3946;
  assign n39440 = ~n39438 & ~n39439;
  assign n39441 = ~n39333 & ~n39440;
  assign po1105 = n39437 | n39441;
  assign n39443 = pi0810 & n39333;
  assign n39444 = pi3414 & po3946;
  assign n39445 = pi0823 & ~po3946;
  assign n39446 = ~n39444 & ~n39445;
  assign n39447 = ~n39333 & ~n39446;
  assign po1106 = n39443 | n39447;
  assign n39449 = pi0811 & n39333;
  assign n39450 = pi3404 & po3946;
  assign n39451 = pi0859 & ~po3946;
  assign n39452 = ~n39450 & ~n39451;
  assign n39453 = ~n39333 & ~n39452;
  assign po1107 = n39449 | n39453;
  assign n39455 = pi0812 & n39333;
  assign n39456 = pi3402 & po3946;
  assign n39457 = pi0730 & ~po3946;
  assign n39458 = ~n39456 & ~n39457;
  assign n39459 = ~n39333 & ~n39458;
  assign po1108 = n39455 | n39459;
  assign n39461 = pi0813 & n39333;
  assign n39462 = pi3403 & po3946;
  assign n39463 = pi0731 & ~po3946;
  assign n39464 = ~n39462 & ~n39463;
  assign n39465 = ~n39333 & ~n39464;
  assign po1109 = n39461 | n39465;
  assign n39467 = pi0814 & n39333;
  assign n39468 = pi3430 & po3946;
  assign n39469 = pi0853 & ~po3946;
  assign n39470 = ~n39468 & ~n39469;
  assign n39471 = ~n39333 & ~n39470;
  assign po1110 = n39467 | n39471;
  assign n39473 = pi0815 & n39333;
  assign n39474 = pi3421 & po3946;
  assign n39475 = pi0854 & ~po3946;
  assign n39476 = ~n39474 & ~n39475;
  assign n39477 = ~n39333 & ~n39476;
  assign po1111 = n39473 | n39477;
  assign n39479 = pi0816 & n39333;
  assign n39480 = pi3422 & po3946;
  assign n39481 = pi0785 & ~po3946;
  assign n39482 = ~n39480 & ~n39481;
  assign n39483 = ~n39333 & ~n39482;
  assign po1112 = n39479 | n39483;
  assign n39485 = pi0817 & n39333;
  assign n39486 = pi3401 & po3946;
  assign n39487 = pi0825 & ~po3946;
  assign n39488 = ~n39486 & ~n39487;
  assign n39489 = ~n39333 & ~n39488;
  assign po1113 = n39485 | n39489;
  assign n39491 = pi0818 & n39333;
  assign n39492 = pi3400 & po3946;
  assign n39493 = pi0938 & ~po3946;
  assign n39494 = ~n39492 & ~n39493;
  assign n39495 = ~n39333 & ~n39494;
  assign po1114 = n39491 | n39495;
  assign n39497 = ~pi0609 & ~pi3579;
  assign n39498 = ~pi1771 & n39497;
  assign n39499 = n9641 & n38277;
  assign n39500 = n9636 & n39499;
  assign n39501 = n38907 & n39500;
  assign n39502 = pi3578 & pi3579;
  assign n39503 = pi3467 & n39502;
  assign n39504 = ~n39501 & ~n39503;
  assign n39505 = ~n39498 & ~n39504;
  assign n39506 = ~pi3579 & ~n10608;
  assign n39507 = ~pi3447 & pi3579;
  assign n39508 = ~n39506 & ~n39507;
  assign n39509 = n39505 & ~n39508;
  assign n39510 = pi0873 & pi0908;
  assign n39511 = pi0907 & n39510;
  assign n39512 = pi0874 & n39511;
  assign n39513 = pi0906 & n39512;
  assign n39514 = pi0905 & n39513;
  assign n39515 = pi0876 & pi0904;
  assign n39516 = n39514 & n39515;
  assign n39517 = pi0902 & pi0903;
  assign n39518 = n39516 & n39517;
  assign n39519 = pi0820 & n39518;
  assign n39520 = pi0910 & n39519;
  assign n39521 = pi0819 & n39520;
  assign n39522 = ~pi0819 & ~n39520;
  assign n39523 = ~n39521 & ~n39522;
  assign n39524 = ~pi0975 & ~pi1422;
  assign n39525 = pi1936 & pi2056;
  assign n39526 = pi1935 & n39525;
  assign n39527 = n39524 & n39526;
  assign n39528 = ~pi3428 & ~n39524;
  assign n39529 = ~n39527 & ~n39528;
  assign n39530 = pi2769 & ~n39529;
  assign n39531 = ~n32788 & ~n39530;
  assign n39532 = ~n39524 & ~n39531;
  assign n39533 = ~n39498 & n39532;
  assign n39534 = ~n39523 & n39533;
  assign n39535 = ~pi0819 & ~n39533;
  assign n39536 = ~n39534 & ~n39535;
  assign n39537 = ~n39505 & n39536;
  assign po1116 = n39509 | n39537;
  assign n39539 = ~pi3579 & ~n15426;
  assign n39540 = ~pi3463 & pi3579;
  assign n39541 = ~n39539 & ~n39540;
  assign n39542 = n39505 & ~n39541;
  assign n39543 = pi0904 & pi0905;
  assign n39544 = n39513 & n39543;
  assign n39545 = n39517 & n39544;
  assign n39546 = pi0876 & n39545;
  assign n39547 = pi0910 & n39546;
  assign n39548 = pi0820 & n39547;
  assign n39549 = ~pi0820 & ~n39547;
  assign n39550 = ~n39548 & ~n39549;
  assign n39551 = n39533 & ~n39550;
  assign n39552 = ~pi0820 & ~n39533;
  assign n39553 = ~n39551 & ~n39552;
  assign n39554 = ~n39505 & n39553;
  assign po1117 = n39542 | n39554;
  assign n39556 = pi0821 & n38745;
  assign n39557 = pi0412 & n38789;
  assign n39558 = pi0385 & n38792;
  assign n39559 = ~n39557 & ~n39558;
  assign n39560 = ~pi3025 & n38760;
  assign n39561 = n39559 & ~n39560;
  assign n39562 = ~pi2973 & n38749;
  assign n39563 = ~pi2818 & n38752;
  assign n39564 = ~pi3001 & n38757;
  assign n39565 = ~n39563 & ~n39564;
  assign n39566 = ~pi3042 & n38770;
  assign n39567 = ~pi3008 & n38772;
  assign n39568 = ~n39566 & ~n39567;
  assign n39569 = ~pi3032 & n38775;
  assign n39570 = n39568 & ~n39569;
  assign n39571 = ~pi3016 & n38766;
  assign n39572 = n39570 & ~n39571;
  assign n39573 = n39565 & n39572;
  assign n39574 = ~n39562 & n39573;
  assign n39575 = n39561 & n39574;
  assign n39576 = ~pi1368 & n38779;
  assign n39577 = ~pi1678 & n38781;
  assign n39578 = ~n39576 & ~n39577;
  assign n39579 = n39575 & n39578;
  assign n39580 = n38798 & ~n39579;
  assign n39581 = ~pi0937 & n38800;
  assign n39582 = pi0852 & ~n38800;
  assign n39583 = ~n39581 & ~n39582;
  assign n39584 = ~n38798 & ~n39583;
  assign n39585 = ~n39580 & ~n39584;
  assign n39586 = ~n38745 & ~n39585;
  assign po1118 = n39556 | n39586;
  assign n39588 = pi0822 & ~n31865;
  assign n39589 = pi0822 & ~n38692;
  assign n39590 = ~n31786 & ~n39589;
  assign n39591 = pi3641 & n39590;
  assign n39592 = ~pi0822 & ~pi3641;
  assign n39593 = ~n39591 & ~n39592;
  assign n39594 = n31865 & n39593;
  assign n39595 = ~n39588 & ~n39594;
  assign n39596 = ~n31777 & ~n39595;
  assign n39597 = pi1719 & n31777;
  assign n39598 = ~n39596 & ~n39597;
  assign n39599 = ~n31779 & ~n39598;
  assign n39600 = ~pi2397 & n31779;
  assign po1119 = n39599 | n39600;
  assign n39602 = pi0823 & n38745;
  assign n39603 = ~pi2792 & n38749;
  assign n39604 = ~pi2899 & n38752;
  assign n39605 = ~n39603 & ~n39604;
  assign n39606 = ~pi2994 & n38757;
  assign n39607 = ~pi3017 & n38760;
  assign n39608 = ~n39606 & ~n39607;
  assign n39609 = pi0810 & n38787;
  assign n39610 = pi0423 & n38789;
  assign n39611 = ~n39609 & ~n39610;
  assign n39612 = pi0377 & n38792;
  assign n39613 = n39611 & ~n39612;
  assign n39614 = ~pi3002 & n38772;
  assign n39615 = ~pi3010 & n38766;
  assign n39616 = ~n39614 & ~n39615;
  assign n39617 = ~n38764 & ~n38769;
  assign n39618 = ~pi1364 & n38779;
  assign n39619 = ~pi1700 & n38781;
  assign n39620 = ~n39618 & ~n39619;
  assign n39621 = ~pi3081 & n38775;
  assign n39622 = ~pi3040 & n38770;
  assign n39623 = ~n39621 & ~n39622;
  assign n39624 = n39620 & n39623;
  assign n39625 = n39617 & n39624;
  assign n39626 = n39616 & n39625;
  assign n39627 = n39613 & n39626;
  assign n39628 = n39608 & n39627;
  assign n39629 = n39605 & n39628;
  assign n39630 = n38798 & ~n39629;
  assign n39631 = pi0859 & n38800;
  assign n39632 = pi0824 & ~n38800;
  assign n39633 = ~n39631 & ~n39632;
  assign n39634 = ~n38798 & ~n39633;
  assign n39635 = ~n39630 & ~n39634;
  assign n39636 = ~n38745 & ~n39635;
  assign po1120 = n39602 | n39636;
  assign n39638 = pi0824 & n38745;
  assign n39639 = ~pi3033 & n38749;
  assign n39640 = ~pi2775 & n38752;
  assign n39641 = ~n39639 & ~n39640;
  assign n39642 = ~pi2954 & n38757;
  assign n39643 = ~pi2815 & n38760;
  assign n39644 = ~n39642 & ~n39643;
  assign n39645 = pi0809 & n38787;
  assign n39646 = pi0422 & n38789;
  assign n39647 = ~n39645 & ~n39646;
  assign n39648 = pi0376 & n38792;
  assign n39649 = n39647 & ~n39648;
  assign n39650 = ~pi2880 & n38772;
  assign n39651 = ~pi3009 & n38766;
  assign n39652 = ~n39650 & ~n39651;
  assign n39653 = ~pi1385 & n38779;
  assign n39654 = ~pi1387 & n38781;
  assign n39655 = ~n39653 & ~n39654;
  assign n39656 = ~pi3026 & n38775;
  assign n39657 = ~pi3061 & n38770;
  assign n39658 = ~n39656 & ~n39657;
  assign n39659 = n39655 & n39658;
  assign n39660 = n39617 & n39659;
  assign n39661 = n39652 & n39660;
  assign n39662 = n39649 & n39661;
  assign n39663 = n39644 & n39662;
  assign n39664 = n39641 & n39663;
  assign n39665 = n38798 & ~n39664;
  assign n39666 = pi0823 & n38800;
  assign n39667 = pi0858 & ~n38800;
  assign n39668 = ~n39666 & ~n39667;
  assign n39669 = ~n38798 & ~n39668;
  assign n39670 = ~n39665 & ~n39669;
  assign n39671 = ~n38745 & ~n39670;
  assign po1121 = n39638 | n39671;
  assign n39673 = pi0825 & n38745;
  assign n39674 = ~pi1005 & n38779;
  assign n39675 = ~pi2972 & n38766;
  assign n39676 = ~n39674 & ~n39675;
  assign n39677 = ~pi3039 & n38749;
  assign n39678 = ~pi2930 & n38752;
  assign n39679 = ~n39677 & ~n39678;
  assign n39680 = ~pi2887 & n38757;
  assign n39681 = ~pi2910 & n38760;
  assign n39682 = ~n39680 & ~n39681;
  assign n39683 = pi0418 & n38789;
  assign n39684 = pi3551 & n39303;
  assign n39685 = ~n39683 & ~n39684;
  assign n39686 = pi0817 & n38787;
  assign n39687 = pi0371 & n38792;
  assign n39688 = ~n39686 & ~n39687;
  assign n39689 = n39685 & n39688;
  assign n39690 = n39682 & n39689;
  assign n39691 = n39679 & n39690;
  assign n39692 = ~pi2857 & n38772;
  assign n39693 = ~pi3044 & n38770;
  assign n39694 = ~n39692 & ~n39693;
  assign n39695 = ~pi3058 & n38775;
  assign n39696 = ~n38764 & ~n39695;
  assign n39697 = n39694 & n39696;
  assign n39698 = n39691 & n39697;
  assign n39699 = pi0565 & n38769;
  assign n39700 = ~pi1073 & n38781;
  assign n39701 = ~n39699 & ~n39700;
  assign n39702 = n39698 & n39701;
  assign n39703 = n39676 & n39702;
  assign n39704 = n38798 & ~n39703;
  assign n39705 = pi0855 & n38800;
  assign n39706 = pi0785 & ~n38800;
  assign n39707 = ~n39705 & ~n39706;
  assign n39708 = ~n38798 & ~n39707;
  assign n39709 = ~n39704 & ~n39708;
  assign n39710 = ~n38745 & ~n39709;
  assign po1122 = n39673 | n39710;
  assign n39712 = ~pi0866 & ~pi3120;
  assign n39713 = ~n9352 & ~n39712;
  assign n39714 = ~n19551 & ~n39713;
  assign n39715 = ~pi3210 & ~n19545;
  assign n39716 = n39712 & n39715;
  assign po1281 = ~n39714 & ~n39716;
  assign n39718 = ~pi1526 & n20345;
  assign n39719 = ~pi1411 & n20347;
  assign n39720 = ~n39718 & ~n39719;
  assign n39721 = ~pi1593 & n20350;
  assign n39722 = ~pi1621 & n20353;
  assign n39723 = ~pi1561 & n20356;
  assign n39724 = ~n39722 & ~n39723;
  assign n39725 = ~pi1507 & n20360;
  assign n39726 = ~pi1489 & n20363;
  assign n39727 = ~n39725 & ~n39726;
  assign n39728 = n39724 & n39727;
  assign n39729 = ~n39721 & n39728;
  assign n39730 = n39720 & n39729;
  assign n39731 = ~pi3120 & ~n39730;
  assign n39732 = pi0826 & ~pi3398;
  assign n39733 = pi3392 & pi3398;
  assign n39734 = ~n39732 & ~n39733;
  assign n39735 = pi3120 & ~n39734;
  assign n39736 = ~n39731 & ~n39735;
  assign n39737 = ~pi0866 & ~n39736;
  assign n39738 = pi0866 & ~n13398;
  assign n39739 = ~n39737 & ~n39738;
  assign n39740 = po1281 & ~n39739;
  assign n39741 = pi0826 & ~po1281;
  assign po1124 = n39740 | n39741;
  assign n39743 = ~pi1421 & n20345;
  assign n39744 = ~pi1545 & n20347;
  assign n39745 = ~n39743 & ~n39744;
  assign n39746 = ~pi1423 & n20350;
  assign n39747 = ~pi1577 & n20353;
  assign n39748 = ~pi1391 & n20356;
  assign n39749 = ~n39747 & ~n39748;
  assign n39750 = ~pi1508 & n20360;
  assign n39751 = ~pi1490 & n20363;
  assign n39752 = ~n39750 & ~n39751;
  assign n39753 = n39749 & n39752;
  assign n39754 = ~n39746 & n39753;
  assign n39755 = n39745 & n39754;
  assign n39756 = ~pi3120 & ~n39755;
  assign n39757 = pi3504 & pi3513;
  assign n39758 = pi0827 & ~pi3513;
  assign n39759 = ~n39757 & ~n39758;
  assign n39760 = pi3120 & ~n39759;
  assign n39761 = ~n39756 & ~n39760;
  assign n39762 = ~pi0866 & ~n39761;
  assign n39763 = pi0866 & ~n13988;
  assign n39764 = ~n39762 & ~n39763;
  assign n39765 = po1281 & ~n39764;
  assign n39766 = pi0827 & ~po1281;
  assign po1125 = n39765 | n39766;
  assign n39768 = ~pi1528 & n20345;
  assign n39769 = ~pi1546 & n20347;
  assign n39770 = ~n39768 & ~n39769;
  assign n39771 = ~pi1401 & n20350;
  assign n39772 = ~pi1509 & n20360;
  assign n39773 = ~pi1390 & n20363;
  assign n39774 = ~n39772 & ~n39773;
  assign n39775 = ~pi1578 & n20353;
  assign n39776 = ~pi1399 & n20356;
  assign n39777 = ~n39775 & ~n39776;
  assign n39778 = n39774 & n39777;
  assign n39779 = ~n39771 & n39778;
  assign n39780 = n39770 & n39779;
  assign n39781 = ~pi3120 & ~n39780;
  assign n39782 = pi3514 & pi3517;
  assign n39783 = pi0828 & ~pi3514;
  assign n39784 = ~n39782 & ~n39783;
  assign n39785 = pi3120 & ~n39784;
  assign n39786 = ~n39781 & ~n39785;
  assign n39787 = ~pi0866 & ~n39786;
  assign n39788 = pi0866 & ~n14816;
  assign n39789 = ~n39787 & ~n39788;
  assign n39790 = po1281 & ~n39789;
  assign n39791 = pi0828 & ~po1281;
  assign po1126 = n39790 | n39791;
  assign n39793 = ~pi1529 & n20345;
  assign n39794 = ~pi1412 & n20347;
  assign n39795 = ~n39793 & ~n39794;
  assign n39796 = ~pi1595 & n20350;
  assign n39797 = ~pi1579 & n20353;
  assign n39798 = ~pi1563 & n20356;
  assign n39799 = ~n39797 & ~n39798;
  assign n39800 = ~pi1510 & n20360;
  assign n39801 = ~pi1492 & n20363;
  assign n39802 = ~n39800 & ~n39801;
  assign n39803 = n39799 & n39802;
  assign n39804 = ~n39796 & n39803;
  assign n39805 = n39795 & n39804;
  assign n39806 = ~pi3120 & ~n39805;
  assign n39807 = pi0829 & ~pi3508;
  assign n39808 = ~n19614 & ~n39807;
  assign n39809 = pi3120 & ~n39808;
  assign n39810 = ~n39806 & ~n39809;
  assign n39811 = ~pi0866 & ~n39810;
  assign n39812 = pi0866 & ~n15115;
  assign n39813 = ~n39811 & ~n39812;
  assign n39814 = po1281 & ~n39813;
  assign n39815 = pi0829 & ~po1281;
  assign po1127 = n39814 | n39815;
  assign n39817 = ~pi1615 & n20345;
  assign n39818 = ~pi1530 & n20347;
  assign n39819 = ~n39817 & ~n39818;
  assign n39820 = ~pi1611 & n20350;
  assign n39821 = ~pi1565 & n20353;
  assign n39822 = ~pi1548 & n20356;
  assign n39823 = ~n39821 & ~n39822;
  assign n39824 = ~pi1494 & n20360;
  assign n39825 = ~pi1476 & n20363;
  assign n39826 = ~n39824 & ~n39825;
  assign n39827 = n39823 & n39826;
  assign n39828 = ~n39820 & n39827;
  assign n39829 = n39819 & n39828;
  assign n39830 = ~pi3120 & ~n39829;
  assign n39831 = pi0830 & ~pi3511;
  assign n39832 = pi3510 & pi3511;
  assign n39833 = ~n39831 & ~n39832;
  assign n39834 = pi3120 & ~n39833;
  assign n39835 = ~n39830 & ~n39834;
  assign n39836 = ~pi0866 & ~n39835;
  assign n39837 = pi0866 & ~n12061;
  assign n39838 = ~n39836 & ~n39837;
  assign n39839 = po1281 & ~n39838;
  assign n39840 = pi0830 & ~po1281;
  assign po1128 = n39839 | n39840;
  assign n39842 = ~n8561 & n36095;
  assign n39843 = n36094 & n39842;
  assign n39844 = ~n36083 & n36096;
  assign n39845 = n39843 & n39844;
  assign n39846 = ~pi0831 & n8561;
  assign n39847 = ~n39845 & ~n39846;
  assign po1129 = po3627 & ~n39847;
  assign n39849 = n36063 & n36069;
  assign n39850 = n9345 & n39849;
  assign n39851 = ~n36083 & n39850;
  assign n39852 = n38864 & n39851;
  assign n39853 = ~pi0832 & n8561;
  assign n39854 = ~n39852 & ~n39853;
  assign po1130 = po3627 & ~n39854;
  assign n39856 = n36096 & n39842;
  assign n39857 = n39851 & n39856;
  assign n39858 = ~pi0833 & n8561;
  assign n39859 = ~n39857 & ~n39858;
  assign po1131 = po3627 & ~n39859;
  assign n39861 = n36083 & n39850;
  assign n39862 = n39856 & n39861;
  assign n39863 = ~pi0834 & n8561;
  assign n39864 = ~n39862 & ~n39863;
  assign po1132 = po3627 & ~n39864;
  assign n39866 = ~n8561 & ~n36099;
  assign n39867 = pi0835 & n8561;
  assign n39868 = ~n39866 & ~n39867;
  assign po1133 = po3627 & n39868;
  assign n39870 = ~n8561 & n36548;
  assign n39871 = pi0836 & n8561;
  assign po1134 = n39870 | n39871;
  assign n39873 = ~n8561 & n36546;
  assign n39874 = pi0837 & n8561;
  assign po1135 = n39873 | n39874;
  assign n39876 = ~n8561 & n36541;
  assign n39877 = pi0838 & n8561;
  assign po1136 = n39876 | n39877;
  assign n39879 = ~n8338 & ~n8354;
  assign n39880 = n8347 & n39879;
  assign n39881 = ~n8332 & n39880;
  assign n39882 = ~pi3099 & n39881;
  assign n39883 = ~n8342 & n39882;
  assign n39884 = pi2986 & ~pi2990;
  assign n39885 = pi2990 & n10778;
  assign n39886 = ~n8585 & ~n16211;
  assign n39887 = ~pi1840 & ~n39886;
  assign n39888 = pi1861 & n39887;
  assign n39889 = ~n39885 & ~n39888;
  assign n39890 = ~n39884 & n39889;
  assign n39891 = n39883 & ~n39890;
  assign n39892 = n8578 & ~n39886;
  assign n39893 = n39883 & n39892;
  assign n39894 = ~n39891 & ~n39893;
  assign n39895 = pi0839 & ~n39894;
  assign n39896 = pi2986 & pi2990;
  assign n39897 = pi2990 & n10771;
  assign n39898 = ~n16213 & ~n39897;
  assign n39899 = ~n39896 & n39898;
  assign n39900 = n39883 & ~n39899;
  assign n39901 = ~n39884 & ~n39900;
  assign n39902 = ~n39896 & n39901;
  assign n39903 = n39896 & ~n39900;
  assign n39904 = ~n39902 & ~n39903;
  assign n39905 = ~n39891 & ~n39904;
  assign n39906 = pi0839 & n39905;
  assign n39907 = ~n39891 & n39900;
  assign n39908 = pi3690 & n39907;
  assign n39909 = ~n39906 & ~n39908;
  assign n39910 = ~n39893 & ~n39909;
  assign po1137 = n39895 | n39910;
  assign n39912 = pi0840 & ~n39894;
  assign n39913 = pi0840 & n39905;
  assign n39914 = pi3689 & n39907;
  assign n39915 = ~n39913 & ~n39914;
  assign n39916 = ~n39893 & ~n39915;
  assign po1138 = n39912 | n39916;
  assign n39918 = pi0841 & ~n39894;
  assign n39919 = pi0841 & n39905;
  assign n39920 = pi3687 & n39907;
  assign n39921 = ~n39919 & ~n39920;
  assign n39922 = ~n39893 & ~n39921;
  assign po1139 = n39918 | n39922;
  assign n39924 = pi0842 & ~n39894;
  assign n39925 = pi0842 & n39905;
  assign n39926 = pi3685 & n39907;
  assign n39927 = ~n39925 & ~n39926;
  assign n39928 = ~n39893 & ~n39927;
  assign po1140 = n39924 | n39928;
  assign n39930 = pi0843 & ~n39894;
  assign n39931 = pi0843 & n39905;
  assign n39932 = pi3684 & n39907;
  assign n39933 = ~n39931 & ~n39932;
  assign n39934 = ~n39893 & ~n39933;
  assign po1141 = n39930 | n39934;
  assign n39936 = pi0844 & ~n39894;
  assign n39937 = pi0844 & n39905;
  assign n39938 = pi3683 & ~n39891;
  assign n39939 = n39900 & n39938;
  assign n39940 = ~n39937 & ~n39939;
  assign n39941 = ~n39893 & ~n39940;
  assign po1142 = n39936 | n39941;
  assign n39943 = ~n12726 & n38962;
  assign n39944 = n38992 & n38997;
  assign n39945 = pi0749 & n39944;
  assign n39946 = pi0845 & n39945;
  assign n39947 = ~pi0845 & ~n39945;
  assign n39948 = ~n39946 & ~n39947;
  assign n39949 = ~n36190 & ~n39948;
  assign n39950 = ~pi0845 & n36190;
  assign n39951 = ~n39949 & ~n39950;
  assign n39952 = ~n38962 & n39951;
  assign po1143 = n39943 | n39952;
  assign n39954 = pi0846 & n39393;
  assign n39955 = ~n15115 & ~n39393;
  assign n39956 = ~n39954 & ~n39955;
  assign po1144 = n39397 | ~n39956;
  assign n39958 = ~pi0847 & ~n38681;
  assign n39959 = pi0847 & n38681;
  assign n39960 = ~n39958 & ~n39959;
  assign n39961 = pi3647 & ~n39960;
  assign n39962 = ~pi0847 & ~pi3647;
  assign n39963 = ~n39961 & ~n39962;
  assign n39964 = n36877 & ~n39963;
  assign n39965 = pi0894 & n36876;
  assign po1145 = n39964 | n39965;
  assign n39967 = ~pi0848 & ~n38380;
  assign n39968 = pi0848 & n38380;
  assign n39969 = ~n39967 & ~n39968;
  assign n39970 = pi3635 & ~n39969;
  assign n39971 = ~pi0848 & ~pi3635;
  assign n39972 = ~n39970 & ~n39971;
  assign n39973 = n36969 & ~n39972;
  assign n39974 = pi0968 & n36968;
  assign po1146 = n39973 | n39974;
  assign n39976 = pi0849 & ~n31865;
  assign n39977 = pi0849 & pi3641;
  assign n39978 = ~pi0849 & ~pi3641;
  assign n39979 = ~n39977 & ~n39978;
  assign n39980 = n31865 & n39979;
  assign n39981 = ~n39976 & ~n39980;
  assign n39982 = ~n31777 & ~n39981;
  assign n39983 = pi1726 & n31777;
  assign n39984 = ~n39982 & ~n39983;
  assign n39985 = ~n31779 & ~n39984;
  assign n39986 = ~pi2098 & n31779;
  assign po1147 = n39985 | n39986;
  assign n39988 = pi0850 & n39393;
  assign n39989 = ~n12415 & ~n39393;
  assign n39990 = ~n39988 & ~n39989;
  assign po1148 = n39397 | ~n39990;
  assign n39992 = pi0851 & n38745;
  assign n39993 = pi0409 & n38789;
  assign n39994 = pi0382 & n38792;
  assign n39995 = ~n39993 & ~n39994;
  assign n39996 = ~pi2790 & n38760;
  assign n39997 = n39995 & ~n39996;
  assign n39998 = ~pi2970 & n38770;
  assign n39999 = ~pi2822 & n38772;
  assign n40000 = ~n39998 & ~n39999;
  assign n40001 = ~pi2971 & n38752;
  assign n40002 = ~pi3067 & n38757;
  assign n40003 = ~n40001 & ~n40002;
  assign n40004 = ~pi3060 & n38775;
  assign n40005 = n40003 & ~n40004;
  assign n40006 = n40000 & n40005;
  assign n40007 = ~pi3036 & n38749;
  assign n40008 = n40006 & ~n40007;
  assign n40009 = ~pi2991 & n38766;
  assign n40010 = n40008 & ~n40009;
  assign n40011 = n39997 & n40010;
  assign n40012 = ~pi1381 & n38779;
  assign n40013 = ~pi1698 & n38781;
  assign n40014 = ~n40012 & ~n40013;
  assign n40015 = n40011 & n40014;
  assign n40016 = n38798 & ~n40015;
  assign n40017 = pi0860 & n38800;
  assign n40018 = pi0938 & ~n38800;
  assign n40019 = ~n40017 & ~n40018;
  assign n40020 = ~n38798 & ~n40019;
  assign n40021 = ~n40016 & ~n40020;
  assign n40022 = ~n38745 & ~n40021;
  assign po1149 = n39992 | n40022;
  assign n40024 = ~pi0860 & ~n38800;
  assign n40025 = ~pi0821 & n38800;
  assign n40026 = ~n40024 & ~n40025;
  assign n40027 = ~n38798 & ~n40026;
  assign n40028 = ~n38745 & ~n40027;
  assign n40029 = ~pi1105 & n38779;
  assign n40030 = ~pi1679 & n38781;
  assign n40031 = ~n40029 & ~n40030;
  assign n40032 = ~pi2977 & n38766;
  assign n40033 = n40031 & ~n40032;
  assign n40034 = ~pi2838 & n38772;
  assign n40035 = n40033 & ~n40034;
  assign n40036 = pi0411 & n38789;
  assign n40037 = pi0384 & n38792;
  assign n40038 = ~n40036 & ~n40037;
  assign n40039 = ~pi3021 & n38760;
  assign n40040 = n40038 & ~n40039;
  assign n40041 = ~pi2907 & n38757;
  assign n40042 = n40040 & ~n40041;
  assign n40043 = ~pi3037 & n38749;
  assign n40044 = ~pi2958 & n38752;
  assign n40045 = ~n40043 & ~n40044;
  assign n40046 = n38798 & n40045;
  assign n40047 = ~pi3028 & n38775;
  assign n40048 = ~pi2811 & n38770;
  assign n40049 = ~n40047 & ~n40048;
  assign n40050 = n40046 & n40049;
  assign n40051 = n40042 & n40050;
  assign n40052 = n40035 & n40051;
  assign n40053 = n40028 & ~n40052;
  assign n40054 = pi0852 & n38745;
  assign po1150 = n40053 | n40054;
  assign n40056 = pi0853 & n38745;
  assign n40057 = pi2813 & n38769;
  assign n40058 = ~pi1074 & n38781;
  assign n40059 = ~n40057 & ~n40058;
  assign n40060 = ~pi3082 & n38749;
  assign n40061 = ~pi3051 & n38752;
  assign n40062 = ~n40060 & ~n40061;
  assign n40063 = ~pi2996 & n38757;
  assign n40064 = ~pi3022 & n38760;
  assign n40065 = ~n40063 & ~n40064;
  assign n40066 = pi0416 & n38789;
  assign n40067 = pi3055 & n39303;
  assign n40068 = ~n40066 & ~n40067;
  assign n40069 = pi0814 & n38787;
  assign n40070 = pi0379 & n38792;
  assign n40071 = ~n40069 & ~n40070;
  assign n40072 = n40068 & n40071;
  assign n40073 = n40065 & n40072;
  assign n40074 = n40062 & n40073;
  assign n40075 = ~pi3005 & n38772;
  assign n40076 = ~pi2902 & n38770;
  assign n40077 = ~n40075 & ~n40076;
  assign n40078 = ~pi3083 & n38775;
  assign n40079 = ~n38764 & ~n40078;
  assign n40080 = n40077 & n40079;
  assign n40081 = n40074 & n40080;
  assign n40082 = ~pi1084 & n38779;
  assign n40083 = ~pi3013 & n38766;
  assign n40084 = ~n40082 & ~n40083;
  assign n40085 = n40081 & n40084;
  assign n40086 = n40059 & n40085;
  assign n40087 = n38798 & ~n40086;
  assign n40088 = pi0854 & n38800;
  assign n40089 = pi3678 & ~n38800;
  assign n40090 = ~n40088 & ~n40089;
  assign n40091 = ~n38798 & ~n40090;
  assign n40092 = ~n40087 & ~n40091;
  assign n40093 = ~n38745 & ~n40092;
  assign po1151 = n40056 | n40093;
  assign n40095 = pi0854 & n38745;
  assign n40096 = ~pi1078 & n38779;
  assign n40097 = ~pi2984 & n38766;
  assign n40098 = ~n40096 & ~n40097;
  assign n40099 = ~pi3038 & n38749;
  assign n40100 = ~pi3052 & n38752;
  assign n40101 = ~n40099 & ~n40100;
  assign n40102 = ~pi2908 & n38757;
  assign n40103 = ~pi2909 & n38760;
  assign n40104 = ~n40102 & ~n40103;
  assign n40105 = pi0417 & n38789;
  assign n40106 = ~pi3188 & n39303;
  assign n40107 = ~n40105 & ~n40106;
  assign n40108 = pi0815 & n38787;
  assign n40109 = pi0380 & n38792;
  assign n40110 = ~n40108 & ~n40109;
  assign n40111 = n40107 & n40110;
  assign n40112 = n40104 & n40111;
  assign n40113 = n40101 & n40112;
  assign n40114 = ~pi2858 & n38772;
  assign n40115 = ~pi3043 & n38770;
  assign n40116 = ~n40114 & ~n40115;
  assign n40117 = ~pi3029 & n38775;
  assign n40118 = ~n38764 & ~n40117;
  assign n40119 = n40116 & n40118;
  assign n40120 = n40113 & n40119;
  assign n40121 = ~pi1610 & n38781;
  assign n40122 = ~pi3145 & n38769;
  assign n40123 = ~n40121 & ~n40122;
  assign n40124 = n40120 & n40123;
  assign n40125 = n40098 & n40124;
  assign n40126 = n38798 & ~n40125;
  assign n40127 = pi0785 & n38800;
  assign n40128 = pi0853 & ~n38800;
  assign n40129 = ~n40127 & ~n40128;
  assign n40130 = ~n38798 & ~n40129;
  assign n40131 = ~n40126 & ~n40130;
  assign n40132 = ~n38745 & ~n40131;
  assign po1152 = n40095 | n40132;
  assign n40134 = pi0855 & n38745;
  assign n40135 = ~pi1077 & n38779;
  assign n40136 = ~pi3015 & n38766;
  assign n40137 = ~n40135 & ~n40136;
  assign n40138 = ~pi3064 & n38749;
  assign n40139 = ~pi3054 & n38752;
  assign n40140 = ~n40138 & ~n40139;
  assign n40141 = ~pi2998 & n38757;
  assign n40142 = ~pi2906 & n38760;
  assign n40143 = ~n40141 & ~n40142;
  assign po3745 = ~pi2860 | pi3573;
  assign n40145 = n39303 & po3745;
  assign n40146 = pi0419 & n38789;
  assign n40147 = ~n40145 & ~n40146;
  assign n40148 = pi0788 & n38787;
  assign n40149 = pi0372 & n38792;
  assign n40150 = ~n40148 & ~n40149;
  assign n40151 = n40147 & n40150;
  assign n40152 = n40143 & n40151;
  assign n40153 = n40140 & n40152;
  assign n40154 = ~pi3007 & n38772;
  assign n40155 = ~pi2904 & n38770;
  assign n40156 = ~n40154 & ~n40155;
  assign n40157 = ~pi3070 & n38775;
  assign n40158 = ~n38764 & ~n40157;
  assign n40159 = n40156 & n40158;
  assign n40160 = n40153 & n40159;
  assign n40161 = pi3452 & n38769;
  assign n40162 = ~pi1604 & n38781;
  assign n40163 = ~n40161 & ~n40162;
  assign n40164 = n40160 & n40163;
  assign n40165 = n40137 & n40164;
  assign n40166 = n38798 & ~n40165;
  assign n40167 = pi0856 & n38800;
  assign n40168 = pi0825 & ~n38800;
  assign n40169 = ~n40167 & ~n40168;
  assign n40170 = ~n38798 & ~n40169;
  assign n40171 = ~n40166 & ~n40170;
  assign n40172 = ~n38745 & ~n40171;
  assign po1153 = n40134 | n40172;
  assign n40174 = pi0856 & n38745;
  assign n40175 = ~pi1076 & n38779;
  assign n40176 = ~pi2886 & n38766;
  assign n40177 = ~n40175 & ~n40176;
  assign n40178 = ~pi3071 & n38749;
  assign n40179 = ~pi3080 & n38752;
  assign n40180 = ~n40178 & ~n40179;
  assign n40181 = ~pi2901 & n38757;
  assign n40182 = ~pi2885 & n38760;
  assign n40183 = ~n40181 & ~n40182;
  assign n40184 = pi0420 & n38789;
  assign n40185 = ~pi3200 & n39303;
  assign n40186 = ~n40184 & ~n40185;
  assign n40187 = pi0806 & n38787;
  assign n40188 = pi0373 & n38792;
  assign n40189 = ~n40187 & ~n40188;
  assign n40190 = n40186 & n40189;
  assign n40191 = n40183 & n40190;
  assign n40192 = n40180 & n40191;
  assign n40193 = ~pi3094 & n38772;
  assign n40194 = ~pi3045 & n38770;
  assign n40195 = ~n40193 & ~n40194;
  assign n40196 = ~pi3030 & n38775;
  assign n40197 = ~n38764 & ~n40196;
  assign n40198 = n40195 & n40197;
  assign n40199 = n40192 & n40198;
  assign n40200 = ~pi1672 & n38781;
  assign n40201 = ~pi3641 & n38769;
  assign n40202 = ~n40200 & ~n40201;
  assign n40203 = n40199 & n40202;
  assign n40204 = n40177 & n40203;
  assign n40205 = n38798 & ~n40204;
  assign n40206 = pi0857 & n38800;
  assign n40207 = pi0855 & ~n38800;
  assign n40208 = ~n40206 & ~n40207;
  assign n40209 = ~n38798 & ~n40208;
  assign n40210 = ~n40205 & ~n40209;
  assign n40211 = ~n38745 & ~n40210;
  assign po1154 = n40174 | n40211;
  assign n40213 = pi0857 & n38745;
  assign n40214 = ~pi2823 & n38749;
  assign n40215 = ~pi2915 & n38752;
  assign n40216 = ~n40214 & ~n40215;
  assign n40217 = ~pi2999 & n38757;
  assign n40218 = ~pi3023 & n38760;
  assign n40219 = ~n40217 & ~n40218;
  assign n40220 = pi0807 & n38787;
  assign n40221 = pi0421 & n38789;
  assign n40222 = ~n40220 & ~n40221;
  assign n40223 = pi0374 & n38792;
  assign n40224 = n40222 & ~n40223;
  assign n40225 = ~pi3077 & n38772;
  assign n40226 = ~pi2959 & n38766;
  assign n40227 = ~n40225 & ~n40226;
  assign n40228 = ~pi1366 & n38779;
  assign n40229 = ~pi1673 & n38781;
  assign n40230 = ~n40228 & ~n40229;
  assign n40231 = ~pi3078 & n38775;
  assign n40232 = ~pi3088 & n38770;
  assign n40233 = ~n40231 & ~n40232;
  assign n40234 = n40230 & n40233;
  assign n40235 = n39617 & n40234;
  assign n40236 = n40227 & n40235;
  assign n40237 = n40224 & n40236;
  assign n40238 = n40219 & n40237;
  assign n40239 = n40216 & n40238;
  assign n40240 = n38798 & ~n40239;
  assign n40241 = pi0858 & n38800;
  assign n40242 = pi0856 & ~n38800;
  assign n40243 = ~n40241 & ~n40242;
  assign n40244 = ~n38798 & ~n40243;
  assign n40245 = ~n40240 & ~n40244;
  assign n40246 = ~n38745 & ~n40245;
  assign po1155 = n40213 | n40246;
  assign n40248 = pi0858 & n38745;
  assign n40249 = ~pi2883 & n38749;
  assign n40250 = ~pi3069 & n38752;
  assign n40251 = ~n40249 & ~n40250;
  assign n40252 = ~pi3000 & n38757;
  assign n40253 = ~pi3024 & n38760;
  assign n40254 = ~n40252 & ~n40253;
  assign n40255 = pi0808 & n38787;
  assign n40256 = pi0405 & n38789;
  assign n40257 = ~n40255 & ~n40256;
  assign n40258 = pi0375 & n38792;
  assign n40259 = n40257 & ~n40258;
  assign n40260 = ~pi3085 & n38772;
  assign n40261 = ~pi2786 & n38766;
  assign n40262 = ~n40260 & ~n40261;
  assign n40263 = ~pi1004 & n38779;
  assign n40264 = ~pi1003 & n38781;
  assign n40265 = ~n40263 & ~n40264;
  assign n40266 = ~pi3031 & n38775;
  assign n40267 = ~pi3046 & n38770;
  assign n40268 = ~n40266 & ~n40267;
  assign n40269 = n40265 & n40268;
  assign n40270 = n39617 & n40269;
  assign n40271 = n40262 & n40270;
  assign n40272 = n40259 & n40271;
  assign n40273 = n40254 & n40272;
  assign n40274 = n40251 & n40273;
  assign n40275 = n38798 & ~n40274;
  assign n40276 = pi0824 & n38800;
  assign n40277 = pi0857 & ~n38800;
  assign n40278 = ~n40276 & ~n40277;
  assign n40279 = ~n38798 & ~n40278;
  assign n40280 = ~n40275 & ~n40279;
  assign n40281 = ~n38745 & ~n40280;
  assign po1156 = n40248 | n40281;
  assign n40283 = pi0859 & n38745;
  assign n40284 = ~pi3034 & n38749;
  assign n40285 = ~pi3048 & n38752;
  assign n40286 = ~n40284 & ~n40285;
  assign n40287 = ~pi2955 & n38757;
  assign n40288 = ~pi3066 & n38760;
  assign n40289 = ~n40287 & ~n40288;
  assign n40290 = pi0811 & n38787;
  assign n40291 = pi0424 & n38789;
  assign n40292 = ~n40290 & ~n40291;
  assign n40293 = pi0378 & n38792;
  assign n40294 = n40292 & ~n40293;
  assign n40295 = ~pi3003 & n38772;
  assign n40296 = ~pi3095 & n38766;
  assign n40297 = ~n40295 & ~n40296;
  assign n40298 = ~pi1365 & n38779;
  assign n40299 = ~pi1671 & n38781;
  assign n40300 = ~n40298 & ~n40299;
  assign n40301 = ~pi3087 & n38775;
  assign n40302 = ~pi3103 & n38770;
  assign n40303 = ~n40301 & ~n40302;
  assign n40304 = n40300 & n40303;
  assign n40305 = n39617 & n40304;
  assign n40306 = n40297 & n40305;
  assign n40307 = n40294 & n40306;
  assign n40308 = n40289 & n40307;
  assign n40309 = n40286 & n40308;
  assign n40310 = n38798 & ~n40309;
  assign n40311 = pi0730 & n38800;
  assign n40312 = pi0823 & ~n38800;
  assign n40313 = ~n40311 & ~n40312;
  assign n40314 = ~n38798 & ~n40313;
  assign n40315 = ~n40310 & ~n40314;
  assign n40316 = ~n38745 & ~n40315;
  assign po1157 = n40283 | n40316;
  assign n40318 = ~pi0852 & n38800;
  assign n40319 = ~pi0851 & ~n38800;
  assign n40320 = ~n40318 & ~n40319;
  assign n40321 = ~n38798 & ~n40320;
  assign n40322 = ~n38745 & ~n40321;
  assign n40323 = ~pi1369 & n38779;
  assign n40324 = ~pi1680 & n38781;
  assign n40325 = ~n40323 & ~n40324;
  assign n40326 = ~pi3012 & n38766;
  assign n40327 = n40325 & ~n40326;
  assign n40328 = ~pi2839 & n38772;
  assign n40329 = n40327 & ~n40328;
  assign n40330 = pi0410 & n38789;
  assign n40331 = pi0383 & n38792;
  assign n40332 = ~n40330 & ~n40331;
  assign n40333 = ~pi3020 & n38760;
  assign n40334 = n40332 & ~n40333;
  assign n40335 = ~pi3073 & n38757;
  assign n40336 = n40334 & ~n40335;
  assign n40337 = ~pi2905 & n38749;
  assign n40338 = ~pi2957 & n38752;
  assign n40339 = ~n40337 & ~n40338;
  assign n40340 = n38798 & n40339;
  assign n40341 = ~pi2859 & n38775;
  assign n40342 = ~pi3041 & n38770;
  assign n40343 = ~n40341 & ~n40342;
  assign n40344 = n40340 & n40343;
  assign n40345 = n40336 & n40344;
  assign n40346 = n40329 & n40345;
  assign n40347 = n40322 & ~n40346;
  assign n40348 = pi0860 & n38745;
  assign po1158 = n40347 | n40348;
  assign n40350 = ~n13121 & n38962;
  assign n40351 = ~pi0861 & ~n39244;
  assign n40352 = pi0861 & n39244;
  assign n40353 = ~n40351 & ~n40352;
  assign n40354 = ~n36190 & ~n40353;
  assign n40355 = ~pi0861 & n36190;
  assign n40356 = ~n40354 & ~n40355;
  assign n40357 = ~n38962 & n40356;
  assign po1159 = n40350 | n40357;
  assign n40359 = ~n13701 & n38962;
  assign n40360 = ~pi0862 & ~n39230;
  assign n40361 = pi0862 & n39230;
  assign n40362 = ~n40360 & ~n40361;
  assign n40363 = ~n36190 & ~n40362;
  assign n40364 = ~pi0862 & n36190;
  assign n40365 = ~n40363 & ~n40364;
  assign n40366 = ~n38962 & n40365;
  assign po1160 = n40359 | n40366;
  assign n40368 = pi3641 & ~n31801;
  assign n40369 = pi0863 & ~pi3641;
  assign n40370 = ~n40368 & ~n40369;
  assign n40371 = n31865 & ~n40370;
  assign n40372 = pi0863 & ~n31865;
  assign n40373 = ~n40371 & ~n40372;
  assign n40374 = ~n31777 & ~n40373;
  assign n40375 = pi1718 & n31777;
  assign n40376 = ~n40374 & ~n40375;
  assign n40377 = ~n31779 & ~n40376;
  assign n40378 = ~pi2093 & n31779;
  assign po1161 = n40377 | n40378;
  assign n40380 = pi0864 & ~n39894;
  assign n40381 = pi0864 & n39905;
  assign n40382 = pi3686 & n39907;
  assign n40383 = ~n40381 & ~n40382;
  assign n40384 = ~n39893 & ~n40383;
  assign po1162 = n40380 | n40384;
  assign n40386 = pi0865 & ~n39894;
  assign n40387 = pi0865 & n39905;
  assign n40388 = pi3688 & n39907;
  assign n40389 = ~n40387 & ~n40388;
  assign n40390 = ~n39893 & ~n40389;
  assign po1163 = n40386 | n40390;
  assign n40392 = pi0866 & n36128;
  assign n40393 = n36060 & n36108;
  assign po1164 = n40392 | n40393;
  assign n40395 = pi0867 & n8561;
  assign n40396 = n36102 & n39842;
  assign n40397 = n36097 & n40396;
  assign n40398 = ~n40395 & ~n40397;
  assign po1165 = po3627 & ~n40398;
  assign n40400 = pi0868 & ~po1281;
  assign n40401 = ~pi1527 & n20345;
  assign n40402 = ~pi1413 & n20347;
  assign n40403 = ~n40401 & ~n40402;
  assign n40404 = ~pi1594 & n20350;
  assign n40405 = ~pi1616 & n20353;
  assign n40406 = ~pi1562 & n20356;
  assign n40407 = ~n40405 & ~n40406;
  assign n40408 = ~pi1617 & n20360;
  assign n40409 = ~pi1491 & n20363;
  assign n40410 = ~n40408 & ~n40409;
  assign n40411 = n40407 & n40410;
  assign n40412 = ~n40404 & n40411;
  assign n40413 = n40403 & n40412;
  assign n40414 = ~pi3120 & ~n40413;
  assign n40415 = pi0868 & ~pi3516;
  assign n40416 = ~n25528 & ~n40415;
  assign n40417 = pi3120 & ~n40416;
  assign n40418 = ~n40414 & ~n40417;
  assign n40419 = ~pi0866 & ~n40418;
  assign n40420 = pi0866 & ~n12415;
  assign n40421 = ~n40419 & ~n40420;
  assign n40422 = po1281 & ~n40421;
  assign po1166 = n40400 | n40422;
  assign n40424 = ~n38903 & ~n38909;
  assign n40425 = ~n12726 & n40424;
  assign n40426 = pi0869 & n38909;
  assign po1167 = n40425 | n40426;
  assign n40428 = ~n9825 & ~n38903;
  assign n40429 = ~n38909 & n40428;
  assign n40430 = pi0870 & n38909;
  assign po1168 = n40429 | n40430;
  assign n40432 = ~n14403 & n40424;
  assign n40433 = pi0871 & n38909;
  assign po1169 = n40432 | n40433;
  assign n40435 = ~n15426 & ~n38903;
  assign n40436 = ~n38909 & n40435;
  assign n40437 = pi0872 & n38909;
  assign po1170 = n40436 | n40437;
  assign n40439 = ~pi3579 & ~n11181;
  assign n40440 = ~pi3464 & pi3579;
  assign n40441 = ~n40439 & ~n40440;
  assign n40442 = n39505 & ~n40441;
  assign n40443 = pi0873 & n39533;
  assign n40444 = ~pi0873 & ~n39533;
  assign n40445 = ~n40443 & ~n40444;
  assign n40446 = ~n39505 & n40445;
  assign po1171 = n40442 | n40446;
  assign n40448 = ~pi3579 & ~n14816;
  assign n40449 = ~pi3446 & pi3579;
  assign n40450 = ~n40448 & ~n40449;
  assign n40451 = n39505 & ~n40450;
  assign n40452 = ~pi0874 & ~n39511;
  assign n40453 = ~n39512 & ~n40452;
  assign n40454 = n39533 & ~n40453;
  assign n40455 = ~pi0874 & ~n39533;
  assign n40456 = ~n40454 & ~n40455;
  assign n40457 = ~n39505 & n40456;
  assign po1172 = n40451 | n40457;
  assign n40459 = ~pi0639 & n10210;
  assign n40460 = ~pi0641 & n40459;
  assign n40461 = ~pi0640 & n40460;
  assign n40462 = ~pi0634 & n40461;
  assign n40463 = ~pi0736 & n40462;
  assign n40464 = ~pi0638 & n40463;
  assign n40465 = ~pi0568 & ~n40464;
  assign n40466 = ~n10296 & n40465;
  assign n40467 = pi3451 & n40466;
  assign n40468 = ~pi0674 & n11532;
  assign n40469 = ~pi0656 & n40468;
  assign n40470 = ~pi0673 & n40469;
  assign n40471 = ~pi0657 & n40470;
  assign n40472 = ~pi0671 & n40471;
  assign n40473 = ~pi0672 & n40472;
  assign n40474 = pi0518 & ~pi3451;
  assign n40475 = ~n40473 & n40474;
  assign n40476 = n11665 & n40475;
  assign n40477 = pi0568 & pi3451;
  assign n40478 = ~n40464 & n40477;
  assign n40479 = n10362 & n40478;
  assign n40480 = ~pi0518 & ~n40473;
  assign n40481 = ~pi3451 & n40480;
  assign n40482 = ~n11615 & n40481;
  assign n40483 = ~n40479 & ~n40482;
  assign n40484 = ~n40476 & n40483;
  assign n40485 = ~n40467 & n40484;
  assign po1173 = pi3427 & ~n40485;
  assign n40487 = ~pi3579 & ~n13121;
  assign n40488 = ~pi3477 & pi3579;
  assign n40489 = ~n40487 & ~n40488;
  assign n40490 = n39505 & ~n40489;
  assign n40491 = ~pi0876 & ~n39544;
  assign n40492 = pi0876 & n39544;
  assign n40493 = ~n40491 & ~n40492;
  assign n40494 = n39533 & ~n40493;
  assign n40495 = ~pi0876 & ~n39533;
  assign n40496 = ~n40494 & ~n40495;
  assign n40497 = ~n39505 & n40496;
  assign po1174 = n40490 | n40497;
  assign po1175 = pi3395 & ~n40485;
  assign po1176 = pi3424 & ~n40485;
  assign po1177 = pi3429 & ~n40485;
  assign n40502 = ~n13121 & ~n38903;
  assign n40503 = ~n38916 & n40502;
  assign n40504 = pi0880 & n38916;
  assign po1178 = n40503 | n40504;
  assign n40506 = ~n13398 & ~n38903;
  assign n40507 = ~n38916 & n40506;
  assign n40508 = pi0881 & n38916;
  assign po1179 = n40507 | n40508;
  assign n40510 = ~n13988 & ~n38903;
  assign n40511 = ~n38916 & n40510;
  assign n40512 = pi0882 & n38916;
  assign po1180 = n40511 | n40512;
  assign n40514 = ~n12415 & ~n38903;
  assign n40515 = ~n38916 & n40514;
  assign n40516 = pi0883 & n38916;
  assign po1181 = n40515 | n40516;
  assign n40518 = ~n38903 & ~n38916;
  assign n40519 = ~n14816 & n40518;
  assign n40520 = pi0884 & n38916;
  assign po1182 = n40519 | n40520;
  assign n40522 = ~n15115 & n40518;
  assign n40523 = pi0885 & n38916;
  assign po1183 = n40522 | n40523;
  assign n40525 = ~n17368 & ~n38903;
  assign n40526 = ~n38916 & n40525;
  assign n40527 = pi0886 & n38916;
  assign po1184 = n40526 | n40527;
  assign n40529 = ~n17199 & ~n38903;
  assign n40530 = ~n38916 & n40529;
  assign n40531 = pi0887 & n38916;
  assign po1185 = n40530 | n40531;
  assign n40533 = ~n38916 & n40428;
  assign n40534 = pi0888 & n38916;
  assign po1186 = n40533 | n40534;
  assign n40536 = ~n10608 & ~n38903;
  assign n40537 = ~n38916 & n40536;
  assign n40538 = pi0889 & n38916;
  assign po1187 = n40537 | n40538;
  assign n40540 = n38901 & n38905;
  assign n40541 = ~n38904 & ~n40540;
  assign n40542 = ~n17199 & ~n40541;
  assign n40543 = pi0890 & n40541;
  assign n40544 = ~n40542 & ~n40543;
  assign n40545 = n38903 & ~n40541;
  assign po1188 = ~n40544 | n40545;
  assign n40547 = ~n14816 & ~n40541;
  assign n40548 = pi0891 & n40541;
  assign n40549 = ~n40547 & ~n40548;
  assign po1189 = n40545 | ~n40549;
  assign n40551 = ~n15115 & ~n40541;
  assign n40552 = pi0892 & n40541;
  assign n40553 = ~n40551 & ~n40552;
  assign po1190 = n40545 | ~n40553;
  assign n40555 = ~n17368 & ~n40541;
  assign n40556 = pi0893 & n40541;
  assign n40557 = ~n40555 & ~n40556;
  assign po1191 = n40545 | ~n40557;
  assign n40559 = ~n13701 & n40424;
  assign n40560 = pi0894 & n38909;
  assign po1192 = n40559 | n40560;
  assign n40562 = ~n38909 & n40525;
  assign n40563 = pi0895 & n38909;
  assign po1193 = n40562 | n40563;
  assign n40565 = ~n38909 & n40529;
  assign n40566 = pi0896 & n38909;
  assign po1194 = n40565 | n40566;
  assign n40568 = ~n38909 & n40536;
  assign n40569 = pi0897 & n38909;
  assign po1195 = n40568 | n40569;
  assign n40571 = ~pi1016 & ~pi1740;
  assign n40572 = ~pi1870 & ~pi1893;
  assign n40573 = ~pi1868 & ~pi1896;
  assign n40574 = ~pi1895 & n40573;
  assign n40575 = ~pi1871 & n40574;
  assign n40576 = n40572 & n40575;
  assign n40577 = ~pi1894 & n40576;
  assign n40578 = ~pi1435 & n40577;
  assign n40579 = ~pi1872 & n40578;
  assign n40580 = n40571 & n40579;
  assign n40581 = ~pi1094 & ~pi1097;
  assign n40582 = n40580 & n40581;
  assign n40583 = ~pi0946 & n40582;
  assign n40584 = ~pi1715 & n40583;
  assign n40585 = ~pi0898 & n40584;
  assign n40586 = pi0898 & ~n40584;
  assign n40587 = ~n40585 & ~n40586;
  assign n40588 = pi1871 & pi1887;
  assign n40589 = ~pi1871 & ~pi1887;
  assign n40590 = ~n40588 & ~n40589;
  assign n40591 = pi1888 & pi1895;
  assign n40592 = ~pi1888 & ~pi1895;
  assign n40593 = ~n40591 & ~n40592;
  assign n40594 = n40590 & n40593;
  assign n40595 = pi1862 & pi1868;
  assign n40596 = ~pi1862 & ~pi1868;
  assign n40597 = ~n40595 & ~n40596;
  assign n40598 = pi1873 & pi1896;
  assign n40599 = ~pi1873 & ~pi1896;
  assign n40600 = ~n40598 & ~n40599;
  assign n40601 = n40597 & n40600;
  assign n40602 = pi1094 & pi1892;
  assign n40603 = ~pi1094 & ~pi1892;
  assign n40604 = ~n40602 & ~n40603;
  assign n40605 = pi1016 & pi1891;
  assign n40606 = ~pi1016 & ~pi1891;
  assign n40607 = ~n40605 & ~n40606;
  assign n40608 = n40604 & n40607;
  assign n40609 = pi1872 & pi1952;
  assign n40610 = ~pi1872 & ~pi1952;
  assign n40611 = ~n40609 & ~n40610;
  assign n40612 = pi1435 & pi1883;
  assign n40613 = ~pi1435 & ~pi1883;
  assign n40614 = ~n40612 & ~n40613;
  assign n40615 = n40611 & n40614;
  assign n40616 = n40608 & n40615;
  assign n40617 = n40601 & n40616;
  assign n40618 = n40594 & n40617;
  assign n40619 = pi0898 & pi1889;
  assign n40620 = ~pi0898 & ~pi1889;
  assign n40621 = ~n40619 & ~n40620;
  assign n40622 = pi0946 & pi1869;
  assign n40623 = ~pi0946 & ~pi1869;
  assign n40624 = ~n40622 & ~n40623;
  assign n40625 = n40621 & n40624;
  assign n40626 = pi1715 & pi1890;
  assign n40627 = ~pi1715 & ~pi1890;
  assign n40628 = ~n40626 & ~n40627;
  assign n40629 = pi1097 & pi1874;
  assign n40630 = ~pi1097 & ~pi1874;
  assign n40631 = ~n40629 & ~n40630;
  assign n40632 = n40628 & n40631;
  assign n40633 = pi1740 & pi1884;
  assign n40634 = ~pi1740 & ~pi1884;
  assign n40635 = ~n40633 & ~n40634;
  assign n40636 = pi1885 & pi1893;
  assign n40637 = ~pi1885 & ~pi1893;
  assign n40638 = ~n40636 & ~n40637;
  assign n40639 = n40635 & n40638;
  assign n40640 = pi1870 & pi1920;
  assign n40641 = ~pi1870 & ~pi1920;
  assign n40642 = ~n40640 & ~n40641;
  assign n40643 = pi1886 & pi1894;
  assign n40644 = ~pi1886 & ~pi1894;
  assign n40645 = ~n40643 & ~n40644;
  assign n40646 = n40642 & n40645;
  assign n40647 = n40639 & n40646;
  assign n40648 = n40632 & n40647;
  assign n40649 = n40625 & n40648;
  assign n40650 = n40618 & n40649;
  assign n40651 = pi3647 & ~n40650;
  assign po1196 = n40587 & n40651;
  assign n40653 = ~pi0899 & n39355;
  assign n40654 = n15426 & ~n39355;
  assign n40655 = ~n40653 & ~n40654;
  assign po1197 = n39359 | n40655;
  assign n40657 = ~n12415 & ~n39351;
  assign n40658 = ~n39374 & n40657;
  assign n40659 = pi0900 & n39374;
  assign po1198 = n40658 | n40659;
  assign n40661 = ~pi1018 & ~pi1748;
  assign n40662 = ~pi1910 & ~pi1916;
  assign n40663 = ~pi1876 & ~pi1912;
  assign n40664 = ~pi1913 & n40663;
  assign n40665 = ~pi1914 & n40664;
  assign n40666 = n40662 & n40665;
  assign n40667 = ~pi1911 & n40666;
  assign n40668 = ~pi1448 & n40667;
  assign n40669 = ~pi1915 & n40668;
  assign n40670 = n40661 & n40669;
  assign n40671 = ~pi1095 & ~pi1098;
  assign n40672 = n40670 & n40671;
  assign n40673 = ~pi0973 & n40672;
  assign n40674 = ~pi1747 & n40673;
  assign n40675 = ~pi0901 & n40674;
  assign n40676 = pi0901 & ~n40674;
  assign n40677 = ~n40675 & ~n40676;
  assign n40678 = pi0901 & pi1903;
  assign n40679 = ~pi0901 & ~pi1903;
  assign n40680 = ~n40678 & ~n40679;
  assign n40681 = pi0973 & pi1904;
  assign n40682 = ~pi0973 & ~pi1904;
  assign n40683 = ~n40681 & ~n40682;
  assign n40684 = n40680 & n40683;
  assign n40685 = pi1747 & pi1905;
  assign n40686 = ~pi1747 & ~pi1905;
  assign n40687 = ~n40685 & ~n40686;
  assign n40688 = pi1098 & pi2053;
  assign n40689 = ~pi1098 & ~pi2053;
  assign n40690 = ~n40688 & ~n40689;
  assign n40691 = n40687 & n40690;
  assign n40692 = pi1901 & pi1914;
  assign n40693 = ~pi1901 & ~pi1914;
  assign n40694 = ~n40692 & ~n40693;
  assign n40695 = pi1902 & pi1913;
  assign n40696 = ~pi1902 & ~pi1913;
  assign n40697 = ~n40695 & ~n40696;
  assign n40698 = n40694 & n40697;
  assign n40699 = pi1912 & pi2052;
  assign n40700 = ~pi1912 & ~pi2052;
  assign n40701 = ~n40699 & ~n40700;
  assign n40702 = pi1876 & pi1907;
  assign n40703 = ~pi1876 & ~pi1907;
  assign n40704 = ~n40702 & ~n40703;
  assign n40705 = n40701 & n40704;
  assign n40706 = n40698 & n40705;
  assign n40707 = n40691 & n40706;
  assign n40708 = n40684 & n40707;
  assign n40709 = pi1748 & pi2055;
  assign n40710 = ~pi1748 & ~pi2055;
  assign n40711 = ~n40709 & ~n40710;
  assign n40712 = pi1899 & pi1910;
  assign n40713 = ~pi1899 & ~pi1910;
  assign n40714 = ~n40712 & ~n40713;
  assign n40715 = n40711 & n40714;
  assign n40716 = pi1916 & pi2054;
  assign n40717 = ~pi1916 & ~pi2054;
  assign n40718 = ~n40716 & ~n40717;
  assign n40719 = pi1900 & pi1911;
  assign n40720 = ~pi1900 & ~pi1911;
  assign n40721 = ~n40719 & ~n40720;
  assign n40722 = n40718 & n40721;
  assign n40723 = pi1095 & pi1906;
  assign n40724 = ~pi1095 & ~pi1906;
  assign n40725 = ~n40723 & ~n40724;
  assign n40726 = pi1018 & pi2051;
  assign n40727 = ~pi1018 & ~pi2051;
  assign n40728 = ~n40726 & ~n40727;
  assign n40729 = n40725 & n40728;
  assign n40730 = pi1915 & pi2057;
  assign n40731 = ~pi1915 & ~pi2057;
  assign n40732 = ~n40730 & ~n40731;
  assign n40733 = pi1448 & pi1898;
  assign n40734 = ~pi1448 & ~pi1898;
  assign n40735 = ~n40733 & ~n40734;
  assign n40736 = n40732 & n40735;
  assign n40737 = n40729 & n40736;
  assign n40738 = n40722 & n40737;
  assign n40739 = n40715 & n40738;
  assign n40740 = n40708 & n40739;
  assign n40741 = pi3635 & ~n40740;
  assign po1199 = n40677 & n40741;
  assign n40743 = ~pi3579 & ~n12726;
  assign n40744 = ~pi3445 & pi3579;
  assign n40745 = ~n40743 & ~n40744;
  assign n40746 = n39505 & ~n40745;
  assign n40747 = pi0876 & n39543;
  assign n40748 = pi0903 & n40747;
  assign n40749 = pi0907 & pi0908;
  assign n40750 = pi0906 & n40749;
  assign n40751 = pi0874 & n40750;
  assign n40752 = n40748 & n40751;
  assign n40753 = pi0873 & n40752;
  assign n40754 = pi0902 & n40753;
  assign n40755 = ~pi0902 & ~n40753;
  assign n40756 = ~n40754 & ~n40755;
  assign n40757 = n39533 & ~n40756;
  assign n40758 = ~pi0902 & ~n39533;
  assign n40759 = ~n40757 & ~n40758;
  assign n40760 = ~n39505 & n40759;
  assign po1200 = n40746 | n40760;
  assign n40762 = ~pi3579 & ~n13701;
  assign n40763 = ~pi3474 & pi3579;
  assign n40764 = ~n40762 & ~n40763;
  assign n40765 = n39505 & ~n40764;
  assign n40766 = ~pi0903 & ~n39516;
  assign n40767 = pi0903 & n39516;
  assign n40768 = ~n40766 & ~n40767;
  assign n40769 = n39533 & ~n40768;
  assign n40770 = ~pi0903 & ~n39533;
  assign n40771 = ~n40769 & ~n40770;
  assign n40772 = ~n39505 & n40771;
  assign po1201 = n40765 | n40772;
  assign n40774 = ~pi3579 & ~n13398;
  assign n40775 = ~pi3476 & pi3579;
  assign n40776 = ~n40774 & ~n40775;
  assign n40777 = n39505 & ~n40776;
  assign n40778 = pi0904 & n39514;
  assign n40779 = ~pi0904 & ~n39514;
  assign n40780 = ~n40778 & ~n40779;
  assign n40781 = n39533 & ~n40780;
  assign n40782 = ~pi0904 & ~n39533;
  assign n40783 = ~n40781 & ~n40782;
  assign n40784 = ~n39505 & n40783;
  assign po1202 = n40777 | n40784;
  assign n40786 = ~pi3579 & ~n13988;
  assign n40787 = ~pi3475 & pi3579;
  assign n40788 = ~n40786 & ~n40787;
  assign n40789 = n39505 & ~n40788;
  assign n40790 = pi0873 & n40751;
  assign n40791 = ~pi0905 & ~n40790;
  assign n40792 = pi0905 & n40790;
  assign n40793 = ~n40791 & ~n40792;
  assign n40794 = n39533 & ~n40793;
  assign n40795 = ~pi0905 & ~n39533;
  assign n40796 = ~n40794 & ~n40795;
  assign n40797 = ~n39505 & n40796;
  assign po1203 = n40789 | n40797;
  assign n40799 = ~pi3579 & ~n12415;
  assign n40800 = ~pi3470 & pi3579;
  assign n40801 = ~n40799 & ~n40800;
  assign n40802 = n39505 & ~n40801;
  assign n40803 = ~pi0906 & ~n39512;
  assign n40804 = ~n39513 & ~n40803;
  assign n40805 = n39533 & ~n40804;
  assign n40806 = ~pi0906 & ~n39533;
  assign n40807 = ~n40805 & ~n40806;
  assign n40808 = ~n39505 & n40807;
  assign po1204 = n40802 | n40808;
  assign n40810 = ~pi3579 & ~n15115;
  assign n40811 = ~pi3462 & pi3579;
  assign n40812 = ~n40810 & ~n40811;
  assign n40813 = n39505 & ~n40812;
  assign n40814 = ~pi0907 & ~n39510;
  assign n40815 = ~n39511 & ~n40814;
  assign n40816 = n39533 & ~n40815;
  assign n40817 = ~pi0907 & ~n39533;
  assign n40818 = ~n40816 & ~n40817;
  assign n40819 = ~n39505 & n40818;
  assign po1205 = n40813 | n40819;
  assign n40821 = ~pi0873 & pi0908;
  assign n40822 = pi0873 & ~pi0908;
  assign n40823 = ~n40821 & ~n40822;
  assign n40824 = n39533 & ~n40823;
  assign n40825 = pi0908 & ~n39533;
  assign n40826 = ~n40824 & ~n40825;
  assign n40827 = ~n39505 & ~n40826;
  assign n40828 = ~pi3579 & ~n12061;
  assign n40829 = ~pi3468 & pi3579;
  assign n40830 = ~n40828 & ~n40829;
  assign n40831 = n39505 & ~n40830;
  assign po1206 = n40827 | n40831;
  assign n40833 = ~pi3579 & ~n9825;
  assign n40834 = ~pi3466 & pi3579;
  assign n40835 = ~n40833 & ~n40834;
  assign n40836 = n39505 & ~n40835;
  assign n40837 = pi0910 & n40790;
  assign n40838 = n40748 & n40837;
  assign n40839 = pi0820 & n40838;
  assign n40840 = pi0902 & n40839;
  assign n40841 = pi0819 & n40840;
  assign n40842 = pi0909 & n40841;
  assign n40843 = ~pi0909 & ~n40841;
  assign n40844 = ~n40842 & ~n40843;
  assign n40845 = n39533 & ~n40844;
  assign n40846 = ~pi0909 & ~n39533;
  assign n40847 = ~n40845 & ~n40846;
  assign n40848 = ~n39505 & n40847;
  assign po1207 = n40836 | n40848;
  assign n40850 = ~pi3579 & ~n14403;
  assign n40851 = ~pi3448 & pi3579;
  assign n40852 = ~n40850 & ~n40851;
  assign n40853 = n39505 & ~n40852;
  assign n40854 = n39515 & n39517;
  assign n40855 = n39514 & n40854;
  assign n40856 = pi0910 & n40855;
  assign n40857 = ~pi0910 & ~n40855;
  assign n40858 = ~n40856 & ~n40857;
  assign n40859 = n39533 & ~n40858;
  assign n40860 = ~pi0910 & ~n39533;
  assign n40861 = ~n40859 & ~n40860;
  assign n40862 = ~n39505 & n40861;
  assign po1208 = n40853 | n40862;
  assign n40864 = ~pi1075 & n38779;
  assign n40865 = ~pi1670 & n38781;
  assign n40866 = ~n40864 & ~n40865;
  assign n40867 = pi0393 & n38792;
  assign n40868 = ~pi0427 & n38789;
  assign n40869 = ~n40867 & ~n40868;
  assign n40870 = n40866 & n40869;
  assign n40871 = ~n38745 & ~n40870;
  assign n40872 = n38798 & n40871;
  assign n40873 = ~pi0911 & n38745;
  assign n40874 = ~n40872 & ~n40873;
  assign n40875 = ~pi1052 & ~n38745;
  assign n40876 = ~n38800 & n40875;
  assign n40877 = ~n38798 & n40876;
  assign po1209 = ~n40874 | n40877;
  assign n40879 = ~pi2017 & ~pi2474;
  assign n40880 = pi3293 & ~n40879;
  assign n40881 = pi1598 & pi3293;
  assign n40882 = ~n38533 & ~n40881;
  assign n40883 = n38538 & n40882;
  assign n40884 = pi1597 & pi3293;
  assign n40885 = pi2019 & pi3293;
  assign n40886 = pi2018 & pi3293;
  assign n40887 = ~n40885 & ~n40886;
  assign n40888 = ~n40884 & n40887;
  assign n40889 = n40883 & n40888;
  assign n40890 = ~n40880 & n40889;
  assign n40891 = pi0912 & ~n40890;
  assign n40892 = n38509 & n40891;
  assign n40893 = ~pi1463 & n20345;
  assign n40894 = ~pi1536 & n20347;
  assign n40895 = ~n40893 & ~n40894;
  assign n40896 = ~pi1464 & n20350;
  assign n40897 = ~pi1571 & n20353;
  assign n40898 = ~pi1408 & n20356;
  assign n40899 = ~n40897 & ~n40898;
  assign n40900 = ~pi1500 & n20360;
  assign n40901 = ~pi1482 & n20363;
  assign n40902 = ~n40900 & ~n40901;
  assign n40903 = n40899 & n40902;
  assign n40904 = ~n40896 & n40903;
  assign n40905 = n40895 & n40904;
  assign n40906 = ~pi1007 & ~n40905;
  assign n40907 = pi1007 & ~n12726;
  assign n40908 = ~n40906 & ~n40907;
  assign n40909 = ~n38527 & n40908;
  assign n40910 = ~pi0912 & n38527;
  assign n40911 = ~n40909 & ~n40910;
  assign n40912 = ~n38509 & n40911;
  assign po1210 = n40892 | n40912;
  assign n40914 = pi2017 & pi3293;
  assign n40915 = n40888 & ~n40914;
  assign n40916 = n40883 & n40915;
  assign n40917 = pi0913 & ~n40916;
  assign n40918 = n38509 & n40917;
  assign n40919 = ~pi1627 & n20360;
  assign n40920 = ~pi1483 & n20363;
  assign n40921 = ~n40919 & ~n40920;
  assign n40922 = ~pi1618 & n20353;
  assign n40923 = ~pi1554 & n20356;
  assign n40924 = ~n40922 & ~n40923;
  assign n40925 = ~pi1518 & n20345;
  assign n40926 = ~pi1537 & n20347;
  assign n40927 = ~n40925 & ~n40926;
  assign n40928 = ~pi1586 & n20350;
  assign n40929 = n40927 & ~n40928;
  assign n40930 = n40924 & n40929;
  assign n40931 = n40921 & n40930;
  assign n40932 = ~pi1007 & ~n40931;
  assign n40933 = pi1007 & ~n13701;
  assign n40934 = ~n40932 & ~n40933;
  assign n40935 = ~n38527 & n40934;
  assign n40936 = ~pi0913 & n38527;
  assign n40937 = ~n40935 & ~n40936;
  assign n40938 = ~n38509 & n40937;
  assign po1211 = n40918 | n40938;
  assign n40940 = ~pi1501 & n20360;
  assign n40941 = ~pi1400 & n20363;
  assign n40942 = ~n40940 & ~n40941;
  assign n40943 = ~pi1572 & n20353;
  assign n40944 = ~pi1404 & n20356;
  assign n40945 = ~n40943 & ~n40944;
  assign n40946 = ~pi1519 & n20345;
  assign n40947 = ~pi1538 & n20347;
  assign n40948 = ~n40946 & ~n40947;
  assign n40949 = ~pi1475 & n20350;
  assign n40950 = n40948 & ~n40949;
  assign n40951 = n40945 & n40950;
  assign n40952 = n40942 & n40951;
  assign n40953 = ~pi1007 & ~n40952;
  assign n40954 = pi1007 & ~n13121;
  assign n40955 = ~n40953 & ~n40954;
  assign n40956 = ~n38527 & n40955;
  assign n40957 = ~pi0914 & n38527;
  assign n40958 = ~n40956 & ~n40957;
  assign n40959 = ~n38509 & n40958;
  assign n40960 = pi0914 & n38509;
  assign n40961 = ~n40889 & n40960;
  assign po1212 = n40959 | n40961;
  assign n40963 = pi0915 & n38509;
  assign n40964 = n40883 & n40887;
  assign n40965 = n40963 & ~n40964;
  assign n40966 = ~pi1520 & n20345;
  assign n40967 = ~pi1416 & n20347;
  assign n40968 = ~n40966 & ~n40967;
  assign n40969 = ~pi1587 & n20350;
  assign n40970 = ~pi1502 & n20360;
  assign n40971 = ~pi1484 & n20363;
  assign n40972 = ~n40970 & ~n40971;
  assign n40973 = ~pi1628 & n20353;
  assign n40974 = ~pi1555 & n20356;
  assign n40975 = ~n40973 & ~n40974;
  assign n40976 = n40972 & n40975;
  assign n40977 = ~n40969 & n40976;
  assign n40978 = n40968 & n40977;
  assign n40979 = ~pi1007 & ~n40978;
  assign n40980 = pi1007 & ~n13398;
  assign n40981 = ~n40979 & ~n40980;
  assign n40982 = ~n38527 & n40981;
  assign n40983 = ~pi0915 & n38527;
  assign n40984 = ~n40982 & ~n40983;
  assign n40985 = ~n38509 & n40984;
  assign po1213 = n40965 | n40985;
  assign n40987 = pi0916 & n38509;
  assign n40988 = n38538 & ~n40885;
  assign n40989 = n40882 & n40988;
  assign n40990 = n40987 & ~n40989;
  assign n40991 = ~pi1395 & n20345;
  assign n40992 = ~pi1539 & n20347;
  assign n40993 = ~n40991 & ~n40992;
  assign n40994 = ~pi1466 & n20350;
  assign n40995 = ~pi1573 & n20353;
  assign n40996 = ~pi1556 & n20356;
  assign n40997 = ~n40995 & ~n40996;
  assign n40998 = ~pi1503 & n20360;
  assign n40999 = ~pi1398 & n20363;
  assign n41000 = ~n40998 & ~n40999;
  assign n41001 = n40997 & n41000;
  assign n41002 = ~n40994 & n41001;
  assign n41003 = n40993 & n41002;
  assign n41004 = ~pi1007 & ~n41003;
  assign n41005 = pi1007 & ~n13988;
  assign n41006 = ~n41004 & ~n41005;
  assign n41007 = ~n38527 & n41006;
  assign n41008 = ~pi0916 & n38527;
  assign n41009 = ~n41007 & ~n41008;
  assign n41010 = ~n38509 & n41009;
  assign po1214 = n40990 | n41010;
  assign n41012 = ~pi1504 & n20360;
  assign n41013 = ~pi1397 & n20363;
  assign n41014 = ~n41012 & ~n41013;
  assign n41015 = ~pi1574 & n20353;
  assign n41016 = ~pi1405 & n20356;
  assign n41017 = ~n41015 & ~n41016;
  assign n41018 = ~pi1522 & n20345;
  assign n41019 = ~pi1541 & n20347;
  assign n41020 = ~n41018 & ~n41019;
  assign n41021 = ~pi1589 & n20350;
  assign n41022 = n41020 & ~n41021;
  assign n41023 = n41017 & n41022;
  assign n41024 = n41014 & n41023;
  assign n41025 = ~pi1007 & ~n41024;
  assign n41026 = pi1007 & ~n12415;
  assign n41027 = ~n41025 & ~n41026;
  assign n41028 = ~n38527 & n41027;
  assign n41029 = ~pi0917 & n38527;
  assign n41030 = ~n41028 & ~n41029;
  assign n41031 = ~n38509 & n41030;
  assign n41032 = pi0917 & n38509;
  assign n41033 = ~n40883 & n41032;
  assign po1215 = n41031 | n41033;
  assign n41035 = ~pi1505 & n20360;
  assign n41036 = ~pi1487 & n20363;
  assign n41037 = ~n41035 & ~n41036;
  assign n41038 = ~pi1575 & n20353;
  assign n41039 = ~pi1559 & n20356;
  assign n41040 = ~n41038 & ~n41039;
  assign n41041 = ~pi1419 & n20345;
  assign n41042 = ~pi1542 & n20347;
  assign n41043 = ~n41041 & ~n41042;
  assign n41044 = ~pi1393 & n20350;
  assign n41045 = n41043 & ~n41044;
  assign n41046 = n41040 & n41045;
  assign n41047 = n41037 & n41046;
  assign n41048 = ~pi1007 & ~n41047;
  assign n41049 = pi1007 & ~n15115;
  assign n41050 = ~n41048 & ~n41049;
  assign n41051 = ~n38527 & n41050;
  assign n41052 = ~pi0918 & n38527;
  assign n41053 = ~n41051 & ~n41052;
  assign n41054 = ~n38509 & n41053;
  assign n41055 = pi0918 & n38509;
  assign n41056 = ~n38538 & n41055;
  assign po1216 = n41054 | n41056;
  assign n41058 = pi0919 & n38509;
  assign n41059 = n38537 & n41058;
  assign n41060 = ~pi1524 & n20345;
  assign n41061 = ~pi1543 & n20347;
  assign n41062 = ~n41060 & ~n41061;
  assign n41063 = ~pi1591 & n20350;
  assign n41064 = ~pi1623 & n20353;
  assign n41065 = ~pi1560 & n20356;
  assign n41066 = ~n41064 & ~n41065;
  assign n41067 = ~pi1622 & n20360;
  assign n41068 = ~pi1488 & n20363;
  assign n41069 = ~n41067 & ~n41068;
  assign n41070 = n41066 & n41069;
  assign n41071 = ~n41063 & n41070;
  assign n41072 = n41062 & n41071;
  assign n41073 = ~pi1007 & ~n41072;
  assign n41074 = pi1007 & ~n12061;
  assign n41075 = ~n41073 & ~n41074;
  assign n41076 = ~n38527 & n41075;
  assign n41077 = ~pi0919 & n38527;
  assign n41078 = ~n41076 & ~n41077;
  assign n41079 = ~n38509 & n41078;
  assign po1217 = n41059 | n41079;
  assign n41081 = ~n8561 & n36084;
  assign n41082 = n36078 & n41081;
  assign n41083 = ~n36063 & n39096;
  assign n41084 = n41082 & n41083;
  assign n41085 = ~pi0920 & n8561;
  assign n41086 = ~n41084 & ~n41085;
  assign po1218 = po3627 & ~n41086;
  assign n41088 = n38864 & n39861;
  assign n41089 = ~pi0921 & n8561;
  assign n41090 = ~n41088 & ~n41089;
  assign po1219 = po3627 & ~n41090;
  assign n41092 = ~pi3252 & n39892;
  assign n41093 = ~pi0445 & n41092;
  assign n41094 = ~pi3252 & ~n39899;
  assign n41095 = ~pi0440 & n41094;
  assign n41096 = pi0922 & ~n41094;
  assign n41097 = ~n41095 & ~n41096;
  assign n41098 = ~pi3252 & ~n39890;
  assign n41099 = ~n41097 & ~n41098;
  assign n41100 = ~pi0453 & n41098;
  assign n41101 = ~n41099 & ~n41100;
  assign n41102 = ~n41092 & ~n41101;
  assign po1220 = n41093 | n41102;
  assign n41104 = ~pi0446 & n41092;
  assign n41105 = ~pi0441 & n41094;
  assign n41106 = pi0923 & ~n41094;
  assign n41107 = ~n41105 & ~n41106;
  assign n41108 = ~n41098 & ~n41107;
  assign n41109 = ~pi0454 & n41098;
  assign n41110 = ~n41108 & ~n41109;
  assign n41111 = ~n41092 & ~n41110;
  assign po1221 = n41104 | n41111;
  assign n41113 = ~pi0447 & n41092;
  assign n41114 = ~pi0442 & n41094;
  assign n41115 = pi0924 & ~n41094;
  assign n41116 = ~n41114 & ~n41115;
  assign n41117 = ~n41098 & ~n41116;
  assign n41118 = ~pi0461 & n41098;
  assign n41119 = ~n41117 & ~n41118;
  assign n41120 = ~n41092 & ~n41119;
  assign po1222 = n41113 | n41120;
  assign n41122 = ~pi0450 & n41092;
  assign n41123 = ~pi0444 & n41094;
  assign n41124 = pi0925 & ~n41094;
  assign n41125 = ~n41123 & ~n41124;
  assign n41126 = ~n41098 & ~n41125;
  assign n41127 = ~pi0456 & n41098;
  assign n41128 = ~n41126 & ~n41127;
  assign n41129 = ~n41092 & ~n41128;
  assign po1223 = n41122 | n41129;
  assign n41131 = ~pi0451 & n41092;
  assign n41132 = ~pi0459 & n41094;
  assign n41133 = pi0926 & ~n41094;
  assign n41134 = ~n41132 & ~n41133;
  assign n41135 = ~n41098 & ~n41134;
  assign n41136 = ~pi0457 & n41098;
  assign n41137 = ~n41135 & ~n41136;
  assign n41138 = ~n41092 & ~n41137;
  assign po1224 = n41131 | n41138;
  assign n41140 = ~pi0462 & n41092;
  assign n41141 = ~pi0449 & n41094;
  assign n41142 = pi0927 & ~n41094;
  assign n41143 = ~n41141 & ~n41142;
  assign n41144 = ~n41098 & ~n41143;
  assign n41145 = ~pi0438 & n41098;
  assign n41146 = ~n41144 & ~n41145;
  assign n41147 = ~n41092 & ~n41146;
  assign po1225 = n41140 | n41147;
  assign n41149 = ~n13701 & n38320;
  assign n41150 = pi0928 & n38310;
  assign n41151 = ~pi0928 & ~n38310;
  assign n41152 = ~n41150 & ~n41151;
  assign n41153 = ~n36181 & ~n41152;
  assign n41154 = ~pi0928 & n36181;
  assign n41155 = ~n41153 & ~n41154;
  assign n41156 = ~n38320 & n41155;
  assign po1226 = n41149 | n41156;
  assign n41158 = ~n9825 & n38320;
  assign n41159 = pi1474 & pi1603;
  assign n41160 = pi1602 & n41159;
  assign n41161 = pi0928 & n41160;
  assign n41162 = pi1090 & n41161;
  assign n41163 = pi2058 & n38304;
  assign n41164 = pi2058 & n38301;
  assign n41165 = ~n41163 & ~n41164;
  assign n41166 = pi1467 & pi1841;
  assign n41167 = ~n41165 & n41166;
  assign n41168 = n41162 & n41167;
  assign n41169 = pi0930 & n41168;
  assign n41170 = pi1066 & n41169;
  assign n41171 = pi0688 & n41170;
  assign n41172 = pi0929 & n41171;
  assign n41173 = ~pi0929 & ~n41171;
  assign n41174 = ~n41172 & ~n41173;
  assign n41175 = ~n36181 & ~n41174;
  assign n41176 = ~pi0929 & n36181;
  assign n41177 = ~n41175 & ~n41176;
  assign n41178 = ~n38320 & n41177;
  assign po1227 = n41158 | n41178;
  assign n41180 = ~n15426 & n38320;
  assign n41181 = n41159 & ~n41165;
  assign n41182 = n41166 & n41181;
  assign n41183 = n38311 & n41182;
  assign n41184 = pi1090 & n41183;
  assign n41185 = pi1602 & n41184;
  assign n41186 = pi0930 & n41185;
  assign n41187 = ~pi0930 & ~n41185;
  assign n41188 = ~n41186 & ~n41187;
  assign n41189 = ~n36181 & ~n41188;
  assign n41190 = ~pi0930 & n36181;
  assign n41191 = ~n41189 & ~n41190;
  assign n41192 = ~n38320 & n41191;
  assign po1228 = n41180 | n41192;
  assign n41194 = pi0931 & pi3647;
  assign n41195 = ~pi0931 & ~pi3647;
  assign n41196 = ~n41194 & ~n41195;
  assign n41197 = n36877 & ~n41196;
  assign n41198 = pi0748 & n36876;
  assign po1229 = n41197 | n41198;
  assign n41200 = pi0932 & n37354;
  assign n41201 = ~pi0932 & ~n37354;
  assign n41202 = ~n41200 & ~n41201;
  assign n41203 = pi3647 & ~n41202;
  assign n41204 = ~pi0932 & ~pi3647;
  assign n41205 = ~n41203 & ~n41204;
  assign n41206 = n36877 & ~n41205;
  assign n41207 = pi0743 & n36876;
  assign po1230 = n41206 | n41207;
  assign n41209 = pi0933 & pi3635;
  assign n41210 = ~pi0933 & ~pi3635;
  assign n41211 = ~n41209 & ~n41210;
  assign n41212 = n36969 & ~n41211;
  assign n41213 = pi0805 & n36968;
  assign po1231 = n41212 | n41213;
  assign n41215 = pi0934 & n37373;
  assign n41216 = ~pi0934 & ~n37373;
  assign n41217 = ~n41215 & ~n41216;
  assign n41218 = pi3635 & ~n41217;
  assign n41219 = ~pi0934 & ~pi3635;
  assign n41220 = ~n41218 & ~n41219;
  assign n41221 = n36969 & ~n41220;
  assign n41222 = pi0801 & n36968;
  assign po1232 = n41221 | n41222;
  assign n41224 = pi0935 & ~pi3635;
  assign n41225 = ~pi0935 & n36887;
  assign n41226 = pi0935 & ~n36887;
  assign n41227 = ~n41225 & ~n41226;
  assign n41228 = pi3635 & ~n41227;
  assign n41229 = ~n41224 & ~n41228;
  assign n41230 = n36969 & n41229;
  assign n41231 = pi0800 & n36968;
  assign po1233 = n41230 | n41231;
  assign po1234 = pi3568 & po0767;
  assign n41234 = pi1668 & pi3681;
  assign n41235 = ~pi1668 & ~pi3681;
  assign n41236 = ~n41234 & ~n41235;
  assign n41237 = ~pi1695 & ~pi3681;
  assign n41238 = pi1695 & pi3681;
  assign n41239 = ~n41237 & ~n41238;
  assign n41240 = ~pi2416 & ~pi3681;
  assign n41241 = pi2416 & pi3681;
  assign n41242 = ~n41240 & ~n41241;
  assign n41243 = ~n41239 & ~n41242;
  assign n41244 = ~pi1851 & n41243;
  assign n41245 = ~n41236 & n41244;
  assign n41246 = ~pi3247 & ~pi3290;
  assign n41247 = ~pi2824 & n41246;
  assign n41248 = ~pi2510 & n41247;
  assign n41249 = n41245 & n41248;
  assign n41250 = pi1380 & pi3681;
  assign n41251 = ~pi1380 & ~pi3681;
  assign n41252 = ~n41250 & ~n41251;
  assign n41253 = ~pi1081 & ~pi3681;
  assign n41254 = pi1081 & pi3681;
  assign n41255 = ~n41253 & ~n41254;
  assign n41256 = ~pi1379 & ~pi3681;
  assign n41257 = pi1379 & pi3681;
  assign n41258 = ~n41256 & ~n41257;
  assign n41259 = ~n41255 & ~n41258;
  assign n41260 = ~n41252 & n41259;
  assign n41261 = n41249 & n41260;
  assign n41262 = pi1908 & pi1917;
  assign n41263 = pi1788 & pi3681;
  assign n41264 = ~pi1788 & ~pi3681;
  assign n41265 = ~n41263 & ~n41264;
  assign n41266 = n41262 & ~n41265;
  assign n41267 = n41261 & n41266;
  assign n41268 = ~pi1006 & ~n41262;
  assign n41269 = ~n41267 & ~n41268;
  assign n41270 = ~pi0936 & n41269;
  assign po1236 = ~pi3583 & ~n41270;
  assign n41272 = ~pi0937 & n38745;
  assign n41273 = ~pi2882 & n38752;
  assign n41274 = ~pi3047 & n38770;
  assign n41275 = ~n41273 & ~n41274;
  assign n41276 = pi0413 & n38789;
  assign n41277 = ~pi1699 & n38781;
  assign n41278 = ~n41276 & ~n41277;
  assign n41279 = pi0386 & n38792;
  assign n41280 = n41278 & ~n41279;
  assign n41281 = n41275 & n41280;
  assign n41282 = ~pi1079 & n38779;
  assign n41283 = n41281 & ~n41282;
  assign n41284 = n38798 & ~n41283;
  assign n41285 = ~pi1045 & n38800;
  assign n41286 = pi0821 & ~n38800;
  assign n41287 = ~n41285 & ~n41286;
  assign n41288 = ~n38798 & ~n41287;
  assign n41289 = ~n41284 & ~n41288;
  assign n41290 = ~n38745 & ~n41289;
  assign po1237 = n41272 | n41290;
  assign n41292 = pi0938 & n38745;
  assign n41293 = ~pi2903 & n38749;
  assign n41294 = ~pi3110 & n38752;
  assign n41295 = ~n41293 & ~n41294;
  assign n41296 = ~pi3072 & n38757;
  assign n41297 = ~pi3019 & n38760;
  assign n41298 = ~n41296 & ~n41297;
  assign n41299 = ~pi1669 & n38781;
  assign n41300 = ~pi1362 & n38779;
  assign n41301 = ~pi2762 & n38764;
  assign n41302 = ~n41300 & ~n41301;
  assign n41303 = ~pi3062 & n38775;
  assign n41304 = ~pi2791 & n38770;
  assign n41305 = ~n41303 & ~n41304;
  assign n41306 = ~n38769 & n41305;
  assign n41307 = n41302 & n41306;
  assign n41308 = ~n41299 & n41307;
  assign n41309 = ~pi2821 & n38772;
  assign n41310 = ~pi3108 & n38766;
  assign n41311 = ~n41309 & ~n41310;
  assign n41312 = n41308 & n41311;
  assign n41313 = pi0818 & n38787;
  assign n41314 = pi0426 & n38789;
  assign n41315 = ~n41313 & ~n41314;
  assign n41316 = pi0392 & n38792;
  assign n41317 = n41315 & ~n41316;
  assign n41318 = n41312 & n41317;
  assign n41319 = n41298 & n41318;
  assign n41320 = n41295 & n41319;
  assign n41321 = n38798 & ~n41320;
  assign n41322 = pi0851 & n38800;
  assign n41323 = pi0731 & ~n38800;
  assign n41324 = ~n41322 & ~n41323;
  assign n41325 = ~n38798 & ~n41324;
  assign n41326 = ~n41321 & ~n41325;
  assign n41327 = ~n38745 & ~n41326;
  assign po1238 = n41292 | n41327;
  assign n41329 = pi3410 & ~pi3416;
  assign po1239 = po1235 & ~n41329;
  assign n41331 = n38259 & ~po3745;
  assign n41332 = pi3330 & ~pi3392;
  assign n41333 = pi3394 & n41332;
  assign n41334 = ~pi3382 & ~n41333;
  assign n41335 = pi3410 & n41334;
  assign n41336 = ~pi0939 & ~n41335;
  assign n41337 = ~pi3416 & n41335;
  assign n41338 = ~n41336 & ~n41337;
  assign po1240 = n41331 & n41338;
  assign n41340 = pi0940 & n36795;
  assign n41341 = ~pi0940 & ~n36795;
  assign n41342 = ~n41340 & ~n41341;
  assign n41343 = pi3647 & ~n41342;
  assign n41344 = ~pi0940 & ~pi3647;
  assign n41345 = ~n41343 & ~n41344;
  assign n41346 = n36877 & ~n41345;
  assign n41347 = pi0742 & n36876;
  assign po1241 = n41346 | n41347;
  assign n41349 = ~pi0941 & n39355;
  assign n41350 = n13701 & ~n39355;
  assign n41351 = ~n41349 & ~n41350;
  assign po1242 = n39359 | n41351;
  assign n41353 = ~pi0452 & n41092;
  assign n41354 = ~pi0460 & n41094;
  assign n41355 = pi0942 & ~n41094;
  assign n41356 = ~n41354 & ~n41355;
  assign n41357 = ~n41098 & ~n41356;
  assign n41358 = ~pi0439 & n41098;
  assign n41359 = ~n41357 & ~n41358;
  assign n41360 = ~n41092 & ~n41359;
  assign po1243 = n41353 | n41360;
  assign n41362 = ~pi0448 & n41092;
  assign n41363 = ~pi0443 & n41094;
  assign n41364 = pi0943 & ~n41094;
  assign n41365 = ~n41363 & ~n41364;
  assign n41366 = ~n41098 & ~n41365;
  assign n41367 = ~pi0455 & n41098;
  assign n41368 = ~n41366 & ~n41367;
  assign n41369 = ~n41092 & ~n41368;
  assign po1244 = n41362 | n41369;
  assign n41371 = ~n8561 & ~n36123;
  assign n41372 = pi0944 & n8561;
  assign n41373 = ~n41371 & ~n41372;
  assign po1245 = po3627 & n41373;
  assign n41375 = n36063 & n39093;
  assign n41376 = n36066 & n36069;
  assign n41377 = n39094 & n41376;
  assign n41378 = n41375 & n41377;
  assign n41379 = ~pi0945 & n8561;
  assign n41380 = ~n41378 & ~n41379;
  assign po1246 = po3627 & ~n41380;
  assign n41382 = ~pi1894 & n40575;
  assign n41383 = ~pi1870 & n41382;
  assign n41384 = ~pi1435 & ~pi1872;
  assign n41385 = n41383 & n41384;
  assign n41386 = ~pi1740 & ~pi1893;
  assign n41387 = n41385 & n41386;
  assign n41388 = ~pi1016 & ~pi1094;
  assign n41389 = n41387 & n41388;
  assign n41390 = ~pi1715 & n41389;
  assign n41391 = ~pi1097 & n41390;
  assign n41392 = ~pi0946 & n41391;
  assign n41393 = pi0946 & ~n41391;
  assign n41394 = ~n41392 & ~n41393;
  assign po1247 = n40651 & n41394;
  assign n41396 = pi0947 & n40541;
  assign n41397 = ~n9825 & ~n40541;
  assign po1248 = n41396 | n41397;
  assign n41399 = pi0948 & n40541;
  assign n41400 = n40502 & ~n40541;
  assign po1249 = n41399 | n41400;
  assign n41402 = pi0949 & n40541;
  assign n41403 = n40506 & ~n40541;
  assign po1250 = n41402 | n41403;
  assign n41405 = pi0950 & n40541;
  assign n41406 = n40510 & ~n40541;
  assign po1251 = n41405 | n41406;
  assign n41408 = pi0951 & n40541;
  assign n41409 = n40514 & ~n40541;
  assign po1252 = n41408 | n41409;
  assign n41411 = ~n12061 & ~n38903;
  assign n41412 = ~n40541 & n41411;
  assign n41413 = pi0952 & n40541;
  assign po1253 = n41412 | n41413;
  assign n41415 = ~n11181 & ~n38903;
  assign n41416 = ~n40541 & n41415;
  assign n41417 = pi0953 & n40541;
  assign po1254 = n41416 | n41417;
  assign n41419 = ~n13398 & ~n39351;
  assign n41420 = ~n39355 & n41419;
  assign n41421 = pi0954 & n39355;
  assign po1255 = n41420 | n41421;
  assign n41423 = ~n13988 & ~n39351;
  assign n41424 = ~n39355 & n41423;
  assign n41425 = pi0955 & n39355;
  assign po1256 = n41424 | n41425;
  assign n41427 = ~n13121 & ~n39351;
  assign n41428 = ~n39355 & n41427;
  assign n41429 = pi0956 & n39355;
  assign po1257 = n41428 | n41429;
  assign n41431 = ~n39351 & ~n39355;
  assign n41432 = ~n14816 & n41431;
  assign n41433 = pi0957 & n39355;
  assign po1258 = n41432 | n41433;
  assign n41435 = ~n17368 & ~n39351;
  assign n41436 = ~n39355 & n41435;
  assign n41437 = pi0958 & n39355;
  assign po1259 = n41436 | n41437;
  assign n41439 = ~n17199 & ~n39351;
  assign n41440 = ~n39355 & n41439;
  assign n41441 = pi0959 & n39355;
  assign po1260 = n41440 | n41441;
  assign n41443 = ~n9825 & ~n39351;
  assign n41444 = ~n39355 & n41443;
  assign n41445 = pi0960 & n39355;
  assign po1261 = n41444 | n41445;
  assign n41447 = ~n10608 & ~n39351;
  assign n41448 = ~n39355 & n41447;
  assign n41449 = pi0961 & n39355;
  assign po1262 = n41448 | n41449;
  assign n41451 = pi0962 & n39374;
  assign n41452 = ~n9825 & ~n39374;
  assign po1263 = n41451 | n41452;
  assign n41454 = pi0963 & n39374;
  assign n41455 = ~n39374 & n41427;
  assign po1264 = n41454 | n41455;
  assign n41457 = pi0964 & n39374;
  assign n41458 = ~n39374 & n41419;
  assign po1265 = n41457 | n41458;
  assign n41460 = pi0965 & n39374;
  assign n41461 = ~n39374 & n41423;
  assign po1266 = n41460 | n41461;
  assign n41463 = ~n12061 & ~n39351;
  assign n41464 = ~n39374 & n41463;
  assign n41465 = pi0966 & n39374;
  assign po1267 = n41464 | n41465;
  assign n41467 = ~n11181 & ~n39351;
  assign n41468 = ~n39374 & n41467;
  assign n41469 = pi0967 & n39374;
  assign po1268 = n41468 | n41469;
  assign n41471 = ~n39351 & ~n39393;
  assign n41472 = ~n13701 & n41471;
  assign n41473 = pi0968 & n39393;
  assign po1269 = n41472 | n41473;
  assign n41475 = ~n39393 & n41435;
  assign n41476 = pi0969 & n39393;
  assign po1270 = n41475 | n41476;
  assign n41478 = ~n39393 & n41439;
  assign n41479 = pi0970 & n39393;
  assign po1271 = n41478 | n41479;
  assign n41481 = ~n15426 & ~n39351;
  assign n41482 = ~n39393 & n41481;
  assign n41483 = pi0971 & n39393;
  assign po1272 = n41482 | n41483;
  assign n41485 = ~n39393 & n41447;
  assign n41486 = pi0972 & n39393;
  assign po1273 = n41485 | n41486;
  assign n41488 = ~pi1911 & n40665;
  assign n41489 = ~pi1916 & n41488;
  assign n41490 = ~pi1448 & ~pi1915;
  assign n41491 = n41489 & n41490;
  assign n41492 = ~pi1748 & ~pi1910;
  assign n41493 = n41491 & n41492;
  assign n41494 = ~pi1018 & ~pi1095;
  assign n41495 = n41493 & n41494;
  assign n41496 = ~pi1747 & n41495;
  assign n41497 = ~pi1098 & n41496;
  assign n41498 = ~pi0973 & n41497;
  assign n41499 = pi0973 & ~n41497;
  assign n41500 = ~n41498 & ~n41499;
  assign po1274 = n40741 & n41500;
  assign n41502 = pi1761 & pi1762;
  assign n41503 = ~pi0609 & n41502;
  assign n41504 = ~pi3243 & ~n41503;
  assign n41505 = ~pi1761 & n41504;
  assign n41506 = ~pi1761 & ~n41503;
  assign n41507 = ~pi1012 & ~pi1033;
  assign n41508 = pi1034 & n41507;
  assign n41509 = pi1039 & n41508;
  assign n41510 = n39500 & n41509;
  assign n41511 = ~n41503 & n41510;
  assign n41512 = ~pi0974 & ~n41511;
  assign n41513 = ~n41506 & ~n41512;
  assign n41514 = n9825 & n41511;
  assign n41515 = n41513 & ~n41514;
  assign po1275 = n41505 | n41515;
  assign n41517 = ~pi1422 & ~n39531;
  assign n41518 = ~pi0975 & ~n41517;
  assign n41519 = n32780 & ~n39531;
  assign n41520 = ~n41518 & ~n41519;
  assign n41521 = ~pi3467 & n39502;
  assign n41522 = n38277 & n38898;
  assign n41523 = n11155 & n41522;
  assign n41524 = ~n41521 & ~n41523;
  assign n41525 = n39504 & n41524;
  assign po1276 = ~n41520 | ~n41525;
  assign n41527 = ~pi2487 & pi3520;
  assign n41528 = pi3211 & ~n41527;
  assign n41529 = ~pi1331 & ~pi3291;
  assign n41530 = ~pi0759 & n41529;
  assign n41531 = ~pi0684 & pi2491;
  assign n41532 = pi3191 & n41531;
  assign n41533 = n41530 & n41532;
  assign n41534 = n41528 & n41533;
  assign n41535 = pi0684 & po3948;
  assign n41536 = ~pi2491 & ~n8670;
  assign n41537 = ~pi0759 & ~n41536;
  assign n41538 = pi3191 & n41537;
  assign n41539 = ~n9352 & ~n41538;
  assign n41540 = ~n41535 & ~n41539;
  assign n41541 = pi1015 & n8738;
  assign n41542 = pi1044 & n41541;
  assign n41543 = ~n41540 & ~n41542;
  assign n41544 = ~n41534 & n41543;
  assign n41545 = pi1015 & ~n41534;
  assign n41546 = ~pi3211 & ~n8670;
  assign n41547 = ~n41527 & ~n41546;
  assign n41548 = ~n16000 & n41547;
  assign n41549 = ~pi1331 & n41548;
  assign n41550 = ~n9352 & ~n41549;
  assign n41551 = n41545 & n41550;
  assign n41552 = ~n41544 & ~n41551;
  assign n41553 = ~pi0976 & ~n41552;
  assign n41554 = pi0976 & n41552;
  assign po1277 = n41553 | n41554;
  assign n41556 = ~n12726 & n41471;
  assign n41557 = pi0977 & n39393;
  assign po1278 = n41556 | n41557;
  assign n41559 = ~n14403 & n41471;
  assign n41560 = pi0978 & n39393;
  assign po1279 = n41559 | n41560;
  assign n41562 = ~pi1512 & n20345;
  assign n41563 = ~pi1531 & n20347;
  assign n41564 = ~n41562 & ~n41563;
  assign n41565 = ~pi1581 & n20350;
  assign n41566 = ~pi1465 & n20360;
  assign n41567 = ~pi1477 & n20363;
  assign n41568 = ~n41566 & ~n41567;
  assign n41569 = ~pi1392 & n20353;
  assign n41570 = ~pi1549 & n20356;
  assign n41571 = ~n41569 & ~n41570;
  assign n41572 = n41568 & n41571;
  assign n41573 = ~n41565 & n41572;
  assign n41574 = n41564 & n41573;
  assign n41575 = ~pi3120 & ~n41574;
  assign n41576 = pi3520 & pi3521;
  assign n41577 = pi0979 & ~pi3521;
  assign n41578 = ~n41576 & ~n41577;
  assign n41579 = pi3120 & ~n41578;
  assign n41580 = ~n41575 & ~n41579;
  assign n41581 = ~pi0866 & ~n41580;
  assign n41582 = pi0866 & ~n11181;
  assign po1282 = n41581 | n41582;
  assign n41584 = ~pi1506 & n20360;
  assign n41585 = ~pi1396 & n20363;
  assign n41586 = ~n41584 & ~n41585;
  assign n41587 = ~pi1576 & n20353;
  assign n41588 = ~pi1403 & n20356;
  assign n41589 = ~n41587 & ~n41588;
  assign n41590 = ~pi1525 & n20345;
  assign n41591 = ~pi1544 & n20347;
  assign n41592 = ~n41590 & ~n41591;
  assign n41593 = ~pi1592 & n20350;
  assign n41594 = n41592 & ~n41593;
  assign n41595 = n41589 & n41594;
  assign n41596 = n41586 & n41595;
  assign n41597 = ~pi1007 & ~n41596;
  assign n41598 = pi1007 & ~n11181;
  assign n41599 = ~n41597 & ~n41598;
  assign n41600 = ~n38527 & n41599;
  assign n41601 = ~pi0980 & n38527;
  assign n41602 = ~n41600 & ~n41601;
  assign po1283 = ~n38509 & n41602;
  assign n41604 = ~n39393 & n41443;
  assign n41605 = pi0981 & n39393;
  assign po1284 = n41604 | n41605;
  assign n41607 = n36095 & n39083;
  assign n41608 = n39844 & n41607;
  assign n41609 = ~pi0982 & n8561;
  assign n41610 = ~n41608 & ~n41609;
  assign po1285 = po3627 & ~n41610;
  assign n41612 = ~pi0983 & n8561;
  assign n41613 = ~n8561 & n36096;
  assign n41614 = ~n36077 & n36080;
  assign n41615 = n36083 & n41614;
  assign n41616 = n41613 & n41615;
  assign n41617 = n36102 & n41616;
  assign n41618 = ~n41612 & ~n41617;
  assign po1286 = po3627 & ~n41618;
  assign n41620 = ~pi0984 & n8561;
  assign n41621 = n39849 & n41616;
  assign n41622 = ~n41620 & ~n41621;
  assign po1287 = po3627 & ~n41622;
  assign n41624 = ~pi0985 & n8561;
  assign n41625 = n36120 & n39094;
  assign n41626 = n41375 & n41625;
  assign n41627 = ~n41624 & ~n41626;
  assign po1288 = po3627 & ~n41627;
  assign n41629 = ~pi0986 & n8561;
  assign n41630 = ~n8561 & n36070;
  assign n41631 = n36078 & n41630;
  assign n41632 = n41375 & n41631;
  assign n41633 = ~n41629 & ~n41632;
  assign po1289 = po3627 & ~n41633;
  assign n41635 = ~pi0987 & n8561;
  assign n41636 = ~n36083 & n41614;
  assign n41637 = n39084 & n41636;
  assign n41638 = ~n41635 & ~n41637;
  assign po1290 = po3627 & ~n41638;
  assign n41640 = ~pi0988 & n8561;
  assign n41641 = n36096 & n39083;
  assign n41642 = n41636 & n41641;
  assign n41643 = ~n41640 & ~n41642;
  assign po1291 = po3627 & ~n41643;
  assign n41645 = ~pi0989 & n8561;
  assign n41646 = n36094 & n38863;
  assign n41647 = n41636 & n41646;
  assign n41648 = ~n41645 & ~n41647;
  assign po1292 = po3627 & ~n41648;
  assign n41650 = ~pi0990 & n8561;
  assign n41651 = ~n36063 & n41082;
  assign n41652 = n36120 & n41651;
  assign n41653 = ~n41650 & ~n41652;
  assign po1293 = po3627 & ~n41653;
  assign n41655 = ~pi0991 & n8561;
  assign n41656 = n41376 & n41651;
  assign n41657 = ~n41655 & ~n41656;
  assign po1294 = po3627 & ~n41657;
  assign n41659 = pi0992 & n8561;
  assign n41660 = n39084 & n41615;
  assign n41661 = ~n41659 & ~n41660;
  assign po1295 = po3627 & ~n41661;
  assign n41663 = pi0993 & n8561;
  assign n41664 = n41615 & n41641;
  assign n41665 = ~n41663 & ~n41664;
  assign po1296 = po3627 & ~n41665;
  assign n41667 = pi0994 & n8561;
  assign n41668 = n41615 & n41646;
  assign n41669 = ~n41667 & ~n41668;
  assign po1297 = po3627 & ~n41669;
  assign n41671 = pi0995 & n8561;
  assign n41672 = ~n8561 & n36094;
  assign n41673 = n36096 & n41672;
  assign n41674 = n41615 & n41673;
  assign n41675 = ~n41671 & ~n41674;
  assign po1298 = po3627 & ~n41675;
  assign n41677 = pi0996 & n8561;
  assign n41678 = ~n36063 & n39093;
  assign n41679 = n41631 & n41678;
  assign n41680 = ~n41677 & ~n41679;
  assign po1299 = po3627 & ~n41680;
  assign n41682 = pi0997 & n8561;
  assign n41683 = n41625 & n41678;
  assign n41684 = ~n41682 & ~n41683;
  assign po1300 = po3627 & ~n41684;
  assign n41686 = pi0998 & n8561;
  assign n41687 = n39095 & n41083;
  assign n41688 = ~n41686 & ~n41687;
  assign po1301 = po3627 & ~n41688;
  assign n41690 = pi0999 & n8561;
  assign n41691 = n41377 & n41678;
  assign n41692 = ~n41690 & ~n41691;
  assign po1302 = po3627 & ~n41692;
  assign n41694 = ~n8561 & n36086;
  assign n41695 = ~pi1000 & n8561;
  assign n41696 = ~n41694 & ~n41695;
  assign po1303 = po3627 & ~n41696;
  assign n41698 = ~pi1001 & ~n36875;
  assign n41699 = pi0739 & pi1067;
  assign n41700 = ~pi0739 & ~pi1067;
  assign n41701 = ~n41699 & ~n41700;
  assign n41702 = pi0741 & pi0931;
  assign n41703 = ~pi0741 & ~pi0931;
  assign n41704 = ~n41702 & ~n41703;
  assign n41705 = pi0884 & pi1069;
  assign n41706 = ~pi0884 & ~pi1069;
  assign n41707 = ~n41705 & ~n41706;
  assign n41708 = pi0885 & pi1088;
  assign n41709 = ~pi0885 & ~pi1088;
  assign n41710 = ~n41708 & ~n41709;
  assign n41711 = n41707 & n41710;
  assign n41712 = n41704 & n41711;
  assign n41713 = n41701 & n41712;
  assign n41714 = ~pi0893 & pi1068;
  assign n41715 = pi0893 & ~pi1068;
  assign n41716 = ~n41714 & ~n41715;
  assign n41717 = n41713 & ~n41716;
  assign n41718 = pi1068 & n36792;
  assign n41719 = pi0890 & n41718;
  assign n41720 = ~n41717 & ~n41719;
  assign n41721 = ~n41698 & n41720;
  assign n41722 = pi0740 & n41721;
  assign n41723 = pi3647 & n41722;
  assign n41724 = ~pi1001 & n36875;
  assign po1304 = n41723 | n41724;
  assign n41726 = ~pi1002 & ~n36967;
  assign n41727 = pi0793 & pi1071;
  assign n41728 = ~pi0793 & ~pi1071;
  assign n41729 = ~n41727 & ~n41728;
  assign n41730 = pi0795 & pi0933;
  assign n41731 = ~pi0795 & ~pi0933;
  assign n41732 = ~n41730 & ~n41731;
  assign n41733 = pi0957 & pi1072;
  assign n41734 = ~pi0957 & ~pi1072;
  assign n41735 = ~n41733 & ~n41734;
  assign n41736 = pi1009 & pi1040;
  assign n41737 = ~pi1009 & ~pi1040;
  assign n41738 = ~n41736 & ~n41737;
  assign n41739 = n41735 & n41738;
  assign n41740 = n41732 & n41739;
  assign n41741 = n41729 & n41740;
  assign n41742 = ~pi0799 & pi1027;
  assign n41743 = pi0799 & ~pi1027;
  assign n41744 = ~n41742 & ~n41743;
  assign n41745 = n41741 & ~n41744;
  assign n41746 = pi1027 & n36885;
  assign n41747 = pi0796 & n41746;
  assign n41748 = ~n41745 & ~n41747;
  assign n41749 = ~n41726 & n41748;
  assign n41750 = pi0794 & n41749;
  assign n41751 = pi3635 & n41750;
  assign n41752 = ~pi1002 & n36967;
  assign po1305 = n41751 | n41752;
  assign po1306 = pi3086 & po0493;
  assign po1307 = pi3559 | ~po3853;
  assign n41756 = ~pi1003 & ~pi1673;
  assign n41757 = ~pi1604 & ~pi1672;
  assign n41758 = n41756 & n41757;
  assign n41759 = ~pi1645 & ~pi1670;
  assign n41760 = ~pi1675 & n41759;
  assign n41761 = ~pi1677 & ~pi1699;
  assign n41762 = ~pi1678 & ~pi1679;
  assign n41763 = n41761 & n41762;
  assign n41764 = n41760 & n41763;
  assign n41765 = ~pi1361 & ~pi1671;
  assign n41766 = ~pi1387 & ~pi1700;
  assign n41767 = n41765 & n41766;
  assign n41768 = ~pi1669 & ~pi1701;
  assign n41769 = ~pi1680 & ~pi1698;
  assign n41770 = n41768 & n41769;
  assign n41771 = ~pi1073 & ~pi1674;
  assign n41772 = n41770 & n41771;
  assign n41773 = ~pi1610 & n41772;
  assign n41774 = ~pi1074 & n41773;
  assign n41775 = n41767 & n41774;
  assign n41776 = n41764 & n41775;
  assign n41777 = ~pi1676 & n41776;
  assign n41778 = n41758 & n41777;
  assign n41779 = pi3641 & ~n41778;
  assign n41780 = ~pi1003 & ~n41779;
  assign n41781 = ~pi1676 & n41760;
  assign n41782 = n41763 & n41781;
  assign n41783 = n41770 & n41782;
  assign n41784 = n41767 & n41783;
  assign n41785 = pi1003 & n41784;
  assign n41786 = ~pi1003 & ~n41784;
  assign n41787 = ~n41785 & ~n41786;
  assign n41788 = n41779 & ~n41787;
  assign po1308 = n41780 | n41788;
  assign n41790 = ~pi1362 & ~pi1363;
  assign n41791 = ~pi1369 & ~pi1381;
  assign n41792 = n41790 & n41791;
  assign n41793 = ~pi1075 & ~pi1382;
  assign n41794 = ~pi1367 & n41793;
  assign n41795 = ~pi1384 & n41794;
  assign n41796 = ~pi1079 & ~pi1383;
  assign n41797 = ~pi1105 & ~pi1368;
  assign n41798 = n41796 & n41797;
  assign n41799 = n41795 & n41798;
  assign n41800 = n41792 & n41799;
  assign n41801 = ~pi1365 & ~pi1386;
  assign n41802 = ~pi1364 & ~pi1385;
  assign n41803 = n41801 & n41802;
  assign n41804 = n41800 & n41803;
  assign n41805 = pi1004 & n41804;
  assign n41806 = ~pi1004 & ~n41804;
  assign n41807 = ~n41805 & ~n41806;
  assign n41808 = po3946 & n41779;
  assign n41809 = ~pi3426 & n41808;
  assign n41810 = ~n41807 & n41809;
  assign n41811 = ~pi1004 & ~n41809;
  assign po1309 = n41810 | n41811;
  assign n41813 = ~pi1005 & ~n41809;
  assign n41814 = ~pi1004 & ~pi1366;
  assign n41815 = ~pi1076 & ~pi1077;
  assign n41816 = n41799 & n41815;
  assign n41817 = n41792 & n41816;
  assign n41818 = n41814 & n41817;
  assign n41819 = n41803 & n41818;
  assign n41820 = ~pi1005 & n41819;
  assign n41821 = pi1005 & ~n41819;
  assign n41822 = ~n41820 & ~n41821;
  assign n41823 = n41809 & n41822;
  assign po1310 = n41813 | n41823;
  assign n41825 = pi1908 & n41248;
  assign n41826 = pi1851 & pi3681;
  assign n41827 = ~pi1851 & ~pi3681;
  assign n41828 = ~n41826 & ~n41827;
  assign n41829 = ~n41239 & ~n41828;
  assign n41830 = ~n41242 & n41829;
  assign n41831 = n41825 & n41830;
  assign n41832 = pi1081 & pi1379;
  assign n41833 = pi1380 & pi1788;
  assign n41834 = pi1668 & pi1695;
  assign n41835 = pi2416 & n41834;
  assign n41836 = pi1851 & pi3247;
  assign n41837 = n41835 & n41836;
  assign n41838 = n41833 & n41837;
  assign n41839 = n41832 & n41838;
  assign n41840 = pi2824 & n41839;
  assign n41841 = pi2510 & pi3290;
  assign n41842 = n41840 & n41841;
  assign n41843 = ~pi1908 & ~n41842;
  assign n41844 = ~n41831 & ~n41843;
  assign n41845 = pi1006 & n41844;
  assign po1311 = ~pi3583 & ~n41845;
  assign n41847 = pi1007 & n36128;
  assign n41848 = n36060 & n36107;
  assign po1312 = n41847 | n41848;
  assign n41850 = n36063 & n41376;
  assign n41851 = n41082 & n41850;
  assign n41852 = ~pi1008 & n8561;
  assign n41853 = ~n41851 & ~n41852;
  assign po1313 = po3627 & ~n41853;
  assign n41855 = ~n15115 & n41431;
  assign n41856 = pi1009 & n39355;
  assign po1314 = n41855 | n41856;
  assign n41858 = n41636 & n41673;
  assign n41859 = ~pi1010 & n8561;
  assign n41860 = ~n41858 & ~n41859;
  assign po1315 = po3627 & ~n41860;
  assign n41862 = ~pi1011 & n8561;
  assign n41863 = n38863 & n41615;
  assign n41864 = n39849 & n41863;
  assign n41865 = ~n41862 & ~n41864;
  assign po1316 = po3627 & ~n41865;
  assign n41867 = ~n10759 & ~n10793;
  assign n41868 = ~n10752 & n41867;
  assign n41869 = n24810 & n41868;
  assign n41870 = ~n8561 & ~n41869;
  assign n41871 = pi1012 & ~n41870;
  assign n41872 = n12114 & n36392;
  assign n41873 = n11795 & ~n36392;
  assign n41874 = ~n41872 & ~n41873;
  assign n41875 = n36403 & ~n41874;
  assign n41876 = pi0413 & n10752;
  assign n41877 = ~n17784 & n36405;
  assign n41878 = ~n41876 & ~n41877;
  assign n41879 = n36392 & ~n41878;
  assign n41880 = ~n17809 & ~n36392;
  assign n41881 = ~n41879 & ~n41880;
  assign n41882 = ~n36403 & n41881;
  assign n41883 = ~n41875 & ~n41882;
  assign n41884 = n36418 & ~n41883;
  assign n41885 = n12061 & n36392;
  assign n41886 = n10608 & ~n36392;
  assign n41887 = ~n41885 & ~n41886;
  assign n41888 = n36403 & ~n41887;
  assign n41889 = n12106 & n36392;
  assign n41890 = n11781 & ~n36392;
  assign n41891 = ~n41889 & ~n41890;
  assign n41892 = ~n36403 & ~n41891;
  assign n41893 = ~n41888 & ~n41892;
  assign n41894 = ~n36418 & ~n41893;
  assign n41895 = ~n41884 & ~n41894;
  assign n41896 = n41870 & n41895;
  assign po1317 = n41871 | n41896;
  assign n41898 = pi1013 & ~n41870;
  assign n41899 = n37158 & n41870;
  assign po1318 = n41898 | n41899;
  assign n41901 = pi0976 & ~pi1014;
  assign n41902 = ~pi0976 & pi1014;
  assign n41903 = ~n41901 & ~n41902;
  assign n41904 = n41543 & ~n41903;
  assign n41905 = ~n15795 & ~n41543;
  assign n41906 = ~n41904 & ~n41905;
  assign n41907 = ~n41552 & ~n41906;
  assign n41908 = pi1014 & n41552;
  assign po1319 = n41907 | n41908;
  assign n41910 = pi1015 & n8745;
  assign n41911 = ~pi1015 & ~n8745;
  assign n41912 = ~n41910 & ~n41911;
  assign n41913 = n41543 & ~n41912;
  assign n41914 = ~pi1015 & n8743;
  assign n41915 = pi1015 & ~n8743;
  assign n41916 = ~n41914 & ~n41915;
  assign n41917 = ~n41543 & n41916;
  assign n41918 = ~n41913 & ~n41917;
  assign n41919 = ~n41552 & ~n41918;
  assign n41920 = ~pi1015 & n41552;
  assign po1320 = n41919 | n41920;
  assign n41922 = pi1016 & ~n41387;
  assign n41923 = ~pi1016 & n41387;
  assign n41924 = ~n41922 & ~n41923;
  assign po1321 = n40651 & n41924;
  assign n41926 = pi1017 & n39355;
  assign n41927 = ~n39355 & n40657;
  assign po1322 = n41926 | n41927;
  assign n41929 = pi1018 & ~n41493;
  assign n41930 = ~pi1018 & n41493;
  assign n41931 = ~n41929 & ~n41930;
  assign po1323 = n40741 & n41931;
  assign n41933 = ~pi3219 & ~n41503;
  assign n41934 = ~pi1762 & n41933;
  assign n41935 = ~pi1762 & ~n41503;
  assign n41936 = n10608 & n41511;
  assign n41937 = ~n41935 & ~n41936;
  assign n41938 = ~pi1019 & ~n41511;
  assign n41939 = n41937 & ~n41938;
  assign po1324 = n41934 | n41939;
  assign n41941 = pi1763 & pi1857;
  assign n41942 = ~pi0609 & n41941;
  assign n41943 = ~pi3241 & ~n41942;
  assign n41944 = ~pi1857 & n41943;
  assign n41945 = ~pi1857 & ~n41942;
  assign n41946 = n41510 & ~n41942;
  assign n41947 = ~pi1020 & ~n41946;
  assign n41948 = ~n41945 & ~n41947;
  assign n41949 = n13121 & n41946;
  assign n41950 = n41948 & ~n41949;
  assign po1325 = n41944 | n41950;
  assign n41952 = pi1764 & pi1765;
  assign n41953 = ~pi0609 & n41952;
  assign n41954 = ~pi3242 & ~n41953;
  assign n41955 = ~pi1764 & n41954;
  assign n41956 = ~pi1764 & ~n41953;
  assign n41957 = n41510 & ~n41953;
  assign n41958 = ~pi1021 & ~n41957;
  assign n41959 = ~n41956 & ~n41958;
  assign n41960 = n13988 & n41957;
  assign n41961 = n41959 & ~n41960;
  assign po1326 = n41955 | n41961;
  assign n41963 = pi1766 & pi1858;
  assign n41964 = ~pi0609 & n41963;
  assign n41965 = ~pi3218 & ~n41964;
  assign n41966 = ~pi1858 & n41965;
  assign n41967 = ~pi1858 & ~n41964;
  assign n41968 = n41510 & ~n41964;
  assign n41969 = ~pi1022 & ~n41968;
  assign n41970 = ~n41967 & ~n41969;
  assign n41971 = n14816 & n41968;
  assign n41972 = n41970 & ~n41971;
  assign po1327 = n41966 | n41972;
  assign n41974 = pi1767 & pi1769;
  assign n41975 = ~pi0609 & n41974;
  assign n41976 = ~pi3223 & ~n41975;
  assign n41977 = ~pi1767 & n41976;
  assign n41978 = ~pi1767 & ~n41975;
  assign n41979 = n41510 & ~n41975;
  assign n41980 = ~pi1023 & ~n41979;
  assign n41981 = ~n41978 & ~n41980;
  assign n41982 = n12061 & n41979;
  assign n41983 = n41981 & ~n41982;
  assign po1328 = n41977 | n41983;
  assign n41985 = pi1768 & pi1854;
  assign n41986 = ~pi0609 & n41985;
  assign n41987 = ~pi3224 & ~n41986;
  assign n41988 = ~pi1768 & n41987;
  assign n41989 = ~pi1768 & ~n41986;
  assign n41990 = n41510 & ~n41986;
  assign n41991 = ~pi1024 & ~n41990;
  assign n41992 = ~n41989 & ~n41991;
  assign n41993 = n17368 & n41990;
  assign n41994 = n41992 & ~n41993;
  assign po1329 = n41988 | n41994;
  assign n41996 = pi1025 & n9352;
  assign n41997 = ~pi1514 & n20345;
  assign n41998 = ~pi1407 & n20347;
  assign n41999 = ~n41997 & ~n41998;
  assign n42000 = ~pi1582 & n20350;
  assign n42001 = ~pi1567 & n20353;
  assign n42002 = ~pi1550 & n20356;
  assign n42003 = ~n42001 & ~n42002;
  assign n42004 = ~pi1496 & n20360;
  assign n42005 = ~pi1478 & n20363;
  assign n42006 = ~n42004 & ~n42005;
  assign n42007 = n42003 & n42006;
  assign n42008 = ~n42000 & n42007;
  assign n42009 = n41999 & n42008;
  assign n42010 = n19550 & ~n42009;
  assign n42011 = ~pi0835 & ~n13398;
  assign n42012 = ~n42010 & ~n42011;
  assign n42013 = ~n9352 & ~n42012;
  assign po1330 = n41996 | n42013;
  assign n42015 = ~pi0933 & ~pi1072;
  assign n42016 = ~pi1027 & ~pi1071;
  assign n42017 = ~pi1040 & n42016;
  assign n42018 = n42015 & n42017;
  assign n42019 = ~pi1026 & ~n42018;
  assign n42020 = pi1026 & n42018;
  assign n42021 = ~n42019 & ~n42020;
  assign n42022 = pi3635 & ~n42021;
  assign n42023 = ~pi1026 & ~pi3635;
  assign n42024 = ~n42022 & ~n42023;
  assign n42025 = n36969 & ~n42024;
  assign n42026 = pi0802 & n36968;
  assign po1331 = n42025 | n42026;
  assign n42028 = pi1027 & ~pi3635;
  assign n42029 = ~pi1027 & ~n36885;
  assign n42030 = ~n41746 & ~n42029;
  assign n42031 = pi3635 & n42030;
  assign n42032 = ~n42028 & ~n42031;
  assign n42033 = n36969 & n42032;
  assign n42034 = pi0850 & n36968;
  assign po1332 = n42033 | n42034;
  assign n42036 = pi1028 & ~n41870;
  assign n42037 = n37110 & n41870;
  assign po1333 = n42036 | n42037;
  assign n42039 = pi1029 & ~n41870;
  assign n42040 = n37183 & n41870;
  assign po1334 = n42039 | n42040;
  assign n42042 = pi1030 & ~n41870;
  assign n42043 = n37134 & n41870;
  assign po1335 = n42042 | n42043;
  assign n42045 = pi1031 & ~n41870;
  assign n42046 = n37207 & n41870;
  assign po1336 = n42045 | n42046;
  assign n42048 = pi1032 & ~n41870;
  assign n42049 = n12493 & n36392;
  assign n42050 = n12138 & ~n36392;
  assign n42051 = ~n42049 & ~n42050;
  assign n42052 = n36403 & ~n42051;
  assign n42053 = ~n17960 & n36405;
  assign n42054 = pi0410 & n10752;
  assign n42055 = ~n42053 & ~n42054;
  assign n42056 = n36392 & ~n42055;
  assign n42057 = ~n17983 & ~n36392;
  assign n42058 = ~n42056 & ~n42057;
  assign n42059 = ~n36403 & n42058;
  assign n42060 = ~n42052 & ~n42059;
  assign n42061 = n36418 & ~n42060;
  assign n42062 = n12415 & n36392;
  assign n42063 = n12726 & ~n36392;
  assign n42064 = ~n42062 & ~n42063;
  assign n42065 = n36403 & ~n42064;
  assign n42066 = n12485 & n36392;
  assign n42067 = n12751 & ~n36392;
  assign n42068 = ~n42066 & ~n42067;
  assign n42069 = ~n36403 & ~n42068;
  assign n42070 = ~n42065 & ~n42069;
  assign n42071 = ~n36418 & ~n42070;
  assign n42072 = ~n42061 & ~n42071;
  assign n42073 = n41870 & n42072;
  assign po1337 = n42048 | n42073;
  assign n42075 = pi1033 & ~n41870;
  assign n42076 = n14545 & n36392;
  assign n42077 = n14475 & ~n36392;
  assign n42078 = ~n42076 & ~n42077;
  assign n42079 = n36403 & ~n42078;
  assign n42080 = ~n17899 & n36405;
  assign n42081 = pi0411 & n10752;
  assign n42082 = ~n42080 & ~n42081;
  assign n42083 = n36392 & ~n42082;
  assign n42084 = ~n17927 & ~n36392;
  assign n42085 = ~n42083 & ~n42084;
  assign n42086 = ~n36403 & n42085;
  assign n42087 = ~n42079 & ~n42086;
  assign n42088 = n36418 & ~n42087;
  assign n42089 = n14816 & n36392;
  assign n42090 = n14403 & ~n36392;
  assign n42091 = ~n42089 & ~n42090;
  assign n42092 = n36403 & ~n42091;
  assign n42093 = n14537 & n36392;
  assign n42094 = n14430 & ~n36392;
  assign n42095 = ~n42093 & ~n42094;
  assign n42096 = ~n36403 & ~n42095;
  assign n42097 = ~n42092 & ~n42096;
  assign n42098 = ~n36418 & ~n42097;
  assign n42099 = ~n42088 & ~n42098;
  assign n42100 = n41870 & n42099;
  assign po1338 = n42075 | n42100;
  assign n42102 = pi1034 & ~n41870;
  assign n42103 = n15195 & n36392;
  assign n42104 = n14832 & ~n36392;
  assign n42105 = ~n42103 & ~n42104;
  assign n42106 = n36403 & ~n42105;
  assign n42107 = ~n17842 & n36405;
  assign n42108 = pi0412 & n10752;
  assign n42109 = ~n42107 & ~n42108;
  assign n42110 = n36392 & ~n42109;
  assign n42111 = ~n17866 & ~n36392;
  assign n42112 = ~n42110 & ~n42111;
  assign n42113 = ~n36403 & n42112;
  assign n42114 = ~n42106 & ~n42113;
  assign n42115 = n36418 & ~n42114;
  assign n42116 = n15115 & n36392;
  assign n42117 = n15426 & ~n36392;
  assign n42118 = ~n42116 & ~n42117;
  assign n42119 = n36403 & ~n42118;
  assign n42120 = n15187 & n36392;
  assign n42121 = n15454 & ~n36392;
  assign n42122 = ~n42120 & ~n42121;
  assign n42123 = ~n36403 & ~n42122;
  assign n42124 = ~n42119 & ~n42123;
  assign n42125 = ~n36418 & ~n42124;
  assign n42126 = ~n42115 & ~n42125;
  assign n42127 = n41870 & n42126;
  assign po1339 = n42102 | n42127;
  assign n42129 = pi1035 & ~n41870;
  assign n42130 = n36430 & n41870;
  assign po1340 = n42129 | n42130;
  assign n42132 = pi1036 & ~n41870;
  assign n42133 = n37085 & n41870;
  assign po1341 = n42132 | n42133;
  assign n42135 = pi1037 & ~n41870;
  assign n42136 = n37235 & n41870;
  assign po1342 = n42135 | n42136;
  assign n42138 = pi1038 & ~n41870;
  assign n42139 = n37061 & n41870;
  assign po1343 = n42138 | n42139;
  assign n42141 = pi1039 & ~n41870;
  assign n42142 = n11682 & n36392;
  assign n42143 = n11200 & ~n36392;
  assign n42144 = ~n42142 & ~n42143;
  assign n42145 = n36403 & ~n42144;
  assign n42146 = ~n17734 & n36405;
  assign n42147 = pi0408 & n10752;
  assign n42148 = ~n42146 & ~n42147;
  assign n42149 = n36392 & ~n42148;
  assign n42150 = ~n17751 & ~n36392;
  assign n42151 = ~n42149 & ~n42150;
  assign n42152 = ~n36403 & n42151;
  assign n42153 = ~n42145 & ~n42152;
  assign n42154 = n36418 & ~n42153;
  assign n42155 = n11181 & n36392;
  assign n42156 = n9825 & ~n36392;
  assign n42157 = ~n42155 & ~n42156;
  assign n42158 = n36403 & ~n42157;
  assign n42159 = n11674 & n36392;
  assign n42160 = n11752 & ~n36392;
  assign n42161 = ~n42159 & ~n42160;
  assign n42162 = ~n36403 & ~n42161;
  assign n42163 = ~n42158 & ~n42162;
  assign n42164 = ~n36418 & ~n42163;
  assign n42165 = ~n42154 & ~n42164;
  assign n42166 = n41870 & n42165;
  assign po1344 = n42141 | n42166;
  assign n42168 = pi1040 & n36883;
  assign n42169 = ~pi1040 & ~n36883;
  assign n42170 = ~n42168 & ~n42169;
  assign n42171 = pi3635 & ~n42170;
  assign n42172 = ~pi1040 & ~pi3635;
  assign n42173 = ~n42171 & ~n42172;
  assign n42174 = n36969 & ~n42173;
  assign n42175 = pi0846 & n36968;
  assign po1345 = n42174 | n42175;
  assign n42177 = pi3394 & n19544;
  assign n42178 = ~pi0684 & ~pi3210;
  assign n42179 = ~n42177 & n42178;
  assign n42180 = ~n19545 & n42179;
  assign n42181 = n19551 & ~n42180;
  assign n42182 = ~n9352 & n42177;
  assign n42183 = ~n41535 & ~n42182;
  assign n42184 = ~n20363 & ~n42183;
  assign n42185 = ~n42180 & n42184;
  assign n42186 = ~n42181 & ~n42185;
  assign n42187 = ~pi1041 & n42186;
  assign n42188 = ~pi1041 & ~n19548;
  assign n42189 = ~n20347 & ~n42188;
  assign n42190 = n42184 & n42189;
  assign n42191 = ~pi1041 & ~n20344;
  assign n42192 = ~n20350 & ~n42191;
  assign n42193 = ~n42184 & n42192;
  assign n42194 = ~n42190 & ~n42193;
  assign n42195 = ~n42186 & n42194;
  assign po1346 = n42187 | n42195;
  assign n42197 = ~pi1042 & n42186;
  assign n42198 = pi1042 & ~n42186;
  assign po1347 = n42197 | n42198;
  assign n42200 = ~n15800 & ~n41543;
  assign n42201 = ~pi1043 & ~n8712;
  assign n42202 = ~n8738 & ~n42201;
  assign n42203 = n41543 & n42202;
  assign n42204 = ~n42200 & ~n42203;
  assign n42205 = ~n41552 & ~n42204;
  assign n42206 = pi1043 & n41552;
  assign po1348 = n42205 | n42206;
  assign n42208 = ~n15798 & ~n41543;
  assign n42209 = ~pi1044 & ~n8738;
  assign n42210 = ~n8745 & ~n42209;
  assign n42211 = n41543 & n42210;
  assign n42212 = ~n42208 & ~n42211;
  assign n42213 = ~n41552 & ~n42212;
  assign n42214 = pi1044 & n41552;
  assign po1349 = n42213 | n42214;
  assign n42216 = ~pi1383 & n38779;
  assign n42217 = ~pi1677 & n38781;
  assign n42218 = ~n42216 & ~n42217;
  assign n42219 = pi0408 & n38789;
  assign n42220 = n42218 & ~n42219;
  assign n42221 = pi0387 & n38792;
  assign n42222 = n42220 & ~n42221;
  assign n42223 = n38798 & ~n42222;
  assign n42224 = ~pi1082 & n38800;
  assign n42225 = ~pi0937 & ~n38800;
  assign n42226 = ~n42224 & ~n42225;
  assign n42227 = ~n38798 & ~n42226;
  assign n42228 = ~n42223 & ~n42227;
  assign n42229 = ~n38745 & ~n42228;
  assign n42230 = ~pi1045 & n38745;
  assign po1350 = n42229 | n42230;
  assign n42232 = ~pi0939 & pi3484;
  assign n42233 = pi3571 & n42232;
  assign po1351 = ~n38259 & n42233;
  assign n42235 = n41540 & ~n41550;
  assign n42236 = ~pi0976 & pi1015;
  assign n42237 = n41550 & n42236;
  assign n42238 = ~pi1014 & n42237;
  assign n42239 = ~pi1044 & n42238;
  assign n42240 = ~pi1043 & n42239;
  assign n42241 = ~pi1015 & n41550;
  assign n42242 = ~n42240 & ~n42241;
  assign n42243 = ~n42235 & ~n42242;
  assign n42244 = pi1047 & n42235;
  assign po1352 = n42243 | n42244;
  assign n42246 = ~n38246 & ~n38248;
  assign n42247 = n38244 & ~n38253;
  assign n42248 = ~n38250 & ~n38252;
  assign n42249 = n42247 & n42248;
  assign n42250 = n38262 & n42249;
  assign n42251 = n38227 & n42250;
  assign n42252 = n42246 & n42251;
  assign n42253 = pi1048 & ~n38262;
  assign po1353 = n42252 | n42253;
  assign n42255 = ~n38248 & ~n38250;
  assign n42256 = ~n38240 & n42255;
  assign n42257 = ~n38227 & n38235;
  assign n42258 = n38254 & n42257;
  assign n42259 = n42256 & n42258;
  assign n42260 = ~n38246 & n42259;
  assign n42261 = n38262 & n42260;
  assign n42262 = ~n38238 & n42261;
  assign n42263 = ~n38242 & n42262;
  assign n42264 = pi1049 & ~n38262;
  assign po1354 = n42263 | n42264;
  assign n42266 = ~pi1050 & n8561;
  assign n42267 = n36102 & n41863;
  assign n42268 = ~n42266 & ~n42267;
  assign po1355 = po3627 & ~n42268;
  assign n42270 = ~pi1051 & n8561;
  assign n42271 = ~n36063 & n36085;
  assign n42272 = n41630 & n42271;
  assign n42273 = ~n42270 & ~n42272;
  assign po1356 = po3627 & ~n42273;
  assign n42275 = ~pi0407 & n38789;
  assign n42276 = ~pi1382 & n38779;
  assign n42277 = ~pi1645 & n38781;
  assign n42278 = ~n42276 & ~n42277;
  assign n42279 = ~n42275 & n42278;
  assign n42280 = pi0390 & n38792;
  assign n42281 = n42279 & ~n42280;
  assign n42282 = n38798 & ~n42281;
  assign n42283 = ~pi0911 & n38800;
  assign n42284 = ~pi1080 & ~n38800;
  assign n42285 = ~n42283 & ~n42284;
  assign n42286 = ~n38798 & ~n42285;
  assign n42287 = ~n42282 & ~n42286;
  assign n42288 = ~n38745 & ~n42287;
  assign n42289 = ~pi1052 & n38745;
  assign po1357 = n42288 | n42289;
  assign n42291 = ~n8561 & n37725;
  assign n42292 = pi1053 & n8561;
  assign po1358 = n42291 | n42292;
  assign n42294 = pi1054 & n8561;
  assign n42295 = ~n8561 & n36021;
  assign po1359 = n42294 | n42295;
  assign n42297 = pi1055 & n8561;
  assign n42298 = ~n8561 & n36023;
  assign po1360 = n42297 | n42298;
  assign n42300 = pi1056 & n8561;
  assign n42301 = ~n8561 & n36042;
  assign po1361 = n42300 | n42301;
  assign n42303 = ~n8561 & n37736;
  assign n42304 = pi1057 & n8561;
  assign po1362 = n42303 | n42304;
  assign n42306 = ~n8561 & n37746;
  assign n42307 = pi1058 & n8561;
  assign po1363 = n42306 | n42307;
  assign n42309 = ~n8561 & n37726;
  assign n42310 = pi1059 & n8561;
  assign po1364 = n42309 | n42310;
  assign n42312 = pi1060 & ~n39903;
  assign n42313 = ~n39891 & ~n42312;
  assign n42314 = ~pi3684 & n39891;
  assign n42315 = ~n42313 & ~n42314;
  assign n42316 = ~n39893 & n42315;
  assign n42317 = pi1060 & n39893;
  assign po1365 = n42316 | n42317;
  assign n42319 = pi1061 & ~n39903;
  assign n42320 = ~n39891 & ~n42319;
  assign n42321 = ~pi3690 & n39891;
  assign n42322 = ~n42320 & ~n42321;
  assign n42323 = ~n39893 & n42322;
  assign n42324 = pi1061 & n39893;
  assign po1366 = n42323 | n42324;
  assign n42326 = pi1062 & ~n39903;
  assign n42327 = ~n39891 & ~n42326;
  assign n42328 = ~pi3689 & n39891;
  assign n42329 = ~n42327 & ~n42328;
  assign n42330 = ~n39893 & n42329;
  assign n42331 = pi1062 & n39893;
  assign po1367 = n42330 | n42331;
  assign n42333 = pi1063 & ~n39903;
  assign n42334 = ~n39891 & ~n42333;
  assign n42335 = ~pi3688 & n39891;
  assign n42336 = ~n42334 & ~n42335;
  assign n42337 = ~n39893 & n42336;
  assign n42338 = pi1063 & n39893;
  assign po1368 = n42337 | n42338;
  assign n42340 = pi1064 & ~n39903;
  assign n42341 = ~n39891 & ~n42340;
  assign n42342 = ~pi3687 & n39891;
  assign n42343 = ~n42341 & ~n42342;
  assign n42344 = ~n39893 & n42343;
  assign n42345 = pi1064 & n39893;
  assign po1369 = n42344 | n42345;
  assign n42347 = pi1065 & ~n39903;
  assign n42348 = ~n39891 & ~n42347;
  assign n42349 = ~pi3686 & n39891;
  assign n42350 = ~n42348 & ~n42349;
  assign n42351 = ~n39893 & n42350;
  assign n42352 = pi1065 & n39893;
  assign po1370 = n42351 | n42352;
  assign n42354 = ~n12726 & n38320;
  assign n42355 = n41161 & n41167;
  assign n42356 = ~pi1066 & ~n42355;
  assign n42357 = pi1066 & n42355;
  assign n42358 = ~n42356 & ~n42357;
  assign n42359 = ~n36181 & ~n42358;
  assign n42360 = ~pi1066 & n36181;
  assign n42361 = ~n42359 & ~n42360;
  assign n42362 = ~n38320 & n42361;
  assign po1371 = n42354 | n42362;
  assign n42364 = ~pi0931 & pi1067;
  assign n42365 = pi0931 & ~pi1067;
  assign n42366 = ~n42364 & ~n42365;
  assign n42367 = pi3647 & ~n42366;
  assign n42368 = ~pi1067 & ~pi3647;
  assign n42369 = ~n42367 & ~n42368;
  assign n42370 = n36877 & ~n42369;
  assign n42371 = pi0747 & n36876;
  assign po1372 = n42370 | n42371;
  assign n42373 = pi1068 & ~pi3647;
  assign n42374 = ~pi1068 & ~n36792;
  assign n42375 = ~n41718 & ~n42374;
  assign n42376 = pi3647 & n42375;
  assign n42377 = ~n42373 & ~n42376;
  assign n42378 = n36877 & n42377;
  assign n42379 = pi0745 & n36876;
  assign po1373 = n42378 | n42379;
  assign n42381 = pi1069 & n36791;
  assign n42382 = ~pi1069 & ~n36791;
  assign n42383 = ~n42381 & ~n42382;
  assign n42384 = pi3647 & ~n42383;
  assign n42385 = ~pi1069 & ~pi3647;
  assign n42386 = ~n42384 & ~n42385;
  assign n42387 = n36877 & ~n42386;
  assign n42388 = pi0746 & n36876;
  assign po1374 = n42387 | n42388;
  assign n42390 = ~pi0848 & n36882;
  assign n42391 = ~pi0935 & n42390;
  assign n42392 = n42018 & n42391;
  assign n42393 = n36892 & n42392;
  assign n42394 = ~pi0690 & n42393;
  assign n42395 = ~pi1091 & n42394;
  assign n42396 = ~pi1070 & ~n42395;
  assign n42397 = pi1070 & n42395;
  assign n42398 = ~n42396 & ~n42397;
  assign n42399 = pi3635 & ~n42398;
  assign n42400 = ~pi1070 & ~pi3635;
  assign n42401 = ~n42399 & ~n42400;
  assign n42402 = n36969 & ~n42401;
  assign n42403 = pi0981 & n36968;
  assign po1375 = n42402 | n42403;
  assign n42405 = pi0933 & ~pi1071;
  assign n42406 = ~pi0933 & pi1071;
  assign n42407 = ~n42405 & ~n42406;
  assign n42408 = pi3635 & ~n42407;
  assign n42409 = ~pi1071 & ~pi3635;
  assign n42410 = ~n42408 & ~n42409;
  assign n42411 = n36969 & ~n42410;
  assign n42412 = pi0804 & n36968;
  assign po1376 = n42411 | n42412;
  assign n42414 = pi1072 & n36884;
  assign n42415 = ~pi1072 & ~n36884;
  assign n42416 = ~n42414 & ~n42415;
  assign n42417 = pi3635 & ~n42416;
  assign n42418 = ~pi1072 & ~pi3635;
  assign n42419 = ~n42417 & ~n42418;
  assign n42420 = n36969 & ~n42419;
  assign n42421 = pi0803 & n36968;
  assign po1377 = n42420 | n42421;
  assign n42423 = ~pi1073 & ~n41779;
  assign n42424 = n41770 & n41781;
  assign n42425 = n41767 & n42424;
  assign n42426 = n41763 & n42425;
  assign n42427 = n41758 & n42426;
  assign n42428 = ~pi1073 & ~n42427;
  assign n42429 = pi1073 & n42427;
  assign n42430 = ~n42428 & ~n42429;
  assign n42431 = n41779 & ~n42430;
  assign po1378 = n42423 | n42431;
  assign n42433 = ~pi1074 & ~n41779;
  assign n42434 = ~pi1073 & ~pi1604;
  assign n42435 = ~pi1671 & ~pi1700;
  assign n42436 = ~pi1361 & n42435;
  assign n42437 = ~pi1701 & n42436;
  assign n42438 = ~pi1679 & n41769;
  assign n42439 = ~pi1669 & n42438;
  assign n42440 = n42437 & n42439;
  assign n42441 = ~pi1003 & ~pi1387;
  assign n42442 = ~pi1672 & ~pi1673;
  assign n42443 = n42441 & n42442;
  assign n42444 = n42440 & n42443;
  assign n42445 = n42434 & n42444;
  assign n42446 = ~pi1678 & ~pi1699;
  assign n42447 = ~pi1676 & ~pi1677;
  assign n42448 = n41760 & n42447;
  assign n42449 = n42446 & n42448;
  assign n42450 = ~pi1610 & n42449;
  assign n42451 = ~pi1674 & n42450;
  assign n42452 = n42445 & n42451;
  assign n42453 = pi1074 & n42452;
  assign n42454 = ~pi1074 & ~n42452;
  assign n42455 = ~n42453 & ~n42454;
  assign n42456 = n41779 & ~n42455;
  assign po1379 = n42433 | n42456;
  assign n42458 = ~pi1075 & ~n41809;
  assign n42459 = pi1075 & n41809;
  assign po1380 = n42458 | n42459;
  assign n42461 = ~pi1076 & ~n41809;
  assign n42462 = n41802 & n41814;
  assign n42463 = ~pi1367 & ~pi1384;
  assign n42464 = n41796 & n42463;
  assign n42465 = n41791 & n41797;
  assign n42466 = n41790 & n41801;
  assign n42467 = n42465 & n42466;
  assign n42468 = n42464 & n42467;
  assign n42469 = n41793 & n42468;
  assign n42470 = n42462 & n42469;
  assign n42471 = ~pi1076 & n42470;
  assign n42472 = pi1076 & ~n42470;
  assign n42473 = ~n42471 & ~n42472;
  assign n42474 = n41809 & n42473;
  assign po1381 = n42461 | n42474;
  assign n42476 = ~pi1077 & ~n41809;
  assign n42477 = ~pi1004 & ~pi1385;
  assign n42478 = ~pi1076 & ~pi1366;
  assign n42479 = n42477 & n42478;
  assign n42480 = ~pi1079 & ~pi1368;
  assign n42481 = ~pi1383 & ~pi1384;
  assign n42482 = n41794 & n42481;
  assign n42483 = n42480 & n42482;
  assign n42484 = ~pi1364 & ~pi1365;
  assign n42485 = ~pi1386 & n42484;
  assign n42486 = ~pi1363 & n42485;
  assign n42487 = ~pi1105 & n41791;
  assign n42488 = ~pi1362 & n42487;
  assign n42489 = n42486 & n42488;
  assign n42490 = n42483 & n42489;
  assign n42491 = n42479 & n42490;
  assign n42492 = ~pi1077 & n42491;
  assign n42493 = pi1077 & ~n42491;
  assign n42494 = ~n42492 & ~n42493;
  assign n42495 = n41809 & n42494;
  assign po1382 = n42476 | n42495;
  assign n42497 = ~pi1078 & ~n41809;
  assign n42498 = n41815 & n42462;
  assign n42499 = n42467 & n42498;
  assign n42500 = n41793 & n42464;
  assign n42501 = n42499 & n42500;
  assign n42502 = ~pi1005 & n42501;
  assign n42503 = ~pi1086 & n42502;
  assign n42504 = ~pi1078 & n42503;
  assign n42505 = pi1078 & ~n42503;
  assign n42506 = ~n42504 & ~n42505;
  assign n42507 = n41809 & n42506;
  assign po1383 = n42497 | n42507;
  assign n42509 = ~pi1079 & ~n41809;
  assign n42510 = ~pi1075 & n42481;
  assign n42511 = ~pi1382 & n42510;
  assign n42512 = ~pi1367 & n42511;
  assign n42513 = ~pi1079 & n42512;
  assign n42514 = pi1079 & ~n42512;
  assign n42515 = ~n42513 & ~n42514;
  assign n42516 = n41809 & n42515;
  assign po1384 = n42509 | n42516;
  assign n42518 = ~pi1367 & n38779;
  assign n42519 = ~pi1675 & n38781;
  assign n42520 = ~n42518 & ~n42519;
  assign n42521 = pi0415 & n38789;
  assign n42522 = n42520 & ~n42521;
  assign n42523 = pi0389 & n38792;
  assign n42524 = n42522 & ~n42523;
  assign n42525 = n38798 & ~n42524;
  assign n42526 = ~pi1052 & n38800;
  assign n42527 = ~pi1082 & ~n38800;
  assign n42528 = ~n42526 & ~n42527;
  assign n42529 = ~n38798 & ~n42528;
  assign n42530 = ~n42525 & ~n42529;
  assign n42531 = ~n38745 & ~n42530;
  assign n42532 = ~pi1080 & n38745;
  assign po1385 = n42531 | n42532;
  assign po1386 = ~pi3583 & po1234;
  assign n42535 = ~pi2492 & pi3397;
  assign n42536 = pi3481 & n42535;
  assign n42537 = ~pi1081 & ~n42536;
  assign n42538 = ~pi1695 & ~pi2416;
  assign n42539 = ~pi1851 & n42538;
  assign n42540 = n41248 & n42539;
  assign n42541 = ~pi1380 & ~pi1788;
  assign n42542 = n42540 & n42541;
  assign n42543 = ~pi1668 & n42542;
  assign n42544 = ~pi1379 & n42543;
  assign n42545 = ~pi1081 & ~n42544;
  assign n42546 = pi1081 & n42544;
  assign n42547 = ~n42545 & ~n42546;
  assign n42548 = n42536 & ~n42547;
  assign po1387 = n42537 | n42548;
  assign n42550 = ~pi1384 & n38779;
  assign n42551 = ~pi1676 & n38781;
  assign n42552 = ~n42550 & ~n42551;
  assign n42553 = pi0414 & n38789;
  assign n42554 = n42552 & ~n42553;
  assign n42555 = pi0388 & n38792;
  assign n42556 = n42554 & ~n42555;
  assign n42557 = n38798 & ~n42556;
  assign n42558 = ~pi1080 & n38800;
  assign n42559 = ~pi1045 & ~n38800;
  assign n42560 = ~n42558 & ~n42559;
  assign n42561 = ~n38798 & ~n42560;
  assign n42562 = ~n42557 & ~n42561;
  assign n42563 = ~n38745 & ~n42562;
  assign n42564 = ~pi1082 & n38745;
  assign po1388 = n42563 | n42564;
  assign n42566 = ~pi1069 & ~pi1088;
  assign n42567 = ~pi0931 & ~pi1068;
  assign n42568 = ~pi1067 & n42567;
  assign n42569 = n42566 & n42568;
  assign n42570 = ~pi1083 & ~n42569;
  assign n42571 = pi1083 & n42569;
  assign n42572 = ~n42570 & ~n42571;
  assign n42573 = pi3647 & ~n42572;
  assign n42574 = ~pi1083 & ~pi3647;
  assign n42575 = ~n42573 & ~n42574;
  assign n42576 = n36877 & ~n42575;
  assign n42577 = pi0744 & n36876;
  assign po1389 = n42576 | n42577;
  assign n42579 = ~pi1084 & ~n41809;
  assign n42580 = ~pi1005 & ~pi1077;
  assign n42581 = ~pi1078 & ~pi1086;
  assign n42582 = n42483 & n42581;
  assign n42583 = n42489 & n42582;
  assign n42584 = n42580 & n42583;
  assign n42585 = n42479 & n42584;
  assign n42586 = ~pi1084 & n42585;
  assign n42587 = pi1084 & ~n42585;
  assign n42588 = ~n42586 & ~n42587;
  assign n42589 = n41809 & n42588;
  assign po1390 = n42579 | n42589;
  assign n42591 = ~pi0847 & n36794;
  assign n42592 = ~pi0940 & n42591;
  assign n42593 = n42569 & n42592;
  assign n42594 = ~pi1085 & ~n42593;
  assign n42595 = pi1085 & n42593;
  assign n42596 = ~n42594 & ~n42595;
  assign n42597 = pi3647 & ~n42596;
  assign n42598 = ~pi1085 & ~pi3647;
  assign n42599 = ~n42597 & ~n42598;
  assign n42600 = n36877 & ~n42599;
  assign n42601 = pi0869 & n36876;
  assign po1391 = n42600 | n42601;
  assign n42603 = ~pi1086 & ~n41809;
  assign n42604 = ~pi1369 & n42480;
  assign n42605 = ~pi1105 & n42604;
  assign n42606 = ~pi1381 & ~pi1386;
  assign n42607 = n41790 & n42606;
  assign n42608 = n42605 & n42607;
  assign n42609 = n42477 & n42608;
  assign n42610 = n42484 & n42609;
  assign n42611 = n42512 & n42580;
  assign n42612 = n42610 & n42611;
  assign n42613 = n42478 & n42612;
  assign n42614 = ~pi1086 & n42613;
  assign n42615 = pi1086 & ~n42613;
  assign n42616 = ~n42614 & ~n42615;
  assign n42617 = n41809 & n42616;
  assign po1392 = n42603 | n42617;
  assign n42619 = n36800 & n42593;
  assign n42620 = ~pi0689 & n42619;
  assign n42621 = ~pi1085 & n42620;
  assign n42622 = ~pi1087 & ~n42621;
  assign n42623 = pi1087 & n42621;
  assign n42624 = ~n42622 & ~n42623;
  assign n42625 = pi3647 & ~n42624;
  assign n42626 = ~pi1087 & ~pi3647;
  assign n42627 = ~n42625 & ~n42626;
  assign n42628 = n36877 & ~n42627;
  assign n42629 = pi0870 & n36876;
  assign po1393 = n42628 | n42629;
  assign n42631 = pi1088 & n36790;
  assign n42632 = ~pi1088 & ~n36790;
  assign n42633 = ~n42631 & ~n42632;
  assign n42634 = pi3647 & ~n42633;
  assign n42635 = ~pi1088 & ~pi3647;
  assign n42636 = ~n42634 & ~n42635;
  assign n42637 = n36877 & ~n42636;
  assign n42638 = pi0737 & n36876;
  assign po1394 = n42637 | n42638;
  assign n42640 = pi1089 & ~n39903;
  assign n42641 = ~n39891 & ~n42640;
  assign n42642 = ~pi3685 & n39891;
  assign n42643 = ~n42641 & ~n42642;
  assign n42644 = ~n39893 & n42643;
  assign n42645 = pi1089 & n39893;
  assign po1395 = n42644 | n42645;
  assign n42647 = ~n14403 & n38320;
  assign n42648 = n38308 & n38311;
  assign n42649 = n38300 & n38307;
  assign n42650 = n42648 & n42649;
  assign n42651 = ~pi1090 & ~n42650;
  assign n42652 = pi1090 & n42650;
  assign n42653 = ~n42651 & ~n42652;
  assign n42654 = ~n36181 & ~n42653;
  assign n42655 = ~pi1090 & n36181;
  assign n42656 = ~n42654 & ~n42655;
  assign n42657 = ~n38320 & n42656;
  assign po1396 = n42647 | n42657;
  assign n42659 = ~pi1091 & ~n42392;
  assign n42660 = pi1091 & n42392;
  assign n42661 = ~n42659 & ~n42660;
  assign n42662 = pi3635 & ~n42661;
  assign n42663 = ~pi1091 & ~pi3635;
  assign n42664 = ~n42662 & ~n42663;
  assign n42665 = n36969 & ~n42664;
  assign n42666 = pi0977 & n36968;
  assign po1397 = n42665 | n42666;
  assign n42668 = pi1092 & ~n39903;
  assign n42669 = ~n39891 & ~n42668;
  assign n42670 = ~pi3683 & n39891;
  assign n42671 = ~n42669 & ~n42670;
  assign n42672 = ~n39893 & n42671;
  assign n42673 = pi1092 & n39893;
  assign po1398 = n42672 | n42673;
  assign n42675 = ~n20352 & ~n20362;
  assign n42676 = n42184 & n42675;
  assign n42677 = ~n19548 & ~n20344;
  assign n42678 = ~n42184 & n42677;
  assign n42679 = ~n42676 & ~n42678;
  assign n42680 = ~n42186 & n42679;
  assign n42681 = ~pi1093 & n42186;
  assign po1399 = n42680 | n42681;
  assign n42683 = ~pi1094 & n40580;
  assign n42684 = pi1094 & ~n40580;
  assign n42685 = ~n42683 & ~n42684;
  assign po1400 = n40651 & n42685;
  assign n42687 = ~pi1095 & n40670;
  assign n42688 = pi1095 & ~n40670;
  assign n42689 = ~n42687 & ~n42688;
  assign po1401 = n40741 & n42689;
  assign n42691 = n41383 & n41386;
  assign n42692 = n41388 & n42691;
  assign n42693 = n41384 & n42692;
  assign n42694 = ~pi1097 & n42693;
  assign n42695 = pi1097 & ~n42693;
  assign n42696 = ~n42694 & ~n42695;
  assign po1403 = n40651 & n42696;
  assign n42698 = n41489 & n41492;
  assign n42699 = n41494 & n42698;
  assign n42700 = n41490 & n42699;
  assign n42701 = ~pi1098 & n42700;
  assign n42702 = pi1098 & ~n42700;
  assign n42703 = ~n42701 & ~n42702;
  assign po1404 = n40741 & n42703;
  assign n42705 = ~pi1763 & ~pi3220;
  assign n42706 = ~n41942 & n42705;
  assign n42707 = ~pi1099 & ~n41946;
  assign n42708 = n13398 & n41946;
  assign n42709 = ~pi1763 & ~n41942;
  assign n42710 = ~n42708 & ~n42709;
  assign n42711 = ~n42707 & n42710;
  assign po1405 = n42706 | n42711;
  assign n42713 = ~pi1765 & ~pi3221;
  assign n42714 = ~n41953 & n42713;
  assign n42715 = ~pi1100 & ~n41957;
  assign n42716 = n12415 & n41957;
  assign n42717 = ~pi1765 & ~n41953;
  assign n42718 = ~n42716 & ~n42717;
  assign n42719 = ~n42715 & n42718;
  assign po1406 = n42714 | n42719;
  assign n42721 = ~pi1766 & ~pi3222;
  assign n42722 = ~n41964 & n42721;
  assign n42723 = ~pi1101 & ~n41968;
  assign n42724 = n15115 & n41968;
  assign n42725 = ~pi1766 & ~n41964;
  assign n42726 = ~n42724 & ~n42725;
  assign n42727 = ~n42723 & n42726;
  assign po1407 = n42722 | n42727;
  assign n42729 = ~pi1854 & ~pi3240;
  assign n42730 = ~n41986 & n42729;
  assign n42731 = ~pi1102 & ~n41990;
  assign n42732 = n17199 & n41990;
  assign n42733 = ~pi1854 & ~n41986;
  assign n42734 = ~n42732 & ~n42733;
  assign n42735 = ~n42731 & n42734;
  assign po1408 = n42730 | n42735;
  assign n42737 = ~pi1769 & ~pi3225;
  assign n42738 = ~n41975 & n42737;
  assign n42739 = ~pi1103 & ~n41979;
  assign n42740 = n11181 & n41979;
  assign n42741 = ~pi1769 & ~n41975;
  assign n42742 = ~n42740 & ~n42741;
  assign n42743 = ~n42739 & n42742;
  assign po1409 = n42738 | n42743;
  assign n42745 = ~pi1104 & pi1373;
  assign n42746 = pi1104 & ~pi1373;
  assign n42747 = ~n42745 & ~n42746;
  assign n42748 = pi2508 & ~pi2992;
  assign n42749 = ~pi3588 & n42748;
  assign n42750 = ~pi2508 & ~pi2992;
  assign n42751 = pi3588 & n42750;
  assign n42752 = ~pi2508 & pi2992;
  assign n42753 = ~pi3588 & n42752;
  assign n42754 = ~n42751 & ~n42753;
  assign n42755 = ~n42749 & n42754;
  assign n42756 = pi0738 & po0038;
  assign n42757 = ~pi0738 & pi3671;
  assign n42758 = ~n42756 & ~n42757;
  assign n42759 = ~pi0880 & ~n42758;
  assign n42760 = pi0880 & n42758;
  assign po3950 = n42759 | n42760;
  assign n42762 = pi3646 & po3950;
  assign po3945 = pi3647 & n42762;
  assign n42764 = n34849 & ~po3945;
  assign n42765 = ~pi3640 & n34859;
  assign n42766 = pi3637 & n34861;
  assign n42767 = pi3634 & ~n34861;
  assign n42768 = ~n42766 & ~n42767;
  assign n42769 = ~n34859 & n42768;
  assign n42770 = ~n42765 & ~n42769;
  assign n42771 = ~n34849 & ~n42770;
  assign n42772 = ~n42764 & ~n42771;
  assign n42773 = n42749 & ~n42772;
  assign n42774 = ~n42755 & ~n42773;
  assign n42775 = ~pi1104 & ~pi1372;
  assign n42776 = ~pi1388 & n42775;
  assign n42777 = ~pi1371 & n42776;
  assign n42778 = ~pi1373 & n42777;
  assign n42779 = n42751 & n42778;
  assign n42780 = ~pi1684 & ~pi1702;
  assign n42781 = ~pi1846 & ~pi1847;
  assign n42782 = pi1607 & pi1703;
  assign n42783 = pi1683 & n42782;
  assign n42784 = pi1682 & n42783;
  assign n42785 = n42781 & n42784;
  assign n42786 = n42780 & n42785;
  assign n42787 = n42779 & n42786;
  assign po2823 = ~n42774 | n42787;
  assign po3310 = n42779 & ~n42786;
  assign n42790 = ~po2823 & ~po3310;
  assign n42791 = ~n42747 & n42790;
  assign n42792 = ~pi0739 & ~n42790;
  assign n42793 = ~n42791 & ~n42792;
  assign po1410 = ~pi1685 | n42793;
  assign n42795 = pi1105 & n42483;
  assign n42796 = ~pi1105 & ~n42483;
  assign n42797 = ~n42795 & ~n42796;
  assign n42798 = n41809 & ~n42797;
  assign n42799 = ~pi1105 & ~n41809;
  assign po1411 = n42798 | n42799;
  assign n42801 = ~pi0976 & n42210;
  assign n42802 = n41903 & ~n42202;
  assign n42803 = n42801 & n42802;
  assign n42804 = ~pi0759 & ~n18968;
  assign n42805 = pi0759 & ~n12726;
  assign n42806 = ~n42804 & ~n42805;
  assign n42807 = ~pi0684 & ~n42806;
  assign n42808 = pi0684 & pi3420;
  assign n42809 = ~n42807 & ~n42808;
  assign n42810 = n42803 & ~n42809;
  assign n42811 = pi1106 & ~n42803;
  assign n42812 = ~n42810 & ~n42811;
  assign n42813 = n41544 & ~n42812;
  assign n42814 = pi1106 & ~n41544;
  assign po1412 = n42813 | n42814;
  assign n42816 = ~pi0759 & n18900;
  assign n42817 = pi0759 & ~n13701;
  assign n42818 = ~n42816 & ~n42817;
  assign n42819 = ~pi0684 & ~n42818;
  assign n42820 = pi0684 & pi3411;
  assign n42821 = ~n42819 & ~n42820;
  assign n42822 = n42803 & ~n42821;
  assign n42823 = pi1107 & ~n42803;
  assign n42824 = ~n42822 & ~n42823;
  assign n42825 = n41544 & ~n42824;
  assign n42826 = pi1107 & ~n41544;
  assign po1413 = n42825 | n42826;
  assign n42828 = ~pi0759 & n18829;
  assign n42829 = pi0759 & ~n13121;
  assign n42830 = ~n42828 & ~n42829;
  assign n42831 = ~pi0684 & ~n42830;
  assign n42832 = pi0684 & pi3406;
  assign n42833 = ~n42831 & ~n42832;
  assign n42834 = n42803 & ~n42833;
  assign n42835 = pi1108 & ~n42803;
  assign n42836 = ~n42834 & ~n42835;
  assign n42837 = n41544 & ~n42836;
  assign n42838 = pi1108 & ~n41544;
  assign po1414 = n42837 | n42838;
  assign n42840 = ~pi0759 & n18755;
  assign n42841 = pi0759 & ~n13398;
  assign n42842 = ~n42840 & ~n42841;
  assign n42843 = ~pi0684 & ~n42842;
  assign n42844 = pi0684 & pi3413;
  assign n42845 = ~n42843 & ~n42844;
  assign n42846 = n42803 & ~n42845;
  assign n42847 = pi1109 & ~n42803;
  assign n42848 = ~n42846 & ~n42847;
  assign n42849 = n41544 & ~n42848;
  assign n42850 = pi1109 & ~n41544;
  assign po1415 = n42849 | n42850;
  assign n42852 = ~pi0759 & n18698;
  assign n42853 = pi0759 & ~n13988;
  assign n42854 = ~n42852 & ~n42853;
  assign n42855 = ~pi0684 & ~n42854;
  assign n42856 = pi0684 & pi3405;
  assign n42857 = ~n42855 & ~n42856;
  assign n42858 = n42803 & ~n42857;
  assign n42859 = pi1110 & ~n42803;
  assign n42860 = ~n42858 & ~n42859;
  assign n42861 = n41544 & ~n42860;
  assign n42862 = pi1110 & ~n41544;
  assign po1416 = n42861 | n42862;
  assign n42864 = ~pi0759 & n18626;
  assign n42865 = pi0759 & ~n12415;
  assign n42866 = ~n42864 & ~n42865;
  assign n42867 = ~pi0684 & ~n42866;
  assign n42868 = pi0684 & pi3414;
  assign n42869 = ~n42867 & ~n42868;
  assign n42870 = n42803 & ~n42869;
  assign n42871 = pi1111 & ~n42803;
  assign n42872 = ~n42870 & ~n42871;
  assign n42873 = n41544 & ~n42872;
  assign n42874 = pi1111 & ~n41544;
  assign po1417 = n42873 | n42874;
  assign n42876 = ~pi0759 & n18593;
  assign n42877 = pi0759 & ~n14816;
  assign n42878 = ~n42876 & ~n42877;
  assign n42879 = ~pi0684 & ~n42878;
  assign n42880 = pi0684 & pi3404;
  assign n42881 = ~n42879 & ~n42880;
  assign n42882 = n42803 & ~n42881;
  assign n42883 = pi1112 & ~n42803;
  assign n42884 = ~n42882 & ~n42883;
  assign n42885 = n41544 & ~n42884;
  assign n42886 = pi1112 & ~n41544;
  assign po1418 = n42885 | n42886;
  assign n42888 = ~pi0759 & n18520;
  assign n42889 = pi0759 & ~n15115;
  assign n42890 = ~n42888 & ~n42889;
  assign n42891 = ~pi0684 & ~n42890;
  assign n42892 = pi0684 & pi3402;
  assign n42893 = ~n42891 & ~n42892;
  assign n42894 = n42803 & ~n42893;
  assign n42895 = pi1113 & ~n42803;
  assign n42896 = ~n42894 & ~n42895;
  assign n42897 = n41544 & ~n42896;
  assign n42898 = pi1113 & ~n41544;
  assign po1419 = n42897 | n42898;
  assign n42900 = ~pi0759 & ~n18402;
  assign n42901 = pi0759 & ~n12061;
  assign n42902 = ~n42900 & ~n42901;
  assign n42903 = ~pi0684 & ~n42902;
  assign n42904 = pi0684 & pi3403;
  assign n42905 = ~n42903 & ~n42904;
  assign n42906 = n42803 & ~n42905;
  assign n42907 = pi1114 & ~n42803;
  assign n42908 = ~n42906 & ~n42907;
  assign n42909 = n41544 & ~n42908;
  assign n42910 = pi1114 & ~n41544;
  assign po1420 = n42909 | n42910;
  assign n42912 = ~pi0759 & n15577;
  assign n42913 = pi0759 & ~n9825;
  assign n42914 = ~n42912 & ~n42913;
  assign n42915 = ~pi0684 & ~n42914;
  assign n42916 = pi0684 & pi3430;
  assign n42917 = ~n42915 & ~n42916;
  assign n42918 = n42803 & ~n42917;
  assign n42919 = pi1115 & ~n42803;
  assign n42920 = ~n42918 & ~n42919;
  assign n42921 = n41544 & ~n42920;
  assign n42922 = pi1115 & ~n41544;
  assign po1421 = n42921 | n42922;
  assign n42924 = ~pi0759 & n16098;
  assign n42925 = pi0759 & ~n10608;
  assign n42926 = ~n42924 & ~n42925;
  assign n42927 = ~pi0684 & ~n42926;
  assign n42928 = pi0684 & pi3421;
  assign n42929 = ~n42927 & ~n42928;
  assign n42930 = n42803 & ~n42929;
  assign n42931 = pi1116 & ~n42803;
  assign n42932 = ~n42930 & ~n42931;
  assign n42933 = n41544 & ~n42932;
  assign n42934 = pi1116 & ~n41544;
  assign po1422 = n42933 | n42934;
  assign n42936 = ~pi0759 & n19148;
  assign n42937 = pi0759 & ~n15426;
  assign n42938 = ~n42936 & ~n42937;
  assign n42939 = ~pi0684 & ~n42938;
  assign n42940 = pi0684 & pi3422;
  assign n42941 = ~n42939 & ~n42940;
  assign n42942 = n42803 & ~n42941;
  assign n42943 = pi1117 & ~n42803;
  assign n42944 = ~n42942 & ~n42943;
  assign n42945 = n41544 & ~n42944;
  assign n42946 = pi1117 & ~n41544;
  assign po1423 = n42945 | n42946;
  assign n42948 = ~pi0759 & n19075;
  assign n42949 = pi0759 & ~n14403;
  assign n42950 = ~n42948 & ~n42949;
  assign n42951 = ~pi0684 & ~n42950;
  assign n42952 = pi0684 & pi3401;
  assign n42953 = ~n42951 & ~n42952;
  assign n42954 = n42803 & ~n42953;
  assign n42955 = pi1118 & ~n42803;
  assign n42956 = ~n42954 & ~n42955;
  assign n42957 = n41544 & ~n42956;
  assign n42958 = pi1118 & ~n41544;
  assign po1424 = n42957 | n42958;
  assign n42960 = ~pi0759 & ~pi3400;
  assign n42961 = pi0759 & ~n11181;
  assign n42962 = ~n42960 & ~n42961;
  assign n42963 = ~pi0684 & ~n42962;
  assign n42964 = pi0684 & pi3400;
  assign n42965 = ~n42963 & ~n42964;
  assign n42966 = n42803 & ~n42965;
  assign n42967 = pi1119 & ~n42803;
  assign n42968 = ~n42966 & ~n42967;
  assign n42969 = n41544 & ~n42968;
  assign n42970 = pi1119 & ~n41544;
  assign po1425 = n42969 | n42970;
  assign n42972 = pi0976 & n42210;
  assign n42973 = n42802 & n42972;
  assign n42974 = ~n42809 & n42973;
  assign n42975 = pi1120 & ~n42973;
  assign n42976 = ~n42974 & ~n42975;
  assign n42977 = n41544 & ~n42976;
  assign n42978 = pi1120 & ~n41544;
  assign po1426 = n42977 | n42978;
  assign n42980 = ~n42821 & n42973;
  assign n42981 = pi1121 & ~n42973;
  assign n42982 = ~n42980 & ~n42981;
  assign n42983 = n41544 & ~n42982;
  assign n42984 = pi1121 & ~n41544;
  assign po1427 = n42983 | n42984;
  assign n42986 = ~n42833 & n42973;
  assign n42987 = pi1122 & ~n42973;
  assign n42988 = ~n42986 & ~n42987;
  assign n42989 = n41544 & ~n42988;
  assign n42990 = pi1122 & ~n41544;
  assign po1428 = n42989 | n42990;
  assign n42992 = ~n42845 & n42973;
  assign n42993 = pi1123 & ~n42973;
  assign n42994 = ~n42992 & ~n42993;
  assign n42995 = n41544 & ~n42994;
  assign n42996 = pi1123 & ~n41544;
  assign po1429 = n42995 | n42996;
  assign n42998 = ~n42857 & n42973;
  assign n42999 = pi1124 & ~n42973;
  assign n43000 = ~n42998 & ~n42999;
  assign n43001 = n41544 & ~n43000;
  assign n43002 = pi1124 & ~n41544;
  assign po1430 = n43001 | n43002;
  assign n43004 = ~n42869 & n42973;
  assign n43005 = pi1125 & ~n42973;
  assign n43006 = ~n43004 & ~n43005;
  assign n43007 = n41544 & ~n43006;
  assign n43008 = pi1125 & ~n41544;
  assign po1431 = n43007 | n43008;
  assign n43010 = ~n42881 & n42973;
  assign n43011 = pi1126 & ~n42973;
  assign n43012 = ~n43010 & ~n43011;
  assign n43013 = n41544 & ~n43012;
  assign n43014 = pi1126 & ~n41544;
  assign po1432 = n43013 | n43014;
  assign n43016 = ~n42893 & n42973;
  assign n43017 = pi1127 & ~n42973;
  assign n43018 = ~n43016 & ~n43017;
  assign n43019 = n41544 & ~n43018;
  assign n43020 = pi1127 & ~n41544;
  assign po1433 = n43019 | n43020;
  assign n43022 = ~n42905 & n42973;
  assign n43023 = pi1128 & ~n42973;
  assign n43024 = ~n43022 & ~n43023;
  assign n43025 = n41544 & ~n43024;
  assign n43026 = pi1128 & ~n41544;
  assign po1434 = n43025 | n43026;
  assign n43028 = ~n42917 & n42973;
  assign n43029 = pi1129 & ~n42973;
  assign n43030 = ~n43028 & ~n43029;
  assign n43031 = n41544 & ~n43030;
  assign n43032 = pi1129 & ~n41544;
  assign po1435 = n43031 | n43032;
  assign n43034 = ~n42929 & n42973;
  assign n43035 = pi1130 & ~n42973;
  assign n43036 = ~n43034 & ~n43035;
  assign n43037 = n41544 & ~n43036;
  assign n43038 = pi1130 & ~n41544;
  assign po1436 = n43037 | n43038;
  assign n43040 = ~n42941 & n42973;
  assign n43041 = pi1131 & ~n42973;
  assign n43042 = ~n43040 & ~n43041;
  assign n43043 = n41544 & ~n43042;
  assign n43044 = pi1131 & ~n41544;
  assign po1437 = n43043 | n43044;
  assign n43046 = ~n42953 & n42973;
  assign n43047 = pi1132 & ~n42973;
  assign n43048 = ~n43046 & ~n43047;
  assign n43049 = n41544 & ~n43048;
  assign n43050 = pi1132 & ~n41544;
  assign po1438 = n43049 | n43050;
  assign n43052 = ~n42965 & n42973;
  assign n43053 = pi1133 & ~n42973;
  assign n43054 = ~n43052 & ~n43053;
  assign n43055 = n41544 & ~n43054;
  assign n43056 = pi1133 & ~n41544;
  assign po1439 = n43055 | n43056;
  assign n43058 = ~pi0976 & ~n42210;
  assign n43059 = ~n41903 & n42202;
  assign n43060 = n43058 & n43059;
  assign n43061 = ~n42809 & n43060;
  assign n43062 = pi1134 & ~n43060;
  assign n43063 = ~n43061 & ~n43062;
  assign n43064 = n41544 & ~n43063;
  assign n43065 = pi1134 & ~n41544;
  assign po1440 = n43064 | n43065;
  assign n43067 = ~n42821 & n43060;
  assign n43068 = pi1135 & ~n43060;
  assign n43069 = ~n43067 & ~n43068;
  assign n43070 = n41544 & ~n43069;
  assign n43071 = pi1135 & ~n41544;
  assign po1441 = n43070 | n43071;
  assign n43073 = ~n42833 & n43060;
  assign n43074 = pi1136 & ~n43060;
  assign n43075 = ~n43073 & ~n43074;
  assign n43076 = n41544 & ~n43075;
  assign n43077 = pi1136 & ~n41544;
  assign po1442 = n43076 | n43077;
  assign n43079 = ~n42845 & n43060;
  assign n43080 = pi1137 & ~n43060;
  assign n43081 = ~n43079 & ~n43080;
  assign n43082 = n41544 & ~n43081;
  assign n43083 = pi1137 & ~n41544;
  assign po1443 = n43082 | n43083;
  assign n43085 = ~n42857 & n43060;
  assign n43086 = pi1138 & ~n43060;
  assign n43087 = ~n43085 & ~n43086;
  assign n43088 = n41544 & ~n43087;
  assign n43089 = pi1138 & ~n41544;
  assign po1444 = n43088 | n43089;
  assign n43091 = ~n42869 & n43060;
  assign n43092 = pi1139 & ~n43060;
  assign n43093 = ~n43091 & ~n43092;
  assign n43094 = n41544 & ~n43093;
  assign n43095 = pi1139 & ~n41544;
  assign po1445 = n43094 | n43095;
  assign n43097 = ~n42881 & n43060;
  assign n43098 = pi1140 & ~n43060;
  assign n43099 = ~n43097 & ~n43098;
  assign n43100 = n41544 & ~n43099;
  assign n43101 = pi1140 & ~n41544;
  assign po1446 = n43100 | n43101;
  assign n43103 = ~n42893 & n43060;
  assign n43104 = pi1141 & ~n43060;
  assign n43105 = ~n43103 & ~n43104;
  assign n43106 = n41544 & ~n43105;
  assign n43107 = pi1141 & ~n41544;
  assign po1447 = n43106 | n43107;
  assign n43109 = ~n42905 & n43060;
  assign n43110 = pi1142 & ~n43060;
  assign n43111 = ~n43109 & ~n43110;
  assign n43112 = n41544 & ~n43111;
  assign n43113 = pi1142 & ~n41544;
  assign po1448 = n43112 | n43113;
  assign n43115 = ~n42917 & n43060;
  assign n43116 = pi1143 & ~n43060;
  assign n43117 = ~n43115 & ~n43116;
  assign n43118 = n41544 & ~n43117;
  assign n43119 = pi1143 & ~n41544;
  assign po1449 = n43118 | n43119;
  assign n43121 = ~n42929 & n43060;
  assign n43122 = pi1144 & ~n43060;
  assign n43123 = ~n43121 & ~n43122;
  assign n43124 = n41544 & ~n43123;
  assign n43125 = pi1144 & ~n41544;
  assign po1450 = n43124 | n43125;
  assign n43127 = ~n42941 & n43060;
  assign n43128 = pi1145 & ~n43060;
  assign n43129 = ~n43127 & ~n43128;
  assign n43130 = n41544 & ~n43129;
  assign n43131 = pi1145 & ~n41544;
  assign po1451 = n43130 | n43131;
  assign n43133 = ~n42953 & n43060;
  assign n43134 = pi1146 & ~n43060;
  assign n43135 = ~n43133 & ~n43134;
  assign n43136 = n41544 & ~n43135;
  assign n43137 = pi1146 & ~n41544;
  assign po1452 = n43136 | n43137;
  assign n43139 = ~n42965 & n43060;
  assign n43140 = pi1147 & ~n43060;
  assign n43141 = ~n43139 & ~n43140;
  assign n43142 = n41544 & ~n43141;
  assign n43143 = pi1147 & ~n41544;
  assign po1453 = n43142 | n43143;
  assign n43145 = pi0976 & ~n42210;
  assign n43146 = n43059 & n43145;
  assign n43147 = ~n42809 & n43146;
  assign n43148 = pi1148 & ~n43146;
  assign n43149 = ~n43147 & ~n43148;
  assign n43150 = n41544 & ~n43149;
  assign n43151 = pi1148 & ~n41544;
  assign po1454 = n43150 | n43151;
  assign n43153 = ~n42821 & n43146;
  assign n43154 = pi1149 & ~n43146;
  assign n43155 = ~n43153 & ~n43154;
  assign n43156 = n41544 & ~n43155;
  assign n43157 = pi1149 & ~n41544;
  assign po1455 = n43156 | n43157;
  assign n43159 = ~n42833 & n43146;
  assign n43160 = pi1150 & ~n43146;
  assign n43161 = ~n43159 & ~n43160;
  assign n43162 = n41544 & ~n43161;
  assign n43163 = pi1150 & ~n41544;
  assign po1456 = n43162 | n43163;
  assign n43165 = ~n42845 & n43146;
  assign n43166 = pi1151 & ~n43146;
  assign n43167 = ~n43165 & ~n43166;
  assign n43168 = n41544 & ~n43167;
  assign n43169 = pi1151 & ~n41544;
  assign po1457 = n43168 | n43169;
  assign n43171 = ~n42857 & n43146;
  assign n43172 = pi1152 & ~n43146;
  assign n43173 = ~n43171 & ~n43172;
  assign n43174 = n41544 & ~n43173;
  assign n43175 = pi1152 & ~n41544;
  assign po1458 = n43174 | n43175;
  assign n43177 = ~n42869 & n43146;
  assign n43178 = pi1153 & ~n43146;
  assign n43179 = ~n43177 & ~n43178;
  assign n43180 = n41544 & ~n43179;
  assign n43181 = pi1153 & ~n41544;
  assign po1459 = n43180 | n43181;
  assign n43183 = ~n42881 & n43146;
  assign n43184 = pi1154 & ~n43146;
  assign n43185 = ~n43183 & ~n43184;
  assign n43186 = n41544 & ~n43185;
  assign n43187 = pi1154 & ~n41544;
  assign po1460 = n43186 | n43187;
  assign n43189 = ~n42893 & n43146;
  assign n43190 = pi1155 & ~n43146;
  assign n43191 = ~n43189 & ~n43190;
  assign n43192 = n41544 & ~n43191;
  assign n43193 = pi1155 & ~n41544;
  assign po1461 = n43192 | n43193;
  assign n43195 = ~n42905 & n43146;
  assign n43196 = pi1156 & ~n43146;
  assign n43197 = ~n43195 & ~n43196;
  assign n43198 = n41544 & ~n43197;
  assign n43199 = pi1156 & ~n41544;
  assign po1462 = n43198 | n43199;
  assign n43201 = ~n42917 & n43146;
  assign n43202 = pi1157 & ~n43146;
  assign n43203 = ~n43201 & ~n43202;
  assign n43204 = n41544 & ~n43203;
  assign n43205 = pi1157 & ~n41544;
  assign po1463 = n43204 | n43205;
  assign n43207 = ~n42929 & n43146;
  assign n43208 = pi1158 & ~n43146;
  assign n43209 = ~n43207 & ~n43208;
  assign n43210 = n41544 & ~n43209;
  assign n43211 = pi1158 & ~n41544;
  assign po1464 = n43210 | n43211;
  assign n43213 = ~n42941 & n43146;
  assign n43214 = pi1159 & ~n43146;
  assign n43215 = ~n43213 & ~n43214;
  assign n43216 = n41544 & ~n43215;
  assign n43217 = pi1159 & ~n41544;
  assign po1465 = n43216 | n43217;
  assign n43219 = ~n42953 & n43146;
  assign n43220 = pi1160 & ~n43146;
  assign n43221 = ~n43219 & ~n43220;
  assign n43222 = n41544 & ~n43221;
  assign n43223 = pi1160 & ~n41544;
  assign po1466 = n43222 | n43223;
  assign n43225 = ~n42965 & n43146;
  assign n43226 = pi1161 & ~n43146;
  assign n43227 = ~n43225 & ~n43226;
  assign n43228 = n41544 & ~n43227;
  assign n43229 = pi1161 & ~n41544;
  assign po1467 = n43228 | n43229;
  assign n43231 = n41903 & n42202;
  assign n43232 = n43058 & n43231;
  assign n43233 = ~n42809 & n43232;
  assign n43234 = pi1162 & ~n43232;
  assign n43235 = ~n43233 & ~n43234;
  assign n43236 = n41544 & ~n43235;
  assign n43237 = pi1162 & ~n41544;
  assign po1468 = n43236 | n43237;
  assign n43239 = ~n42821 & n43232;
  assign n43240 = pi1163 & ~n43232;
  assign n43241 = ~n43239 & ~n43240;
  assign n43242 = n41544 & ~n43241;
  assign n43243 = pi1163 & ~n41544;
  assign po1469 = n43242 | n43243;
  assign n43245 = ~n42833 & n43232;
  assign n43246 = pi1164 & ~n43232;
  assign n43247 = ~n43245 & ~n43246;
  assign n43248 = n41544 & ~n43247;
  assign n43249 = pi1164 & ~n41544;
  assign po1470 = n43248 | n43249;
  assign n43251 = ~n42845 & n43232;
  assign n43252 = pi1165 & ~n43232;
  assign n43253 = ~n43251 & ~n43252;
  assign n43254 = n41544 & ~n43253;
  assign n43255 = pi1165 & ~n41544;
  assign po1471 = n43254 | n43255;
  assign n43257 = ~n42857 & n43232;
  assign n43258 = pi1166 & ~n43232;
  assign n43259 = ~n43257 & ~n43258;
  assign n43260 = n41544 & ~n43259;
  assign n43261 = pi1166 & ~n41544;
  assign po1472 = n43260 | n43261;
  assign n43263 = ~n42869 & n43232;
  assign n43264 = pi1167 & ~n43232;
  assign n43265 = ~n43263 & ~n43264;
  assign n43266 = n41544 & ~n43265;
  assign n43267 = pi1167 & ~n41544;
  assign po1473 = n43266 | n43267;
  assign n43269 = ~n42881 & n43232;
  assign n43270 = pi1168 & ~n43232;
  assign n43271 = ~n43269 & ~n43270;
  assign n43272 = n41544 & ~n43271;
  assign n43273 = pi1168 & ~n41544;
  assign po1474 = n43272 | n43273;
  assign n43275 = ~n42893 & n43232;
  assign n43276 = pi1169 & ~n43232;
  assign n43277 = ~n43275 & ~n43276;
  assign n43278 = n41544 & ~n43277;
  assign n43279 = pi1169 & ~n41544;
  assign po1475 = n43278 | n43279;
  assign n43281 = ~n42905 & n43232;
  assign n43282 = pi1170 & ~n43232;
  assign n43283 = ~n43281 & ~n43282;
  assign n43284 = n41544 & ~n43283;
  assign n43285 = pi1170 & ~n41544;
  assign po1476 = n43284 | n43285;
  assign n43287 = ~n42917 & n43232;
  assign n43288 = pi1171 & ~n43232;
  assign n43289 = ~n43287 & ~n43288;
  assign n43290 = n41544 & ~n43289;
  assign n43291 = pi1171 & ~n41544;
  assign po1477 = n43290 | n43291;
  assign n43293 = ~n42929 & n43232;
  assign n43294 = pi1172 & ~n43232;
  assign n43295 = ~n43293 & ~n43294;
  assign n43296 = n41544 & ~n43295;
  assign n43297 = pi1172 & ~n41544;
  assign po1478 = n43296 | n43297;
  assign n43299 = ~n42941 & n43232;
  assign n43300 = pi1173 & ~n43232;
  assign n43301 = ~n43299 & ~n43300;
  assign n43302 = n41544 & ~n43301;
  assign n43303 = pi1173 & ~n41544;
  assign po1479 = n43302 | n43303;
  assign n43305 = ~n42953 & n43232;
  assign n43306 = pi1174 & ~n43232;
  assign n43307 = ~n43305 & ~n43306;
  assign n43308 = n41544 & ~n43307;
  assign n43309 = pi1174 & ~n41544;
  assign po1480 = n43308 | n43309;
  assign n43311 = ~n42965 & n43232;
  assign n43312 = pi1175 & ~n43232;
  assign n43313 = ~n43311 & ~n43312;
  assign n43314 = n41544 & ~n43313;
  assign n43315 = pi1175 & ~n41544;
  assign po1481 = n43314 | n43315;
  assign n43317 = n43145 & n43231;
  assign n43318 = ~n42809 & n43317;
  assign n43319 = pi1176 & ~n43317;
  assign n43320 = ~n43318 & ~n43319;
  assign n43321 = n41544 & ~n43320;
  assign n43322 = pi1176 & ~n41544;
  assign po1482 = n43321 | n43322;
  assign n43324 = ~n42821 & n43317;
  assign n43325 = pi1177 & ~n43317;
  assign n43326 = ~n43324 & ~n43325;
  assign n43327 = n41544 & ~n43326;
  assign n43328 = pi1177 & ~n41544;
  assign po1483 = n43327 | n43328;
  assign n43330 = ~n42833 & n43317;
  assign n43331 = pi1178 & ~n43317;
  assign n43332 = ~n43330 & ~n43331;
  assign n43333 = n41544 & ~n43332;
  assign n43334 = pi1178 & ~n41544;
  assign po1484 = n43333 | n43334;
  assign n43336 = ~n42845 & n43317;
  assign n43337 = pi1179 & ~n43317;
  assign n43338 = ~n43336 & ~n43337;
  assign n43339 = n41544 & ~n43338;
  assign n43340 = pi1179 & ~n41544;
  assign po1485 = n43339 | n43340;
  assign n43342 = ~n42857 & n43317;
  assign n43343 = pi1180 & ~n43317;
  assign n43344 = ~n43342 & ~n43343;
  assign n43345 = n41544 & ~n43344;
  assign n43346 = pi1180 & ~n41544;
  assign po1486 = n43345 | n43346;
  assign n43348 = ~n42869 & n43317;
  assign n43349 = pi1181 & ~n43317;
  assign n43350 = ~n43348 & ~n43349;
  assign n43351 = n41544 & ~n43350;
  assign n43352 = pi1181 & ~n41544;
  assign po1487 = n43351 | n43352;
  assign n43354 = ~n42881 & n43317;
  assign n43355 = pi1182 & ~n43317;
  assign n43356 = ~n43354 & ~n43355;
  assign n43357 = n41544 & ~n43356;
  assign n43358 = pi1182 & ~n41544;
  assign po1488 = n43357 | n43358;
  assign n43360 = ~n42893 & n43317;
  assign n43361 = pi1183 & ~n43317;
  assign n43362 = ~n43360 & ~n43361;
  assign n43363 = n41544 & ~n43362;
  assign n43364 = pi1183 & ~n41544;
  assign po1489 = n43363 | n43364;
  assign n43366 = ~n42905 & n43317;
  assign n43367 = pi1184 & ~n43317;
  assign n43368 = ~n43366 & ~n43367;
  assign n43369 = n41544 & ~n43368;
  assign n43370 = pi1184 & ~n41544;
  assign po1490 = n43369 | n43370;
  assign n43372 = ~n42917 & n43317;
  assign n43373 = pi1185 & ~n43317;
  assign n43374 = ~n43372 & ~n43373;
  assign n43375 = n41544 & ~n43374;
  assign n43376 = pi1185 & ~n41544;
  assign po1491 = n43375 | n43376;
  assign n43378 = ~n42929 & n43317;
  assign n43379 = pi1186 & ~n43317;
  assign n43380 = ~n43378 & ~n43379;
  assign n43381 = n41544 & ~n43380;
  assign n43382 = pi1186 & ~n41544;
  assign po1492 = n43381 | n43382;
  assign n43384 = ~n42941 & n43317;
  assign n43385 = pi1187 & ~n43317;
  assign n43386 = ~n43384 & ~n43385;
  assign n43387 = n41544 & ~n43386;
  assign n43388 = pi1187 & ~n41544;
  assign po1493 = n43387 | n43388;
  assign n43390 = ~n42953 & n43317;
  assign n43391 = pi1188 & ~n43317;
  assign n43392 = ~n43390 & ~n43391;
  assign n43393 = n41544 & ~n43392;
  assign n43394 = pi1188 & ~n41544;
  assign po1494 = n43393 | n43394;
  assign n43396 = ~n42965 & n43317;
  assign n43397 = pi1189 & ~n43317;
  assign n43398 = ~n43396 & ~n43397;
  assign n43399 = n41544 & ~n43398;
  assign n43400 = pi1189 & ~n41544;
  assign po1495 = n43399 | n43400;
  assign n43402 = ~n41903 & ~n42202;
  assign n43403 = n43058 & n43402;
  assign n43404 = ~n42809 & n43403;
  assign n43405 = pi1190 & ~n43403;
  assign n43406 = ~n43404 & ~n43405;
  assign n43407 = n41544 & ~n43406;
  assign n43408 = pi1190 & ~n41544;
  assign po1496 = n43407 | n43408;
  assign n43410 = ~n42821 & n43403;
  assign n43411 = pi1191 & ~n43403;
  assign n43412 = ~n43410 & ~n43411;
  assign n43413 = n41544 & ~n43412;
  assign n43414 = pi1191 & ~n41544;
  assign po1497 = n43413 | n43414;
  assign n43416 = ~n42833 & n43403;
  assign n43417 = pi1192 & ~n43403;
  assign n43418 = ~n43416 & ~n43417;
  assign n43419 = n41544 & ~n43418;
  assign n43420 = pi1192 & ~n41544;
  assign po1498 = n43419 | n43420;
  assign n43422 = ~n42845 & n43403;
  assign n43423 = pi1193 & ~n43403;
  assign n43424 = ~n43422 & ~n43423;
  assign n43425 = n41544 & ~n43424;
  assign n43426 = pi1193 & ~n41544;
  assign po1499 = n43425 | n43426;
  assign n43428 = ~n42857 & n43403;
  assign n43429 = pi1194 & ~n43403;
  assign n43430 = ~n43428 & ~n43429;
  assign n43431 = n41544 & ~n43430;
  assign n43432 = pi1194 & ~n41544;
  assign po1500 = n43431 | n43432;
  assign n43434 = ~n42869 & n43403;
  assign n43435 = pi1195 & ~n43403;
  assign n43436 = ~n43434 & ~n43435;
  assign n43437 = n41544 & ~n43436;
  assign n43438 = pi1195 & ~n41544;
  assign po1501 = n43437 | n43438;
  assign n43440 = ~n42881 & n43403;
  assign n43441 = pi1196 & ~n43403;
  assign n43442 = ~n43440 & ~n43441;
  assign n43443 = n41544 & ~n43442;
  assign n43444 = pi1196 & ~n41544;
  assign po1502 = n43443 | n43444;
  assign n43446 = ~n42893 & n43403;
  assign n43447 = pi1197 & ~n43403;
  assign n43448 = ~n43446 & ~n43447;
  assign n43449 = n41544 & ~n43448;
  assign n43450 = pi1197 & ~n41544;
  assign po1503 = n43449 | n43450;
  assign n43452 = ~n42905 & n43403;
  assign n43453 = pi1198 & ~n43403;
  assign n43454 = ~n43452 & ~n43453;
  assign n43455 = n41544 & ~n43454;
  assign n43456 = pi1198 & ~n41544;
  assign po1504 = n43455 | n43456;
  assign n43458 = ~n42917 & n43403;
  assign n43459 = pi1199 & ~n43403;
  assign n43460 = ~n43458 & ~n43459;
  assign n43461 = n41544 & ~n43460;
  assign n43462 = pi1199 & ~n41544;
  assign po1505 = n43461 | n43462;
  assign n43464 = ~n42929 & n43403;
  assign n43465 = pi1200 & ~n43403;
  assign n43466 = ~n43464 & ~n43465;
  assign n43467 = n41544 & ~n43466;
  assign n43468 = pi1200 & ~n41544;
  assign po1506 = n43467 | n43468;
  assign n43470 = ~n42941 & n43403;
  assign n43471 = pi1201 & ~n43403;
  assign n43472 = ~n43470 & ~n43471;
  assign n43473 = n41544 & ~n43472;
  assign n43474 = pi1201 & ~n41544;
  assign po1507 = n43473 | n43474;
  assign n43476 = ~n42953 & n43403;
  assign n43477 = pi1202 & ~n43403;
  assign n43478 = ~n43476 & ~n43477;
  assign n43479 = n41544 & ~n43478;
  assign n43480 = pi1202 & ~n41544;
  assign po1508 = n43479 | n43480;
  assign n43482 = ~n42965 & n43403;
  assign n43483 = pi1203 & ~n43403;
  assign n43484 = ~n43482 & ~n43483;
  assign n43485 = n41544 & ~n43484;
  assign n43486 = pi1203 & ~n41544;
  assign po1509 = n43485 | n43486;
  assign n43488 = n43145 & n43402;
  assign n43489 = ~n42809 & n43488;
  assign n43490 = pi1204 & ~n43488;
  assign n43491 = ~n43489 & ~n43490;
  assign n43492 = n41544 & ~n43491;
  assign n43493 = pi1204 & ~n41544;
  assign po1510 = n43492 | n43493;
  assign n43495 = ~n42821 & n43488;
  assign n43496 = pi1205 & ~n43488;
  assign n43497 = ~n43495 & ~n43496;
  assign n43498 = n41544 & ~n43497;
  assign n43499 = pi1205 & ~n41544;
  assign po1511 = n43498 | n43499;
  assign n43501 = ~n42833 & n43488;
  assign n43502 = pi1206 & ~n43488;
  assign n43503 = ~n43501 & ~n43502;
  assign n43504 = n41544 & ~n43503;
  assign n43505 = pi1206 & ~n41544;
  assign po1512 = n43504 | n43505;
  assign n43507 = ~n42845 & n43488;
  assign n43508 = pi1207 & ~n43488;
  assign n43509 = ~n43507 & ~n43508;
  assign n43510 = n41544 & ~n43509;
  assign n43511 = pi1207 & ~n41544;
  assign po1513 = n43510 | n43511;
  assign n43513 = ~n42857 & n43488;
  assign n43514 = pi1208 & ~n43488;
  assign n43515 = ~n43513 & ~n43514;
  assign n43516 = n41544 & ~n43515;
  assign n43517 = pi1208 & ~n41544;
  assign po1514 = n43516 | n43517;
  assign n43519 = ~n42869 & n43488;
  assign n43520 = pi1209 & ~n43488;
  assign n43521 = ~n43519 & ~n43520;
  assign n43522 = n41544 & ~n43521;
  assign n43523 = pi1209 & ~n41544;
  assign po1515 = n43522 | n43523;
  assign n43525 = ~n42881 & n43488;
  assign n43526 = pi1210 & ~n43488;
  assign n43527 = ~n43525 & ~n43526;
  assign n43528 = n41544 & ~n43527;
  assign n43529 = pi1210 & ~n41544;
  assign po1516 = n43528 | n43529;
  assign n43531 = ~n42893 & n43488;
  assign n43532 = pi1211 & ~n43488;
  assign n43533 = ~n43531 & ~n43532;
  assign n43534 = n41544 & ~n43533;
  assign n43535 = pi1211 & ~n41544;
  assign po1517 = n43534 | n43535;
  assign n43537 = ~n42905 & n43488;
  assign n43538 = pi1212 & ~n43488;
  assign n43539 = ~n43537 & ~n43538;
  assign n43540 = n41544 & ~n43539;
  assign n43541 = pi1212 & ~n41544;
  assign po1518 = n43540 | n43541;
  assign n43543 = ~n42917 & n43488;
  assign n43544 = pi1213 & ~n43488;
  assign n43545 = ~n43543 & ~n43544;
  assign n43546 = n41544 & ~n43545;
  assign n43547 = pi1213 & ~n41544;
  assign po1519 = n43546 | n43547;
  assign n43549 = ~n42929 & n43488;
  assign n43550 = pi1214 & ~n43488;
  assign n43551 = ~n43549 & ~n43550;
  assign n43552 = n41544 & ~n43551;
  assign n43553 = pi1214 & ~n41544;
  assign po1520 = n43552 | n43553;
  assign n43555 = ~n42941 & n43488;
  assign n43556 = pi1215 & ~n43488;
  assign n43557 = ~n43555 & ~n43556;
  assign n43558 = n41544 & ~n43557;
  assign n43559 = pi1215 & ~n41544;
  assign po1521 = n43558 | n43559;
  assign n43561 = ~n42953 & n43488;
  assign n43562 = pi1216 & ~n43488;
  assign n43563 = ~n43561 & ~n43562;
  assign n43564 = n41544 & ~n43563;
  assign n43565 = pi1216 & ~n41544;
  assign po1522 = n43564 | n43565;
  assign n43567 = ~n42965 & n43488;
  assign n43568 = pi1217 & ~n43488;
  assign n43569 = ~n43567 & ~n43568;
  assign n43570 = n41544 & ~n43569;
  assign n43571 = pi1217 & ~n41544;
  assign po1523 = n43570 | n43571;
  assign n43573 = n42802 & n43058;
  assign n43574 = ~n42809 & n43573;
  assign n43575 = pi1218 & ~n43573;
  assign n43576 = ~n43574 & ~n43575;
  assign n43577 = n41544 & ~n43576;
  assign n43578 = pi1218 & ~n41544;
  assign po1524 = n43577 | n43578;
  assign n43580 = ~n42821 & n43573;
  assign n43581 = pi1219 & ~n43573;
  assign n43582 = ~n43580 & ~n43581;
  assign n43583 = n41544 & ~n43582;
  assign n43584 = pi1219 & ~n41544;
  assign po1525 = n43583 | n43584;
  assign n43586 = ~n42833 & n43573;
  assign n43587 = pi1220 & ~n43573;
  assign n43588 = ~n43586 & ~n43587;
  assign n43589 = n41544 & ~n43588;
  assign n43590 = pi1220 & ~n41544;
  assign po1526 = n43589 | n43590;
  assign n43592 = ~n42845 & n43573;
  assign n43593 = pi1221 & ~n43573;
  assign n43594 = ~n43592 & ~n43593;
  assign n43595 = n41544 & ~n43594;
  assign n43596 = pi1221 & ~n41544;
  assign po1527 = n43595 | n43596;
  assign n43598 = ~n42857 & n43573;
  assign n43599 = pi1222 & ~n43573;
  assign n43600 = ~n43598 & ~n43599;
  assign n43601 = n41544 & ~n43600;
  assign n43602 = pi1222 & ~n41544;
  assign po1528 = n43601 | n43602;
  assign n43604 = ~n42869 & n43573;
  assign n43605 = pi1223 & ~n43573;
  assign n43606 = ~n43604 & ~n43605;
  assign n43607 = n41544 & ~n43606;
  assign n43608 = pi1223 & ~n41544;
  assign po1529 = n43607 | n43608;
  assign n43610 = ~n42881 & n43573;
  assign n43611 = pi1224 & ~n43573;
  assign n43612 = ~n43610 & ~n43611;
  assign n43613 = n41544 & ~n43612;
  assign n43614 = pi1224 & ~n41544;
  assign po1530 = n43613 | n43614;
  assign n43616 = ~n42893 & n43573;
  assign n43617 = pi1225 & ~n43573;
  assign n43618 = ~n43616 & ~n43617;
  assign n43619 = n41544 & ~n43618;
  assign n43620 = pi1225 & ~n41544;
  assign po1531 = n43619 | n43620;
  assign n43622 = ~n42905 & n43573;
  assign n43623 = pi1226 & ~n43573;
  assign n43624 = ~n43622 & ~n43623;
  assign n43625 = n41544 & ~n43624;
  assign n43626 = pi1226 & ~n41544;
  assign po1532 = n43625 | n43626;
  assign n43628 = ~n42917 & n43573;
  assign n43629 = pi1227 & ~n43573;
  assign n43630 = ~n43628 & ~n43629;
  assign n43631 = n41544 & ~n43630;
  assign n43632 = pi1227 & ~n41544;
  assign po1533 = n43631 | n43632;
  assign n43634 = ~n42929 & n43573;
  assign n43635 = pi1228 & ~n43573;
  assign n43636 = ~n43634 & ~n43635;
  assign n43637 = n41544 & ~n43636;
  assign n43638 = pi1228 & ~n41544;
  assign po1534 = n43637 | n43638;
  assign n43640 = ~n42941 & n43573;
  assign n43641 = pi1229 & ~n43573;
  assign n43642 = ~n43640 & ~n43641;
  assign n43643 = n41544 & ~n43642;
  assign n43644 = pi1229 & ~n41544;
  assign po1535 = n43643 | n43644;
  assign n43646 = ~n42953 & n43573;
  assign n43647 = pi1230 & ~n43573;
  assign n43648 = ~n43646 & ~n43647;
  assign n43649 = n41544 & ~n43648;
  assign n43650 = pi1230 & ~n41544;
  assign po1536 = n43649 | n43650;
  assign n43652 = ~n42965 & n43573;
  assign n43653 = pi1231 & ~n43573;
  assign n43654 = ~n43652 & ~n43653;
  assign n43655 = n41544 & ~n43654;
  assign n43656 = pi1231 & ~n41544;
  assign po1537 = n43655 | n43656;
  assign n43658 = n42801 & n43059;
  assign n43659 = ~n42809 & n43658;
  assign n43660 = pi1232 & ~n43658;
  assign n43661 = ~n43659 & ~n43660;
  assign n43662 = n41544 & ~n43661;
  assign n43663 = pi1232 & ~n41544;
  assign po1538 = n43662 | n43663;
  assign n43665 = ~n42821 & n43658;
  assign n43666 = pi1233 & ~n43658;
  assign n43667 = ~n43665 & ~n43666;
  assign n43668 = n41544 & ~n43667;
  assign n43669 = pi1233 & ~n41544;
  assign po1539 = n43668 | n43669;
  assign n43671 = ~n42833 & n43658;
  assign n43672 = pi1234 & ~n43658;
  assign n43673 = ~n43671 & ~n43672;
  assign n43674 = n41544 & ~n43673;
  assign n43675 = pi1234 & ~n41544;
  assign po1540 = n43674 | n43675;
  assign n43677 = ~n42845 & n43658;
  assign n43678 = pi1235 & ~n43658;
  assign n43679 = ~n43677 & ~n43678;
  assign n43680 = n41544 & ~n43679;
  assign n43681 = pi1235 & ~n41544;
  assign po1541 = n43680 | n43681;
  assign n43683 = ~n42857 & n43658;
  assign n43684 = pi1236 & ~n43658;
  assign n43685 = ~n43683 & ~n43684;
  assign n43686 = n41544 & ~n43685;
  assign n43687 = pi1236 & ~n41544;
  assign po1542 = n43686 | n43687;
  assign n43689 = ~n42869 & n43658;
  assign n43690 = pi1237 & ~n43658;
  assign n43691 = ~n43689 & ~n43690;
  assign n43692 = n41544 & ~n43691;
  assign n43693 = pi1237 & ~n41544;
  assign po1543 = n43692 | n43693;
  assign n43695 = ~n42881 & n43658;
  assign n43696 = pi1238 & ~n43658;
  assign n43697 = ~n43695 & ~n43696;
  assign n43698 = n41544 & ~n43697;
  assign n43699 = pi1238 & ~n41544;
  assign po1544 = n43698 | n43699;
  assign n43701 = ~n42893 & n43658;
  assign n43702 = pi1239 & ~n43658;
  assign n43703 = ~n43701 & ~n43702;
  assign n43704 = n41544 & ~n43703;
  assign n43705 = pi1239 & ~n41544;
  assign po1545 = n43704 | n43705;
  assign n43707 = ~n42905 & n43658;
  assign n43708 = pi1240 & ~n43658;
  assign n43709 = ~n43707 & ~n43708;
  assign n43710 = n41544 & ~n43709;
  assign n43711 = pi1240 & ~n41544;
  assign po1546 = n43710 | n43711;
  assign n43713 = ~n42917 & n43658;
  assign n43714 = pi1241 & ~n43658;
  assign n43715 = ~n43713 & ~n43714;
  assign n43716 = n41544 & ~n43715;
  assign n43717 = pi1241 & ~n41544;
  assign po1547 = n43716 | n43717;
  assign n43719 = ~n42929 & n43658;
  assign n43720 = pi1242 & ~n43658;
  assign n43721 = ~n43719 & ~n43720;
  assign n43722 = n41544 & ~n43721;
  assign n43723 = pi1242 & ~n41544;
  assign po1548 = n43722 | n43723;
  assign n43725 = ~n42941 & n43658;
  assign n43726 = pi1243 & ~n43658;
  assign n43727 = ~n43725 & ~n43726;
  assign n43728 = n41544 & ~n43727;
  assign n43729 = pi1243 & ~n41544;
  assign po1549 = n43728 | n43729;
  assign n43731 = ~n42953 & n43658;
  assign n43732 = pi1244 & ~n43658;
  assign n43733 = ~n43731 & ~n43732;
  assign n43734 = n41544 & ~n43733;
  assign n43735 = pi1244 & ~n41544;
  assign po1550 = n43734 | n43735;
  assign n43737 = ~n42965 & n43658;
  assign n43738 = pi1245 & ~n43658;
  assign n43739 = ~n43737 & ~n43738;
  assign n43740 = n41544 & ~n43739;
  assign n43741 = pi1245 & ~n41544;
  assign po1551 = n43740 | n43741;
  assign n43743 = n42972 & n43059;
  assign n43744 = ~n42809 & n43743;
  assign n43745 = pi1246 & ~n43743;
  assign n43746 = ~n43744 & ~n43745;
  assign n43747 = n41544 & ~n43746;
  assign n43748 = pi1246 & ~n41544;
  assign po1552 = n43747 | n43748;
  assign n43750 = ~n42821 & n43743;
  assign n43751 = pi1247 & ~n43743;
  assign n43752 = ~n43750 & ~n43751;
  assign n43753 = n41544 & ~n43752;
  assign n43754 = pi1247 & ~n41544;
  assign po1553 = n43753 | n43754;
  assign n43756 = ~n42833 & n43743;
  assign n43757 = pi1248 & ~n43743;
  assign n43758 = ~n43756 & ~n43757;
  assign n43759 = n41544 & ~n43758;
  assign n43760 = pi1248 & ~n41544;
  assign po1554 = n43759 | n43760;
  assign n43762 = ~n42845 & n43743;
  assign n43763 = pi1249 & ~n43743;
  assign n43764 = ~n43762 & ~n43763;
  assign n43765 = n41544 & ~n43764;
  assign n43766 = pi1249 & ~n41544;
  assign po1555 = n43765 | n43766;
  assign n43768 = ~n42857 & n43743;
  assign n43769 = pi1250 & ~n43743;
  assign n43770 = ~n43768 & ~n43769;
  assign n43771 = n41544 & ~n43770;
  assign n43772 = pi1250 & ~n41544;
  assign po1556 = n43771 | n43772;
  assign n43774 = ~n42869 & n43743;
  assign n43775 = pi1251 & ~n43743;
  assign n43776 = ~n43774 & ~n43775;
  assign n43777 = n41544 & ~n43776;
  assign n43778 = pi1251 & ~n41544;
  assign po1557 = n43777 | n43778;
  assign n43780 = ~n42881 & n43743;
  assign n43781 = pi1252 & ~n43743;
  assign n43782 = ~n43780 & ~n43781;
  assign n43783 = n41544 & ~n43782;
  assign n43784 = pi1252 & ~n41544;
  assign po1558 = n43783 | n43784;
  assign n43786 = ~n42893 & n43743;
  assign n43787 = pi1253 & ~n43743;
  assign n43788 = ~n43786 & ~n43787;
  assign n43789 = n41544 & ~n43788;
  assign n43790 = pi1253 & ~n41544;
  assign po1559 = n43789 | n43790;
  assign n43792 = ~n42905 & n43743;
  assign n43793 = pi1254 & ~n43743;
  assign n43794 = ~n43792 & ~n43793;
  assign n43795 = n41544 & ~n43794;
  assign n43796 = pi1254 & ~n41544;
  assign po1560 = n43795 | n43796;
  assign n43798 = ~n42917 & n43743;
  assign n43799 = pi1255 & ~n43743;
  assign n43800 = ~n43798 & ~n43799;
  assign n43801 = n41544 & ~n43800;
  assign n43802 = pi1255 & ~n41544;
  assign po1561 = n43801 | n43802;
  assign n43804 = ~n42929 & n43743;
  assign n43805 = pi1256 & ~n43743;
  assign n43806 = ~n43804 & ~n43805;
  assign n43807 = n41544 & ~n43806;
  assign n43808 = pi1256 & ~n41544;
  assign po1562 = n43807 | n43808;
  assign n43810 = ~n42941 & n43743;
  assign n43811 = pi1257 & ~n43743;
  assign n43812 = ~n43810 & ~n43811;
  assign n43813 = n41544 & ~n43812;
  assign n43814 = pi1257 & ~n41544;
  assign po1563 = n43813 | n43814;
  assign n43816 = ~n42953 & n43743;
  assign n43817 = pi1258 & ~n43743;
  assign n43818 = ~n43816 & ~n43817;
  assign n43819 = n41544 & ~n43818;
  assign n43820 = pi1258 & ~n41544;
  assign po1564 = n43819 | n43820;
  assign n43822 = ~n42965 & n43743;
  assign n43823 = pi1259 & ~n43743;
  assign n43824 = ~n43822 & ~n43823;
  assign n43825 = n41544 & ~n43824;
  assign n43826 = pi1259 & ~n41544;
  assign po1565 = n43825 | n43826;
  assign n43828 = n42801 & n43231;
  assign n43829 = ~n42809 & n43828;
  assign n43830 = pi1260 & ~n43828;
  assign n43831 = ~n43829 & ~n43830;
  assign n43832 = n41544 & ~n43831;
  assign n43833 = pi1260 & ~n41544;
  assign po1566 = n43832 | n43833;
  assign n43835 = ~n42821 & n43828;
  assign n43836 = pi1261 & ~n43828;
  assign n43837 = ~n43835 & ~n43836;
  assign n43838 = n41544 & ~n43837;
  assign n43839 = pi1261 & ~n41544;
  assign po1567 = n43838 | n43839;
  assign n43841 = ~n42833 & n43828;
  assign n43842 = pi1262 & ~n43828;
  assign n43843 = ~n43841 & ~n43842;
  assign n43844 = n41544 & ~n43843;
  assign n43845 = pi1262 & ~n41544;
  assign po1568 = n43844 | n43845;
  assign n43847 = ~n42845 & n43828;
  assign n43848 = pi1263 & ~n43828;
  assign n43849 = ~n43847 & ~n43848;
  assign n43850 = n41544 & ~n43849;
  assign n43851 = pi1263 & ~n41544;
  assign po1569 = n43850 | n43851;
  assign n43853 = ~n42857 & n43828;
  assign n43854 = pi1264 & ~n43828;
  assign n43855 = ~n43853 & ~n43854;
  assign n43856 = n41544 & ~n43855;
  assign n43857 = pi1264 & ~n41544;
  assign po1570 = n43856 | n43857;
  assign n43859 = ~n42869 & n43828;
  assign n43860 = pi1265 & ~n43828;
  assign n43861 = ~n43859 & ~n43860;
  assign n43862 = n41544 & ~n43861;
  assign n43863 = pi1265 & ~n41544;
  assign po1571 = n43862 | n43863;
  assign n43865 = ~n42881 & n43828;
  assign n43866 = pi1266 & ~n43828;
  assign n43867 = ~n43865 & ~n43866;
  assign n43868 = n41544 & ~n43867;
  assign n43869 = pi1266 & ~n41544;
  assign po1572 = n43868 | n43869;
  assign n43871 = ~n42893 & n43828;
  assign n43872 = pi1267 & ~n43828;
  assign n43873 = ~n43871 & ~n43872;
  assign n43874 = n41544 & ~n43873;
  assign n43875 = pi1267 & ~n41544;
  assign po1573 = n43874 | n43875;
  assign n43877 = ~n42905 & n43828;
  assign n43878 = pi1268 & ~n43828;
  assign n43879 = ~n43877 & ~n43878;
  assign n43880 = n41544 & ~n43879;
  assign n43881 = pi1268 & ~n41544;
  assign po1574 = n43880 | n43881;
  assign n43883 = ~n42917 & n43828;
  assign n43884 = pi1269 & ~n43828;
  assign n43885 = ~n43883 & ~n43884;
  assign n43886 = n41544 & ~n43885;
  assign n43887 = pi1269 & ~n41544;
  assign po1575 = n43886 | n43887;
  assign n43889 = ~n42929 & n43828;
  assign n43890 = pi1270 & ~n43828;
  assign n43891 = ~n43889 & ~n43890;
  assign n43892 = n41544 & ~n43891;
  assign n43893 = pi1270 & ~n41544;
  assign po1576 = n43892 | n43893;
  assign n43895 = ~n42941 & n43828;
  assign n43896 = pi1271 & ~n43828;
  assign n43897 = ~n43895 & ~n43896;
  assign n43898 = n41544 & ~n43897;
  assign n43899 = pi1271 & ~n41544;
  assign po1577 = n43898 | n43899;
  assign n43901 = ~n42953 & n43828;
  assign n43902 = pi1272 & ~n43828;
  assign n43903 = ~n43901 & ~n43902;
  assign n43904 = n41544 & ~n43903;
  assign n43905 = pi1272 & ~n41544;
  assign po1578 = n43904 | n43905;
  assign n43907 = ~n42965 & n43828;
  assign n43908 = pi1273 & ~n43828;
  assign n43909 = ~n43907 & ~n43908;
  assign n43910 = n41544 & ~n43909;
  assign n43911 = pi1273 & ~n41544;
  assign po1579 = n43910 | n43911;
  assign n43913 = n42972 & n43231;
  assign n43914 = ~n42809 & n43913;
  assign n43915 = pi1274 & ~n43913;
  assign n43916 = ~n43914 & ~n43915;
  assign n43917 = n41544 & ~n43916;
  assign n43918 = pi1274 & ~n41544;
  assign po1580 = n43917 | n43918;
  assign n43920 = ~n42821 & n43913;
  assign n43921 = pi1275 & ~n43913;
  assign n43922 = ~n43920 & ~n43921;
  assign n43923 = n41544 & ~n43922;
  assign n43924 = pi1275 & ~n41544;
  assign po1581 = n43923 | n43924;
  assign n43926 = ~n42833 & n43913;
  assign n43927 = pi1276 & ~n43913;
  assign n43928 = ~n43926 & ~n43927;
  assign n43929 = n41544 & ~n43928;
  assign n43930 = pi1276 & ~n41544;
  assign po1582 = n43929 | n43930;
  assign n43932 = ~n42845 & n43913;
  assign n43933 = pi1277 & ~n43913;
  assign n43934 = ~n43932 & ~n43933;
  assign n43935 = n41544 & ~n43934;
  assign n43936 = pi1277 & ~n41544;
  assign po1583 = n43935 | n43936;
  assign n43938 = ~n42857 & n43913;
  assign n43939 = pi1278 & ~n43913;
  assign n43940 = ~n43938 & ~n43939;
  assign n43941 = n41544 & ~n43940;
  assign n43942 = pi1278 & ~n41544;
  assign po1584 = n43941 | n43942;
  assign n43944 = ~n42869 & n43913;
  assign n43945 = pi1279 & ~n43913;
  assign n43946 = ~n43944 & ~n43945;
  assign n43947 = n41544 & ~n43946;
  assign n43948 = pi1279 & ~n41544;
  assign po1585 = n43947 | n43948;
  assign n43950 = ~n42881 & n43913;
  assign n43951 = pi1280 & ~n43913;
  assign n43952 = ~n43950 & ~n43951;
  assign n43953 = n41544 & ~n43952;
  assign n43954 = pi1280 & ~n41544;
  assign po1586 = n43953 | n43954;
  assign n43956 = ~n42893 & n43913;
  assign n43957 = pi1281 & ~n43913;
  assign n43958 = ~n43956 & ~n43957;
  assign n43959 = n41544 & ~n43958;
  assign n43960 = pi1281 & ~n41544;
  assign po1587 = n43959 | n43960;
  assign n43962 = ~n42905 & n43913;
  assign n43963 = pi1282 & ~n43913;
  assign n43964 = ~n43962 & ~n43963;
  assign n43965 = n41544 & ~n43964;
  assign n43966 = pi1282 & ~n41544;
  assign po1588 = n43965 | n43966;
  assign n43968 = ~n42917 & n43913;
  assign n43969 = pi1283 & ~n43913;
  assign n43970 = ~n43968 & ~n43969;
  assign n43971 = n41544 & ~n43970;
  assign n43972 = pi1283 & ~n41544;
  assign po1589 = n43971 | n43972;
  assign n43974 = ~n42929 & n43913;
  assign n43975 = pi1284 & ~n43913;
  assign n43976 = ~n43974 & ~n43975;
  assign n43977 = n41544 & ~n43976;
  assign n43978 = pi1284 & ~n41544;
  assign po1590 = n43977 | n43978;
  assign n43980 = ~n42941 & n43913;
  assign n43981 = pi1285 & ~n43913;
  assign n43982 = ~n43980 & ~n43981;
  assign n43983 = n41544 & ~n43982;
  assign n43984 = pi1285 & ~n41544;
  assign po1591 = n43983 | n43984;
  assign n43986 = ~n42953 & n43913;
  assign n43987 = pi1286 & ~n43913;
  assign n43988 = ~n43986 & ~n43987;
  assign n43989 = n41544 & ~n43988;
  assign n43990 = pi1286 & ~n41544;
  assign po1592 = n43989 | n43990;
  assign n43992 = ~n42965 & n43913;
  assign n43993 = pi1287 & ~n43913;
  assign n43994 = ~n43992 & ~n43993;
  assign n43995 = n41544 & ~n43994;
  assign n43996 = pi1287 & ~n41544;
  assign po1593 = n43995 | n43996;
  assign n43998 = n42801 & n43402;
  assign n43999 = ~n42809 & n43998;
  assign n44000 = pi1288 & ~n43998;
  assign n44001 = ~n43999 & ~n44000;
  assign n44002 = n41544 & ~n44001;
  assign n44003 = pi1288 & ~n41544;
  assign po1594 = n44002 | n44003;
  assign n44005 = ~n42821 & n43998;
  assign n44006 = pi1289 & ~n43998;
  assign n44007 = ~n44005 & ~n44006;
  assign n44008 = n41544 & ~n44007;
  assign n44009 = pi1289 & ~n41544;
  assign po1595 = n44008 | n44009;
  assign n44011 = ~n42833 & n43998;
  assign n44012 = pi1290 & ~n43998;
  assign n44013 = ~n44011 & ~n44012;
  assign n44014 = n41544 & ~n44013;
  assign n44015 = pi1290 & ~n41544;
  assign po1596 = n44014 | n44015;
  assign n44017 = ~n42845 & n43998;
  assign n44018 = pi1291 & ~n43998;
  assign n44019 = ~n44017 & ~n44018;
  assign n44020 = n41544 & ~n44019;
  assign n44021 = pi1291 & ~n41544;
  assign po1597 = n44020 | n44021;
  assign n44023 = ~n42857 & n43998;
  assign n44024 = pi1292 & ~n43998;
  assign n44025 = ~n44023 & ~n44024;
  assign n44026 = n41544 & ~n44025;
  assign n44027 = pi1292 & ~n41544;
  assign po1598 = n44026 | n44027;
  assign n44029 = ~n42869 & n43998;
  assign n44030 = pi1293 & ~n43998;
  assign n44031 = ~n44029 & ~n44030;
  assign n44032 = n41544 & ~n44031;
  assign n44033 = pi1293 & ~n41544;
  assign po1599 = n44032 | n44033;
  assign n44035 = ~n42881 & n43998;
  assign n44036 = pi1294 & ~n43998;
  assign n44037 = ~n44035 & ~n44036;
  assign n44038 = n41544 & ~n44037;
  assign n44039 = pi1294 & ~n41544;
  assign po1600 = n44038 | n44039;
  assign n44041 = ~n42893 & n43998;
  assign n44042 = pi1295 & ~n43998;
  assign n44043 = ~n44041 & ~n44042;
  assign n44044 = n41544 & ~n44043;
  assign n44045 = pi1295 & ~n41544;
  assign po1601 = n44044 | n44045;
  assign n44047 = ~n42905 & n43998;
  assign n44048 = pi1296 & ~n43998;
  assign n44049 = ~n44047 & ~n44048;
  assign n44050 = n41544 & ~n44049;
  assign n44051 = pi1296 & ~n41544;
  assign po1602 = n44050 | n44051;
  assign n44053 = ~n42917 & n43998;
  assign n44054 = pi1297 & ~n43998;
  assign n44055 = ~n44053 & ~n44054;
  assign n44056 = n41544 & ~n44055;
  assign n44057 = pi1297 & ~n41544;
  assign po1603 = n44056 | n44057;
  assign n44059 = ~n42929 & n43998;
  assign n44060 = pi1298 & ~n43998;
  assign n44061 = ~n44059 & ~n44060;
  assign n44062 = n41544 & ~n44061;
  assign n44063 = pi1298 & ~n41544;
  assign po1604 = n44062 | n44063;
  assign n44065 = ~n42941 & n43998;
  assign n44066 = pi1299 & ~n43998;
  assign n44067 = ~n44065 & ~n44066;
  assign n44068 = n41544 & ~n44067;
  assign n44069 = pi1299 & ~n41544;
  assign po1605 = n44068 | n44069;
  assign n44071 = ~n42953 & n43998;
  assign n44072 = pi1300 & ~n43998;
  assign n44073 = ~n44071 & ~n44072;
  assign n44074 = n41544 & ~n44073;
  assign n44075 = pi1300 & ~n41544;
  assign po1606 = n44074 | n44075;
  assign n44077 = ~n42965 & n43998;
  assign n44078 = pi1301 & ~n43998;
  assign n44079 = ~n44077 & ~n44078;
  assign n44080 = n41544 & ~n44079;
  assign n44081 = pi1301 & ~n41544;
  assign po1607 = n44080 | n44081;
  assign n44083 = n42972 & n43402;
  assign n44084 = ~n42809 & n44083;
  assign n44085 = pi1302 & ~n44083;
  assign n44086 = ~n44084 & ~n44085;
  assign n44087 = n41544 & ~n44086;
  assign n44088 = pi1302 & ~n41544;
  assign po1608 = n44087 | n44088;
  assign n44090 = ~n42821 & n44083;
  assign n44091 = pi1303 & ~n44083;
  assign n44092 = ~n44090 & ~n44091;
  assign n44093 = n41544 & ~n44092;
  assign n44094 = pi1303 & ~n41544;
  assign po1609 = n44093 | n44094;
  assign n44096 = ~n42833 & n44083;
  assign n44097 = pi1304 & ~n44083;
  assign n44098 = ~n44096 & ~n44097;
  assign n44099 = n41544 & ~n44098;
  assign n44100 = pi1304 & ~n41544;
  assign po1610 = n44099 | n44100;
  assign n44102 = ~n42845 & n44083;
  assign n44103 = pi1305 & ~n44083;
  assign n44104 = ~n44102 & ~n44103;
  assign n44105 = n41544 & ~n44104;
  assign n44106 = pi1305 & ~n41544;
  assign po1611 = n44105 | n44106;
  assign n44108 = ~n42857 & n44083;
  assign n44109 = pi1306 & ~n44083;
  assign n44110 = ~n44108 & ~n44109;
  assign n44111 = n41544 & ~n44110;
  assign n44112 = pi1306 & ~n41544;
  assign po1612 = n44111 | n44112;
  assign n44114 = ~n42869 & n44083;
  assign n44115 = pi1307 & ~n44083;
  assign n44116 = ~n44114 & ~n44115;
  assign n44117 = n41544 & ~n44116;
  assign n44118 = pi1307 & ~n41544;
  assign po1613 = n44117 | n44118;
  assign n44120 = ~n42881 & n44083;
  assign n44121 = pi1308 & ~n44083;
  assign n44122 = ~n44120 & ~n44121;
  assign n44123 = n41544 & ~n44122;
  assign n44124 = pi1308 & ~n41544;
  assign po1614 = n44123 | n44124;
  assign n44126 = ~n42893 & n44083;
  assign n44127 = pi1309 & ~n44083;
  assign n44128 = ~n44126 & ~n44127;
  assign n44129 = n41544 & ~n44128;
  assign n44130 = pi1309 & ~n41544;
  assign po1615 = n44129 | n44130;
  assign n44132 = ~n42905 & n44083;
  assign n44133 = pi1310 & ~n44083;
  assign n44134 = ~n44132 & ~n44133;
  assign n44135 = n41544 & ~n44134;
  assign n44136 = pi1310 & ~n41544;
  assign po1616 = n44135 | n44136;
  assign n44138 = ~n42917 & n44083;
  assign n44139 = pi1311 & ~n44083;
  assign n44140 = ~n44138 & ~n44139;
  assign n44141 = n41544 & ~n44140;
  assign n44142 = pi1311 & ~n41544;
  assign po1617 = n44141 | n44142;
  assign n44144 = ~n42929 & n44083;
  assign n44145 = pi1312 & ~n44083;
  assign n44146 = ~n44144 & ~n44145;
  assign n44147 = n41544 & ~n44146;
  assign n44148 = pi1312 & ~n41544;
  assign po1618 = n44147 | n44148;
  assign n44150 = ~n42941 & n44083;
  assign n44151 = pi1313 & ~n44083;
  assign n44152 = ~n44150 & ~n44151;
  assign n44153 = n41544 & ~n44152;
  assign n44154 = pi1313 & ~n41544;
  assign po1619 = n44153 | n44154;
  assign n44156 = ~n42953 & n44083;
  assign n44157 = pi1314 & ~n44083;
  assign n44158 = ~n44156 & ~n44157;
  assign n44159 = n41544 & ~n44158;
  assign n44160 = pi1314 & ~n41544;
  assign po1620 = n44159 | n44160;
  assign n44162 = ~n42965 & n44083;
  assign n44163 = pi1315 & ~n44083;
  assign n44164 = ~n44162 & ~n44163;
  assign n44165 = n41544 & ~n44164;
  assign n44166 = pi1315 & ~n41544;
  assign po1621 = n44165 | n44166;
  assign n44168 = n42802 & n43145;
  assign n44169 = ~n42809 & n44168;
  assign n44170 = pi1316 & ~n44168;
  assign n44171 = ~n44169 & ~n44170;
  assign n44172 = n41544 & ~n44171;
  assign n44173 = pi1316 & ~n41544;
  assign po1622 = n44172 | n44173;
  assign n44175 = ~n42821 & n44168;
  assign n44176 = pi1317 & ~n44168;
  assign n44177 = ~n44175 & ~n44176;
  assign n44178 = n41544 & ~n44177;
  assign n44179 = pi1317 & ~n41544;
  assign po1623 = n44178 | n44179;
  assign n44181 = ~n42833 & n44168;
  assign n44182 = pi1318 & ~n44168;
  assign n44183 = ~n44181 & ~n44182;
  assign n44184 = n41544 & ~n44183;
  assign n44185 = pi1318 & ~n41544;
  assign po1624 = n44184 | n44185;
  assign n44187 = ~n42845 & n44168;
  assign n44188 = pi1319 & ~n44168;
  assign n44189 = ~n44187 & ~n44188;
  assign n44190 = n41544 & ~n44189;
  assign n44191 = pi1319 & ~n41544;
  assign po1625 = n44190 | n44191;
  assign n44193 = ~n42857 & n44168;
  assign n44194 = pi1320 & ~n44168;
  assign n44195 = ~n44193 & ~n44194;
  assign n44196 = n41544 & ~n44195;
  assign n44197 = pi1320 & ~n41544;
  assign po1626 = n44196 | n44197;
  assign n44199 = ~n42869 & n44168;
  assign n44200 = pi1321 & ~n44168;
  assign n44201 = ~n44199 & ~n44200;
  assign n44202 = n41544 & ~n44201;
  assign n44203 = pi1321 & ~n41544;
  assign po1627 = n44202 | n44203;
  assign n44205 = ~n42881 & n44168;
  assign n44206 = pi1322 & ~n44168;
  assign n44207 = ~n44205 & ~n44206;
  assign n44208 = n41544 & ~n44207;
  assign n44209 = pi1322 & ~n41544;
  assign po1628 = n44208 | n44209;
  assign n44211 = ~n42893 & n44168;
  assign n44212 = pi1323 & ~n44168;
  assign n44213 = ~n44211 & ~n44212;
  assign n44214 = n41544 & ~n44213;
  assign n44215 = pi1323 & ~n41544;
  assign po1629 = n44214 | n44215;
  assign n44217 = ~n42905 & n44168;
  assign n44218 = pi1324 & ~n44168;
  assign n44219 = ~n44217 & ~n44218;
  assign n44220 = n41544 & ~n44219;
  assign n44221 = pi1324 & ~n41544;
  assign po1630 = n44220 | n44221;
  assign n44223 = ~n42917 & n44168;
  assign n44224 = pi1325 & ~n44168;
  assign n44225 = ~n44223 & ~n44224;
  assign n44226 = n41544 & ~n44225;
  assign n44227 = pi1325 & ~n41544;
  assign po1631 = n44226 | n44227;
  assign n44229 = ~n42929 & n44168;
  assign n44230 = pi1326 & ~n44168;
  assign n44231 = ~n44229 & ~n44230;
  assign n44232 = n41544 & ~n44231;
  assign n44233 = pi1326 & ~n41544;
  assign po1632 = n44232 | n44233;
  assign n44235 = ~n42941 & n44168;
  assign n44236 = pi1327 & ~n44168;
  assign n44237 = ~n44235 & ~n44236;
  assign n44238 = n41544 & ~n44237;
  assign n44239 = pi1327 & ~n41544;
  assign po1633 = n44238 | n44239;
  assign n44241 = ~n42953 & n44168;
  assign n44242 = pi1328 & ~n44168;
  assign n44243 = ~n44241 & ~n44242;
  assign n44244 = n41544 & ~n44243;
  assign n44245 = pi1328 & ~n41544;
  assign po1634 = n44244 | n44245;
  assign n44247 = ~n42965 & n44168;
  assign n44248 = pi1329 & ~n44168;
  assign n44249 = ~n44247 & ~n44248;
  assign n44250 = n41544 & ~n44249;
  assign n44251 = pi1329 & ~n41544;
  assign po1635 = n44250 | n44251;
  assign n44253 = ~n38238 & ~n38248;
  assign n44254 = ~n38227 & ~n38235;
  assign n44255 = ~n38246 & n44254;
  assign n44256 = n44253 & n44255;
  assign n44257 = n38229 & n44256;
  assign n44258 = n38262 & n44257;
  assign n44259 = n38243 & n44258;
  assign n44260 = n38255 & n44259;
  assign n44261 = pi1330 & ~n38262;
  assign po1636 = n44260 | n44261;
  assign n44263 = n36060 & n36114;
  assign n44264 = pi1331 & n36128;
  assign po1637 = n44263 | n44264;
  assign n44266 = pi1332 & n8561;
  assign n44267 = ~n8561 & n39108;
  assign po1638 = n44266 | n44267;
  assign n44269 = pi1333 & n8561;
  assign n44270 = ~n8561 & n39109;
  assign po1639 = n44269 | n44270;
  assign n44272 = pi1334 & n8561;
  assign n44273 = ~n8561 & n37748;
  assign po1640 = n44272 | n44273;
  assign n44275 = ~n8561 & n39106;
  assign n44276 = pi1335 & n8561;
  assign po1641 = n44275 | n44276;
  assign n44278 = ~n8561 & n39107;
  assign n44279 = pi1336 & n8561;
  assign po1642 = n44278 | n44279;
  assign n44281 = pi1337 & n8561;
  assign n44282 = ~n8561 & n38600;
  assign po1643 = n44281 | n44282;
  assign n44284 = pi1338 & n8561;
  assign n44285 = ~n8561 & n38603;
  assign po1644 = n44284 | n44285;
  assign n44287 = pi1339 & n8561;
  assign n44288 = ~n8561 & n38598;
  assign po1645 = n44287 | n44288;
  assign n44290 = pi1340 & n8561;
  assign n44291 = ~n8561 & n36026;
  assign po1646 = n44290 | n44291;
  assign n44293 = pi1341 & n8561;
  assign n44294 = ~n8561 & n36025;
  assign po1647 = n44293 | n44294;
  assign n44296 = pi1342 & n8561;
  assign n44297 = ~n8561 & n36029;
  assign po1648 = n44296 | n44297;
  assign n44299 = pi1343 & n8561;
  assign n44300 = ~n8561 & n36033;
  assign po1649 = n44299 | n44300;
  assign n44302 = ~n8561 & n37742;
  assign n44303 = pi1344 & n8561;
  assign po1650 = n44302 | n44303;
  assign n44305 = pi1345 & n8561;
  assign n44306 = ~n8561 & n38621;
  assign po1651 = n44305 | n44306;
  assign n44308 = ~n8561 & n38623;
  assign n44309 = pi1346 & n8561;
  assign po1652 = n44308 | n44309;
  assign n44311 = pi1347 & n8561;
  assign n44312 = ~n8561 & n38620;
  assign po1653 = n44311 | n44312;
  assign n44314 = ~n8561 & n38624;
  assign n44315 = pi1348 & n8561;
  assign po1654 = n44314 | n44315;
  assign n44317 = ~n8561 & n36038;
  assign n44318 = pi1349 & n8561;
  assign po1655 = n44317 | n44318;
  assign n44320 = pi1350 & n8561;
  assign n44321 = ~n8561 & n38610;
  assign po1656 = n44320 | n44321;
  assign n44323 = pi1351 & n8561;
  assign n44324 = ~n8561 & n38611;
  assign po1657 = n44323 | n44324;
  assign n44326 = pi1352 & n8561;
  assign n44327 = ~n8561 & n38615;
  assign po1658 = n44326 | n44327;
  assign n44329 = ~n8561 & n38613;
  assign n44330 = pi1353 & n8561;
  assign po1659 = n44329 | n44330;
  assign n44332 = pi1354 & n8561;
  assign n44333 = ~n8561 & n36014;
  assign po1660 = n44332 | n44333;
  assign n44335 = pi1355 & n8561;
  assign n44336 = ~n8561 & n36017;
  assign po1661 = n44335 | n44336;
  assign n44338 = pi1356 & n8561;
  assign n44339 = ~n8561 & n36050;
  assign po1662 = n44338 | n44339;
  assign n44341 = pi1357 & n8561;
  assign n44342 = ~n8561 & n36051;
  assign po1663 = n44341 | n44342;
  assign n44344 = ~n8561 & n37744;
  assign n44345 = pi1358 & n8561;
  assign po1664 = n44344 | n44345;
  assign n44347 = ~n8561 & n37730;
  assign n44348 = pi1359 & n8561;
  assign po1665 = n44347 | n44348;
  assign n44350 = pi1360 & n8561;
  assign n44351 = ~n8561 & n36539;
  assign po1666 = n44350 | n44351;
  assign n44353 = ~pi1361 & ~n41779;
  assign n44354 = pi1361 & n41783;
  assign n44355 = ~pi1361 & ~n41783;
  assign n44356 = ~n44354 & ~n44355;
  assign n44357 = n41779 & ~n44356;
  assign po1667 = n44353 | n44357;
  assign n44359 = n42465 & n42500;
  assign n44360 = pi1362 & n44359;
  assign n44361 = ~pi1362 & ~n44359;
  assign n44362 = ~n44360 & ~n44361;
  assign n44363 = n41809 & ~n44362;
  assign n44364 = ~pi1362 & ~n41809;
  assign po1668 = n44363 | n44364;
  assign n44366 = n42483 & n42488;
  assign n44367 = ~pi1363 & ~n44366;
  assign n44368 = pi1363 & n44366;
  assign n44369 = ~n44367 & ~n44368;
  assign n44370 = n41809 & ~n44369;
  assign n44371 = ~pi1363 & ~n41809;
  assign po1669 = n44370 | n44371;
  assign n44373 = n42466 & n44359;
  assign n44374 = pi1364 & n44373;
  assign n44375 = ~pi1364 & ~n44373;
  assign n44376 = ~n44374 & ~n44375;
  assign n44377 = n41809 & ~n44376;
  assign n44378 = ~pi1364 & ~n41809;
  assign po1670 = n44377 | n44378;
  assign n44380 = n42512 & n42605;
  assign n44381 = n42607 & n44380;
  assign n44382 = pi1365 & n44381;
  assign n44383 = ~pi1365 & ~n44381;
  assign n44384 = ~n44382 & ~n44383;
  assign n44385 = n41809 & ~n44384;
  assign n44386 = ~pi1365 & ~n41809;
  assign po1671 = n44385 | n44386;
  assign n44388 = n42512 & n42610;
  assign n44389 = ~pi1366 & ~n44388;
  assign n44390 = pi1366 & n44388;
  assign n44391 = ~n44389 & ~n44390;
  assign n44392 = n41809 & ~n44391;
  assign n44393 = ~pi1366 & ~n41809;
  assign po1672 = n44392 | n44393;
  assign n44395 = ~pi1367 & ~n41793;
  assign n44396 = pi1367 & n41793;
  assign n44397 = ~n44395 & ~n44396;
  assign n44398 = n41809 & ~n44397;
  assign n44399 = ~pi1367 & ~n41809;
  assign po1673 = n44398 | n44399;
  assign n44401 = ~pi1368 & ~n42500;
  assign n44402 = pi1368 & n42500;
  assign n44403 = ~n44401 & ~n44402;
  assign n44404 = n41809 & ~n44403;
  assign n44405 = ~pi1368 & ~n41809;
  assign po1674 = n44404 | n44405;
  assign n44407 = pi1369 & n41799;
  assign n44408 = ~pi1369 & ~n41799;
  assign n44409 = ~n44407 & ~n44408;
  assign n44410 = n41809 & ~n44409;
  assign n44411 = ~pi1369 & ~n41809;
  assign po1675 = n44410 | n44411;
  assign n44413 = ~pi1370 & ~pi3641;
  assign n44414 = pi3641 & ~n37404;
  assign n44415 = ~n44413 & ~n44414;
  assign n44416 = n37393 & ~n44415;
  assign n44417 = pi1430 & ~n37393;
  assign po1676 = n44416 | n44417;
  assign n44419 = ~pi1104 & ~pi1373;
  assign n44420 = ~pi1372 & n44419;
  assign n44421 = ~pi1388 & n44420;
  assign n44422 = ~pi1371 & ~n44421;
  assign n44423 = pi1371 & n44421;
  assign n44424 = ~n44422 & ~n44423;
  assign n44425 = n42790 & ~n44424;
  assign n44426 = ~pi0893 & ~n42790;
  assign n44427 = ~n44425 & ~n44426;
  assign po1677 = pi1685 & n44427;
  assign n44429 = pi1372 & ~n44419;
  assign n44430 = ~n44420 & ~n44429;
  assign n44431 = n42790 & n44430;
  assign n44432 = ~pi0885 & ~n42790;
  assign n44433 = ~n44431 & ~n44432;
  assign po1678 = ~pi1685 | n44433;
  assign n44435 = pi1373 & n42790;
  assign n44436 = ~pi0741 & ~n42790;
  assign n44437 = ~n44435 & ~n44436;
  assign po1679 = ~pi1685 | n44437;
  assign n44439 = ~pi1377 & ~pi1389;
  assign n44440 = ~pi1376 & n44439;
  assign n44441 = ~pi1375 & n44440;
  assign n44442 = ~pi1374 & ~n44441;
  assign n44443 = pi1374 & n44441;
  assign n44444 = ~n44442 & ~n44443;
  assign n44445 = pi2509 & ~pi2993;
  assign n44446 = ~pi3554 & n44445;
  assign n44447 = ~pi2509 & ~pi2993;
  assign n44448 = pi3554 & n44447;
  assign n44449 = ~pi2509 & pi2993;
  assign n44450 = ~pi3554 & n44449;
  assign n44451 = ~n44448 & ~n44450;
  assign n44452 = ~n44446 & n44451;
  assign n44453 = pi0792 & po0034;
  assign n44454 = ~pi0792 & pi3669;
  assign n44455 = ~n44453 & ~n44454;
  assign n44456 = ~pi0956 & ~n44455;
  assign n44457 = pi0956 & n44455;
  assign po3943 = n44456 | n44457;
  assign n44459 = pi3636 & po3943;
  assign po3937 = pi3635 & n44459;
  assign n44461 = n35387 & ~po3937;
  assign n44462 = ~pi3630 & n35397;
  assign n44463 = pi3629 & n35399;
  assign n44464 = pi3628 & ~n35399;
  assign n44465 = ~n44463 & ~n44464;
  assign n44466 = ~n35397 & n44465;
  assign n44467 = ~n44462 & ~n44466;
  assign n44468 = ~n35387 & ~n44467;
  assign n44469 = ~n44461 & ~n44468;
  assign n44470 = n44446 & ~n44469;
  assign n44471 = ~n44452 & ~n44470;
  assign n44472 = ~pi1376 & ~pi1389;
  assign n44473 = ~pi1375 & n44472;
  assign n44474 = ~pi1374 & n44473;
  assign n44475 = ~pi1377 & n44474;
  assign n44476 = n44448 & n44475;
  assign n44477 = ~pi1629 & ~pi1687;
  assign n44478 = ~pi1848 & ~pi1849;
  assign n44479 = pi1608 & pi1644;
  assign n44480 = pi1648 & n44479;
  assign n44481 = pi1686 & n44480;
  assign n44482 = n44478 & n44481;
  assign n44483 = n44477 & n44482;
  assign n44484 = n44476 & n44483;
  assign po2824 = ~n44471 | n44484;
  assign po3311 = n44476 & ~n44483;
  assign n44487 = ~po2824 & ~po3311;
  assign n44488 = ~n44444 & n44487;
  assign n44489 = ~pi0799 & ~n44487;
  assign n44490 = ~n44488 & ~n44489;
  assign po1680 = pi1688 & n44490;
  assign n44492 = pi1375 & ~n44440;
  assign n44493 = ~n44441 & ~n44492;
  assign n44494 = n44487 & n44493;
  assign n44495 = ~pi0957 & ~n44487;
  assign n44496 = ~n44494 & ~n44495;
  assign po1681 = ~pi1688 | n44496;
  assign n44498 = pi1376 & ~n44439;
  assign n44499 = ~n44440 & ~n44498;
  assign n44500 = n44487 & n44499;
  assign n44501 = ~pi1009 & ~n44487;
  assign n44502 = ~n44500 & ~n44501;
  assign po1682 = ~pi1688 | n44502;
  assign n44504 = pi1377 & n44487;
  assign n44505 = ~pi0795 & ~n44487;
  assign n44506 = ~n44504 & ~n44505;
  assign po1683 = ~pi1688 | n44506;
  assign n44508 = ~pi1689 & ~pi1690;
  assign n44509 = ~pi1646 & ~pi1850;
  assign n44510 = ~pi1694 & n44509;
  assign n44511 = ~pi1643 & n44510;
  assign n44512 = ~pi1691 & n44511;
  assign n44513 = ~pi1692 & n44512;
  assign n44514 = ~pi1693 & n44513;
  assign n44515 = ~pi1649 & n44514;
  assign n44516 = n44508 & n44515;
  assign n44517 = ~pi1378 & n44516;
  assign n44518 = pi1378 & ~n44516;
  assign n44519 = ~n44517 & ~n44518;
  assign n44520 = pi1691 & pi1834;
  assign n44521 = ~pi1691 & ~pi1834;
  assign n44522 = ~n44520 & ~n44521;
  assign n44523 = pi1643 & pi1839;
  assign n44524 = ~pi1643 & ~pi1839;
  assign n44525 = ~n44523 & ~n44524;
  assign n44526 = pi1692 & pi1853;
  assign n44527 = ~pi1692 & ~pi1853;
  assign n44528 = ~n44526 & ~n44527;
  assign n44529 = pi1693 & pi1852;
  assign n44530 = ~pi1693 & ~pi1852;
  assign n44531 = ~n44529 & ~n44530;
  assign n44532 = n44528 & n44531;
  assign n44533 = n44525 & n44532;
  assign n44534 = n44522 & n44533;
  assign n44535 = pi1690 & pi1832;
  assign n44536 = ~pi1690 & ~pi1832;
  assign n44537 = ~n44535 & ~n44536;
  assign n44538 = n44534 & n44537;
  assign n44539 = ~pi1649 & ~pi1833;
  assign n44540 = pi1649 & pi1833;
  assign n44541 = ~n44539 & ~n44540;
  assign n44542 = ~pi1689 & ~pi1831;
  assign n44543 = pi1689 & pi1831;
  assign n44544 = ~n44542 & ~n44543;
  assign n44545 = pi1378 & ~pi1830;
  assign n44546 = ~pi1378 & pi1830;
  assign n44547 = ~n44545 & ~n44546;
  assign n44548 = n44544 & ~n44547;
  assign n44549 = n44541 & n44548;
  assign n44550 = n44538 & n44549;
  assign po1684 = n44519 & ~n44550;
  assign n44552 = ~pi1379 & ~n42536;
  assign n44553 = ~pi1668 & ~pi1695;
  assign n44554 = n42541 & n44553;
  assign n44555 = ~pi1851 & ~pi2416;
  assign n44556 = n41248 & n44555;
  assign n44557 = n44554 & n44556;
  assign n44558 = pi1379 & n44557;
  assign n44559 = ~pi1379 & ~n44557;
  assign n44560 = ~n44558 & ~n44559;
  assign n44561 = n42536 & ~n44560;
  assign po1685 = n44552 | n44561;
  assign n44563 = ~pi1380 & ~n42536;
  assign n44564 = n41248 & n44553;
  assign n44565 = n44555 & n44564;
  assign n44566 = pi1380 & n44565;
  assign n44567 = ~pi1380 & ~n44565;
  assign n44568 = ~n44566 & ~n44567;
  assign n44569 = n42536 & ~n44568;
  assign po1686 = n44563 | n44569;
  assign n44571 = ~pi1381 & ~n44380;
  assign n44572 = pi1381 & n44380;
  assign n44573 = ~n44571 & ~n44572;
  assign n44574 = n41809 & ~n44573;
  assign n44575 = ~pi1381 & ~n41809;
  assign po1687 = n44574 | n44575;
  assign n44577 = pi1075 & ~pi1382;
  assign n44578 = ~pi1075 & pi1382;
  assign n44579 = ~n44577 & ~n44578;
  assign n44580 = n41809 & ~n44579;
  assign n44581 = ~pi1382 & ~n41809;
  assign po1688 = n44580 | n44581;
  assign n44583 = pi1383 & n41795;
  assign n44584 = ~pi1383 & ~n41795;
  assign n44585 = ~n44583 & ~n44584;
  assign n44586 = n41809 & ~n44585;
  assign n44587 = ~pi1383 & ~n41809;
  assign po1689 = n44586 | n44587;
  assign n44589 = pi1384 & n41794;
  assign n44590 = ~pi1384 & ~n41794;
  assign n44591 = ~n44589 & ~n44590;
  assign n44592 = n41809 & ~n44591;
  assign n44593 = ~pi1384 & ~n41809;
  assign po1690 = n44592 | n44593;
  assign n44595 = n42486 & n44366;
  assign n44596 = pi1385 & n44595;
  assign n44597 = ~pi1385 & ~n44595;
  assign n44598 = ~n44596 & ~n44597;
  assign n44599 = n41809 & ~n44598;
  assign n44600 = ~pi1385 & ~n41809;
  assign po1691 = n44599 | n44600;
  assign n44602 = pi1386 & n41800;
  assign n44603 = ~pi1386 & ~n41800;
  assign n44604 = ~n44602 & ~n44603;
  assign n44605 = n41809 & ~n44604;
  assign n44606 = ~pi1386 & ~n41809;
  assign po1692 = n44605 | n44606;
  assign n44608 = ~pi1387 & ~n41779;
  assign n44609 = n42439 & n42449;
  assign n44610 = n42437 & n44609;
  assign n44611 = pi1387 & n44610;
  assign n44612 = ~pi1387 & ~n44610;
  assign n44613 = ~n44611 & ~n44612;
  assign n44614 = n41779 & ~n44613;
  assign po1693 = n44608 | n44614;
  assign n44616 = pi1388 & ~n44420;
  assign n44617 = ~n44421 & ~n44616;
  assign n44618 = n42790 & n44617;
  assign n44619 = ~pi0884 & ~n42790;
  assign n44620 = ~n44618 & ~n44619;
  assign po1694 = ~pi1685 | n44620;
  assign n44622 = pi1377 & ~pi1389;
  assign n44623 = ~pi1377 & pi1389;
  assign n44624 = ~n44622 & ~n44623;
  assign n44625 = n44487 & ~n44624;
  assign n44626 = ~pi0793 & ~n44487;
  assign n44627 = ~n44625 & ~n44626;
  assign po1695 = ~pi1688 | n44627;
  assign n44629 = ~pi1390 & ~n42185;
  assign n44630 = ~pi1042 & ~n42675;
  assign n44631 = ~n42189 & n44630;
  assign n44632 = pi1390 & ~n44631;
  assign n44633 = ~pi0828 & n44631;
  assign n44634 = ~n44632 & ~n44633;
  assign n44635 = n42185 & n44634;
  assign po1696 = n44629 | n44635;
  assign n44637 = ~pi1391 & ~n42185;
  assign n44638 = n42189 & n44630;
  assign n44639 = pi0827 & n44638;
  assign n44640 = ~pi1391 & ~n44638;
  assign n44641 = ~n44639 & ~n44640;
  assign n44642 = n42185 & ~n44641;
  assign po1697 = n44637 | n44642;
  assign n44644 = ~pi1392 & ~n42185;
  assign n44645 = pi1042 & n42675;
  assign n44646 = n42189 & n44645;
  assign n44647 = pi0979 & n44646;
  assign n44648 = ~pi1392 & ~n44646;
  assign n44649 = ~n44647 & ~n44648;
  assign n44650 = n42185 & ~n44649;
  assign po1698 = n44644 | n44650;
  assign n44652 = ~pi1393 & ~n42185;
  assign n44653 = ~pi1042 & n42675;
  assign n44654 = n42189 & n44653;
  assign n44655 = pi0918 & n44654;
  assign n44656 = ~pi1393 & ~n44654;
  assign n44657 = ~n44655 & ~n44656;
  assign n44658 = n42185 & ~n44657;
  assign po1699 = n44652 | n44658;
  assign n44660 = ~pi1394 & ~n42185;
  assign n44661 = pi0659 & n44646;
  assign n44662 = ~pi1394 & ~n44646;
  assign n44663 = ~n44661 & ~n44662;
  assign n44664 = n42185 & ~n44663;
  assign po1700 = n44660 | n44664;
  assign n44666 = ~pi1395 & ~n42185;
  assign n44667 = ~n42189 & n44653;
  assign n44668 = pi1395 & ~n44667;
  assign n44669 = ~pi0916 & n44667;
  assign n44670 = ~n44668 & ~n44669;
  assign n44671 = n42185 & n44670;
  assign po1701 = n44666 | n44671;
  assign n44673 = ~pi1396 & ~n42185;
  assign n44674 = pi1396 & ~n44631;
  assign n44675 = ~pi0980 & n44631;
  assign n44676 = ~n44674 & ~n44675;
  assign n44677 = n42185 & n44676;
  assign po1702 = n44673 | n44677;
  assign n44679 = ~pi1397 & ~n42185;
  assign n44680 = pi1397 & ~n44631;
  assign n44681 = ~pi0917 & n44631;
  assign n44682 = ~n44680 & ~n44681;
  assign n44683 = n42185 & n44682;
  assign po1703 = n44679 | n44683;
  assign n44685 = ~pi1398 & ~n42185;
  assign n44686 = pi1398 & ~n44631;
  assign n44687 = ~pi0916 & n44631;
  assign n44688 = ~n44686 & ~n44687;
  assign n44689 = n42185 & n44688;
  assign po1704 = n44685 | n44689;
  assign n44691 = ~pi1399 & ~n42185;
  assign n44692 = pi0828 & n44638;
  assign n44693 = ~pi1399 & ~n44638;
  assign n44694 = ~n44692 & ~n44693;
  assign n44695 = n42185 & ~n44694;
  assign po1705 = n44691 | n44695;
  assign n44697 = ~pi1400 & ~n42185;
  assign n44698 = pi1400 & ~n44631;
  assign n44699 = ~pi0914 & n44631;
  assign n44700 = ~n44698 & ~n44699;
  assign n44701 = n42185 & n44700;
  assign po1706 = n44697 | n44701;
  assign n44703 = ~pi1401 & ~n42185;
  assign n44704 = pi0828 & n44654;
  assign n44705 = ~pi1401 & ~n44654;
  assign n44706 = ~n44704 & ~n44705;
  assign n44707 = n42185 & ~n44706;
  assign po1707 = n44703 | n44707;
  assign n44709 = ~pi1402 & ~n42185;
  assign n44710 = pi1402 & ~n44631;
  assign n44711 = ~pi0586 & n44631;
  assign n44712 = ~n44710 & ~n44711;
  assign n44713 = n42185 & n44712;
  assign po1708 = n44709 | n44713;
  assign n44715 = ~pi1403 & ~n42185;
  assign n44716 = pi0980 & n44638;
  assign n44717 = ~pi1403 & ~n44638;
  assign n44718 = ~n44716 & ~n44717;
  assign n44719 = n42185 & ~n44718;
  assign po1709 = n44715 | n44719;
  assign n44721 = ~pi1404 & ~n42185;
  assign n44722 = pi0914 & n44638;
  assign n44723 = ~pi1404 & ~n44638;
  assign n44724 = ~n44722 & ~n44723;
  assign n44725 = n42185 & ~n44724;
  assign po1710 = n44721 | n44725;
  assign n44727 = ~pi1405 & ~n42185;
  assign n44728 = pi0917 & n44638;
  assign n44729 = ~pi1405 & ~n44638;
  assign n44730 = ~n44728 & ~n44729;
  assign n44731 = n42185 & ~n44730;
  assign po1711 = n44727 | n44731;
  assign n44733 = ~pi1406 & ~n42185;
  assign n44734 = pi1406 & ~n44631;
  assign n44735 = ~pi0196 & n44631;
  assign n44736 = ~n44734 & ~n44735;
  assign n44737 = n42185 & n44736;
  assign po1712 = n44733 | n44737;
  assign n44739 = ~pi1407 & ~n42185;
  assign n44740 = n42189 & ~n42675;
  assign n44741 = pi1042 & n44740;
  assign n44742 = ~pi3633 & n44741;
  assign n44743 = ~pi1407 & ~n44741;
  assign n44744 = ~n44742 & ~n44743;
  assign n44745 = n42185 & ~n44744;
  assign po1713 = n44739 | n44745;
  assign n44747 = ~pi1408 & ~n42185;
  assign n44748 = pi0912 & n44638;
  assign n44749 = ~pi1408 & ~n44638;
  assign n44750 = ~n44748 & ~n44749;
  assign n44751 = n42185 & ~n44750;
  assign po1714 = n44747 | n44751;
  assign n44753 = ~pi1409 & ~n42185;
  assign n44754 = pi0196 & n44638;
  assign n44755 = ~pi1409 & ~n44638;
  assign n44756 = ~n44754 & ~n44755;
  assign n44757 = n42185 & ~n44756;
  assign po1715 = n44753 | n44757;
  assign n44759 = ~pi1410 & ~n42185;
  assign n44760 = pi0586 & n44638;
  assign n44761 = ~pi1410 & ~n44638;
  assign n44762 = ~n44760 & ~n44761;
  assign n44763 = n42185 & ~n44762;
  assign po1716 = n44759 | n44763;
  assign n44765 = ~pi1411 & ~n42185;
  assign n44766 = pi0826 & n44741;
  assign n44767 = ~pi1411 & ~n44741;
  assign n44768 = ~n44766 & ~n44767;
  assign n44769 = n42185 & ~n44768;
  assign po1717 = n44765 | n44769;
  assign n44771 = ~pi1412 & ~n42185;
  assign n44772 = pi0829 & n44741;
  assign n44773 = ~pi1412 & ~n44741;
  assign n44774 = ~n44772 & ~n44773;
  assign n44775 = n42185 & ~n44774;
  assign po1718 = n44771 | n44775;
  assign n44777 = ~pi1413 & ~n42185;
  assign n44778 = pi0868 & n44741;
  assign n44779 = ~pi1413 & ~n44741;
  assign n44780 = ~n44778 & ~n44779;
  assign n44781 = n42185 & ~n44780;
  assign po1719 = n44777 | n44781;
  assign n44783 = ~pi1414 & ~n42185;
  assign n44784 = pi0149 & n44654;
  assign n44785 = ~pi1414 & ~n44654;
  assign n44786 = ~n44784 & ~n44785;
  assign n44787 = n42185 & ~n44786;
  assign po1720 = n44783 | n44787;
  assign n44789 = ~pi1415 & ~n42185;
  assign n44790 = pi0708 & n44741;
  assign n44791 = ~pi1415 & ~n44741;
  assign n44792 = ~n44790 & ~n44791;
  assign n44793 = n42185 & ~n44792;
  assign po1721 = n44789 | n44793;
  assign n44795 = ~pi1416 & ~n42185;
  assign n44796 = pi0915 & n44741;
  assign n44797 = ~pi1416 & ~n44741;
  assign n44798 = ~n44796 & ~n44797;
  assign n44799 = n42185 & ~n44798;
  assign po1722 = n44795 | n44799;
  assign n44801 = ~pi1417 & ~n42185;
  assign n44802 = pi0152 & n44741;
  assign n44803 = ~pi1417 & ~n44741;
  assign n44804 = ~n44802 & ~n44803;
  assign n44805 = n42185 & ~n44804;
  assign po1723 = n44801 | n44805;
  assign n44807 = ~pi1418 & ~n25623;
  assign n44808 = pi0405 & pi0422;
  assign n44809 = n25623 & n44808;
  assign n44810 = n24807 & n25623;
  assign n44811 = pi0423 & pi0424;
  assign n44812 = n44810 & n44811;
  assign n44813 = ~n44809 & ~n44812;
  assign po1724 = n44807 | ~n44813;
  assign n44815 = ~pi1419 & ~n42185;
  assign n44816 = pi1419 & ~n44667;
  assign n44817 = ~pi0918 & n44667;
  assign n44818 = ~n44816 & ~n44817;
  assign n44819 = n42185 & n44818;
  assign po1725 = n44815 | n44819;
  assign n44821 = ~pi1420 & ~n42185;
  assign n44822 = pi1420 & ~n44667;
  assign n44823 = ~pi0149 & n44667;
  assign n44824 = ~n44822 & ~n44823;
  assign n44825 = n42185 & n44824;
  assign po1726 = n44821 | n44825;
  assign n44827 = ~pi1421 & ~n42185;
  assign n44828 = pi1421 & ~n44667;
  assign n44829 = ~pi0827 & n44667;
  assign n44830 = ~n44828 & ~n44829;
  assign n44831 = n42185 & n44830;
  assign po1727 = n44827 | n44831;
  assign n44833 = ~pi3579 & ~n17199;
  assign n44834 = ~pi3465 & pi3579;
  assign n44835 = ~n44833 & ~n44834;
  assign n44836 = n39505 & ~n44835;
  assign n44837 = pi1422 & ~n39505;
  assign po1728 = n44836 | n44837;
  assign n44839 = ~pi1423 & ~n42185;
  assign n44840 = pi0827 & n44654;
  assign n44841 = ~pi1423 & ~n44654;
  assign n44842 = ~n44840 & ~n44841;
  assign n44843 = n42185 & ~n44842;
  assign po1729 = n44839 | n44843;
  assign n44845 = ~pi1424 & ~n25623;
  assign po1730 = ~n44813 | n44845;
  assign n44847 = ~pi1425 & ~n25623;
  assign po1731 = ~n44813 | n44847;
  assign n44849 = pi1012 & pi1033;
  assign n44850 = ~pi1034 & n44849;
  assign n44851 = pi1039 & n44850;
  assign po3132 = n41522 & n44851;
  assign n44853 = pi0609 & po3132;
  assign n44854 = ~n17368 & n44853;
  assign n44855 = pi1426 & ~n44853;
  assign po1732 = n44854 | n44855;
  assign n44857 = ~n13121 & n44853;
  assign n44858 = pi1427 & ~n44853;
  assign po1733 = n44857 | n44858;
  assign n44860 = ~n13398 & n44853;
  assign n44861 = pi1428 & ~n44853;
  assign po1734 = n44860 | n44861;
  assign n44863 = ~n13988 & n44853;
  assign n44864 = pi1429 & ~n44853;
  assign po1735 = n44863 | n44864;
  assign n44866 = ~n12415 & n44853;
  assign n44867 = pi1430 & ~n44853;
  assign po1736 = n44866 | n44867;
  assign n44869 = ~n14816 & n44853;
  assign n44870 = pi1431 & ~n44853;
  assign po1737 = n44869 | n44870;
  assign n44872 = ~n15115 & n44853;
  assign n44873 = pi1432 & ~n44853;
  assign po1738 = n44872 | n44873;
  assign n44875 = ~n12061 & n44853;
  assign n44876 = pi1433 & ~n44853;
  assign po1739 = n44875 | n44876;
  assign n44878 = ~n11181 & n44853;
  assign n44879 = pi1434 & ~n44853;
  assign po1740 = n44878 | n44879;
  assign n44881 = pi1435 & ~n42691;
  assign n44882 = ~pi1435 & n42691;
  assign n44883 = ~n44881 & ~n44882;
  assign po1741 = n40651 & n44883;
  assign n44885 = n9644 & n41522;
  assign n44886 = pi0609 & n44885;
  assign n44887 = pi1436 & ~n44886;
  assign n44888 = ~n12726 & n44886;
  assign po1742 = n44887 | n44888;
  assign n44890 = pi1437 & ~n44886;
  assign n44891 = ~n13701 & n44886;
  assign po1743 = n44890 | n44891;
  assign n44893 = ~n13121 & n44886;
  assign n44894 = pi1438 & ~n44886;
  assign po1744 = n44893 | n44894;
  assign n44896 = ~n13398 & n44886;
  assign n44897 = pi1439 & ~n44886;
  assign po1745 = n44896 | n44897;
  assign n44899 = ~n13988 & n44886;
  assign n44900 = pi1440 & ~n44886;
  assign po1746 = n44899 | n44900;
  assign n44902 = ~n12415 & n44886;
  assign n44903 = pi1441 & ~n44886;
  assign po1747 = n44902 | n44903;
  assign n44905 = ~n14816 & n44886;
  assign n44906 = pi1442 & ~n44886;
  assign po1748 = n44905 | n44906;
  assign n44908 = ~n15115 & n44886;
  assign n44909 = pi1443 & ~n44886;
  assign po1749 = n44908 | n44909;
  assign n44911 = ~n12061 & n44886;
  assign n44912 = pi1444 & ~n44886;
  assign po1750 = n44911 | n44912;
  assign n44914 = pi1445 & ~n44886;
  assign n44915 = ~n15426 & n44886;
  assign po1751 = n44914 | n44915;
  assign n44917 = pi1446 & ~n44886;
  assign n44918 = ~n14403 & n44886;
  assign po1752 = n44917 | n44918;
  assign n44920 = ~n11181 & n44886;
  assign n44921 = pi1447 & ~n44886;
  assign po1753 = n44920 | n44921;
  assign n44923 = pi1448 & ~n42698;
  assign n44924 = ~pi1448 & n42698;
  assign n44925 = ~n44923 & ~n44924;
  assign po1754 = n40741 & n44925;
  assign n44927 = pi3651 & ~pi3652;
  assign po1755 = ~pi3529 | n44927;
  assign po1756 = ~pi3529 | ~n44927;
  assign n44930 = ~pi0876 & ~pi0904;
  assign n44931 = ~pi0902 & ~pi0903;
  assign n44932 = ~pi0820 & ~pi0910;
  assign n44933 = ~pi0819 & ~pi0909;
  assign n44934 = n44932 & n44933;
  assign n44935 = n44931 & n44934;
  assign n44936 = n44930 & n44935;
  assign n44937 = ~pi0908 & n44936;
  assign n44938 = ~pi0907 & n44937;
  assign n44939 = ~pi0873 & n44938;
  assign n44940 = ~pi0874 & n44939;
  assign n44941 = ~pi0905 & ~pi0906;
  assign n44942 = n32780 & n39530;
  assign n44943 = n44941 & n44942;
  assign n44944 = n44940 & n44943;
  assign po1757 = pi1449 & ~n44944;
  assign n44946 = ~n39498 & ~n41524;
  assign n44947 = ~n40745 & n44946;
  assign n44948 = pi1450 & ~n44946;
  assign po1758 = n44947 | n44948;
  assign n44950 = ~n40764 & n44946;
  assign n44951 = pi1451 & ~n44946;
  assign po1759 = n44950 | n44951;
  assign n44953 = ~n40489 & n44946;
  assign n44954 = pi1452 & ~n44946;
  assign po1760 = n44953 | n44954;
  assign n44956 = ~n40776 & n44946;
  assign n44957 = pi1453 & ~n44946;
  assign po1761 = n44956 | n44957;
  assign n44959 = ~n40788 & n44946;
  assign n44960 = pi1454 & ~n44946;
  assign po1762 = n44959 | n44960;
  assign n44962 = ~n40801 & n44946;
  assign n44963 = pi1455 & ~n44946;
  assign po1763 = n44962 | n44963;
  assign n44965 = ~n40450 & n44946;
  assign n44966 = pi1456 & ~n44946;
  assign po1764 = n44965 | n44966;
  assign n44968 = ~n40812 & n44946;
  assign n44969 = pi1457 & ~n44946;
  assign po1765 = n44968 | n44969;
  assign n44971 = ~n40830 & n44946;
  assign n44972 = pi1458 & ~n44946;
  assign po1766 = n44971 | n44972;
  assign n44974 = ~n39541 & n44946;
  assign n44975 = pi1459 & ~n44946;
  assign po1767 = n44974 | n44975;
  assign n44977 = ~n40852 & n44946;
  assign n44978 = pi1460 & ~n44946;
  assign po1768 = n44977 | n44978;
  assign n44980 = ~n40441 & n44946;
  assign n44981 = pi1461 & ~n44946;
  assign po1769 = n44980 | n44981;
  assign n44983 = ~pi0565 & pi3582;
  assign n44984 = pi3641 & po3852;
  assign n44985 = pi0565 & ~pi3641;
  assign n44986 = ~n44984 & ~n44985;
  assign n44987 = ~pi3631 & ~n44986;
  assign n44988 = pi2409 & pi3344;
  assign n44989 = pi2529 & ~pi3680;
  assign n44990 = ~pi3680 & ~n44989;
  assign n44991 = pi2647 & ~n44990;
  assign n44992 = n44988 & n44991;
  assign n44993 = n44987 & ~n44992;
  assign n44994 = ~n44983 & n44993;
  assign n44995 = ~po3616 & ~n44983;
  assign n44996 = n8312 & n44992;
  assign n44997 = po3646 & n44996;
  assign n44998 = n44995 & n44997;
  assign n44999 = ~n44994 & ~n44998;
  assign n45000 = ~pi2789 & ~pi3257;
  assign n45001 = ~n44999 & ~n45000;
  assign n45002 = pi0565 & n8358;
  assign n45003 = n45001 & n45002;
  assign n45004 = n8193 & ~n44983;
  assign n45005 = pi1462 & ~n45004;
  assign n45006 = n44999 & n45005;
  assign po1771 = n45003 | n45006;
  assign n45008 = ~pi1463 & ~n42185;
  assign n45009 = pi1463 & ~n44667;
  assign n45010 = ~pi0912 & n44667;
  assign n45011 = ~n45009 & ~n45010;
  assign n45012 = n42185 & n45011;
  assign po1772 = n45008 | n45012;
  assign n45014 = ~pi1464 & ~n42185;
  assign n45015 = pi0912 & n44654;
  assign n45016 = ~pi1464 & ~n44654;
  assign n45017 = ~n45015 & ~n45016;
  assign n45018 = n42185 & ~n45017;
  assign po1773 = n45014 | n45018;
  assign n45020 = ~pi1465 & ~n42185;
  assign n45021 = ~n42189 & n44645;
  assign n45022 = pi1465 & ~n45021;
  assign n45023 = ~pi0979 & n45021;
  assign n45024 = ~n45022 & ~n45023;
  assign n45025 = n42185 & n45024;
  assign po1774 = n45020 | n45025;
  assign n45027 = ~pi1466 & ~n42185;
  assign n45028 = pi0916 & n44654;
  assign n45029 = ~pi1466 & ~n44654;
  assign n45030 = ~n45028 & ~n45029;
  assign n45031 = n42185 & ~n45030;
  assign po1775 = n45027 | n45031;
  assign n45033 = ~n12415 & n38320;
  assign n45034 = pi1467 & n38307;
  assign n45035 = ~pi1467 & ~n38307;
  assign n45036 = ~n45034 & ~n45035;
  assign n45037 = ~n36181 & ~n45036;
  assign n45038 = ~pi1467 & n36181;
  assign n45039 = ~n45037 & ~n45038;
  assign n45040 = ~n38320 & n45039;
  assign po1776 = n45033 | n45040;
  assign n45042 = ~pi1468 & ~n25623;
  assign po1777 = ~n44813 | n45042;
  assign n45044 = ~pi1469 & ~n25623;
  assign po1778 = ~n44813 | n45044;
  assign n45046 = ~pi1470 & ~n25623;
  assign po1779 = ~n44813 | n45046;
  assign n45048 = ~pi1471 & ~n25623;
  assign po1780 = ~n44813 | n45048;
  assign n45050 = ~pi0423 & n44810;
  assign n45051 = pi0424 & n45050;
  assign n45052 = ~pi1472 & ~n25623;
  assign n45053 = ~pi0405 & pi0422;
  assign n45054 = n25623 & n45053;
  assign n45055 = ~n45052 & ~n45054;
  assign po1781 = n45051 | ~n45055;
  assign n45057 = ~pi1473 & ~n25623;
  assign po1782 = ~n44813 | n45057;
  assign n45059 = ~n13398 & n38320;
  assign n45060 = pi1474 & n42649;
  assign n45061 = ~pi1474 & ~n42649;
  assign n45062 = ~n45060 & ~n45061;
  assign n45063 = ~n36181 & ~n45062;
  assign n45064 = ~pi1474 & n36181;
  assign n45065 = ~n45063 & ~n45064;
  assign n45066 = ~n38320 & n45065;
  assign po1783 = n45059 | n45066;
  assign n45068 = ~pi1475 & ~n42185;
  assign n45069 = pi0914 & n44654;
  assign n45070 = ~pi1475 & ~n44654;
  assign n45071 = ~n45069 & ~n45070;
  assign n45072 = n42185 & ~n45071;
  assign po1784 = n45068 | n45072;
  assign n45074 = ~pi1476 & ~n42185;
  assign n45075 = pi1476 & ~n44631;
  assign n45076 = ~pi0830 & n44631;
  assign n45077 = ~n45075 & ~n45076;
  assign n45078 = n42185 & n45077;
  assign po1785 = n45074 | n45078;
  assign n45080 = ~pi1477 & ~n42185;
  assign n45081 = pi1477 & ~n44631;
  assign n45082 = ~pi0979 & n44631;
  assign n45083 = ~n45081 & ~n45082;
  assign n45084 = n42185 & n45083;
  assign po1786 = n45080 | n45084;
  assign n45086 = ~pi1478 & ~n42185;
  assign n45087 = pi1478 & ~n44631;
  assign n45088 = pi3633 & n44631;
  assign n45089 = ~n45087 & ~n45088;
  assign n45090 = n42185 & n45089;
  assign po1787 = n45086 | n45090;
  assign n45092 = ~pi1479 & ~n42185;
  assign n45093 = pi1479 & ~n44631;
  assign n45094 = ~pi0143 & n44631;
  assign n45095 = ~n45093 & ~n45094;
  assign n45096 = n42185 & n45095;
  assign po1788 = n45092 | n45096;
  assign n45098 = ~pi1480 & ~n42185;
  assign n45099 = pi1480 & ~n44631;
  assign n45100 = ~pi0659 & n44631;
  assign n45101 = ~n45099 & ~n45100;
  assign n45102 = n42185 & n45101;
  assign po1789 = n45098 | n45102;
  assign n45104 = ~pi1481 & ~n42185;
  assign n45105 = pi1481 & ~n44631;
  assign n45106 = ~pi0152 & n44631;
  assign n45107 = ~n45105 & ~n45106;
  assign n45108 = n42185 & n45107;
  assign po1790 = n45104 | n45108;
  assign n45110 = ~pi1482 & ~n42185;
  assign n45111 = pi1482 & ~n44631;
  assign n45112 = ~pi0912 & n44631;
  assign n45113 = ~n45111 & ~n45112;
  assign n45114 = n42185 & n45113;
  assign po1791 = n45110 | n45114;
  assign n45116 = ~pi1483 & ~n42185;
  assign n45117 = pi1483 & ~n44631;
  assign n45118 = ~pi0913 & n44631;
  assign n45119 = ~n45117 & ~n45118;
  assign n45120 = n42185 & n45119;
  assign po1792 = n45116 | n45120;
  assign n45122 = ~pi1484 & ~n42185;
  assign n45123 = pi1484 & ~n44631;
  assign n45124 = ~pi0915 & n44631;
  assign n45125 = ~n45123 & ~n45124;
  assign n45126 = n42185 & n45125;
  assign po1793 = n45122 | n45126;
  assign n45128 = ~pi1485 & ~n42185;
  assign n45129 = pi1485 & ~n44631;
  assign n45130 = ~pi0134 & n44631;
  assign n45131 = ~n45129 & ~n45130;
  assign n45132 = n42185 & n45131;
  assign po1794 = n45128 | n45132;
  assign n45134 = ~pi1486 & ~n42185;
  assign n45135 = pi1486 & ~n44631;
  assign n45136 = ~pi0708 & n44631;
  assign n45137 = ~n45135 & ~n45136;
  assign n45138 = n42185 & n45137;
  assign po1795 = n45134 | n45138;
  assign n45140 = ~pi1487 & ~n42185;
  assign n45141 = pi1487 & ~n44631;
  assign n45142 = ~pi0918 & n44631;
  assign n45143 = ~n45141 & ~n45142;
  assign n45144 = n42185 & n45143;
  assign po1796 = n45140 | n45144;
  assign n45146 = ~pi1488 & ~n42185;
  assign n45147 = pi1488 & ~n44631;
  assign n45148 = ~pi0919 & n44631;
  assign n45149 = ~n45147 & ~n45148;
  assign n45150 = n42185 & n45149;
  assign po1797 = n45146 | n45150;
  assign n45152 = ~pi1489 & ~n42185;
  assign n45153 = pi1489 & ~n44631;
  assign n45154 = ~pi0826 & n44631;
  assign n45155 = ~n45153 & ~n45154;
  assign n45156 = n42185 & n45155;
  assign po1798 = n45152 | n45156;
  assign n45158 = ~pi1490 & ~n42185;
  assign n45159 = pi1490 & ~n44631;
  assign n45160 = ~pi0827 & n44631;
  assign n45161 = ~n45159 & ~n45160;
  assign n45162 = n42185 & n45161;
  assign po1799 = n45158 | n45162;
  assign n45164 = ~pi1491 & ~n42185;
  assign n45165 = pi1491 & ~n44631;
  assign n45166 = ~pi0868 & n44631;
  assign n45167 = ~n45165 & ~n45166;
  assign n45168 = n42185 & n45167;
  assign po1800 = n45164 | n45168;
  assign n45170 = ~pi1492 & ~n42185;
  assign n45171 = pi1492 & ~n44631;
  assign n45172 = ~pi0829 & n44631;
  assign n45173 = ~n45171 & ~n45172;
  assign n45174 = n42185 & n45173;
  assign po1801 = n45170 | n45174;
  assign n45176 = ~pi1493 & ~n42185;
  assign n45177 = pi1493 & ~n44631;
  assign n45178 = ~pi0149 & n44631;
  assign n45179 = ~n45177 & ~n45178;
  assign n45180 = n42185 & n45179;
  assign po1802 = n45176 | n45180;
  assign n45182 = ~pi1494 & ~n42185;
  assign n45183 = pi1494 & ~n45021;
  assign n45184 = ~pi0830 & n45021;
  assign n45185 = ~n45183 & ~n45184;
  assign n45186 = n42185 & n45185;
  assign po1803 = n45182 | n45186;
  assign n45188 = ~pi1495 & ~n42185;
  assign n45189 = pi1495 & ~n45021;
  assign n45190 = ~pi0586 & n45021;
  assign n45191 = ~n45189 & ~n45190;
  assign n45192 = n42185 & n45191;
  assign po1804 = n45188 | n45192;
  assign n45194 = ~pi1496 & ~n42185;
  assign n45195 = pi1496 & ~n45021;
  assign n45196 = pi3633 & n45021;
  assign n45197 = ~n45195 & ~n45196;
  assign n45198 = n42185 & n45197;
  assign po1805 = n45194 | n45198;
  assign n45200 = ~pi1497 & ~n42185;
  assign n45201 = pi1497 & ~n45021;
  assign n45202 = ~pi0143 & n45021;
  assign n45203 = ~n45201 & ~n45202;
  assign n45204 = n42185 & n45203;
  assign po1806 = n45200 | n45204;
  assign n45206 = ~pi1498 & ~n42185;
  assign n45207 = pi1498 & ~n45021;
  assign n45208 = ~pi0196 & n45021;
  assign n45209 = ~n45207 & ~n45208;
  assign n45210 = n42185 & n45209;
  assign po1807 = n45206 | n45210;
  assign n45212 = ~pi1499 & ~n42185;
  assign n45213 = pi1499 & ~n45021;
  assign n45214 = ~pi0152 & n45021;
  assign n45215 = ~n45213 & ~n45214;
  assign n45216 = n42185 & n45215;
  assign po1808 = n45212 | n45216;
  assign n45218 = ~pi1500 & ~n42185;
  assign n45219 = pi1500 & ~n45021;
  assign n45220 = ~pi0912 & n45021;
  assign n45221 = ~n45219 & ~n45220;
  assign n45222 = n42185 & n45221;
  assign po1809 = n45218 | n45222;
  assign n45224 = ~pi1501 & ~n42185;
  assign n45225 = pi1501 & ~n45021;
  assign n45226 = ~pi0914 & n45021;
  assign n45227 = ~n45225 & ~n45226;
  assign n45228 = n42185 & n45227;
  assign po1810 = n45224 | n45228;
  assign n45230 = ~pi1502 & ~n42185;
  assign n45231 = pi1502 & ~n45021;
  assign n45232 = ~pi0915 & n45021;
  assign n45233 = ~n45231 & ~n45232;
  assign n45234 = n42185 & n45233;
  assign po1811 = n45230 | n45234;
  assign n45236 = ~pi1503 & ~n42185;
  assign n45237 = pi1503 & ~n45021;
  assign n45238 = ~pi0916 & n45021;
  assign n45239 = ~n45237 & ~n45238;
  assign n45240 = n42185 & n45239;
  assign po1812 = n45236 | n45240;
  assign n45242 = ~pi1504 & ~n42185;
  assign n45243 = pi1504 & ~n45021;
  assign n45244 = ~pi0917 & n45021;
  assign n45245 = ~n45243 & ~n45244;
  assign n45246 = n42185 & n45245;
  assign po1813 = n45242 | n45246;
  assign n45248 = ~pi1505 & ~n42185;
  assign n45249 = pi1505 & ~n45021;
  assign n45250 = ~pi0918 & n45021;
  assign n45251 = ~n45249 & ~n45250;
  assign n45252 = n42185 & n45251;
  assign po1814 = n45248 | n45252;
  assign n45254 = ~pi1506 & ~n42185;
  assign n45255 = pi1506 & ~n45021;
  assign n45256 = ~pi0980 & n45021;
  assign n45257 = ~n45255 & ~n45256;
  assign n45258 = n42185 & n45257;
  assign po1815 = n45254 | n45258;
  assign n45260 = ~pi1507 & ~n42185;
  assign n45261 = pi1507 & ~n45021;
  assign n45262 = ~pi0826 & n45021;
  assign n45263 = ~n45261 & ~n45262;
  assign n45264 = n42185 & n45263;
  assign po1816 = n45260 | n45264;
  assign n45266 = ~pi1508 & ~n42185;
  assign n45267 = pi1508 & ~n45021;
  assign n45268 = ~pi0827 & n45021;
  assign n45269 = ~n45267 & ~n45268;
  assign n45270 = n42185 & n45269;
  assign po1817 = n45266 | n45270;
  assign n45272 = ~pi1509 & ~n42185;
  assign n45273 = pi1509 & ~n45021;
  assign n45274 = ~pi0828 & n45021;
  assign n45275 = ~n45273 & ~n45274;
  assign n45276 = n42185 & n45275;
  assign po1818 = n45272 | n45276;
  assign n45278 = ~pi1510 & ~n42185;
  assign n45279 = pi1510 & ~n45021;
  assign n45280 = ~pi0829 & n45021;
  assign n45281 = ~n45279 & ~n45280;
  assign n45282 = n42185 & n45281;
  assign po1819 = n45278 | n45282;
  assign n45284 = ~pi1511 & ~n42185;
  assign n45285 = pi1511 & ~n45021;
  assign n45286 = ~pi0149 & n45021;
  assign n45287 = ~n45285 & ~n45286;
  assign n45288 = n42185 & n45287;
  assign po1820 = n45284 | n45288;
  assign n45290 = ~pi1512 & ~n42185;
  assign n45291 = pi1512 & ~n44667;
  assign n45292 = ~pi0979 & n44667;
  assign n45293 = ~n45291 & ~n45292;
  assign n45294 = n42185 & n45293;
  assign po1821 = n45290 | n45294;
  assign n45296 = ~pi1513 & ~n42185;
  assign n45297 = pi1513 & ~n44667;
  assign n45298 = ~pi0586 & n44667;
  assign n45299 = ~n45297 & ~n45298;
  assign n45300 = n42185 & n45299;
  assign po1822 = n45296 | n45300;
  assign n45302 = ~pi1514 & ~n42185;
  assign n45303 = pi1514 & ~n44667;
  assign n45304 = pi3633 & n44667;
  assign n45305 = ~n45303 & ~n45304;
  assign n45306 = n42185 & n45305;
  assign po1823 = n45302 | n45306;
  assign n45308 = ~pi1515 & ~n42185;
  assign n45309 = pi1515 & ~n44667;
  assign n45310 = ~pi0659 & n44667;
  assign n45311 = ~n45309 & ~n45310;
  assign n45312 = n42185 & n45311;
  assign po1824 = n45308 | n45312;
  assign n45314 = ~pi1516 & ~n42185;
  assign n45315 = pi1516 & ~n44667;
  assign n45316 = ~pi0196 & n44667;
  assign n45317 = ~n45315 & ~n45316;
  assign n45318 = n42185 & n45317;
  assign po1825 = n45314 | n45318;
  assign n45320 = ~pi1517 & ~n42185;
  assign n45321 = pi1517 & ~n44667;
  assign n45322 = ~pi0152 & n44667;
  assign n45323 = ~n45321 & ~n45322;
  assign n45324 = n42185 & n45323;
  assign po1826 = n45320 | n45324;
  assign n45326 = ~pi1518 & ~n42185;
  assign n45327 = pi1518 & ~n44667;
  assign n45328 = ~pi0913 & n44667;
  assign n45329 = ~n45327 & ~n45328;
  assign n45330 = n42185 & n45329;
  assign po1827 = n45326 | n45330;
  assign n45332 = ~pi1519 & ~n42185;
  assign n45333 = pi1519 & ~n44667;
  assign n45334 = ~pi0914 & n44667;
  assign n45335 = ~n45333 & ~n45334;
  assign n45336 = n42185 & n45335;
  assign po1828 = n45332 | n45336;
  assign n45338 = ~pi1520 & ~n42185;
  assign n45339 = pi1520 & ~n44667;
  assign n45340 = ~pi0915 & n44667;
  assign n45341 = ~n45339 & ~n45340;
  assign n45342 = n42185 & n45341;
  assign po1829 = n45338 | n45342;
  assign n45344 = ~pi1521 & ~n42185;
  assign n45345 = pi1521 & ~n44667;
  assign n45346 = ~pi0134 & n44667;
  assign n45347 = ~n45345 & ~n45346;
  assign n45348 = n42185 & n45347;
  assign po1830 = n45344 | n45348;
  assign n45350 = ~pi1522 & ~n42185;
  assign n45351 = pi1522 & ~n44667;
  assign n45352 = ~pi0917 & n44667;
  assign n45353 = ~n45351 & ~n45352;
  assign n45354 = n42185 & n45353;
  assign po1831 = n45350 | n45354;
  assign n45356 = ~pi1523 & ~n42185;
  assign n45357 = pi1523 & ~n44667;
  assign n45358 = ~pi0708 & n44667;
  assign n45359 = ~n45357 & ~n45358;
  assign n45360 = n42185 & n45359;
  assign po1832 = n45356 | n45360;
  assign n45362 = ~pi1524 & ~n42185;
  assign n45363 = pi1524 & ~n44667;
  assign n45364 = ~pi0919 & n44667;
  assign n45365 = ~n45363 & ~n45364;
  assign n45366 = n42185 & n45365;
  assign po1833 = n45362 | n45366;
  assign n45368 = ~pi1525 & ~n42185;
  assign n45369 = pi1525 & ~n44667;
  assign n45370 = ~pi0980 & n44667;
  assign n45371 = ~n45369 & ~n45370;
  assign n45372 = n42185 & n45371;
  assign po1834 = n45368 | n45372;
  assign n45374 = ~pi1526 & ~n42185;
  assign n45375 = pi1526 & ~n44667;
  assign n45376 = ~pi0826 & n44667;
  assign n45377 = ~n45375 & ~n45376;
  assign n45378 = n42185 & n45377;
  assign po1835 = n45374 | n45378;
  assign n45380 = ~pi1527 & ~n42185;
  assign n45381 = pi1527 & ~n44667;
  assign n45382 = ~pi0868 & n44667;
  assign n45383 = ~n45381 & ~n45382;
  assign n45384 = n42185 & n45383;
  assign po1836 = n45380 | n45384;
  assign n45386 = ~pi1528 & ~n42185;
  assign n45387 = pi1528 & ~n44667;
  assign n45388 = ~pi0828 & n44667;
  assign n45389 = ~n45387 & ~n45388;
  assign n45390 = n42185 & n45389;
  assign po1837 = n45386 | n45390;
  assign n45392 = ~pi1529 & ~n42185;
  assign n45393 = pi1529 & ~n44667;
  assign n45394 = ~pi0829 & n44667;
  assign n45395 = ~n45393 & ~n45394;
  assign n45396 = n42185 & n45395;
  assign po1838 = n45392 | n45396;
  assign n45398 = ~pi1530 & ~n42185;
  assign n45399 = pi0830 & n44741;
  assign n45400 = ~pi1530 & ~n44741;
  assign n45401 = ~n45399 & ~n45400;
  assign n45402 = n42185 & ~n45401;
  assign po1839 = n45398 | n45402;
  assign n45404 = ~pi1531 & ~n42185;
  assign n45405 = pi0979 & n44741;
  assign n45406 = ~pi1531 & ~n44741;
  assign n45407 = ~n45405 & ~n45406;
  assign n45408 = n42185 & ~n45407;
  assign po1840 = n45404 | n45408;
  assign n45410 = ~pi1532 & ~n42185;
  assign n45411 = pi0586 & n44741;
  assign n45412 = ~pi1532 & ~n44741;
  assign n45413 = ~n45411 & ~n45412;
  assign n45414 = n42185 & ~n45413;
  assign po1841 = n45410 | n45414;
  assign n45416 = ~pi1533 & ~n42185;
  assign n45417 = pi0143 & n44741;
  assign n45418 = ~pi1533 & ~n44741;
  assign n45419 = ~n45417 & ~n45418;
  assign n45420 = n42185 & ~n45419;
  assign po1842 = n45416 | n45420;
  assign n45422 = ~pi1534 & ~n42185;
  assign n45423 = pi0659 & n44741;
  assign n45424 = ~pi1534 & ~n44741;
  assign n45425 = ~n45423 & ~n45424;
  assign n45426 = n42185 & ~n45425;
  assign po1843 = n45422 | n45426;
  assign n45428 = ~pi1535 & ~n42185;
  assign n45429 = pi0196 & n44741;
  assign n45430 = ~pi1535 & ~n44741;
  assign n45431 = ~n45429 & ~n45430;
  assign n45432 = n42185 & ~n45431;
  assign po1844 = n45428 | n45432;
  assign n45434 = ~pi1536 & ~n42185;
  assign n45435 = pi0912 & n44741;
  assign n45436 = ~pi1536 & ~n44741;
  assign n45437 = ~n45435 & ~n45436;
  assign n45438 = n42185 & ~n45437;
  assign po1845 = n45434 | n45438;
  assign n45440 = ~pi1537 & ~n42185;
  assign n45441 = pi0913 & n44741;
  assign n45442 = ~pi1537 & ~n44741;
  assign n45443 = ~n45441 & ~n45442;
  assign n45444 = n42185 & ~n45443;
  assign po1846 = n45440 | n45444;
  assign n45446 = ~pi1538 & ~n42185;
  assign n45447 = pi0914 & n44741;
  assign n45448 = ~pi1538 & ~n44741;
  assign n45449 = ~n45447 & ~n45448;
  assign n45450 = n42185 & ~n45449;
  assign po1847 = n45446 | n45450;
  assign n45452 = ~pi1539 & ~n42185;
  assign n45453 = pi0916 & n44741;
  assign n45454 = ~pi1539 & ~n44741;
  assign n45455 = ~n45453 & ~n45454;
  assign n45456 = n42185 & ~n45455;
  assign po1848 = n45452 | n45456;
  assign n45458 = ~pi1540 & ~n42185;
  assign n45459 = pi0134 & n44741;
  assign n45460 = ~pi1540 & ~n44741;
  assign n45461 = ~n45459 & ~n45460;
  assign n45462 = n42185 & ~n45461;
  assign po1849 = n45458 | n45462;
  assign n45464 = ~pi1541 & ~n42185;
  assign n45465 = pi0917 & n44741;
  assign n45466 = ~pi1541 & ~n44741;
  assign n45467 = ~n45465 & ~n45466;
  assign n45468 = n42185 & ~n45467;
  assign po1850 = n45464 | n45468;
  assign n45470 = ~pi1542 & ~n42185;
  assign n45471 = pi0918 & n44741;
  assign n45472 = ~pi1542 & ~n44741;
  assign n45473 = ~n45471 & ~n45472;
  assign n45474 = n42185 & ~n45473;
  assign po1851 = n45470 | n45474;
  assign n45476 = ~pi1543 & ~n42185;
  assign n45477 = pi0919 & n44741;
  assign n45478 = ~pi1543 & ~n44741;
  assign n45479 = ~n45477 & ~n45478;
  assign n45480 = n42185 & ~n45479;
  assign po1852 = n45476 | n45480;
  assign n45482 = ~pi1544 & ~n42185;
  assign n45483 = pi0980 & n44741;
  assign n45484 = ~pi1544 & ~n44741;
  assign n45485 = ~n45483 & ~n45484;
  assign n45486 = n42185 & ~n45485;
  assign po1853 = n45482 | n45486;
  assign n45488 = ~pi1545 & ~n42185;
  assign n45489 = pi0827 & n44741;
  assign n45490 = ~pi1545 & ~n44741;
  assign n45491 = ~n45489 & ~n45490;
  assign n45492 = n42185 & ~n45491;
  assign po1854 = n45488 | n45492;
  assign n45494 = ~pi1546 & ~n42185;
  assign n45495 = pi0828 & n44741;
  assign n45496 = ~pi1546 & ~n44741;
  assign n45497 = ~n45495 & ~n45496;
  assign n45498 = n42185 & ~n45497;
  assign po1855 = n45494 | n45498;
  assign n45500 = ~pi1547 & ~n42185;
  assign n45501 = pi0149 & n44741;
  assign n45502 = ~pi1547 & ~n44741;
  assign n45503 = ~n45501 & ~n45502;
  assign n45504 = n42185 & ~n45503;
  assign po1856 = n45500 | n45504;
  assign n45506 = ~pi1548 & ~n42185;
  assign n45507 = pi0830 & n44638;
  assign n45508 = ~pi1548 & ~n44638;
  assign n45509 = ~n45507 & ~n45508;
  assign n45510 = n42185 & ~n45509;
  assign po1857 = n45506 | n45510;
  assign n45512 = ~pi1549 & ~n42185;
  assign n45513 = pi0979 & n44638;
  assign n45514 = ~pi1549 & ~n44638;
  assign n45515 = ~n45513 & ~n45514;
  assign n45516 = n42185 & ~n45515;
  assign po1858 = n45512 | n45516;
  assign n45518 = ~pi1550 & ~n42185;
  assign n45519 = ~pi3633 & n44638;
  assign n45520 = ~pi1550 & ~n44638;
  assign n45521 = ~n45519 & ~n45520;
  assign n45522 = n42185 & ~n45521;
  assign po1859 = n45518 | n45522;
  assign n45524 = ~pi1551 & ~n42185;
  assign n45525 = pi0143 & n44638;
  assign n45526 = ~pi1551 & ~n44638;
  assign n45527 = ~n45525 & ~n45526;
  assign n45528 = n42185 & ~n45527;
  assign po1860 = n45524 | n45528;
  assign n45530 = ~pi1552 & ~n42185;
  assign n45531 = pi0659 & n44638;
  assign n45532 = ~pi1552 & ~n44638;
  assign n45533 = ~n45531 & ~n45532;
  assign n45534 = n42185 & ~n45533;
  assign po1861 = n45530 | n45534;
  assign n45536 = ~pi1553 & ~n42185;
  assign n45537 = pi0152 & n44638;
  assign n45538 = ~pi1553 & ~n44638;
  assign n45539 = ~n45537 & ~n45538;
  assign n45540 = n42185 & ~n45539;
  assign po1862 = n45536 | n45540;
  assign n45542 = ~pi1554 & ~n42185;
  assign n45543 = pi0913 & n44638;
  assign n45544 = ~pi1554 & ~n44638;
  assign n45545 = ~n45543 & ~n45544;
  assign n45546 = n42185 & ~n45545;
  assign po1863 = n45542 | n45546;
  assign n45548 = ~pi1555 & ~n42185;
  assign n45549 = pi0915 & n44638;
  assign n45550 = ~pi1555 & ~n44638;
  assign n45551 = ~n45549 & ~n45550;
  assign n45552 = n42185 & ~n45551;
  assign po1864 = n45548 | n45552;
  assign n45554 = ~pi1556 & ~n42185;
  assign n45555 = pi0916 & n44638;
  assign n45556 = ~pi1556 & ~n44638;
  assign n45557 = ~n45555 & ~n45556;
  assign n45558 = n42185 & ~n45557;
  assign po1865 = n45554 | n45558;
  assign n45560 = ~pi1557 & ~n42185;
  assign n45561 = pi0134 & n44638;
  assign n45562 = ~pi1557 & ~n44638;
  assign n45563 = ~n45561 & ~n45562;
  assign n45564 = n42185 & ~n45563;
  assign po1866 = n45560 | n45564;
  assign n45566 = ~pi1558 & ~n42185;
  assign n45567 = pi0708 & n44638;
  assign n45568 = ~pi1558 & ~n44638;
  assign n45569 = ~n45567 & ~n45568;
  assign n45570 = n42185 & ~n45569;
  assign po1867 = n45566 | n45570;
  assign n45572 = ~pi1559 & ~n42185;
  assign n45573 = pi0918 & n44638;
  assign n45574 = ~pi1559 & ~n44638;
  assign n45575 = ~n45573 & ~n45574;
  assign n45576 = n42185 & ~n45575;
  assign po1868 = n45572 | n45576;
  assign n45578 = ~pi1560 & ~n42185;
  assign n45579 = pi0919 & n44638;
  assign n45580 = ~pi1560 & ~n44638;
  assign n45581 = ~n45579 & ~n45580;
  assign n45582 = n42185 & ~n45581;
  assign po1869 = n45578 | n45582;
  assign n45584 = ~pi1561 & ~n42185;
  assign n45585 = pi0826 & n44638;
  assign n45586 = ~pi1561 & ~n44638;
  assign n45587 = ~n45585 & ~n45586;
  assign n45588 = n42185 & ~n45587;
  assign po1870 = n45584 | n45588;
  assign n45590 = ~pi1562 & ~n42185;
  assign n45591 = pi0868 & n44638;
  assign n45592 = ~pi1562 & ~n44638;
  assign n45593 = ~n45591 & ~n45592;
  assign n45594 = n42185 & ~n45593;
  assign po1871 = n45590 | n45594;
  assign n45596 = ~pi1563 & ~n42185;
  assign n45597 = pi0829 & n44638;
  assign n45598 = ~pi1563 & ~n44638;
  assign n45599 = ~n45597 & ~n45598;
  assign n45600 = n42185 & ~n45599;
  assign po1872 = n45596 | n45600;
  assign n45602 = ~pi1564 & ~n42185;
  assign n45603 = pi0149 & n44638;
  assign n45604 = ~pi1564 & ~n44638;
  assign n45605 = ~n45603 & ~n45604;
  assign n45606 = n42185 & ~n45605;
  assign po1873 = n45602 | n45606;
  assign n45608 = ~pi1565 & ~n42185;
  assign n45609 = pi0830 & n44646;
  assign n45610 = ~pi1565 & ~n44646;
  assign n45611 = ~n45609 & ~n45610;
  assign n45612 = n42185 & ~n45611;
  assign po1874 = n45608 | n45612;
  assign n45614 = ~pi1566 & ~n42185;
  assign n45615 = pi0586 & n44646;
  assign n45616 = ~pi1566 & ~n44646;
  assign n45617 = ~n45615 & ~n45616;
  assign n45618 = n42185 & ~n45617;
  assign po1875 = n45614 | n45618;
  assign n45620 = ~pi1567 & ~n42185;
  assign n45621 = ~pi3633 & n44646;
  assign n45622 = ~pi1567 & ~n44646;
  assign n45623 = ~n45621 & ~n45622;
  assign n45624 = n42185 & ~n45623;
  assign po1876 = n45620 | n45624;
  assign n45626 = ~pi1568 & ~n42185;
  assign n45627 = pi0143 & n44646;
  assign n45628 = ~pi1568 & ~n44646;
  assign n45629 = ~n45627 & ~n45628;
  assign n45630 = n42185 & ~n45629;
  assign po1877 = n45626 | n45630;
  assign n45632 = ~pi1569 & ~n42185;
  assign n45633 = pi0196 & n44646;
  assign n45634 = ~pi1569 & ~n44646;
  assign n45635 = ~n45633 & ~n45634;
  assign n45636 = n42185 & ~n45635;
  assign po1878 = n45632 | n45636;
  assign n45638 = ~pi1570 & ~n42185;
  assign n45639 = pi0152 & n44646;
  assign n45640 = ~pi1570 & ~n44646;
  assign n45641 = ~n45639 & ~n45640;
  assign n45642 = n42185 & ~n45641;
  assign po1879 = n45638 | n45642;
  assign n45644 = ~pi1571 & ~n42185;
  assign n45645 = pi0912 & n44646;
  assign n45646 = ~pi1571 & ~n44646;
  assign n45647 = ~n45645 & ~n45646;
  assign n45648 = n42185 & ~n45647;
  assign po1880 = n45644 | n45648;
  assign n45650 = ~pi1572 & ~n42185;
  assign n45651 = pi0914 & n44646;
  assign n45652 = ~pi1572 & ~n44646;
  assign n45653 = ~n45651 & ~n45652;
  assign n45654 = n42185 & ~n45653;
  assign po1881 = n45650 | n45654;
  assign n45656 = ~pi1573 & ~n42185;
  assign n45657 = pi0916 & n44646;
  assign n45658 = ~pi1573 & ~n44646;
  assign n45659 = ~n45657 & ~n45658;
  assign n45660 = n42185 & ~n45659;
  assign po1882 = n45656 | n45660;
  assign n45662 = ~pi1574 & ~n42185;
  assign n45663 = pi0917 & n44646;
  assign n45664 = ~pi1574 & ~n44646;
  assign n45665 = ~n45663 & ~n45664;
  assign n45666 = n42185 & ~n45665;
  assign po1883 = n45662 | n45666;
  assign n45668 = ~pi1575 & ~n42185;
  assign n45669 = pi0918 & n44646;
  assign n45670 = ~pi1575 & ~n44646;
  assign n45671 = ~n45669 & ~n45670;
  assign n45672 = n42185 & ~n45671;
  assign po1884 = n45668 | n45672;
  assign n45674 = ~pi1576 & ~n42185;
  assign n45675 = pi0980 & n44646;
  assign n45676 = ~pi1576 & ~n44646;
  assign n45677 = ~n45675 & ~n45676;
  assign n45678 = n42185 & ~n45677;
  assign po1885 = n45674 | n45678;
  assign n45680 = ~pi1577 & ~n42185;
  assign n45681 = pi0827 & n44646;
  assign n45682 = ~pi1577 & ~n44646;
  assign n45683 = ~n45681 & ~n45682;
  assign n45684 = n42185 & ~n45683;
  assign po1886 = n45680 | n45684;
  assign n45686 = ~pi1578 & ~n42185;
  assign n45687 = pi0828 & n44646;
  assign n45688 = ~pi1578 & ~n44646;
  assign n45689 = ~n45687 & ~n45688;
  assign n45690 = n42185 & ~n45689;
  assign po1887 = n45686 | n45690;
  assign n45692 = ~pi1579 & ~n42185;
  assign n45693 = pi0829 & n44646;
  assign n45694 = ~pi1579 & ~n44646;
  assign n45695 = ~n45693 & ~n45694;
  assign n45696 = n42185 & ~n45695;
  assign po1888 = n45692 | n45696;
  assign n45698 = ~pi1580 & ~n42185;
  assign n45699 = pi0149 & n44646;
  assign n45700 = ~pi1580 & ~n44646;
  assign n45701 = ~n45699 & ~n45700;
  assign n45702 = n42185 & ~n45701;
  assign po1889 = n45698 | n45702;
  assign n45704 = ~pi1581 & ~n42185;
  assign n45705 = pi0979 & n44654;
  assign n45706 = ~pi1581 & ~n44654;
  assign n45707 = ~n45705 & ~n45706;
  assign n45708 = n42185 & ~n45707;
  assign po1890 = n45704 | n45708;
  assign n45710 = ~pi1582 & ~n42185;
  assign n45711 = ~pi3633 & n44654;
  assign n45712 = ~pi1582 & ~n44654;
  assign n45713 = ~n45711 & ~n45712;
  assign n45714 = n42185 & ~n45713;
  assign po1891 = n45710 | n45714;
  assign n45716 = ~pi1583 & ~n42185;
  assign n45717 = pi0659 & n44654;
  assign n45718 = ~pi1583 & ~n44654;
  assign n45719 = ~n45717 & ~n45718;
  assign n45720 = n42185 & ~n45719;
  assign po1892 = n45716 | n45720;
  assign n45722 = ~pi1584 & ~n42185;
  assign n45723 = pi0196 & n44654;
  assign n45724 = ~pi1584 & ~n44654;
  assign n45725 = ~n45723 & ~n45724;
  assign n45726 = n42185 & ~n45725;
  assign po1893 = n45722 | n45726;
  assign n45728 = ~pi1585 & ~n42185;
  assign n45729 = pi0152 & n44654;
  assign n45730 = ~pi1585 & ~n44654;
  assign n45731 = ~n45729 & ~n45730;
  assign n45732 = n42185 & ~n45731;
  assign po1894 = n45728 | n45732;
  assign n45734 = ~pi1586 & ~n42185;
  assign n45735 = pi0913 & n44654;
  assign n45736 = ~pi1586 & ~n44654;
  assign n45737 = ~n45735 & ~n45736;
  assign n45738 = n42185 & ~n45737;
  assign po1895 = n45734 | n45738;
  assign n45740 = ~pi1587 & ~n42185;
  assign n45741 = pi0915 & n44654;
  assign n45742 = ~pi1587 & ~n44654;
  assign n45743 = ~n45741 & ~n45742;
  assign n45744 = n42185 & ~n45743;
  assign po1896 = n45740 | n45744;
  assign n45746 = ~pi1588 & ~n42185;
  assign n45747 = pi0134 & n44654;
  assign n45748 = ~pi1588 & ~n44654;
  assign n45749 = ~n45747 & ~n45748;
  assign n45750 = n42185 & ~n45749;
  assign po1897 = n45746 | n45750;
  assign n45752 = ~pi1589 & ~n42185;
  assign n45753 = pi0917 & n44654;
  assign n45754 = ~pi1589 & ~n44654;
  assign n45755 = ~n45753 & ~n45754;
  assign n45756 = n42185 & ~n45755;
  assign po1898 = n45752 | n45756;
  assign n45758 = ~pi1590 & ~n42185;
  assign n45759 = pi0708 & n44654;
  assign n45760 = ~pi1590 & ~n44654;
  assign n45761 = ~n45759 & ~n45760;
  assign n45762 = n42185 & ~n45761;
  assign po1899 = n45758 | n45762;
  assign n45764 = ~pi1591 & ~n42185;
  assign n45765 = pi0919 & n44654;
  assign n45766 = ~pi1591 & ~n44654;
  assign n45767 = ~n45765 & ~n45766;
  assign n45768 = n42185 & ~n45767;
  assign po1900 = n45764 | n45768;
  assign n45770 = ~pi1592 & ~n42185;
  assign n45771 = pi0980 & n44654;
  assign n45772 = ~pi1592 & ~n44654;
  assign n45773 = ~n45771 & ~n45772;
  assign n45774 = n42185 & ~n45773;
  assign po1901 = n45770 | n45774;
  assign n45776 = ~pi1593 & ~n42185;
  assign n45777 = pi0826 & n44654;
  assign n45778 = ~pi1593 & ~n44654;
  assign n45779 = ~n45777 & ~n45778;
  assign n45780 = n42185 & ~n45779;
  assign po1902 = n45776 | n45780;
  assign n45782 = ~pi1594 & ~n42185;
  assign n45783 = pi0868 & n44654;
  assign n45784 = ~pi1594 & ~n44654;
  assign n45785 = ~n45783 & ~n45784;
  assign n45786 = n42185 & ~n45785;
  assign po1903 = n45782 | n45786;
  assign n45788 = ~pi1595 & ~n42185;
  assign n45789 = pi0829 & n44654;
  assign n45790 = ~pi1595 & ~n44654;
  assign n45791 = ~n45789 & ~n45790;
  assign n45792 = n42185 & ~n45791;
  assign po1904 = n45788 | n45792;
  assign n45794 = pi1596 & ~pi3137;
  assign n45795 = ~pi2564 & ~n45794;
  assign n45796 = ~pi1596 & pi3137;
  assign po1905 = n45795 | n45796;
  assign n45798 = n38240 & n38262;
  assign n45799 = n38256 & n45798;
  assign n45800 = pi1597 & ~n38262;
  assign po1906 = n45799 | n45800;
  assign n45802 = n38243 & ~n38253;
  assign n45803 = n42248 & n45802;
  assign n45804 = n38262 & n45803;
  assign n45805 = n38246 & n45804;
  assign n45806 = n44253 & n45805;
  assign n45807 = pi1598 & ~n38262;
  assign po1907 = n45806 | n45807;
  assign n45809 = ~n8561 & n35999;
  assign n45810 = pi1599 & n8561;
  assign po1908 = n45809 | n45810;
  assign n45812 = ~n8561 & n38602;
  assign n45813 = pi1600 & n8561;
  assign po1909 = n45812 | n45813;
  assign n45815 = pi1601 & pi3252;
  assign n45816 = ~pi2505 & ~pi2522;
  assign n45817 = ~pi2503 & pi2504;
  assign n45818 = ~n45816 & n45817;
  assign n45819 = pi2504 & ~n45816;
  assign n45820 = pi2503 & ~n45819;
  assign n45821 = ~n45818 & ~n45820;
  assign n45822 = ~pi2759 & ~n45821;
  assign n45823 = pi2759 & n45821;
  assign n45824 = ~n45822 & ~n45823;
  assign n45825 = ~pi2504 & n45816;
  assign n45826 = ~n45819 & ~n45825;
  assign n45827 = ~pi3199 & n45826;
  assign n45828 = pi3199 & ~n45826;
  assign n45829 = ~n45827 & ~n45828;
  assign n45830 = n45824 & n45829;
  assign n45831 = pi2505 & pi2522;
  assign n45832 = ~n45816 & ~n45831;
  assign n45833 = pi3281 & n45832;
  assign n45834 = ~pi3281 & ~n45832;
  assign n45835 = ~n45833 & ~n45834;
  assign n45836 = ~pi2505 & pi3343;
  assign n45837 = pi2505 & ~pi3343;
  assign n45838 = ~n45836 & ~n45837;
  assign n45839 = pi3099 & ~n45838;
  assign n45840 = pi2503 & n45819;
  assign n45841 = ~pi2049 & ~n45840;
  assign n45842 = pi2049 & n45840;
  assign n45843 = ~n45841 & ~n45842;
  assign n45844 = n45839 & ~n45843;
  assign n45845 = n45835 & n45844;
  assign n45846 = n45830 & n45845;
  assign po1910 = n45815 | n45846;
  assign n45848 = ~n13121 & n38320;
  assign n45849 = pi1602 & n41182;
  assign n45850 = ~pi1602 & ~n41182;
  assign n45851 = ~n45849 & ~n45850;
  assign n45852 = ~n36181 & ~n45851;
  assign n45853 = ~pi1602 & n36181;
  assign n45854 = ~n45852 & ~n45853;
  assign n45855 = ~n38320 & n45854;
  assign po1911 = n45848 | n45855;
  assign n45857 = ~n13988 & n38320;
  assign n45858 = pi1603 & n41167;
  assign n45859 = ~pi1603 & ~n41167;
  assign n45860 = ~n45858 & ~n45859;
  assign n45861 = ~n36181 & ~n45860;
  assign n45862 = ~pi1603 & n36181;
  assign n45863 = ~n45861 & ~n45862;
  assign n45864 = ~n38320 & n45863;
  assign po1912 = n45857 | n45864;
  assign n45866 = ~pi1604 & ~n41779;
  assign n45867 = n42444 & n42449;
  assign n45868 = pi1604 & n45867;
  assign n45869 = ~pi1604 & ~n45867;
  assign n45870 = ~n45868 & ~n45869;
  assign n45871 = n41779 & ~n45870;
  assign po1913 = n45866 | n45871;
  assign n45873 = pi1605 & pi3641;
  assign n45874 = ~pi1605 & ~pi3641;
  assign n45875 = ~n45873 & ~n45874;
  assign n45876 = n37393 & ~n45875;
  assign n45877 = pi1434 & ~n37393;
  assign po1914 = n45876 | n45877;
  assign n45879 = ~pi1606 & ~n31859;
  assign n45880 = ~n31860 & ~n45879;
  assign n45881 = pi3641 & ~n45880;
  assign n45882 = ~pi1606 & ~pi3641;
  assign n45883 = ~n45881 & ~n45882;
  assign n45884 = n37390 & ~n45883;
  assign n45885 = ~n37392 & n45884;
  assign n45886 = pi1431 & ~n37393;
  assign po1915 = n45885 | n45886;
  assign n45888 = pi0950 & po2823;
  assign n45889 = pi1607 & ~pi1847;
  assign n45890 = ~pi1846 & n42780;
  assign n45891 = pi1703 & n45890;
  assign n45892 = n45889 & n45891;
  assign n45893 = ~pi1847 & n45891;
  assign n45894 = ~pi1607 & ~n45893;
  assign n45895 = ~n45892 & ~n45894;
  assign n45896 = po3310 & ~n45895;
  assign n45897 = ~pi1607 & ~po3310;
  assign n45898 = ~n45896 & ~n45897;
  assign n45899 = ~po2823 & ~n45898;
  assign po1916 = n45888 | n45899;
  assign n45901 = pi0965 & po2824;
  assign n45902 = pi1608 & ~pi1848;
  assign n45903 = ~pi1849 & n44477;
  assign n45904 = pi1644 & n45903;
  assign n45905 = n45902 & n45904;
  assign n45906 = ~pi1848 & n45904;
  assign n45907 = ~pi1608 & ~n45906;
  assign n45908 = ~n45905 & ~n45907;
  assign n45909 = po3311 & ~n45908;
  assign n45910 = ~pi1608 & ~po3311;
  assign n45911 = ~n45909 & ~n45910;
  assign n45912 = ~po2824 & ~n45911;
  assign po1917 = n45901 | n45912;
  assign n45914 = ~pi1609 & n44550;
  assign n45915 = pi1609 & ~n44550;
  assign po1918 = n45914 | n45915;
  assign n45917 = ~pi1610 & ~n41779;
  assign n45918 = n41757 & n41771;
  assign n45919 = ~pi1675 & ~pi1676;
  assign n45920 = n41761 & n45919;
  assign n45921 = n41759 & n45920;
  assign n45922 = n41762 & n41769;
  assign n45923 = n41765 & n41768;
  assign n45924 = n45922 & n45923;
  assign n45925 = n41756 & n41766;
  assign n45926 = n45924 & n45925;
  assign n45927 = n45921 & n45926;
  assign n45928 = n45918 & n45927;
  assign n45929 = ~pi1610 & ~n45928;
  assign n45930 = pi1610 & n45928;
  assign n45931 = ~n45929 & ~n45930;
  assign n45932 = n41779 & ~n45931;
  assign po1919 = n45917 | n45932;
  assign n45934 = ~pi1611 & ~n42185;
  assign n45935 = pi0830 & n44654;
  assign n45936 = ~pi1611 & ~n44654;
  assign n45937 = ~n45935 & ~n45936;
  assign n45938 = n42185 & ~n45937;
  assign po1920 = n45934 | n45938;
  assign n45940 = ~pi1612 & ~n42185;
  assign n45941 = pi1612 & ~n44667;
  assign n45942 = ~pi0143 & n44667;
  assign n45943 = ~n45941 & ~n45942;
  assign n45944 = n42185 & n45943;
  assign po1921 = n45940 | n45944;
  assign n45946 = ~pi1613 & ~n42185;
  assign n45947 = pi0143 & n44654;
  assign n45948 = ~pi1613 & ~n44654;
  assign n45949 = ~n45947 & ~n45948;
  assign n45950 = n42185 & ~n45949;
  assign po1922 = n45946 | n45950;
  assign n45952 = ~pi1614 & ~n42185;
  assign n45953 = pi0586 & n44654;
  assign n45954 = ~pi1614 & ~n44654;
  assign n45955 = ~n45953 & ~n45954;
  assign n45956 = n42185 & ~n45955;
  assign po1923 = n45952 | n45956;
  assign n45958 = ~pi1615 & ~n42185;
  assign n45959 = pi1615 & ~n44667;
  assign n45960 = ~pi0830 & n44667;
  assign n45961 = ~n45959 & ~n45960;
  assign n45962 = n42185 & n45961;
  assign po1924 = n45958 | n45962;
  assign n45964 = ~pi1616 & ~n42185;
  assign n45965 = pi0868 & n44646;
  assign n45966 = ~pi1616 & ~n44646;
  assign n45967 = ~n45965 & ~n45966;
  assign n45968 = n42185 & ~n45967;
  assign po1925 = n45964 | n45968;
  assign n45970 = ~pi1617 & ~n42185;
  assign n45971 = pi1617 & ~n45021;
  assign n45972 = ~pi0868 & n45021;
  assign n45973 = ~n45971 & ~n45972;
  assign n45974 = n42185 & n45973;
  assign po1926 = n45970 | n45974;
  assign n45976 = ~pi1618 & ~n42185;
  assign n45977 = pi0913 & n44646;
  assign n45978 = ~pi1618 & ~n44646;
  assign n45979 = ~n45977 & ~n45978;
  assign n45980 = n42185 & ~n45979;
  assign po1927 = n45976 | n45980;
  assign n45982 = ~pi1619 & ~n42185;
  assign n45983 = pi0708 & n44646;
  assign n45984 = ~pi1619 & ~n44646;
  assign n45985 = ~n45983 & ~n45984;
  assign n45986 = n42185 & ~n45985;
  assign po1928 = n45982 | n45986;
  assign n45988 = ~pi1620 & ~n42185;
  assign n45989 = pi1620 & ~n45021;
  assign n45990 = ~pi0134 & n45021;
  assign n45991 = ~n45989 & ~n45990;
  assign n45992 = n42185 & n45991;
  assign po1929 = n45988 | n45992;
  assign n45994 = ~pi1621 & ~n42185;
  assign n45995 = pi0826 & n44646;
  assign n45996 = ~pi1621 & ~n44646;
  assign n45997 = ~n45995 & ~n45996;
  assign n45998 = n42185 & ~n45997;
  assign po1930 = n45994 | n45998;
  assign n46000 = ~pi1622 & ~n42185;
  assign n46001 = pi1622 & ~n45021;
  assign n46002 = ~pi0919 & n45021;
  assign n46003 = ~n46001 & ~n46002;
  assign n46004 = n42185 & n46003;
  assign po1931 = n46000 | n46004;
  assign n46006 = ~pi1623 & ~n42185;
  assign n46007 = pi0919 & n44646;
  assign n46008 = ~pi1623 & ~n44646;
  assign n46009 = ~n46007 & ~n46008;
  assign n46010 = n42185 & ~n46009;
  assign po1932 = n46006 | n46010;
  assign n46012 = ~pi1624 & ~n42185;
  assign n46013 = pi1624 & ~n45021;
  assign n46014 = ~pi0708 & n45021;
  assign n46015 = ~n46013 & ~n46014;
  assign n46016 = n42185 & n46015;
  assign po1933 = n46012 | n46016;
  assign n46018 = ~pi1625 & ~n42185;
  assign n46019 = pi0134 & n44646;
  assign n46020 = ~pi1625 & ~n44646;
  assign n46021 = ~n46019 & ~n46020;
  assign n46022 = n42185 & ~n46021;
  assign po1934 = n46018 | n46022;
  assign n46024 = ~pi1626 & ~n42185;
  assign n46025 = pi1626 & ~n45021;
  assign n46026 = ~pi0659 & n45021;
  assign n46027 = ~n46025 & ~n46026;
  assign n46028 = n42185 & n46027;
  assign po1935 = n46024 | n46028;
  assign n46030 = ~pi1627 & ~n42185;
  assign n46031 = pi1627 & ~n45021;
  assign n46032 = ~pi0913 & n45021;
  assign n46033 = ~n46031 & ~n46032;
  assign n46034 = n42185 & n46033;
  assign po1936 = n46030 | n46034;
  assign n46036 = ~pi1628 & ~n42185;
  assign n46037 = pi0915 & n44646;
  assign n46038 = ~pi1628 & ~n44646;
  assign n46039 = ~n46037 & ~n46038;
  assign n46040 = n42185 & ~n46039;
  assign po1937 = n46036 | n46040;
  assign n46042 = pi0798 & po2824;
  assign n46043 = ~pi1629 & ~n44478;
  assign n46044 = pi1629 & n44478;
  assign n46045 = ~n46043 & ~n46044;
  assign n46046 = po3311 & ~n46045;
  assign n46047 = ~pi1629 & ~po3311;
  assign n46048 = ~n46046 & ~n46047;
  assign n46049 = ~po2824 & n46048;
  assign po1938 = n46042 | n46049;
  assign n46051 = ~pi1630 & ~n37331;
  assign n46052 = pi0616 & n37700;
  assign n46053 = pi0632 & n46052;
  assign n46054 = ~pi1630 & ~n46052;
  assign n46055 = ~n46053 & ~n46054;
  assign n46056 = n37331 & ~n46055;
  assign po1939 = n46051 | n46056;
  assign n46058 = ~pi1631 & ~n37331;
  assign n46059 = pi0593 & n46052;
  assign n46060 = ~pi1631 & ~n46052;
  assign n46061 = ~n46059 & ~n46060;
  assign n46062 = n37331 & ~n46061;
  assign po1940 = n46058 | n46062;
  assign n46064 = ~pi1632 & ~n37331;
  assign n46065 = pi0594 & n46052;
  assign n46066 = ~pi1632 & ~n46052;
  assign n46067 = ~n46065 & ~n46066;
  assign n46068 = n37331 & ~n46067;
  assign po1941 = n46064 | n46068;
  assign n46070 = ~pi1633 & ~n37331;
  assign n46071 = pi0571 & n46052;
  assign n46072 = ~pi1633 & ~n46052;
  assign n46073 = ~n46071 & ~n46072;
  assign n46074 = n37331 & ~n46073;
  assign po1942 = n46070 | n46074;
  assign n46076 = ~pi1634 & ~n37331;
  assign n46077 = ~pi0616 & ~n37700;
  assign n46078 = ~pi1634 & ~n46077;
  assign n46079 = pi0594 & n46077;
  assign n46080 = ~n46078 & ~n46079;
  assign n46081 = n37331 & ~n46080;
  assign po1943 = n46076 | n46081;
  assign n46083 = ~pi1635 & ~n37331;
  assign n46084 = pi0590 & n46052;
  assign n46085 = ~pi1635 & ~n46052;
  assign n46086 = ~n46084 & ~n46085;
  assign n46087 = n37331 & ~n46086;
  assign po1944 = n46083 | n46087;
  assign n46089 = ~pi1636 & ~n37331;
  assign n46090 = ~pi1636 & ~n46077;
  assign n46091 = pi0593 & n46077;
  assign n46092 = ~n46090 & ~n46091;
  assign n46093 = n37331 & ~n46092;
  assign po1945 = n46089 | n46093;
  assign n46095 = ~pi1637 & ~n37331;
  assign n46096 = ~pi1637 & ~n46077;
  assign n46097 = pi0603 & n46077;
  assign n46098 = ~n46096 & ~n46097;
  assign n46099 = n37331 & ~n46098;
  assign po1946 = n46095 | n46099;
  assign n46101 = ~pi1638 & ~n37331;
  assign n46102 = ~pi1638 & ~n46077;
  assign n46103 = pi0632 & n46077;
  assign n46104 = ~n46102 & ~n46103;
  assign n46105 = n37331 & ~n46104;
  assign po1947 = n46101 | n46105;
  assign n46107 = ~pi1639 & ~n37331;
  assign n46108 = ~pi1639 & ~n46077;
  assign n46109 = pi0571 & n46077;
  assign n46110 = ~n46108 & ~n46109;
  assign n46111 = n37331 & ~n46110;
  assign po1948 = n46107 | n46111;
  assign n46113 = pi0423 & n25623;
  assign n46114 = ~n24807 & n46113;
  assign n46115 = ~pi1640 & ~n25623;
  assign po1949 = n46114 | n46115;
  assign po1951 = ~pi3395 & ~pi3638;
  assign n46118 = ~pi0955 & po3448;
  assign n46119 = ~n31887 & ~n46118;
  assign n46120 = pi1447 & ~n46119;
  assign n46121 = pi3635 & n46120;
  assign po1952 = pi1642 | n46121;
  assign n46123 = pi1643 & ~n44510;
  assign n46124 = ~n44511 & ~n46123;
  assign po1953 = ~n44550 & n46124;
  assign n46126 = pi0900 & po2824;
  assign n46127 = ~pi1629 & n44478;
  assign n46128 = ~pi1687 & n46127;
  assign n46129 = pi1644 & ~n46128;
  assign n46130 = ~pi1644 & n46128;
  assign n46131 = ~n46129 & ~n46130;
  assign n46132 = po3311 & n46131;
  assign n46133 = ~pi1644 & ~po3311;
  assign n46134 = ~n46132 & ~n46133;
  assign n46135 = ~po2824 & ~n46134;
  assign po1954 = n46126 | n46135;
  assign n46137 = ~pi1645 & ~n41779;
  assign n46138 = ~pi1645 & pi1670;
  assign n46139 = pi1645 & ~pi1670;
  assign n46140 = ~n46138 & ~n46139;
  assign n46141 = n41779 & ~n46140;
  assign po1955 = n46137 | n46141;
  assign po1956 = pi1646 & ~n44550;
  assign n46144 = pi0424 & n25623;
  assign n46145 = ~n24807 & n46144;
  assign n46146 = ~pi1647 & ~n25623;
  assign po1957 = n46145 | n46146;
  assign n46148 = pi0964 & po2824;
  assign n46149 = n44478 & n44479;
  assign n46150 = n44477 & n46149;
  assign n46151 = ~pi1648 & n46150;
  assign n46152 = pi1648 & ~n46150;
  assign n46153 = ~n46151 & ~n46152;
  assign n46154 = po3311 & n46153;
  assign n46155 = ~pi1648 & ~po3311;
  assign n46156 = ~n46154 & ~n46155;
  assign n46157 = ~po2824 & ~n46156;
  assign po1958 = n46148 | n46157;
  assign n46159 = ~pi1691 & ~pi1693;
  assign n46160 = ~pi1643 & ~pi1692;
  assign n46161 = n46159 & n46160;
  assign n46162 = n44510 & n46161;
  assign n46163 = ~pi1649 & n46162;
  assign n46164 = pi1649 & ~n46162;
  assign n46165 = ~n46163 & ~n46164;
  assign po1959 = ~n44550 & n46165;
  assign n46167 = ~pi1650 & ~n37331;
  assign n46168 = ~pi1650 & ~n46077;
  assign n46169 = pi0590 & n46077;
  assign n46170 = ~n46168 & ~n46169;
  assign n46171 = n37331 & ~n46170;
  assign po1960 = n46167 | n46171;
  assign n46173 = ~pi1651 & ~n37331;
  assign n46174 = ~pi1651 & ~n46077;
  assign n46175 = pi0602 & n46077;
  assign n46176 = ~n46174 & ~n46175;
  assign n46177 = n37331 & ~n46176;
  assign po1961 = n46173 | n46177;
  assign n46179 = ~pi1652 & ~n37331;
  assign n46180 = ~pi1652 & ~n46077;
  assign n46181 = pi0572 & n46077;
  assign n46182 = ~n46180 & ~n46181;
  assign n46183 = n37331 & ~n46182;
  assign po1962 = n46179 | n46183;
  assign n46185 = ~pi1653 & ~n37331;
  assign n46186 = ~pi1653 & ~n46077;
  assign n46187 = pi0591 & n46077;
  assign n46188 = ~n46186 & ~n46187;
  assign n46189 = n37331 & ~n46188;
  assign po1963 = n46185 | n46189;
  assign n46191 = ~pi1654 & ~n37331;
  assign n46192 = ~pi1654 & ~n46077;
  assign n46193 = pi0592 & n46077;
  assign n46194 = ~n46192 & ~n46193;
  assign n46195 = n37331 & ~n46194;
  assign po1964 = n46191 | n46195;
  assign n46197 = ~pi1655 & ~n37331;
  assign n46198 = ~pi1655 & ~n46077;
  assign n46199 = pi0573 & n46077;
  assign n46200 = ~n46198 & ~n46199;
  assign n46201 = n37331 & ~n46200;
  assign po1965 = n46197 | n46201;
  assign n46203 = ~pi1656 & ~n37331;
  assign n46204 = ~pi1656 & ~n46077;
  assign n46205 = pi0595 & n46077;
  assign n46206 = ~n46204 & ~n46205;
  assign n46207 = n37331 & ~n46206;
  assign po1966 = n46203 | n46207;
  assign n46209 = ~pi1657 & ~n37331;
  assign n46210 = ~pi1657 & ~n46077;
  assign n46211 = pi0585 & n46077;
  assign n46212 = ~n46210 & ~n46211;
  assign n46213 = n37331 & ~n46212;
  assign po1967 = n46209 | n46213;
  assign n46215 = ~pi1658 & ~n37331;
  assign n46216 = pi0602 & n46052;
  assign n46217 = ~pi1658 & ~n46052;
  assign n46218 = ~n46216 & ~n46217;
  assign n46219 = n37331 & ~n46218;
  assign po1968 = n46215 | n46219;
  assign n46221 = ~pi1659 & ~n37331;
  assign n46222 = pi0572 & n46052;
  assign n46223 = ~pi1659 & ~n46052;
  assign n46224 = ~n46222 & ~n46223;
  assign n46225 = n37331 & ~n46224;
  assign po1969 = n46221 | n46225;
  assign n46227 = ~pi1660 & ~n37331;
  assign n46228 = pi0591 & n46052;
  assign n46229 = ~pi1660 & ~n46052;
  assign n46230 = ~n46228 & ~n46229;
  assign n46231 = n37331 & ~n46230;
  assign po1970 = n46227 | n46231;
  assign n46233 = ~pi1661 & ~n37331;
  assign n46234 = pi0603 & n46052;
  assign n46235 = ~pi1661 & ~n46052;
  assign n46236 = ~n46234 & ~n46235;
  assign n46237 = n37331 & ~n46236;
  assign po1971 = n46233 | n46237;
  assign n46239 = ~pi1662 & ~n37331;
  assign n46240 = pi0592 & n46052;
  assign n46241 = ~pi1662 & ~n46052;
  assign n46242 = ~n46240 & ~n46241;
  assign n46243 = n37331 & ~n46242;
  assign po1972 = n46239 | n46243;
  assign n46245 = ~pi1663 & ~n37331;
  assign n46246 = pi0573 & n46052;
  assign n46247 = ~pi1663 & ~n46052;
  assign n46248 = ~n46246 & ~n46247;
  assign n46249 = n37331 & ~n46248;
  assign po1973 = n46245 | n46249;
  assign n46251 = ~pi1664 & ~n37331;
  assign n46252 = pi0595 & n46052;
  assign n46253 = ~pi1664 & ~n46052;
  assign n46254 = ~n46252 & ~n46253;
  assign n46255 = n37331 & ~n46254;
  assign po1974 = n46251 | n46255;
  assign n46257 = ~pi1665 & ~n37331;
  assign n46258 = pi0585 & n46052;
  assign n46259 = ~pi1665 & ~n46052;
  assign n46260 = ~n46258 & ~n46259;
  assign n46261 = n37331 & ~n46260;
  assign po1975 = n46257 | n46261;
  assign n46263 = po3627 & n25623;
  assign n46264 = pi0420 & ~n8615;
  assign n46265 = n46263 & ~n46264;
  assign n46266 = ~pi1666 & n36128;
  assign po1976 = n46265 | n46266;
  assign n46268 = pi0420 & po3627;
  assign n46269 = n25623 & n46268;
  assign n46270 = ~n8615 & n46269;
  assign n46271 = ~pi1667 & n36128;
  assign po1977 = n46270 | n46271;
  assign n46273 = ~pi1668 & ~n42536;
  assign n46274 = ~pi1668 & ~n42540;
  assign n46275 = pi1668 & n42540;
  assign n46276 = ~n46274 & ~n46275;
  assign n46277 = n42536 & ~n46276;
  assign po1978 = n46273 | n46277;
  assign n46279 = ~pi1669 & ~n41779;
  assign n46280 = n45921 & n45922;
  assign n46281 = pi1669 & n46280;
  assign n46282 = ~pi1669 & ~n46280;
  assign n46283 = ~n46281 & ~n46282;
  assign n46284 = n41779 & ~n46283;
  assign po1979 = n46279 | n46284;
  assign n46286 = ~pi1670 & ~n41779;
  assign n46287 = pi1670 & n41779;
  assign po1980 = n46286 | n46287;
  assign n46289 = ~pi1671 & ~n41779;
  assign n46290 = ~pi1361 & ~pi1698;
  assign n46291 = n41768 & n46290;
  assign n46292 = ~pi1680 & n42446;
  assign n46293 = ~pi1679 & n46292;
  assign n46294 = ~pi1670 & n42447;
  assign n46295 = ~pi1645 & n46294;
  assign n46296 = ~pi1675 & n46295;
  assign n46297 = n46293 & n46296;
  assign n46298 = n46291 & n46297;
  assign n46299 = pi1671 & n46298;
  assign n46300 = ~pi1671 & ~n46298;
  assign n46301 = ~n46299 & ~n46300;
  assign n46302 = n41779 & ~n46301;
  assign po1981 = n46289 | n46302;
  assign n46304 = ~pi1672 & ~n41779;
  assign n46305 = n45920 & n45924;
  assign n46306 = n41759 & n46305;
  assign n46307 = n45925 & n46306;
  assign n46308 = ~pi1672 & ~n46307;
  assign n46309 = pi1672 & n46307;
  assign n46310 = ~n46308 & ~n46309;
  assign n46311 = n41779 & ~n46310;
  assign po1982 = n46304 | n46311;
  assign n46313 = ~pi1673 & ~n41779;
  assign n46314 = n46291 & n46293;
  assign n46315 = n42441 & n46314;
  assign n46316 = n42435 & n46315;
  assign n46317 = n46296 & n46316;
  assign n46318 = ~pi1673 & ~n46317;
  assign n46319 = pi1673 & n46317;
  assign n46320 = ~n46318 & ~n46319;
  assign n46321 = n41779 & ~n46320;
  assign po1983 = n46313 | n46321;
  assign n46323 = ~pi1674 & ~n41779;
  assign n46324 = n42434 & n46296;
  assign n46325 = n42442 & n46324;
  assign n46326 = n46316 & n46325;
  assign n46327 = pi1674 & n46326;
  assign n46328 = ~pi1674 & ~n46326;
  assign n46329 = ~n46327 & ~n46328;
  assign n46330 = n41779 & ~n46329;
  assign po1984 = n46323 | n46330;
  assign n46332 = ~pi1675 & ~n41779;
  assign n46333 = ~pi1675 & ~n41759;
  assign n46334 = pi1675 & n41759;
  assign n46335 = ~n46333 & ~n46334;
  assign n46336 = n41779 & ~n46335;
  assign po1985 = n46332 | n46336;
  assign n46338 = ~pi1676 & ~n41779;
  assign n46339 = pi1676 & n41760;
  assign n46340 = ~pi1676 & ~n41760;
  assign n46341 = ~n46339 & ~n46340;
  assign n46342 = n41779 & ~n46341;
  assign po1986 = n46338 | n46342;
  assign n46344 = ~pi1677 & ~n41779;
  assign n46345 = ~pi1677 & ~n41781;
  assign n46346 = pi1677 & n41781;
  assign n46347 = ~n46345 & ~n46346;
  assign n46348 = n41779 & ~n46347;
  assign po1987 = n46344 | n46348;
  assign n46350 = ~pi1678 & ~n41779;
  assign n46351 = ~pi1678 & ~n45921;
  assign n46352 = pi1678 & n45921;
  assign n46353 = ~n46351 & ~n46352;
  assign n46354 = n41779 & ~n46353;
  assign po1988 = n46350 | n46354;
  assign n46356 = ~pi1679 & ~n41779;
  assign n46357 = pi1679 & n42449;
  assign n46358 = ~pi1679 & ~n42449;
  assign n46359 = ~n46357 & ~n46358;
  assign n46360 = n41779 & ~n46359;
  assign po1989 = n46356 | n46360;
  assign n46362 = ~pi1680 & ~n41779;
  assign n46363 = pi1680 & n41782;
  assign n46364 = ~pi1680 & ~n41782;
  assign n46365 = ~n46363 & ~n46364;
  assign n46366 = n41779 & ~n46365;
  assign po1990 = n46362 | n46366;
  assign n46368 = pi1433 & ~n37393;
  assign n46369 = ~pi1605 & ~pi1681;
  assign n46370 = ~n31858 & ~n46369;
  assign n46371 = pi3641 & ~n46370;
  assign n46372 = ~pi1681 & ~pi3641;
  assign n46373 = ~n46371 & ~n46372;
  assign n46374 = n37390 & ~n46373;
  assign n46375 = ~n37392 & n46374;
  assign po1991 = n46368 | n46375;
  assign n46377 = pi0948 & po2823;
  assign n46378 = pi1683 & ~pi1684;
  assign n46379 = ~pi1702 & n42781;
  assign n46380 = pi1703 & n46379;
  assign n46381 = pi1607 & n46380;
  assign n46382 = n46378 & n46381;
  assign n46383 = ~pi1682 & n46382;
  assign n46384 = pi1682 & ~n46382;
  assign n46385 = ~n46383 & ~n46384;
  assign n46386 = po3310 & n46385;
  assign n46387 = ~pi1682 & ~po3310;
  assign n46388 = ~n46386 & ~n46387;
  assign n46389 = ~po2823 & ~n46388;
  assign po1992 = n46377 | n46389;
  assign n46391 = pi0949 & po2823;
  assign n46392 = n42781 & n42782;
  assign n46393 = n42780 & n46392;
  assign n46394 = ~pi1683 & n46393;
  assign n46395 = pi1683 & ~n46393;
  assign n46396 = ~n46394 & ~n46395;
  assign n46397 = po3310 & n46396;
  assign n46398 = ~pi1683 & ~po3310;
  assign n46399 = ~n46397 & ~n46398;
  assign n46400 = ~po2823 & ~n46399;
  assign po1993 = n46391 | n46400;
  assign n46402 = pi0891 & po2823;
  assign n46403 = pi1684 & n46379;
  assign n46404 = ~pi1684 & ~n46379;
  assign n46405 = ~n46403 & ~n46404;
  assign n46406 = po3310 & ~n46405;
  assign n46407 = ~pi1684 & ~po3310;
  assign n46408 = ~n46406 & ~n46407;
  assign n46409 = ~po2823 & n46408;
  assign po1994 = n46402 | n46409;
  assign po1995 = pi0890 & n36875;
  assign n46412 = pi0963 & po2824;
  assign n46413 = pi1648 & ~pi1687;
  assign n46414 = pi1644 & n46127;
  assign n46415 = pi1608 & n46414;
  assign n46416 = n46413 & n46415;
  assign n46417 = ~pi1686 & n46416;
  assign n46418 = pi1686 & ~n46416;
  assign n46419 = ~n46417 & ~n46418;
  assign n46420 = po3311 & n46419;
  assign n46421 = ~pi1686 & ~po3311;
  assign n46422 = ~n46420 & ~n46421;
  assign n46423 = ~po2824 & ~n46422;
  assign po1996 = n46412 | n46423;
  assign n46425 = pi0797 & po2824;
  assign n46426 = pi1687 & n46127;
  assign n46427 = ~pi1687 & ~n46127;
  assign n46428 = ~n46426 & ~n46427;
  assign n46429 = po3311 & ~n46428;
  assign n46430 = ~pi1687 & ~po3311;
  assign n46431 = ~n46429 & ~n46430;
  assign n46432 = ~po2824 & n46431;
  assign po1997 = n46425 | n46432;
  assign po1998 = pi0796 & n36967;
  assign n46435 = ~pi1850 & n46160;
  assign n46436 = ~pi1694 & n46435;
  assign n46437 = n46159 & n46436;
  assign n46438 = ~pi1646 & n46437;
  assign n46439 = ~pi1690 & n46438;
  assign n46440 = ~pi1649 & n46439;
  assign n46441 = ~pi1689 & n46440;
  assign n46442 = pi1689 & ~n46440;
  assign n46443 = ~n46441 & ~n46442;
  assign po1999 = ~n44550 & n46443;
  assign n46445 = n44511 & n46159;
  assign n46446 = ~pi1649 & n46445;
  assign n46447 = ~pi1692 & n46446;
  assign n46448 = ~pi1690 & n46447;
  assign n46449 = pi1690 & ~n46447;
  assign n46450 = ~n46448 & ~n46449;
  assign po2000 = ~n44550 & n46450;
  assign n46452 = ~pi1646 & n46436;
  assign n46453 = pi1691 & ~n46452;
  assign n46454 = ~pi1691 & n46452;
  assign n46455 = ~n46453 & ~n46454;
  assign po2001 = ~n44550 & n46455;
  assign n46457 = ~pi1692 & n44511;
  assign n46458 = pi1692 & ~n44511;
  assign n46459 = ~n46457 & ~n46458;
  assign po2002 = ~n44550 & n46459;
  assign n46461 = pi1693 & ~n44513;
  assign n46462 = ~n44514 & ~n46461;
  assign po2003 = ~n44550 & n46462;
  assign n46464 = pi1694 & ~n44509;
  assign n46465 = ~n44510 & ~n46464;
  assign po2004 = ~n44550 & n46465;
  assign n46467 = ~pi1695 & ~n42536;
  assign n46468 = ~pi1695 & ~n44556;
  assign n46469 = pi1695 & n44556;
  assign n46470 = ~n46468 & ~n46469;
  assign n46471 = n42536 & ~n46470;
  assign po2005 = n46467 | n46471;
  assign n46473 = ~pi1698 & ~n41779;
  assign n46474 = ~pi1698 & ~n46297;
  assign n46475 = pi1698 & n46297;
  assign n46476 = ~n46474 & ~n46475;
  assign n46477 = n41779 & ~n46476;
  assign po2006 = n46473 | n46477;
  assign n46479 = ~pi1699 & ~n41779;
  assign n46480 = ~pi1699 & ~n46296;
  assign n46481 = pi1699 & n46296;
  assign n46482 = ~n46480 & ~n46481;
  assign n46483 = n41779 & ~n46482;
  assign po2007 = n46479 | n46483;
  assign n46485 = ~pi1700 & ~n41779;
  assign n46486 = n45923 & n46280;
  assign n46487 = pi1700 & n46486;
  assign n46488 = ~pi1700 & ~n46486;
  assign n46489 = ~n46487 & ~n46488;
  assign n46490 = n41779 & ~n46489;
  assign po2008 = n46485 | n46490;
  assign n46492 = ~pi1701 & ~n41779;
  assign n46493 = ~pi1701 & ~n44609;
  assign n46494 = pi1701 & n44609;
  assign n46495 = ~n46493 & ~n46494;
  assign n46496 = n41779 & ~n46495;
  assign po2009 = n46492 | n46496;
  assign n46498 = pi0892 & po2823;
  assign n46499 = ~pi1702 & ~n42781;
  assign n46500 = pi1702 & n42781;
  assign n46501 = ~n46499 & ~n46500;
  assign n46502 = po3310 & ~n46501;
  assign n46503 = ~pi1702 & ~po3310;
  assign n46504 = ~n46502 & ~n46503;
  assign n46505 = ~po2823 & n46504;
  assign po2010 = n46498 | n46505;
  assign n46507 = pi0951 & po2823;
  assign n46508 = ~pi1684 & n46379;
  assign n46509 = pi1703 & ~n46508;
  assign n46510 = ~pi1703 & n46508;
  assign n46511 = ~n46509 & ~n46510;
  assign n46512 = po3310 & n46511;
  assign n46513 = ~pi1703 & ~po3310;
  assign n46514 = ~n46512 & ~n46513;
  assign n46515 = ~po2823 & ~n46514;
  assign po2011 = n46507 | n46515;
  assign n46517 = pi1432 & ~n37393;
  assign n46518 = ~pi1704 & ~n31858;
  assign n46519 = ~n31859 & ~n46518;
  assign n46520 = pi3641 & ~n46519;
  assign n46521 = ~pi1704 & ~pi3641;
  assign n46522 = ~n46520 & ~n46521;
  assign n46523 = n37390 & ~n46522;
  assign n46524 = ~n37392 & n46523;
  assign po2012 = n46517 | n46524;
  assign n46526 = n38906 & n44849;
  assign n46527 = ~pi1039 & n46526;
  assign n46528 = ~pi1034 & n46527;
  assign n46529 = ~n14403 & n46528;
  assign n46530 = pi1705 & ~n46528;
  assign po2013 = n46529 | n46530;
  assign n46532 = ~pi1012 & n11105;
  assign n46533 = pi1039 & n46532;
  assign n46534 = n38906 & n46533;
  assign n46535 = ~n13121 & n46534;
  assign n46536 = pi1706 & ~n46534;
  assign po2014 = n46535 | n46536;
  assign n46538 = ~pi1707 & ~n37331;
  assign n46539 = ~pi0616 & n37700;
  assign n46540 = ~pi1707 & ~n46539;
  assign n46541 = pi0603 & n46539;
  assign n46542 = ~n46540 & ~n46541;
  assign n46543 = n37331 & ~n46542;
  assign po2015 = n46538 | n46543;
  assign n46545 = ~pi1708 & ~n37331;
  assign n46546 = ~pi1708 & ~n46539;
  assign n46547 = pi0571 & n46539;
  assign n46548 = ~n46546 & ~n46547;
  assign n46549 = n37331 & ~n46548;
  assign po2016 = n46545 | n46549;
  assign n46551 = ~pi1709 & ~n37331;
  assign n46552 = ~pi1709 & ~n46052;
  assign n46553 = pi0578 & n46052;
  assign n46554 = ~n46552 & ~n46553;
  assign n46555 = n37331 & ~n46554;
  assign po2017 = n46551 | n46555;
  assign n46557 = ~pi1710 & ~n37331;
  assign n46558 = pi0616 & ~n37700;
  assign n46559 = pi0594 & n46558;
  assign n46560 = ~pi1710 & ~n46558;
  assign n46561 = ~n46559 & ~n46560;
  assign n46562 = n37331 & ~n46561;
  assign po2018 = n46557 | n46562;
  assign n46564 = ~pi1711 & ~n37331;
  assign n46565 = pi0632 & n46558;
  assign n46566 = ~pi1711 & ~n46558;
  assign n46567 = ~n46565 & ~n46566;
  assign n46568 = n37331 & ~n46567;
  assign po2019 = n46564 | n46568;
  assign n46570 = ~pi1712 & ~n37331;
  assign n46571 = pi0590 & n46558;
  assign n46572 = ~pi1712 & ~n46558;
  assign n46573 = ~n46571 & ~n46572;
  assign n46574 = n37331 & ~n46573;
  assign po2020 = n46570 | n46574;
  assign n46576 = ~pi1797 & n15594;
  assign n46577 = ~pi3191 & ~n9352;
  assign n46578 = ~n46576 & n46577;
  assign n46579 = ~n15594 & ~n15599;
  assign n46580 = ~n46578 & ~n46579;
  assign n46581 = ~n15592 & ~n15597;
  assign n46582 = n46578 & ~n46581;
  assign n46583 = ~n46580 & ~n46582;
  assign n46584 = pi3191 & ~pi3291;
  assign n46585 = pi2383 & n46584;
  assign n46586 = n46578 & ~n46585;
  assign n46587 = pi2383 & ~n16000;
  assign n46588 = ~n9352 & ~n46587;
  assign n46589 = ~pi1797 & n46588;
  assign n46590 = ~n46585 & n46589;
  assign n46591 = ~n46586 & ~n46590;
  assign n46592 = ~n46583 & ~n46591;
  assign n46593 = pi1713 & n46591;
  assign po2021 = n46592 | n46593;
  assign n46595 = ~pi2555 & ~n15426;
  assign n46596 = ~n26062 & n46595;
  assign n46597 = pi1714 & n26062;
  assign n46598 = ~n46596 & ~n46597;
  assign n46599 = pi2555 & ~n26062;
  assign n46600 = ~pi1897 & n46599;
  assign po2022 = ~n46598 | n46600;
  assign n46602 = ~pi1868 & ~pi1894;
  assign n46603 = ~pi1896 & n46602;
  assign n46604 = ~pi1871 & n46603;
  assign n46605 = ~pi1895 & n46604;
  assign n46606 = n40572 & n46605;
  assign n46607 = ~pi1740 & n46606;
  assign n46608 = ~pi1435 & n46607;
  assign n46609 = n40581 & n46608;
  assign n46610 = ~pi1016 & n46609;
  assign n46611 = ~pi1872 & n46610;
  assign n46612 = ~pi1715 & n46611;
  assign n46613 = pi1715 & ~n46611;
  assign n46614 = ~n46612 & ~n46613;
  assign po2023 = n40651 & n46614;
  assign n46616 = ~n13398 & n46534;
  assign n46617 = pi1716 & ~n46534;
  assign po2024 = n46616 | n46617;
  assign n46619 = ~n13988 & n46534;
  assign n46620 = pi1717 & ~n46534;
  assign po2025 = n46619 | n46620;
  assign n46622 = ~n12415 & n46534;
  assign n46623 = pi1718 & ~n46534;
  assign po2026 = n46622 | n46623;
  assign n46625 = ~n14816 & n46534;
  assign n46626 = pi1719 & ~n46534;
  assign po2027 = n46625 | n46626;
  assign n46628 = ~n15115 & n46534;
  assign n46629 = pi1720 & ~n46534;
  assign po2028 = n46628 | n46629;
  assign n46631 = ~n12061 & n46534;
  assign n46632 = pi1721 & ~n46534;
  assign po2029 = n46631 | n46632;
  assign n46634 = ~n17368 & n46534;
  assign n46635 = pi1722 & ~n46534;
  assign po2030 = n46634 | n46635;
  assign n46637 = ~n17199 & n46534;
  assign n46638 = pi1723 & ~n46534;
  assign po2031 = n46637 | n46638;
  assign n46640 = ~n15426 & n46534;
  assign n46641 = pi1724 & ~n46534;
  assign po2032 = n46640 | n46641;
  assign n46643 = ~n14403 & n46534;
  assign n46644 = pi1725 & ~n46534;
  assign po2033 = n46643 | n46644;
  assign n46646 = ~n11181 & n46534;
  assign n46647 = pi1726 & ~n46534;
  assign po2034 = n46646 | n46647;
  assign n46649 = pi0609 & n9636;
  assign n46650 = n39499 & n46649;
  assign n46651 = pi1039 & n11105;
  assign n46652 = pi1012 & n46651;
  assign n46653 = n46650 & n46652;
  assign n46654 = ~n12726 & n46653;
  assign n46655 = pi1727 & ~n46653;
  assign po2035 = n46654 | n46655;
  assign n46657 = ~n13701 & n46653;
  assign n46658 = pi1728 & ~n46653;
  assign po2036 = n46657 | n46658;
  assign n46660 = ~n13121 & n46653;
  assign n46661 = pi1729 & ~n46653;
  assign po2037 = n46660 | n46661;
  assign n46663 = ~n13398 & n46653;
  assign n46664 = pi1730 & ~n46653;
  assign po2038 = n46663 | n46664;
  assign n46666 = ~n13988 & n46653;
  assign n46667 = pi1731 & ~n46653;
  assign po2039 = n46666 | n46667;
  assign n46669 = ~n12415 & n46653;
  assign n46670 = pi1732 & ~n46653;
  assign po2040 = n46669 | n46670;
  assign n46672 = ~n14816 & n46653;
  assign n46673 = pi1733 & ~n46653;
  assign po2041 = n46672 | n46673;
  assign n46675 = ~n15115 & n46653;
  assign n46676 = pi1734 & ~n46653;
  assign po2042 = n46675 | n46676;
  assign n46678 = ~n12061 & n46653;
  assign n46679 = pi1735 & ~n46653;
  assign po2043 = n46678 | n46679;
  assign n46681 = ~n15426 & n46653;
  assign n46682 = pi1736 & ~n46653;
  assign po2044 = n46681 | n46682;
  assign n46684 = ~n14403 & n46653;
  assign n46685 = pi1737 & ~n46653;
  assign po2045 = n46684 | n46685;
  assign n46687 = ~n11181 & n46653;
  assign n46688 = pi1738 & ~n46653;
  assign po2046 = n46687 | n46688;
  assign n46690 = ~pi1739 & ~n40651;
  assign n46691 = pi1739 & n40651;
  assign po2047 = n46690 | n46691;
  assign n46693 = ~pi1740 & n40577;
  assign n46694 = pi1740 & ~n40577;
  assign n46695 = ~n46693 & ~n46694;
  assign po2048 = n40651 & n46695;
  assign n46697 = ~pi2555 & ~n13701;
  assign n46698 = ~n26062 & n46697;
  assign n46699 = pi1741 & n26062;
  assign n46700 = ~n46698 & ~n46699;
  assign po2049 = n46600 | ~n46700;
  assign n46702 = ~pi2555 & ~n12726;
  assign n46703 = ~n26062 & n46702;
  assign n46704 = pi1742 & n26062;
  assign n46705 = ~n46703 & ~n46704;
  assign po2050 = n46600 | ~n46705;
  assign n46707 = ~pi2555 & ~n9825;
  assign n46708 = ~n26062 & n46707;
  assign n46709 = pi1743 & n26062;
  assign n46710 = ~n46708 & ~n46709;
  assign po2051 = n46600 | ~n46710;
  assign n46712 = ~pi2555 & ~n10608;
  assign n46713 = ~n26062 & n46712;
  assign n46714 = pi1744 & n26062;
  assign n46715 = ~n46713 & ~n46714;
  assign po2052 = n46600 | ~n46715;
  assign n46717 = ~pi2555 & ~n14403;
  assign n46718 = ~n26062 & n46717;
  assign n46719 = pi1745 & n26062;
  assign n46720 = ~n46718 & ~n46719;
  assign po2053 = n46600 | ~n46720;
  assign n46722 = ~pi1746 & ~n40741;
  assign n46723 = pi1746 & n40741;
  assign po2054 = n46722 | n46723;
  assign n46725 = ~pi1911 & ~pi1912;
  assign n46726 = ~pi1876 & n46725;
  assign n46727 = ~pi1914 & n46726;
  assign n46728 = ~pi1913 & n46727;
  assign n46729 = n40662 & n46728;
  assign n46730 = ~pi1748 & n46729;
  assign n46731 = ~pi1448 & n46730;
  assign n46732 = n40671 & n46731;
  assign n46733 = ~pi1018 & n46732;
  assign n46734 = ~pi1915 & n46733;
  assign n46735 = ~pi1747 & n46734;
  assign n46736 = pi1747 & ~n46734;
  assign n46737 = ~n46735 & ~n46736;
  assign po2055 = n40741 & n46737;
  assign n46739 = ~pi1748 & n40667;
  assign n46740 = pi1748 & ~n40667;
  assign n46741 = ~n46739 & ~n46740;
  assign po2056 = n40741 & n46741;
  assign n46743 = n39349 & n46650;
  assign n46744 = ~n9825 & n46743;
  assign n46745 = pi1749 & ~n46743;
  assign po2057 = n46744 | n46745;
  assign n46747 = ~n10608 & n46743;
  assign n46748 = pi1750 & ~n46743;
  assign po2058 = n46747 | n46748;
  assign n46750 = ~n13121 & n46743;
  assign n46751 = pi1751 & ~n46743;
  assign po2059 = n46750 | n46751;
  assign n46753 = ~n13398 & n46743;
  assign n46754 = pi1752 & ~n46743;
  assign po2060 = n46753 | n46754;
  assign n46756 = ~n13988 & n46743;
  assign n46757 = pi1753 & ~n46743;
  assign po2061 = n46756 | n46757;
  assign n46759 = ~n12415 & n46743;
  assign n46760 = pi1754 & ~n46743;
  assign po2062 = n46759 | n46760;
  assign n46762 = ~n14816 & n46743;
  assign n46763 = pi1755 & ~n46743;
  assign po2063 = n46762 | n46763;
  assign n46765 = ~n15115 & n46743;
  assign n46766 = pi1756 & ~n46743;
  assign po2064 = n46765 | n46766;
  assign n46768 = ~n12061 & n46743;
  assign n46769 = pi1757 & ~n46743;
  assign po2065 = n46768 | n46769;
  assign n46771 = ~n17368 & n46743;
  assign n46772 = pi1758 & ~n46743;
  assign po2066 = n46771 | n46772;
  assign n46774 = ~n17199 & n46743;
  assign n46775 = pi1759 & ~n46743;
  assign po2067 = n46774 | n46775;
  assign n46777 = ~n11181 & n46743;
  assign n46778 = pi1760 & ~n46743;
  assign po2068 = n46777 | n46778;
  assign n46780 = n39353 & n46650;
  assign n46781 = ~n9825 & n46780;
  assign n46782 = pi1761 & ~n46780;
  assign po2069 = n46781 | n46782;
  assign n46784 = ~n10608 & n46780;
  assign n46785 = pi1762 & ~n46780;
  assign po2070 = n46784 | n46785;
  assign n46787 = ~n13398 & n46780;
  assign n46788 = pi1763 & ~n46780;
  assign po2071 = n46787 | n46788;
  assign n46790 = ~n13988 & n46780;
  assign n46791 = pi1764 & ~n46780;
  assign po2072 = n46790 | n46791;
  assign n46793 = ~n12415 & n46780;
  assign n46794 = pi1765 & ~n46780;
  assign po2073 = n46793 | n46794;
  assign n46796 = ~n15115 & n46780;
  assign n46797 = pi1766 & ~n46780;
  assign po2074 = n46796 | n46797;
  assign n46799 = ~n12061 & n46780;
  assign n46800 = pi1767 & ~n46780;
  assign po2075 = n46799 | n46800;
  assign n46802 = ~n17368 & n46780;
  assign n46803 = pi1768 & ~n46780;
  assign po2076 = n46802 | n46803;
  assign n46805 = ~n11181 & n46780;
  assign n46806 = pi1769 & ~n46780;
  assign po2077 = n46805 | n46806;
  assign n46808 = pi3572 & pi3645;
  assign n46809 = n32780 & ~n34595;
  assign n46810 = n46808 & n46809;
  assign n46811 = pi0975 & n8592;
  assign n46812 = ~n34595 & n46811;
  assign n46813 = ~pi1770 & ~n46812;
  assign n46814 = ~pi1770 & ~pi1855;
  assign n46815 = ~n32784 & ~n46814;
  assign n46816 = n46812 & ~n46815;
  assign n46817 = ~n46813 & ~n46816;
  assign n46818 = ~n46810 & ~n46817;
  assign n46819 = pi1923 & n46810;
  assign po2078 = n46818 | n46819;
  assign n46821 = ~pi1771 & ~n46808;
  assign n46822 = pi3440 & pi3507;
  assign n46823 = n46821 & ~n46822;
  assign po2079 = n39531 & ~n46823;
  assign n46825 = n11105 & n38906;
  assign n46826 = pi1012 & n46825;
  assign n46827 = ~pi1039 & n46826;
  assign n46828 = ~n12726 & n46827;
  assign n46829 = pi1772 & ~n46827;
  assign po2081 = n46828 | n46829;
  assign n46831 = ~n13701 & n46827;
  assign n46832 = pi1773 & ~n46827;
  assign po2082 = n46831 | n46832;
  assign n46834 = ~n13121 & n46827;
  assign n46835 = pi1774 & ~n46827;
  assign po2083 = n46834 | n46835;
  assign n46837 = ~n13398 & n46827;
  assign n46838 = pi1775 & ~n46827;
  assign po2084 = n46837 | n46838;
  assign n46840 = ~n13988 & n46827;
  assign n46841 = pi1776 & ~n46827;
  assign po2085 = n46840 | n46841;
  assign n46843 = ~n12415 & n46827;
  assign n46844 = pi1777 & ~n46827;
  assign po2086 = n46843 | n46844;
  assign n46846 = ~n14816 & n46827;
  assign n46847 = pi1778 & ~n46827;
  assign po2087 = n46846 | n46847;
  assign n46849 = ~n15115 & n46827;
  assign n46850 = pi1779 & ~n46827;
  assign po2088 = n46849 | n46850;
  assign n46852 = ~n12061 & n46827;
  assign n46853 = pi1780 & ~n46827;
  assign po2089 = n46852 | n46853;
  assign n46855 = ~n17199 & n46827;
  assign n46856 = pi1781 & ~n46827;
  assign po2090 = n46855 | n46856;
  assign n46858 = ~n9825 & n46827;
  assign n46859 = pi1782 & ~n46827;
  assign po2091 = n46858 | n46859;
  assign n46861 = ~n10608 & n46827;
  assign n46862 = pi1783 & ~n46827;
  assign po2092 = n46861 | n46862;
  assign n46864 = ~n15426 & n46827;
  assign n46865 = pi1784 & ~n46827;
  assign po2093 = n46864 | n46865;
  assign n46867 = ~n14403 & n46827;
  assign n46868 = pi1785 & ~n46827;
  assign po2094 = n46867 | n46868;
  assign n46870 = ~n11181 & n46827;
  assign n46871 = pi1786 & ~n46827;
  assign po2095 = n46870 | n46871;
  assign n46873 = ~n8561 & ~n44983;
  assign n46874 = pi1787 & ~n46873;
  assign n46875 = n44999 & n46874;
  assign n46876 = pi3257 & n8358;
  assign n46877 = ~pi2779 & ~n46876;
  assign n46878 = ~n44999 & ~n46877;
  assign po2096 = n46875 | n46878;
  assign n46880 = ~pi1788 & ~n42536;
  assign n46881 = ~pi2824 & ~pi3247;
  assign n46882 = ~pi1851 & n46881;
  assign n46883 = ~pi2510 & n46882;
  assign n46884 = n42538 & n46883;
  assign n46885 = ~pi3290 & n46884;
  assign n46886 = ~pi1668 & n46885;
  assign n46887 = ~pi1380 & n46886;
  assign n46888 = ~pi1788 & ~n46887;
  assign n46889 = pi1788 & n46887;
  assign n46890 = ~n46888 & ~n46889;
  assign n46891 = n42536 & ~n46890;
  assign po2097 = n46880 | n46891;
  assign n46893 = ~pi1789 & ~n25623;
  assign po2098 = n44810 | n46893;
  assign n46895 = ~n12061 & n25547;
  assign n46896 = ~n16568 & ~n25547;
  assign n46897 = ~n46895 & ~n46896;
  assign n46898 = ~n30537 & ~n46897;
  assign n46899 = ~n11006 & n30537;
  assign n46900 = ~n46898 & ~n46899;
  assign n46901 = n30536 & ~n46900;
  assign n46902 = pi1790 & ~n30536;
  assign po2099 = n46901 | n46902;
  assign n46904 = ~n17105 & ~n25547;
  assign n46905 = ~n17199 & n25547;
  assign n46906 = ~n46904 & ~n46905;
  assign n46907 = ~n30537 & n46906;
  assign n46908 = n9556 & n30537;
  assign n46909 = ~n46907 & ~n46908;
  assign n46910 = n30536 & n46909;
  assign n46911 = pi1791 & ~n30536;
  assign po2100 = n46910 | n46911;
  assign n46913 = ~n17199 & n46528;
  assign n46914 = pi1792 & ~n46528;
  assign po2101 = n46913 | n46914;
  assign n46916 = ~pi0411 & ~pi0412;
  assign n46917 = ~pi0408 & n46916;
  assign n46918 = ~pi0413 & n46917;
  assign n46919 = n16037 & ~n46918;
  assign n46920 = n24813 & n46919;
  assign n46921 = pi0408 & n46920;
  assign n46922 = pi0413 & ~n25526;
  assign n46923 = ~pi0411 & pi0413;
  assign n46924 = ~n46922 & ~n46923;
  assign n46925 = pi0411 & n25526;
  assign n46926 = pi0412 & ~pi0413;
  assign n46927 = n46925 & n46926;
  assign n46928 = n46924 & ~n46927;
  assign n46929 = ~pi0412 & pi0413;
  assign n46930 = n46928 & ~n46929;
  assign n46931 = n46921 & ~n46930;
  assign n46932 = ~pi1793 & ~n46920;
  assign po2102 = n46931 | n46932;
  assign n46934 = ~pi0412 & ~pi0413;
  assign n46935 = n46925 & n46934;
  assign n46936 = n46924 & ~n46935;
  assign n46937 = pi0412 & pi0413;
  assign n46938 = n46936 & ~n46937;
  assign n46939 = n46921 & ~n46938;
  assign n46940 = ~pi1794 & ~n46920;
  assign po2103 = n46939 | n46940;
  assign n46942 = pi0411 & pi0413;
  assign n46943 = ~n46922 & ~n46942;
  assign n46944 = ~pi0411 & pi0425;
  assign n46945 = pi0406 & n46944;
  assign n46946 = n46926 & n46945;
  assign n46947 = n46943 & ~n46946;
  assign n46948 = ~n46929 & n46947;
  assign n46949 = n46921 & ~n46948;
  assign n46950 = ~pi1795 & ~n46920;
  assign po2104 = n46949 | n46950;
  assign n46952 = n46934 & n46945;
  assign n46953 = n46943 & ~n46952;
  assign n46954 = ~n46937 & n46953;
  assign n46955 = n46921 & ~n46954;
  assign n46956 = ~pi1796 & ~n46920;
  assign po2105 = n46955 | n46956;
  assign n46958 = pi1797 & n46591;
  assign n46959 = pi1797 & n15599;
  assign n46960 = ~pi1797 & ~n15599;
  assign n46961 = ~n46959 & ~n46960;
  assign n46962 = ~n46578 & ~n46961;
  assign n46963 = pi1797 & ~n15594;
  assign n46964 = ~n46576 & ~n46963;
  assign n46965 = n46578 & n46964;
  assign n46966 = ~n46962 & ~n46965;
  assign n46967 = ~n46591 & n46966;
  assign po2106 = n46958 | n46967;
  assign n46969 = pi1798 & n46591;
  assign n46970 = ~pi1798 & ~n46591;
  assign po2107 = n46969 | n46970;
  assign n46972 = ~pi1798 & ~n46581;
  assign n46973 = ~pi3330 & n46972;
  assign n46974 = pi1799 & ~n46972;
  assign n46975 = ~n46973 & ~n46974;
  assign n46976 = n46586 & ~n46975;
  assign n46977 = pi1799 & ~n46586;
  assign po2108 = n46976 | n46977;
  assign n46979 = ~pi1798 & n46581;
  assign n46980 = ~pi3330 & n46979;
  assign n46981 = pi1800 & ~n46979;
  assign n46982 = ~n46980 & ~n46981;
  assign n46983 = n46586 & ~n46982;
  assign n46984 = pi1800 & ~n46586;
  assign po2109 = n46983 | n46984;
  assign n46986 = ~pi1801 & ~n37331;
  assign n46987 = pi0602 & n46558;
  assign n46988 = ~pi1801 & ~n46558;
  assign n46989 = ~n46987 & ~n46988;
  assign n46990 = n37331 & ~n46989;
  assign po2110 = n46986 | n46990;
  assign n46992 = ~pi1802 & ~n37331;
  assign n46993 = pi0571 & n46558;
  assign n46994 = ~pi1802 & ~n46558;
  assign n46995 = ~n46993 & ~n46994;
  assign n46996 = n37331 & ~n46995;
  assign po2111 = n46992 | n46996;
  assign n46998 = ~pi1803 & ~n37331;
  assign n46999 = pi0572 & n46558;
  assign n47000 = ~pi1803 & ~n46558;
  assign n47001 = ~n46999 & ~n47000;
  assign n47002 = n37331 & ~n47001;
  assign po2112 = n46998 | n47002;
  assign n47004 = ~pi1804 & ~n37331;
  assign n47005 = pi0591 & n46558;
  assign n47006 = ~pi1804 & ~n46558;
  assign n47007 = ~n47005 & ~n47006;
  assign n47008 = n37331 & ~n47007;
  assign po2113 = n47004 | n47008;
  assign n47010 = ~pi1805 & ~n37331;
  assign n47011 = pi0603 & n46558;
  assign n47012 = ~pi1805 & ~n46558;
  assign n47013 = ~n47011 & ~n47012;
  assign n47014 = n37331 & ~n47013;
  assign po2114 = n47010 | n47014;
  assign n47016 = ~pi1806 & ~n37331;
  assign n47017 = pi0592 & n46558;
  assign n47018 = ~pi1806 & ~n46558;
  assign n47019 = ~n47017 & ~n47018;
  assign n47020 = n37331 & ~n47019;
  assign po2115 = n47016 | n47020;
  assign n47022 = ~pi1807 & ~n37331;
  assign n47023 = pi0573 & n46558;
  assign n47024 = ~pi1807 & ~n46558;
  assign n47025 = ~n47023 & ~n47024;
  assign n47026 = n37331 & ~n47025;
  assign po2116 = n47022 | n47026;
  assign n47028 = ~pi1808 & ~n37331;
  assign n47029 = pi0593 & n46558;
  assign n47030 = ~pi1808 & ~n46558;
  assign n47031 = ~n47029 & ~n47030;
  assign n47032 = n37331 & ~n47031;
  assign po2117 = n47028 | n47032;
  assign n47034 = ~pi1809 & ~n37331;
  assign n47035 = pi0595 & n46558;
  assign n47036 = ~pi1809 & ~n46558;
  assign n47037 = ~n47035 & ~n47036;
  assign n47038 = n37331 & ~n47037;
  assign po2118 = n47034 | n47038;
  assign n47040 = ~pi1810 & ~n37331;
  assign n47041 = pi0585 & n46558;
  assign n47042 = ~pi1810 & ~n46558;
  assign n47043 = ~n47041 & ~n47042;
  assign n47044 = n37331 & ~n47043;
  assign po2119 = n47040 | n47044;
  assign n47046 = ~pi1811 & ~n37331;
  assign n47047 = pi0578 & n46077;
  assign n47048 = ~pi1811 & ~n46077;
  assign n47049 = ~n47047 & ~n47048;
  assign n47050 = n37331 & ~n47049;
  assign po2120 = n47046 | n47050;
  assign n47052 = ~pi1812 & ~n37331;
  assign n47053 = ~pi1812 & ~n46539;
  assign n47054 = pi0590 & n46539;
  assign n47055 = ~n47053 & ~n47054;
  assign n47056 = n37331 & ~n47055;
  assign po2121 = n47052 | n47056;
  assign n47058 = ~pi1813 & ~n37331;
  assign n47059 = ~pi1813 & ~n46539;
  assign n47060 = pi0602 & n46539;
  assign n47061 = ~n47059 & ~n47060;
  assign n47062 = n37331 & ~n47061;
  assign po2122 = n47058 | n47062;
  assign n47064 = ~pi1814 & ~n37331;
  assign n47065 = ~pi1814 & ~n46539;
  assign n47066 = pi0572 & n46539;
  assign n47067 = ~n47065 & ~n47066;
  assign n47068 = n37331 & ~n47067;
  assign po2123 = n47064 | n47068;
  assign n47070 = ~pi1815 & ~n37331;
  assign n47071 = ~pi1815 & ~n46539;
  assign n47072 = pi0591 & n46539;
  assign n47073 = ~n47071 & ~n47072;
  assign n47074 = n37331 & ~n47073;
  assign po2124 = n47070 | n47074;
  assign n47076 = ~pi1816 & ~n37331;
  assign n47077 = ~pi1816 & ~n46539;
  assign n47078 = pi0592 & n46539;
  assign n47079 = ~n47077 & ~n47078;
  assign n47080 = n37331 & ~n47079;
  assign po2125 = n47076 | n47080;
  assign n47082 = ~pi1817 & ~n37331;
  assign n47083 = ~pi1817 & ~n46539;
  assign n47084 = pi0632 & n46539;
  assign n47085 = ~n47083 & ~n47084;
  assign n47086 = n37331 & ~n47085;
  assign po2126 = n47082 | n47086;
  assign n47088 = ~pi1818 & ~n37331;
  assign n47089 = ~pi1818 & ~n46539;
  assign n47090 = pi0573 & n46539;
  assign n47091 = ~n47089 & ~n47090;
  assign n47092 = n37331 & ~n47091;
  assign po2127 = n47088 | n47092;
  assign n47094 = ~pi1819 & ~n37331;
  assign n47095 = ~pi1819 & ~n46539;
  assign n47096 = pi0595 & n46539;
  assign n47097 = ~n47095 & ~n47096;
  assign n47098 = n37331 & ~n47097;
  assign po2128 = n47094 | n47098;
  assign n47100 = ~pi1820 & ~n37331;
  assign n47101 = ~pi1820 & ~n46539;
  assign n47102 = pi0594 & n46539;
  assign n47103 = ~n47101 & ~n47102;
  assign n47104 = n37331 & ~n47103;
  assign po2129 = n47100 | n47104;
  assign n47106 = ~pi1821 & ~n37331;
  assign n47107 = ~pi1821 & ~n46539;
  assign n47108 = pi0585 & n46539;
  assign n47109 = ~n47107 & ~n47108;
  assign n47110 = n37331 & ~n47109;
  assign po2130 = n47106 | n47110;
  assign n47112 = ~pi3443 & ~pi3536;
  assign n47113 = pi3374 & ~n47112;
  assign n47114 = pi1822 & n47113;
  assign n47115 = pi3217 & ~n47114;
  assign n47116 = pi2019 & ~po3627;
  assign po2131 = n47115 & ~n47116;
  assign n47118 = n15793 & ~n33813;
  assign n47119 = ~pi1823 & n33813;
  assign n47120 = ~n47118 & ~n47119;
  assign po2132 = po3627 & ~n47120;
  assign n47122 = n9373 & n35814;
  assign n47123 = pi0405 & n47122;
  assign n47124 = ~pi0421 & n47123;
  assign n47125 = pi0405 & ~pi0421;
  assign n47126 = n34038 & n47125;
  assign n47127 = ~n47124 & ~n47126;
  assign n47128 = ~n24813 & n47127;
  assign n47129 = ~pi0419 & n8609;
  assign n47130 = pi0418 & n47129;
  assign n47131 = pi0420 & n47130;
  assign n47132 = n47128 & ~n47131;
  assign n47133 = ~n15589 & n47132;
  assign n47134 = ~n9377 & n47133;
  assign n47135 = ~n8561 & ~n47134;
  assign n47136 = ~pi1824 & n8561;
  assign n47137 = ~n47135 & ~n47136;
  assign po2133 = po3627 & ~n47137;
  assign n47139 = pi1930 & ~n33813;
  assign n47140 = ~n15929 & n47139;
  assign n47141 = pi1825 & ~n47139;
  assign n47142 = ~n47140 & ~n47141;
  assign po2134 = po3627 & n47142;
  assign n47144 = ~n15991 & n47139;
  assign n47145 = pi1826 & ~n47139;
  assign n47146 = ~n47144 & ~n47145;
  assign po2135 = po3627 & n47146;
  assign n47148 = ~n15992 & n47139;
  assign n47149 = pi1827 & ~n47139;
  assign n47150 = ~n47148 & ~n47149;
  assign po2136 = po3627 & n47150;
  assign n47152 = ~n12726 & n46528;
  assign n47153 = pi1828 & ~n46528;
  assign po2137 = n47152 | n47153;
  assign n47155 = ~n13701 & n46528;
  assign n47156 = pi1829 & ~n46528;
  assign po2138 = n47155 | n47156;
  assign n47158 = ~n13121 & n46528;
  assign n47159 = pi1830 & ~n46528;
  assign po2139 = n47158 | n47159;
  assign n47161 = ~n13398 & n46528;
  assign n47162 = pi1831 & ~n46528;
  assign po2140 = n47161 | n47162;
  assign n47164 = ~n13988 & n46528;
  assign n47165 = pi1832 & ~n46528;
  assign po2141 = n47164 | n47165;
  assign n47167 = ~n12415 & n46528;
  assign n47168 = pi1833 & ~n46528;
  assign po2142 = n47167 | n47168;
  assign n47170 = ~n15115 & n46528;
  assign n47171 = pi1834 & ~n46528;
  assign po2143 = n47170 | n47171;
  assign n47173 = ~n17368 & n46528;
  assign n47174 = pi1835 & ~n46528;
  assign po2144 = n47173 | n47174;
  assign n47176 = ~n9825 & n46528;
  assign n47177 = pi1836 & ~n46528;
  assign po2145 = n47176 | n47177;
  assign n47179 = ~n10608 & n46528;
  assign n47180 = pi1837 & ~n46528;
  assign po2146 = n47179 | n47180;
  assign n47182 = ~n15426 & n46528;
  assign n47183 = pi1838 & ~n46528;
  assign po2147 = n47182 | n47183;
  assign n47185 = ~n11181 & n46528;
  assign n47186 = pi1839 & ~n46528;
  assign po2148 = n47185 | n47186;
  assign n47188 = pi1840 & ~pi1861;
  assign n47189 = ~n8596 & ~n47188;
  assign n47190 = ~n36181 & ~n39886;
  assign n47191 = n47189 & n47190;
  assign n47192 = ~pi1840 & ~n47190;
  assign n47193 = ~n47191 & ~n47192;
  assign po2149 = ~n36189 & n47193;
  assign n47195 = ~n14816 & n38320;
  assign n47196 = ~pi1841 & n41165;
  assign n47197 = pi1841 & ~n41165;
  assign n47198 = ~n47196 & ~n47197;
  assign n47199 = ~n36181 & ~n47198;
  assign n47200 = ~pi1841 & n36181;
  assign n47201 = ~n47199 & ~n47200;
  assign n47202 = ~n38320 & n47201;
  assign po2150 = n47195 | n47202;
  assign n47204 = pi0498 & n35314;
  assign n47205 = pi0551 & ~pi0563;
  assign n47206 = pi0497 & n35322;
  assign n47207 = ~pi0553 & n47206;
  assign n47208 = ~pi0504 & n47207;
  assign n47209 = ~pi0552 & n47208;
  assign n47210 = n47205 & n47209;
  assign n47211 = n47204 & n47210;
  assign n47212 = ~n38373 & n47211;
  assign n47213 = pi1842 & ~n47211;
  assign po2151 = n47212 | n47213;
  assign n47215 = ~pi0498 & n35314;
  assign n47216 = n47210 & n47215;
  assign n47217 = ~n38373 & n47216;
  assign n47218 = pi1843 & ~n47216;
  assign po2152 = n47217 | n47218;
  assign n47220 = ~pi0559 & pi0560;
  assign n47221 = pi0501 & n35425;
  assign n47222 = ~pi0561 & n47221;
  assign n47223 = ~pi0502 & n47222;
  assign n47224 = ~pi0564 & n47223;
  assign n47225 = n47220 & n47224;
  assign n47226 = n35417 & n47225;
  assign n47227 = pi0503 & n47226;
  assign n47228 = ~n38357 & n47227;
  assign n47229 = pi1844 & ~n47227;
  assign po2153 = n47228 | n47229;
  assign n47231 = ~pi0503 & n35417;
  assign n47232 = n47225 & n47231;
  assign n47233 = ~n38357 & n47232;
  assign n47234 = pi1845 & ~n47232;
  assign po2154 = n47233 | n47234;
  assign n47236 = pi0952 & po2823;
  assign n47237 = pi1846 & pi1847;
  assign n47238 = ~n42781 & ~n47237;
  assign n47239 = po3310 & n47238;
  assign n47240 = ~pi1846 & ~po3310;
  assign n47241 = ~n47239 & ~n47240;
  assign n47242 = ~po2823 & n47241;
  assign po2155 = n47236 | n47242;
  assign n47244 = pi0953 & po2823;
  assign n47245 = pi1847 & po3310;
  assign n47246 = ~pi1847 & ~po3310;
  assign n47247 = ~n47245 & ~n47246;
  assign n47248 = ~po2823 & n47247;
  assign po2156 = n47244 | n47248;
  assign n47250 = pi0967 & po2824;
  assign n47251 = pi1848 & po3311;
  assign n47252 = ~pi1848 & ~po3311;
  assign n47253 = ~n47251 & ~n47252;
  assign n47254 = ~po2824 & n47253;
  assign po2157 = n47250 | n47254;
  assign n47256 = pi0966 & po2824;
  assign n47257 = pi1848 & pi1849;
  assign n47258 = ~n44478 & ~n47257;
  assign n47259 = po3311 & n47258;
  assign n47260 = ~pi1849 & ~po3311;
  assign n47261 = ~n47259 & ~n47260;
  assign n47262 = ~po2824 & n47261;
  assign po2158 = n47256 | n47262;
  assign n47264 = pi1646 & ~pi1850;
  assign n47265 = ~pi1646 & pi1850;
  assign n47266 = ~n47264 & ~n47265;
  assign po2159 = ~n44550 & ~n47266;
  assign n47268 = ~pi1851 & ~n42536;
  assign n47269 = pi1851 & n41248;
  assign n47270 = ~pi1851 & ~n41248;
  assign n47271 = ~n47269 & ~n47270;
  assign n47272 = n42536 & ~n47271;
  assign po2160 = n47268 | n47272;
  assign n47274 = ~n14816 & n46528;
  assign n47275 = pi1852 & ~n46528;
  assign po2161 = n47274 | n47275;
  assign n47277 = ~n12061 & n46528;
  assign n47278 = pi1853 & ~n46528;
  assign po2162 = n47277 | n47278;
  assign n47280 = ~n17199 & n46780;
  assign n47281 = pi1854 & ~n46780;
  assign po2163 = n47280 | n47281;
  assign n47283 = ~pi1855 & ~n46812;
  assign n47284 = pi1855 & n46812;
  assign n47285 = ~n47283 & ~n47284;
  assign n47286 = ~n46810 & ~n47285;
  assign n47287 = pi1924 & n46810;
  assign po2164 = n47286 | n47287;
  assign n47289 = ~pi1422 & ~pi3645;
  assign n47290 = ~pi3572 & n47289;
  assign n47291 = ~pi1856 & ~n47290;
  assign n47292 = pi1856 & n47290;
  assign n47293 = ~n47291 & ~n47292;
  assign po2165 = ~n41525 | n47293;
  assign n47295 = ~n13121 & n46780;
  assign n47296 = pi1857 & ~n46780;
  assign po2166 = n47295 | n47296;
  assign n47298 = ~n14816 & n46780;
  assign n47299 = pi1858 & ~n46780;
  assign po2167 = n47298 | n47299;
  assign n47301 = ~pi1859 & ~n37331;
  assign n47302 = ~pi1859 & ~n46539;
  assign n47303 = pi0593 & n46539;
  assign n47304 = ~n47302 & ~n47303;
  assign n47305 = n37331 & ~n47304;
  assign po2168 = n47301 | n47305;
  assign po2169 = ~pi3419 & pi3562;
  assign n47308 = pi0783 & pi3099;
  assign n47309 = n39883 & ~n47308;
  assign n47310 = ~n8599 & ~n16214;
  assign n47311 = ~pi1860 & n47310;
  assign n47312 = ~n10780 & n47311;
  assign n47313 = n47309 & ~n47312;
  assign n47314 = ~n10773 & ~n34654;
  assign n47315 = ~n8586 & n47314;
  assign n47316 = pi3590 & ~n47315;
  assign n47317 = pi3585 & n47316;
  assign n47318 = n47308 & n47317;
  assign n47319 = ~n47313 & ~n47318;
  assign po2170 = pi1860 | ~n47319;
  assign n47321 = pi1861 & n47190;
  assign n47322 = ~pi1861 & ~n47190;
  assign n47323 = ~n47321 & ~n47322;
  assign po2171 = ~n36189 & n47323;
  assign n47325 = n9667 & n38906;
  assign n47326 = ~n12061 & n47325;
  assign n47327 = pi1862 & ~n47325;
  assign po2172 = n47326 | n47327;
  assign n47329 = ~pi1863 & ~n47139;
  assign n47330 = pi0036 & n47139;
  assign po2173 = n47329 | n47330;
  assign n47332 = ~pi1864 & ~n37331;
  assign n47333 = pi0578 & n46539;
  assign n47334 = ~pi1864 & ~n46539;
  assign n47335 = ~n47333 & ~n47334;
  assign n47336 = n37331 & ~n47335;
  assign po2174 = n47332 | n47336;
  assign n47338 = ~pi1865 & ~n37331;
  assign n47339 = ~pi1865 & ~n46558;
  assign n47340 = pi0578 & n46558;
  assign n47341 = ~n47339 & ~n47340;
  assign n47342 = n37331 & ~n47341;
  assign po2175 = n47338 | n47342;
  assign n47344 = ~n17199 & n30466;
  assign n47345 = pi1866 & n26062;
  assign n47346 = ~n46600 & ~n47345;
  assign po2176 = n47344 | ~n47346;
  assign n47348 = ~n13121 & n30466;
  assign n47349 = pi1867 & n26062;
  assign n47350 = ~n46600 & ~n47349;
  assign po2177 = n47348 | ~n47350;
  assign n47352 = pi1868 & pi1896;
  assign n47353 = ~n40573 & ~n47352;
  assign po2178 = n40651 & n47353;
  assign n47355 = ~n17199 & n47325;
  assign n47356 = pi1869 & ~n47325;
  assign po2179 = n47355 | n47356;
  assign n47358 = ~pi1870 & n46605;
  assign n47359 = pi1870 & ~n46605;
  assign n47360 = ~n47358 & ~n47359;
  assign po2180 = n40651 & n47360;
  assign n47362 = pi1871 & ~n40574;
  assign n47363 = ~n40575 & ~n47362;
  assign po2181 = n40651 & n47363;
  assign n47365 = ~pi1872 & n46608;
  assign n47366 = pi1872 & ~n46608;
  assign n47367 = ~n47365 & ~n47366;
  assign po2182 = n40651 & n47367;
  assign n47369 = ~n11181 & n47325;
  assign n47370 = pi1873 & ~n47325;
  assign po2183 = n47369 | n47370;
  assign n47372 = ~n10608 & n47325;
  assign n47373 = pi1874 & ~n47325;
  assign po2184 = n47372 | n47373;
  assign n47375 = n31776 & ~n37392;
  assign n47376 = pi3444 & ~n31779;
  assign po2185 = n47375 & n47376;
  assign po2186 = pi1876 & n40741;
  assign n47379 = ~n12726 & n46534;
  assign n47380 = pi1877 & ~n46534;
  assign po2187 = n47379 | n47380;
  assign n47382 = ~n13701 & n46534;
  assign n47383 = pi1878 & ~n46534;
  assign po2188 = n47382 | n47383;
  assign n47385 = ~n9825 & n46534;
  assign n47386 = pi1879 & ~n46534;
  assign po2189 = n47385 | n47386;
  assign n47388 = ~n10608 & n46534;
  assign n47389 = pi1880 & ~n46534;
  assign po2190 = n47388 | n47389;
  assign n47391 = n38277 & n38897;
  assign n47392 = n9641 & n47391;
  assign n47393 = n9649 & n47392;
  assign po3455 = n11105 & n47393;
  assign n47395 = pi0609 & po3455;
  assign n47396 = ~n15426 & n47395;
  assign n47397 = ~pi1881 & ~n47395;
  assign po2191 = n47396 | n47397;
  assign po2192 = po0493 & ~n37392;
  assign po2193 = ~pi1882 | pi2814;
  assign n47401 = ~n13701 & n47325;
  assign n47402 = pi1883 & ~n47325;
  assign po2194 = n47401 | n47402;
  assign n47404 = ~n13121 & n47325;
  assign n47405 = pi1884 & ~n47325;
  assign po2195 = n47404 | n47405;
  assign n47407 = ~n13398 & n47325;
  assign n47408 = pi1885 & ~n47325;
  assign po2196 = n47407 | n47408;
  assign n47410 = ~n12415 & n47325;
  assign n47411 = pi1886 & ~n47325;
  assign po2197 = n47410 | n47411;
  assign n47413 = ~n14816 & n47325;
  assign n47414 = pi1887 & ~n47325;
  assign po2198 = n47413 | n47414;
  assign n47416 = ~n15115 & n47325;
  assign n47417 = pi1888 & ~n47325;
  assign po2199 = n47416 | n47417;
  assign n47419 = ~n17368 & n47325;
  assign n47420 = pi1889 & ~n47325;
  assign po2200 = n47419 | n47420;
  assign n47422 = ~n9825 & n47325;
  assign n47423 = pi1890 & ~n47325;
  assign po2201 = n47422 | n47423;
  assign n47425 = ~n14403 & n47325;
  assign n47426 = pi1891 & ~n47325;
  assign po2202 = n47425 | n47426;
  assign n47428 = ~n15426 & n47325;
  assign n47429 = pi1892 & ~n47325;
  assign po2203 = n47428 | n47429;
  assign n47431 = ~pi1893 & n41383;
  assign n47432 = pi1893 & ~n41383;
  assign n47433 = ~n47431 & ~n47432;
  assign po2204 = n40651 & n47433;
  assign n47435 = pi1894 & ~n40575;
  assign n47436 = ~n41382 & ~n47435;
  assign po2205 = n40651 & n47436;
  assign n47438 = pi1895 & ~n40573;
  assign n47439 = ~n40574 & ~n47438;
  assign po2206 = n40651 & n47439;
  assign po2207 = pi1896 & n40651;
  assign n47442 = ~n17368 & n30466;
  assign n47443 = pi1897 & n26062;
  assign n47444 = ~n46600 & ~n47443;
  assign po2208 = n47442 | ~n47444;
  assign n47446 = n38906 & n41509;
  assign n47447 = ~n13701 & n47446;
  assign n47448 = pi1898 & ~n47446;
  assign po2209 = n47447 | n47448;
  assign n47450 = ~n13398 & n47446;
  assign n47451 = pi1899 & ~n47446;
  assign po2210 = n47450 | n47451;
  assign n47453 = ~n12415 & n47446;
  assign n47454 = pi1900 & ~n47446;
  assign po2211 = n47453 | n47454;
  assign n47456 = ~n14816 & n47446;
  assign n47457 = pi1901 & ~n47446;
  assign po2212 = n47456 | n47457;
  assign n47459 = ~n15115 & n47446;
  assign n47460 = pi1902 & ~n47446;
  assign po2213 = n47459 | n47460;
  assign n47462 = ~n17368 & n47446;
  assign n47463 = pi1903 & ~n47446;
  assign po2214 = n47462 | n47463;
  assign n47465 = ~n17199 & n47446;
  assign n47466 = pi1904 & ~n47446;
  assign po2215 = n47465 | n47466;
  assign n47468 = ~n9825 & n47446;
  assign n47469 = pi1905 & ~n47446;
  assign po2216 = n47468 | n47469;
  assign n47471 = ~n15426 & n47446;
  assign n47472 = pi1906 & ~n47446;
  assign po2217 = n47471 | n47472;
  assign n47474 = ~n11181 & n47446;
  assign n47475 = pi1907 & ~n47446;
  assign po2218 = n47474 | n47475;
  assign n47477 = ~n17368 & n44885;
  assign n47478 = pi1908 & ~n44885;
  assign po2219 = n47477 | n47478;
  assign n47480 = ~n10608 & n44885;
  assign n47481 = pi1909 & ~n44885;
  assign po2220 = n47480 | n47481;
  assign n47483 = ~pi1910 & n41489;
  assign n47484 = pi1910 & ~n41489;
  assign n47485 = ~n47483 & ~n47484;
  assign po2221 = n40741 & n47485;
  assign n47487 = pi1911 & ~n40665;
  assign n47488 = ~n41488 & ~n47487;
  assign po2222 = n40741 & n47488;
  assign n47490 = pi1876 & pi1912;
  assign n47491 = ~n40663 & ~n47490;
  assign po2223 = n40741 & n47491;
  assign n47493 = pi1913 & ~n40663;
  assign n47494 = ~n40664 & ~n47493;
  assign po2224 = n40741 & n47494;
  assign n47496 = pi1914 & ~n40664;
  assign n47497 = ~n40665 & ~n47496;
  assign po2225 = n40741 & n47497;
  assign n47499 = ~pi1915 & n46731;
  assign n47500 = pi1915 & ~n46731;
  assign n47501 = ~n47499 & ~n47500;
  assign po2226 = n40741 & n47501;
  assign n47503 = ~pi1916 & n46728;
  assign n47504 = pi1916 & ~n46728;
  assign n47505 = ~n47503 & ~n47504;
  assign po2227 = n40741 & n47505;
  assign n47507 = ~n17199 & n44885;
  assign n47508 = pi1917 & ~n44885;
  assign po2228 = n47507 | n47508;
  assign n47510 = n38906 & n46652;
  assign n47511 = ~n12726 & n47510;
  assign n47512 = pi1918 & ~n47510;
  assign po2229 = n47511 | n47512;
  assign n47514 = ~n13701 & n47510;
  assign n47515 = pi1919 & ~n47510;
  assign po2230 = n47514 | n47515;
  assign n47517 = ~n13988 & n47325;
  assign n47518 = pi1920 & ~n47325;
  assign po2231 = n47517 | n47518;
  assign n47520 = ~n13121 & n47510;
  assign n47521 = pi1921 & ~n47510;
  assign po2232 = n47520 | n47521;
  assign n47523 = ~n13398 & n47510;
  assign n47524 = pi1922 & ~n47510;
  assign po2233 = n47523 | n47524;
  assign n47526 = ~n13988 & n47510;
  assign n47527 = pi1923 & ~n47510;
  assign po2234 = n47526 | n47527;
  assign n47529 = ~n12415 & n47510;
  assign n47530 = pi1924 & ~n47510;
  assign po2235 = n47529 | n47530;
  assign n47532 = ~n14816 & n47510;
  assign n47533 = pi1925 & ~n47510;
  assign po2236 = n47532 | n47533;
  assign n47535 = ~n15115 & n47510;
  assign n47536 = pi1926 & ~n47510;
  assign po2237 = n47535 | n47536;
  assign n47538 = ~n12061 & n47510;
  assign n47539 = pi1927 & ~n47510;
  assign po2238 = n47538 | n47539;
  assign n47541 = ~n17368 & n47510;
  assign n47542 = pi1928 & ~n47510;
  assign po2239 = n47541 | n47542;
  assign n47544 = ~n17199 & n47510;
  assign n47545 = pi1929 & ~n47510;
  assign po2240 = n47544 | n47545;
  assign n47547 = ~n9825 & n47510;
  assign n47548 = pi1930 & ~n47510;
  assign po2241 = n47547 | n47548;
  assign n47550 = ~n15426 & n47510;
  assign n47551 = pi1931 & ~n47510;
  assign po2242 = n47550 | n47551;
  assign n47553 = ~n14403 & n47510;
  assign n47554 = pi1932 & ~n47510;
  assign po2243 = n47553 | n47554;
  assign n47556 = ~n11181 & n47510;
  assign n47557 = pi1933 & ~n47510;
  assign po2244 = n47556 | n47557;
  assign n47559 = n10767 & ~n10769;
  assign n47560 = ~po3855 & n25532;
  assign n47561 = ~n9881 & n47560;
  assign n47562 = n15462 & ~n47561;
  assign n47563 = ~n47559 & n47562;
  assign n47564 = pi1934 & n47561;
  assign po2245 = n47563 | n47564;
  assign n47566 = ~n34595 & n46822;
  assign n47567 = pi1918 & n47566;
  assign n47568 = ~pi3147 & ~n34595;
  assign n47569 = ~pi1935 & ~n39525;
  assign n47570 = ~n39526 & ~n47569;
  assign n47571 = n47568 & ~n47570;
  assign n47572 = ~pi1935 & ~n47568;
  assign n47573 = ~n47571 & ~n47572;
  assign n47574 = ~n47566 & ~n47573;
  assign po2246 = n47567 | n47574;
  assign n47576 = pi1921 & n47566;
  assign n47577 = ~pi1936 & n47568;
  assign n47578 = pi1936 & ~n47568;
  assign n47579 = ~n47577 & ~n47578;
  assign n47580 = ~n47566 & n47579;
  assign po2247 = n47576 | n47580;
  assign n47582 = ~pi1937 & ~n32784;
  assign n47583 = pi1937 & n32784;
  assign n47584 = ~n47582 & ~n47583;
  assign n47585 = n46812 & ~n47584;
  assign n47586 = ~pi1937 & ~n46812;
  assign n47587 = ~n47585 & ~n47586;
  assign n47588 = ~n46810 & ~n47587;
  assign n47589 = pi1922 & n46810;
  assign po2248 = n47588 | n47589;
  assign n47591 = n39499 & n44851;
  assign n47592 = n46649 & n47591;
  assign n47593 = ~n13121 & n47592;
  assign n47594 = pi1938 & ~n47592;
  assign po2249 = n47593 | n47594;
  assign n47596 = ~n13398 & n47592;
  assign n47597 = pi1939 & ~n47592;
  assign po2250 = n47596 | n47597;
  assign n47599 = ~n13988 & n47592;
  assign n47600 = pi1940 & ~n47592;
  assign po2251 = n47599 | n47600;
  assign n47602 = ~n12415 & n47592;
  assign n47603 = pi1941 & ~n47592;
  assign po2252 = n47602 | n47603;
  assign n47605 = ~n14816 & n47592;
  assign n47606 = pi1942 & ~n47592;
  assign po2253 = n47605 | n47606;
  assign n47608 = ~n15115 & n47592;
  assign n47609 = pi1943 & ~n47592;
  assign po2254 = n47608 | n47609;
  assign n47611 = ~n12061 & n47592;
  assign n47612 = pi1944 & ~n47592;
  assign po2255 = n47611 | n47612;
  assign n47614 = ~n11181 & n47592;
  assign n47615 = pi1945 & ~n47592;
  assign po2256 = n47614 | n47615;
  assign n47617 = ~n8307 & ~n44983;
  assign n47618 = n8232 & ~po0014;
  assign n47619 = pi3256 & n47618;
  assign n47620 = n47617 & n47619;
  assign n47621 = pi3698 & n47620;
  assign n47622 = pi1946 & ~n47620;
  assign po2257 = n47621 | n47622;
  assign n47624 = pi3697 & n47620;
  assign n47625 = pi1947 & ~n47620;
  assign po2258 = n47624 | n47625;
  assign n47627 = pi3696 & n47620;
  assign n47628 = pi1948 & ~n47620;
  assign po2259 = n47627 | n47628;
  assign n47630 = pi3695 & n47620;
  assign n47631 = pi1949 & ~n47620;
  assign po2260 = n47630 | n47631;
  assign n47633 = pi3694 & n47620;
  assign n47634 = pi1950 & ~n47620;
  assign po2261 = n47633 | n47634;
  assign n47636 = pi3693 & n47620;
  assign n47637 = pi1951 & ~n47620;
  assign po2262 = n47636 | n47637;
  assign n47639 = ~n12726 & n47325;
  assign n47640 = pi1952 & ~n47325;
  assign po2263 = n47639 | n47640;
  assign n47642 = n16037 & ~n24818;
  assign n47643 = n46268 & n47642;
  assign n47644 = ~n8615 & n47643;
  assign n47645 = ~pi1953 & n36128;
  assign po2264 = n47644 | n47645;
  assign n47647 = ~pi1954 & ~n47139;
  assign n47648 = pi0007 & n47139;
  assign po2265 = n47647 | n47648;
  assign n47650 = ~n12726 & n25547;
  assign n47651 = ~n16855 & ~n25547;
  assign n47652 = ~n47650 & ~n47651;
  assign n47653 = ~n30537 & n47652;
  assign n47654 = n13578 & n30537;
  assign n47655 = ~n47653 & ~n47654;
  assign n47656 = n30536 & n47655;
  assign n47657 = pi1955 & ~n30536;
  assign po2266 = n47656 | n47657;
  assign n47659 = ~n13701 & n25547;
  assign n47660 = ~n16819 & ~n25547;
  assign n47661 = ~n47659 & ~n47660;
  assign n47662 = ~n30537 & n47661;
  assign n47663 = n12984 & n30537;
  assign n47664 = ~n47662 & ~n47663;
  assign n47665 = n30536 & n47664;
  assign n47666 = pi1956 & ~n30536;
  assign po2267 = n47665 | n47666;
  assign n47668 = ~n13121 & n25547;
  assign n47669 = ~n16784 & ~n25547;
  assign n47670 = ~n47668 & ~n47669;
  assign n47671 = ~n30537 & n47670;
  assign n47672 = n13168 & n30537;
  assign n47673 = ~n47671 & ~n47672;
  assign n47674 = n30536 & n47673;
  assign n47675 = pi1957 & ~n30536;
  assign po2268 = n47674 | n47675;
  assign n47677 = ~n13398 & n25547;
  assign n47678 = ~n16748 & ~n25547;
  assign n47679 = ~n47677 & ~n47678;
  assign n47680 = ~n30537 & n47679;
  assign n47681 = n13816 & n30537;
  assign n47682 = ~n47680 & ~n47681;
  assign n47683 = n30536 & n47682;
  assign n47684 = pi1958 & ~n30536;
  assign po2269 = n47683 | n47684;
  assign n47686 = ~n13988 & n25547;
  assign n47687 = ~n16712 & ~n25547;
  assign n47688 = ~n47686 & ~n47687;
  assign n47689 = ~n30537 & n47688;
  assign n47690 = n12243 & n30537;
  assign n47691 = ~n47689 & ~n47690;
  assign n47692 = n30536 & n47691;
  assign n47693 = pi1959 & ~n30536;
  assign po2270 = n47692 | n47693;
  assign n47695 = ~n12415 & n25547;
  assign n47696 = ~n16676 & ~n25547;
  assign n47697 = ~n47695 & ~n47696;
  assign n47698 = ~n30537 & n47697;
  assign n47699 = n14644 & n30537;
  assign n47700 = ~n47698 & ~n47699;
  assign n47701 = n30536 & n47700;
  assign n47702 = pi1960 & ~n30536;
  assign po2271 = n47701 | n47702;
  assign n47704 = ~n14816 & n25547;
  assign n47705 = ~n16640 & ~n25547;
  assign n47706 = ~n47704 & ~n47705;
  assign n47707 = ~n30537 & n47706;
  assign n47708 = n14877 & n30537;
  assign n47709 = ~n47707 & ~n47708;
  assign n47710 = n30536 & n47709;
  assign n47711 = pi1961 & ~n30536;
  assign po2272 = n47710 | n47711;
  assign n47713 = ~n15115 & n25547;
  assign n47714 = ~n16604 & ~n25547;
  assign n47715 = ~n47713 & ~n47714;
  assign n47716 = ~n30537 & n47715;
  assign n47717 = n11829 & n30537;
  assign n47718 = ~n47716 & ~n47717;
  assign n47719 = n30536 & n47718;
  assign n47720 = pi1962 & ~n30536;
  assign po2273 = n47719 | n47720;
  assign n47722 = ~n17368 & n25547;
  assign n47723 = ~n17397 & ~n25547;
  assign n47724 = ~n47722 & ~n47723;
  assign n47725 = ~n30537 & n47724;
  assign n47726 = n17031 & n30537;
  assign n47727 = ~n47725 & ~n47726;
  assign n47728 = n30536 & n47727;
  assign n47729 = pi1963 & ~n30536;
  assign po2274 = n47728 | n47729;
  assign n47731 = ~n9825 & n25547;
  assign n47732 = ~n16999 & ~n25547;
  assign n47733 = ~n47731 & ~n47732;
  assign n47734 = ~n30537 & n47733;
  assign n47735 = n10482 & n30537;
  assign n47736 = ~n47734 & ~n47735;
  assign n47737 = n30536 & n47736;
  assign n47738 = pi1964 & ~n30536;
  assign po2275 = n47737 | n47738;
  assign n47740 = ~n10608 & n25547;
  assign n47741 = ~n16963 & ~n25547;
  assign n47742 = ~n47740 & ~n47741;
  assign n47743 = ~n30537 & n47742;
  assign n47744 = n15294 & n30537;
  assign n47745 = ~n47743 & ~n47744;
  assign n47746 = n30536 & n47745;
  assign n47747 = pi1965 & ~n30536;
  assign po2276 = n47746 | n47747;
  assign n47749 = ~n15426 & n25547;
  assign n47750 = ~n16927 & ~n25547;
  assign n47751 = ~n47749 & ~n47750;
  assign n47752 = ~n30537 & n47751;
  assign n47753 = n14277 & n30537;
  assign n47754 = ~n47752 & ~n47753;
  assign n47755 = n30536 & n47754;
  assign n47756 = pi1966 & ~n30536;
  assign po2277 = n47755 | n47756;
  assign n47758 = ~n14403 & n25547;
  assign n47759 = ~n16891 & ~n25547;
  assign n47760 = ~n47758 & ~n47759;
  assign n47761 = ~n30537 & n47760;
  assign n47762 = n12542 & n30537;
  assign n47763 = ~n47761 & ~n47762;
  assign n47764 = n30536 & n47763;
  assign n47765 = pi1967 & ~n30536;
  assign po2278 = n47764 | n47765;
  assign n47767 = ~pi1968 & ~n47139;
  assign n47768 = pi0034 & n47139;
  assign po2279 = n47767 | n47768;
  assign n47770 = ~pi1969 & ~n47139;
  assign n47771 = pi0005 & n47139;
  assign po2280 = n47770 | n47771;
  assign n47773 = ~pi1970 & ~n47139;
  assign n47774 = pi0003 & n47139;
  assign po2281 = n47773 | n47774;
  assign n47776 = ~n8561 & n9373;
  assign n47777 = ~pi0420 & n47776;
  assign n47778 = ~pi0421 & n47777;
  assign n47779 = pi0419 & n47778;
  assign n47780 = ~pi0405 & n47779;
  assign n47781 = ~pi0419 & ~n8561;
  assign n47782 = n9373 & n47781;
  assign n47783 = ~pi0421 & n47782;
  assign n47784 = pi0420 & n47783;
  assign n47785 = pi0405 & n47784;
  assign n47786 = ~n47780 & ~n47785;
  assign n47787 = ~n47642 & n47786;
  assign n47788 = ~pi1971 & n47787;
  assign n47789 = pi0421 & ~n47787;
  assign po2282 = n47788 | n47789;
  assign n47791 = ~pi1972 & n47787;
  assign n47792 = pi0405 & ~n47787;
  assign po2283 = n47791 | n47792;
  assign n47794 = ~pi1973 & n47787;
  assign n47795 = pi0422 & ~n47787;
  assign po2284 = n47794 | n47795;
  assign n47797 = ~pi1974 & n47787;
  assign n47798 = pi0423 & ~n47787;
  assign po2285 = n47797 | n47798;
  assign n47800 = ~pi1975 & n47787;
  assign n47801 = pi0424 & ~n47787;
  assign po2286 = n47800 | n47801;
  assign n47803 = pi0995 & ~pi3426;
  assign n47804 = ~n9399 & ~n47803;
  assign n47805 = ~n9403 & n47804;
  assign n47806 = ~n9404 & ~n47805;
  assign n47807 = ~n37833 & n47806;
  assign n47808 = pi1976 & ~n47806;
  assign po2287 = n47807 | n47808;
  assign n47810 = ~n37586 & n47806;
  assign n47811 = pi1977 & ~n47806;
  assign po2288 = n47810 | n47811;
  assign n47813 = ~n37850 & n47806;
  assign n47814 = pi1978 & ~n47806;
  assign po2289 = n47813 | n47814;
  assign n47816 = ~n37867 & n47806;
  assign n47817 = pi1979 & ~n47806;
  assign po2290 = n47816 | n47817;
  assign n47819 = ~n37884 & n47806;
  assign n47820 = pi1980 & ~n47806;
  assign po2291 = n47819 | n47820;
  assign n47822 = ~n37901 & n47806;
  assign n47823 = pi1981 & ~n47806;
  assign po2292 = n47822 | n47823;
  assign n47825 = ~n37918 & n47806;
  assign n47826 = pi1982 & ~n47806;
  assign po2293 = n47825 | n47826;
  assign n47828 = ~n37935 & n47806;
  assign n47829 = pi1983 & ~n47806;
  assign po2294 = n47828 | n47829;
  assign n47831 = ~n37613 & n47806;
  assign n47832 = pi1984 & ~n47806;
  assign po2295 = n47831 | n47832;
  assign n47834 = ~n37952 & n47806;
  assign n47835 = pi1985 & ~n47806;
  assign po2296 = n47834 | n47835;
  assign n47837 = pi3398 & n46972;
  assign n47838 = pi1986 & ~n46972;
  assign n47839 = ~n47837 & ~n47838;
  assign n47840 = n46586 & ~n47839;
  assign n47841 = pi1986 & ~n46586;
  assign po2297 = n47840 | n47841;
  assign n47843 = pi3520 & n46972;
  assign n47844 = pi1987 & ~n46972;
  assign n47845 = ~n47843 & ~n47844;
  assign n47846 = n46586 & ~n47845;
  assign n47847 = pi1987 & ~n46586;
  assign po2298 = n47846 | n47847;
  assign n47849 = pi3392 & n46972;
  assign n47850 = pi1988 & ~n46972;
  assign n47851 = ~n47849 & ~n47850;
  assign n47852 = n46586 & ~n47851;
  assign n47853 = pi1988 & ~n46586;
  assign po2299 = n47852 | n47853;
  assign n47855 = ~pi3394 & n46972;
  assign n47856 = pi1989 & ~n46972;
  assign n47857 = ~n47855 & ~n47856;
  assign n47858 = n46586 & ~n47857;
  assign n47859 = pi1989 & ~n46586;
  assign po2300 = n47858 | n47859;
  assign n47861 = ~pi1990 & ~n46586;
  assign n47862 = pi2514 & n46972;
  assign n47863 = ~pi1990 & ~n46972;
  assign n47864 = ~n47862 & ~n47863;
  assign n47865 = n46586 & ~n47864;
  assign po2301 = n47861 | n47865;
  assign n47867 = pi3512 & n46972;
  assign n47868 = pi1991 & ~n46972;
  assign n47869 = ~n47867 & ~n47868;
  assign n47870 = n46586 & ~n47869;
  assign n47871 = pi1991 & ~n46586;
  assign po2302 = n47870 | n47871;
  assign n47873 = pi3513 & n46972;
  assign n47874 = pi1992 & ~n46972;
  assign n47875 = ~n47873 & ~n47874;
  assign n47876 = n46586 & ~n47875;
  assign n47877 = pi1992 & ~n46586;
  assign po2303 = n47876 | n47877;
  assign n47879 = pi3514 & n46972;
  assign n47880 = pi1993 & ~n46972;
  assign n47881 = ~n47879 & ~n47880;
  assign n47882 = n46586 & ~n47881;
  assign n47883 = pi1993 & ~n46586;
  assign po2304 = n47882 | n47883;
  assign n47885 = pi3518 & n46972;
  assign n47886 = pi1994 & ~n46972;
  assign n47887 = ~n47885 & ~n47886;
  assign n47888 = n46586 & ~n47887;
  assign n47889 = pi1994 & ~n46586;
  assign po2305 = n47888 | n47889;
  assign n47891 = pi3516 & n46972;
  assign n47892 = pi1995 & ~n46972;
  assign n47893 = ~n47891 & ~n47892;
  assign n47894 = n46586 & ~n47893;
  assign n47895 = pi1995 & ~n46586;
  assign po2306 = n47894 | n47895;
  assign n47897 = pi1798 & ~n46581;
  assign n47898 = ~pi3330 & n47897;
  assign n47899 = pi1996 & ~n47897;
  assign n47900 = ~n47898 & ~n47899;
  assign n47901 = n46586 & ~n47900;
  assign n47902 = pi1996 & ~n46586;
  assign po2307 = n47901 | n47902;
  assign n47904 = ~pi3394 & n47897;
  assign n47905 = pi1997 & ~n47897;
  assign n47906 = ~n47904 & ~n47905;
  assign n47907 = n46586 & ~n47906;
  assign n47908 = pi1997 & ~n46586;
  assign po2308 = n47907 | n47908;
  assign n47910 = pi3511 & n46979;
  assign n47911 = pi1998 & ~n46979;
  assign n47912 = ~n47910 & ~n47911;
  assign n47913 = n46586 & ~n47912;
  assign n47914 = pi1998 & ~n46586;
  assign po2309 = n47913 | n47914;
  assign n47916 = pi3392 & n46979;
  assign n47917 = pi1999 & ~n46979;
  assign n47918 = ~n47916 & ~n47917;
  assign n47919 = n46586 & ~n47918;
  assign n47920 = pi1999 & ~n46586;
  assign po2310 = n47919 | n47920;
  assign n47922 = ~pi3394 & n46979;
  assign n47923 = pi2000 & ~n46979;
  assign n47924 = ~n47922 & ~n47923;
  assign n47925 = n46586 & ~n47924;
  assign n47926 = pi2000 & ~n46586;
  assign po2311 = n47925 | n47926;
  assign n47928 = ~pi2001 & ~n46586;
  assign n47929 = pi2514 & n46979;
  assign n47930 = ~pi2001 & ~n46979;
  assign n47931 = ~n47929 & ~n47930;
  assign n47932 = n46586 & ~n47931;
  assign po2312 = n47928 | n47932;
  assign n47934 = pi3512 & n46979;
  assign n47935 = pi2002 & ~n46979;
  assign n47936 = ~n47934 & ~n47935;
  assign n47937 = n46586 & ~n47936;
  assign n47938 = pi2002 & ~n46586;
  assign po2313 = n47937 | n47938;
  assign n47940 = pi3514 & n46979;
  assign n47941 = pi2003 & ~n46979;
  assign n47942 = ~n47940 & ~n47941;
  assign n47943 = n46586 & ~n47942;
  assign n47944 = pi2003 & ~n46586;
  assign po2314 = n47943 | n47944;
  assign n47946 = pi3516 & n46979;
  assign n47947 = pi2004 & ~n46979;
  assign n47948 = ~n47946 & ~n47947;
  assign n47949 = n46586 & ~n47948;
  assign n47950 = pi2004 & ~n46586;
  assign po2315 = n47949 | n47950;
  assign n47952 = pi3517 & n46979;
  assign n47953 = pi2005 & ~n46979;
  assign n47954 = ~n47952 & ~n47953;
  assign n47955 = n46586 & ~n47954;
  assign n47956 = pi2005 & ~n46586;
  assign po2316 = n47955 | n47956;
  assign n47958 = pi3509 & n46979;
  assign n47959 = pi2006 & ~n46979;
  assign n47960 = ~n47958 & ~n47959;
  assign n47961 = n46586 & ~n47960;
  assign n47962 = pi2006 & ~n46586;
  assign po2317 = n47961 | n47962;
  assign n47964 = pi3521 & n46979;
  assign n47965 = pi2007 & ~n46979;
  assign n47966 = ~n47964 & ~n47965;
  assign n47967 = n46586 & ~n47966;
  assign n47968 = pi2007 & ~n46586;
  assign po2318 = n47967 | n47968;
  assign n47970 = pi1798 & n46581;
  assign n47971 = ~pi3330 & n47970;
  assign n47972 = pi2008 & ~n47970;
  assign n47973 = ~n47971 & ~n47972;
  assign n47974 = n46586 & ~n47973;
  assign n47975 = pi2008 & ~n46586;
  assign po2319 = n47974 | n47975;
  assign n47977 = ~pi3394 & n47970;
  assign n47978 = pi2009 & ~n47970;
  assign n47979 = ~n47977 & ~n47978;
  assign n47980 = n46586 & ~n47979;
  assign n47981 = pi2009 & ~n46586;
  assign po2320 = n47980 | n47981;
  assign n47983 = n9415 & ~n12801;
  assign n47984 = ~n9415 & ~n13121;
  assign n47985 = ~n47983 & ~n47984;
  assign n47986 = n9361 & n47985;
  assign n47987 = ~n9415 & ~n12785;
  assign n47988 = ~n47983 & ~n47987;
  assign n47989 = ~n9361 & n47988;
  assign n47990 = ~n47986 & ~n47989;
  assign n47991 = n9377 & n47990;
  assign n47992 = pi0425 & n47131;
  assign n47993 = ~n47991 & ~n47992;
  assign n47994 = po3831 & ~n47993;
  assign n47995 = pi2010 & ~po3831;
  assign po2321 = n47994 | n47995;
  assign n47997 = n9415 & ~n13735;
  assign n47998 = ~n9415 & ~n13988;
  assign n47999 = ~n47997 & ~n47998;
  assign n48000 = n9361 & n47999;
  assign n48001 = ~n9415 & ~n14046;
  assign n48002 = ~n47997 & ~n48001;
  assign n48003 = ~n9361 & n48002;
  assign n48004 = ~n48000 & ~n48003;
  assign n48005 = n9377 & n48004;
  assign n48006 = pi0409 & n47131;
  assign n48007 = ~n48005 & ~n48006;
  assign n48008 = po3831 & ~n48007;
  assign n48009 = pi2011 & ~po3831;
  assign po2322 = n48008 | n48009;
  assign n48011 = n9415 & ~n17960;
  assign n48012 = ~n9415 & ~n12415;
  assign n48013 = ~n48011 & ~n48012;
  assign n48014 = n9361 & n48013;
  assign n48015 = ~n9415 & ~n17983;
  assign n48016 = ~n48011 & ~n48015;
  assign n48017 = ~n9361 & n48016;
  assign n48018 = ~n48014 & ~n48017;
  assign n48019 = n9377 & n48018;
  assign n48020 = pi0410 & n47131;
  assign n48021 = ~n48019 & ~n48020;
  assign n48022 = po3831 & ~n48021;
  assign n48023 = pi2012 & ~po3831;
  assign po2323 = n48022 | n48023;
  assign n48025 = n9415 & ~n17899;
  assign n48026 = ~n9415 & ~n14816;
  assign n48027 = ~n48025 & ~n48026;
  assign n48028 = n9361 & n48027;
  assign n48029 = ~n9415 & ~n17927;
  assign n48030 = ~n48025 & ~n48029;
  assign n48031 = ~n9361 & n48030;
  assign n48032 = ~n48028 & ~n48031;
  assign n48033 = n9377 & n48032;
  assign n48034 = pi0411 & n47131;
  assign n48035 = ~n48033 & ~n48034;
  assign n48036 = po3831 & ~n48035;
  assign n48037 = pi2013 & ~po3831;
  assign po2324 = n48036 | n48037;
  assign n48039 = n9415 & ~n17842;
  assign n48040 = ~n9415 & ~n15115;
  assign n48041 = ~n48039 & ~n48040;
  assign n48042 = n9361 & n48041;
  assign n48043 = ~n9415 & ~n17866;
  assign n48044 = ~n48039 & ~n48043;
  assign n48045 = ~n9361 & n48044;
  assign n48046 = ~n48042 & ~n48045;
  assign n48047 = n9377 & n48046;
  assign n48048 = pi0412 & n47131;
  assign n48049 = ~n48047 & ~n48048;
  assign n48050 = po3831 & ~n48049;
  assign n48051 = pi2014 & ~po3831;
  assign po2325 = n48050 | n48051;
  assign n48053 = n9415 & ~n17784;
  assign n48054 = ~n9415 & ~n12061;
  assign n48055 = ~n48053 & ~n48054;
  assign n48056 = n9361 & n48055;
  assign n48057 = ~n9415 & ~n17809;
  assign n48058 = ~n48053 & ~n48057;
  assign n48059 = ~n9361 & n48058;
  assign n48060 = ~n48056 & ~n48059;
  assign n48061 = n9377 & n48060;
  assign n48062 = pi0413 & n47131;
  assign n48063 = ~n48061 & ~n48062;
  assign n48064 = po3831 & ~n48063;
  assign n48065 = pi2015 & ~po3831;
  assign po2326 = n48064 | n48065;
  assign n48067 = n9415 & ~n17734;
  assign n48068 = ~n9415 & ~n11181;
  assign n48069 = ~n48067 & ~n48068;
  assign n48070 = n9361 & n48069;
  assign n48071 = ~n9415 & ~n17751;
  assign n48072 = ~n48067 & ~n48071;
  assign n48073 = ~n9361 & n48072;
  assign n48074 = ~n48070 & ~n48073;
  assign n48075 = n9377 & n48074;
  assign n48076 = pi0408 & n47131;
  assign n48077 = ~n48075 & ~n48076;
  assign n48078 = po3831 & ~n48077;
  assign n48079 = pi2016 & ~po3831;
  assign po2327 = n48078 | n48079;
  assign n48081 = n38248 & n38262;
  assign n48082 = n38255 & n48081;
  assign n48083 = pi2017 & ~n38262;
  assign po2328 = n48082 | n48083;
  assign n48085 = n38242 & n42256;
  assign n48086 = n38254 & n38262;
  assign n48087 = n48085 & n48086;
  assign n48088 = pi2018 & ~n38262;
  assign po2329 = n48087 | n48088;
  assign n48090 = n38238 & n42255;
  assign n48091 = n38262 & n48090;
  assign n48092 = n38243 & n48091;
  assign n48093 = n38254 & n48092;
  assign n48094 = pi2019 & ~n38262;
  assign po2330 = n48093 | n48094;
  assign n48096 = po3627 & n47642;
  assign n48097 = ~n46264 & n48096;
  assign n48098 = ~pi2020 & n36128;
  assign po2331 = n48097 | n48098;
  assign n48100 = pi0418 & n8607;
  assign n48101 = n34039 & n48100;
  assign n48102 = n8609 & n48101;
  assign n48103 = ~n47124 & ~n48102;
  assign n48104 = n35838 & n48103;
  assign n48105 = ~n35828 & n48104;
  assign n48106 = ~n8561 & ~n48105;
  assign n48107 = ~pi2021 & n8561;
  assign n48108 = ~n48106 & ~n48107;
  assign po2332 = po3627 & ~n48108;
  assign n48110 = ~pi2022 & ~n47139;
  assign n48111 = pi0002 & n47139;
  assign po2333 = n48110 | n48111;
  assign n48113 = ~pi2023 & ~n47139;
  assign n48114 = pi0011 & n47139;
  assign po2334 = n48113 | n48114;
  assign n48116 = ~pi2024 & ~n47139;
  assign n48117 = pi0010 & n47139;
  assign po2335 = n48116 | n48117;
  assign n48119 = ~pi2025 & ~n47139;
  assign n48120 = pi0009 & n47139;
  assign po2336 = n48119 | n48120;
  assign n48122 = ~pi2026 & ~n47139;
  assign n48123 = pi0008 & n47139;
  assign po2337 = n48122 | n48123;
  assign n48125 = ~pi2027 & ~n47139;
  assign n48126 = pi0006 & n47139;
  assign po2338 = n48125 | n48126;
  assign n48128 = ~pi2028 & ~n47139;
  assign n48129 = pi0004 & n47139;
  assign po2339 = n48128 | n48129;
  assign n48131 = ~pi2029 & ~n47139;
  assign n48132 = ~n15935 & n47139;
  assign po2340 = n48131 | n48132;
  assign n48134 = ~pi2030 & ~n47139;
  assign n48135 = ~n15932 & n47139;
  assign po2341 = n48134 | n48135;
  assign n48137 = ~pi2031 & ~n47139;
  assign n48138 = pi0028 & n47139;
  assign po2342 = n48137 | n48138;
  assign n48140 = ~pi2032 & ~n47139;
  assign n48141 = pi0037 & n47139;
  assign po2343 = n48140 | n48141;
  assign n48143 = ~pi2033 & ~n47139;
  assign n48144 = pi0035 & n47139;
  assign po2344 = n48143 | n48144;
  assign n48146 = ~pi2034 & ~n47139;
  assign n48147 = pi0033 & n47139;
  assign po2345 = n48146 | n48147;
  assign n48149 = ~pi2035 & ~n47139;
  assign n48150 = pi0031 & n47139;
  assign po2346 = n48149 | n48150;
  assign n48152 = ~pi2036 & ~n47139;
  assign n48153 = pi0029 & n47139;
  assign po2347 = n48152 | n48153;
  assign n48155 = ~pi2037 & ~n47139;
  assign n48156 = pi0022 & n47139;
  assign po2348 = n48155 | n48156;
  assign n48158 = ~pi2038 & ~n47139;
  assign n48159 = pi0021 & n47139;
  assign po2349 = n48158 | n48159;
  assign n48161 = ~pi2039 & ~n47139;
  assign n48162 = pi0020 & n47139;
  assign po2350 = n48161 | n48162;
  assign n48164 = ~pi2040 & ~n47139;
  assign n48165 = pi0018 & n47139;
  assign po2351 = n48164 | n48165;
  assign n48167 = ~pi2041 & ~n47139;
  assign n48168 = pi0017 & n47139;
  assign po2352 = n48167 | n48168;
  assign n48170 = ~pi2042 & ~n47139;
  assign n48171 = pi0016 & n47139;
  assign po2353 = n48170 | n48171;
  assign n48173 = ~pi2043 & ~n47139;
  assign n48174 = pi0027 & n47139;
  assign po2354 = n48173 | n48174;
  assign n48176 = ~pi2044 & ~n47139;
  assign n48177 = pi0026 & n47139;
  assign po2355 = n48176 | n48177;
  assign n48179 = ~pi2045 & ~n47139;
  assign n48180 = pi0025 & n47139;
  assign po2356 = n48179 | n48180;
  assign n48182 = ~pi2046 & ~n47139;
  assign n48183 = ~n15953 & n47139;
  assign po2357 = n48182 | n48183;
  assign n48185 = ~pi2047 & ~n47139;
  assign n48186 = ~n15951 & n47139;
  assign po2358 = n48185 | n48186;
  assign n48188 = n10770 & ~n36181;
  assign n48189 = ~pi2048 & n48188;
  assign n48190 = pi2048 & ~n48188;
  assign po2359 = n48189 | n48190;
  assign n48192 = ~pi1860 & n8201;
  assign n48193 = ~pi2049 & ~n48192;
  assign n48194 = pi3281 & pi3343;
  assign n48195 = pi3199 & n48194;
  assign n48196 = pi2759 & n48195;
  assign n48197 = pi2049 & n48196;
  assign n48198 = ~pi2049 & ~n48196;
  assign n48199 = ~n48197 & ~n48198;
  assign n48200 = n48192 & ~n48199;
  assign n48201 = ~n48193 & ~n48200;
  assign po2360 = ~n36174 & n48201;
  assign n48203 = ~pi2050 & ~n47139;
  assign n48204 = pi0014 & n47139;
  assign po2361 = n48203 | n48204;
  assign n48206 = ~n14403 & n47446;
  assign n48207 = pi2051 & ~n47446;
  assign po2362 = n48206 | n48207;
  assign n48209 = ~n12061 & n47446;
  assign n48210 = pi2052 & ~n47446;
  assign po2363 = n48209 | n48210;
  assign n48212 = ~n10608 & n47446;
  assign n48213 = pi2053 & ~n47446;
  assign po2364 = n48212 | n48213;
  assign n48215 = ~n13988 & n47446;
  assign n48216 = pi2054 & ~n47446;
  assign po2365 = n48215 | n48216;
  assign n48218 = ~n13121 & n47446;
  assign n48219 = pi2055 & ~n47446;
  assign po2366 = n48218 | n48219;
  assign n48221 = pi1919 & n47566;
  assign n48222 = ~pi1936 & ~pi2056;
  assign n48223 = ~n39525 & ~n48222;
  assign n48224 = n47568 & ~n48223;
  assign n48225 = ~pi2056 & ~n47568;
  assign n48226 = ~n48224 & ~n48225;
  assign n48227 = ~n47566 & ~n48226;
  assign po2367 = n48221 | n48227;
  assign n48229 = ~n12726 & n47446;
  assign n48230 = pi2057 & ~n47446;
  assign po2368 = n48229 | n48230;
  assign n48232 = ~n15115 & n38320;
  assign n48233 = ~pi2058 & n38305;
  assign n48234 = ~n38306 & ~n48233;
  assign n48235 = ~n36181 & ~n48234;
  assign n48236 = ~pi2058 & n36181;
  assign n48237 = ~n48235 & ~n48236;
  assign n48238 = ~n38320 & n48237;
  assign po2369 = n48232 | n48238;
  assign n48240 = ~n11181 & n38320;
  assign n48241 = ~pi2059 & n8598;
  assign n48242 = ~n38302 & ~n48241;
  assign n48243 = ~n36181 & ~n48242;
  assign n48244 = ~pi2059 & n36181;
  assign n48245 = ~n48243 & ~n48244;
  assign n48246 = ~n38320 & n48245;
  assign po2370 = n48240 | n48246;
  assign n48248 = ~pi2060 & ~n47139;
  assign n48249 = pi0024 & n47139;
  assign po2371 = n48248 | n48249;
  assign n48251 = ~n12061 & n38320;
  assign n48252 = ~n38301 & ~n38303;
  assign n48253 = ~n38302 & ~n48252;
  assign n48254 = n38302 & n48252;
  assign n48255 = ~n48253 & ~n48254;
  assign n48256 = ~n36181 & ~n48255;
  assign n48257 = ~pi2061 & n36181;
  assign n48258 = ~n48256 & ~n48257;
  assign n48259 = ~n38320 & n48258;
  assign po2372 = n48251 | n48259;
  assign n48261 = ~pi2062 & ~n47139;
  assign n48262 = pi0015 & n47139;
  assign po2373 = n48261 | n48262;
  assign n48264 = ~pi2063 & ~n47139;
  assign n48265 = pi0030 & n47139;
  assign po2374 = n48264 | n48265;
  assign n48267 = ~pi2064 & ~n47139;
  assign n48268 = pi0019 & n47139;
  assign po2375 = n48267 | n48268;
  assign n48270 = ~pi2065 & ~n47139;
  assign n48271 = pi0023 & n47139;
  assign po2376 = n48270 | n48271;
  assign n48273 = ~pi2066 & ~n47139;
  assign n48274 = pi0032 & n47139;
  assign po2377 = n48273 | n48274;
  assign n48276 = ~pi0985 & n35623;
  assign n48277 = ~pi3426 & n48276;
  assign n48278 = ~n13701 & n48277;
  assign n48279 = pi2067 & ~n48277;
  assign po2378 = n48278 | n48279;
  assign n48281 = ~pi0986 & n35625;
  assign n48282 = ~pi3426 & n48281;
  assign n48283 = ~n12061 & n48282;
  assign n48284 = pi2068 & ~n48282;
  assign po2379 = n48283 | n48284;
  assign n48286 = pi3516 & n47970;
  assign n48287 = pi2069 & ~n47970;
  assign n48288 = ~n48286 & ~n48287;
  assign n48289 = n46586 & ~n48288;
  assign n48290 = pi2069 & ~n46586;
  assign po2380 = n48289 | n48290;
  assign n48292 = pi3519 & n47897;
  assign n48293 = pi2070 & ~n47897;
  assign n48294 = ~n48292 & ~n48293;
  assign n48295 = n46586 & ~n48294;
  assign n48296 = pi2070 & ~n46586;
  assign po2381 = n48295 | n48296;
  assign n48298 = pi3392 & n47897;
  assign n48299 = pi2071 & ~n47897;
  assign n48300 = ~n48298 & ~n48299;
  assign n48301 = n46586 & ~n48300;
  assign n48302 = pi2071 & ~n46586;
  assign po2382 = n48301 | n48302;
  assign n48304 = pi3504 & n47970;
  assign n48305 = pi2072 & ~n47970;
  assign n48306 = ~n48304 & ~n48305;
  assign n48307 = n46586 & ~n48306;
  assign n48308 = pi2072 & ~n46586;
  assign po2383 = n48307 | n48308;
  assign n48310 = pi3511 & n47897;
  assign n48311 = pi2073 & ~n47897;
  assign n48312 = ~n48310 & ~n48311;
  assign n48313 = n46586 & ~n48312;
  assign n48314 = pi2073 & ~n46586;
  assign po2384 = n48313 | n48314;
  assign n48316 = pi3504 & n46972;
  assign n48317 = pi2074 & ~n46972;
  assign n48318 = ~n48316 & ~n48317;
  assign n48319 = n46586 & ~n48318;
  assign n48320 = pi2074 & ~n46586;
  assign po2385 = n48319 | n48320;
  assign n48322 = pi3511 & n46972;
  assign n48323 = pi2075 & ~n46972;
  assign n48324 = ~n48322 & ~n48323;
  assign n48325 = n46586 & ~n48324;
  assign n48326 = pi2075 & ~n46586;
  assign po2386 = n48325 | n48326;
  assign n48328 = pi2076 & ~n47970;
  assign n48329 = pi3519 & n47970;
  assign n48330 = ~n48328 & ~n48329;
  assign n48331 = n46586 & ~n48330;
  assign n48332 = pi2076 & ~n46586;
  assign po2387 = n48331 | n48332;
  assign n48334 = pi3519 & n46972;
  assign n48335 = pi2077 & ~n46972;
  assign n48336 = ~n48334 & ~n48335;
  assign n48337 = n46586 & ~n48336;
  assign n48338 = pi2077 & ~n46586;
  assign po2388 = n48337 | n48338;
  assign n48340 = pi3688 & n47620;
  assign n48341 = pi2078 & ~n47620;
  assign po2389 = n48340 | n48341;
  assign n48343 = ~pi2079 & ~n46920;
  assign n48344 = pi0406 & pi0413;
  assign n48345 = ~n46942 & ~n48344;
  assign n48346 = pi0413 & ~pi0425;
  assign n48347 = n48345 & ~n48346;
  assign n48348 = pi0408 & ~n48347;
  assign n48349 = pi0408 & n46937;
  assign n48350 = ~n48348 & ~n48349;
  assign n48351 = pi0408 & n46934;
  assign n48352 = ~pi0406 & ~pi0411;
  assign n48353 = pi0425 & n48352;
  assign n48354 = n48351 & n48353;
  assign n48355 = n48350 & ~n48354;
  assign n48356 = n46920 & ~n48355;
  assign po2390 = n48343 | n48356;
  assign n48358 = ~pi2080 & ~n46920;
  assign n48359 = ~pi0406 & pi0413;
  assign n48360 = pi0413 & pi0425;
  assign n48361 = ~n48359 & ~n48360;
  assign n48362 = ~n46923 & n48361;
  assign n48363 = pi0408 & ~n48362;
  assign n48364 = ~n48349 & ~n48363;
  assign n48365 = pi0406 & ~pi0425;
  assign n48366 = pi0411 & n48365;
  assign n48367 = n48351 & n48366;
  assign n48368 = n48364 & ~n48367;
  assign n48369 = n46920 & ~n48368;
  assign po2391 = n48358 | n48369;
  assign n48371 = ~pi2081 & ~n46920;
  assign n48372 = pi0408 & n46929;
  assign n48373 = ~n48363 & ~n48372;
  assign n48374 = pi0408 & ~pi0413;
  assign n48375 = pi0412 & n48374;
  assign n48376 = n48366 & n48375;
  assign n48377 = n48373 & ~n48376;
  assign n48378 = n46920 & ~n48377;
  assign po2392 = n48371 | n48378;
  assign n48380 = ~n8199 & ~n8209;
  assign n48381 = ~n8232 & n48380;
  assign n48382 = ~n8196 & n48381;
  assign n48383 = ~n8211 & n48382;
  assign n48384 = ~pi2082 & n48383;
  assign n48385 = pi2798 & pi2825;
  assign n48386 = pi2799 & n48385;
  assign n48387 = pi2600 & n48386;
  assign n48388 = pi2082 & n48387;
  assign n48389 = ~pi2082 & ~n48387;
  assign n48390 = ~n48388 & ~n48389;
  assign n48391 = ~n48383 & ~n48390;
  assign n48392 = ~n48384 & ~n48391;
  assign n48393 = ~po3646 & po3616;
  assign n48394 = ~po3645 & po3647;
  assign n48395 = n48393 & n48394;
  assign n48396 = ~n8199 & n48393;
  assign n48397 = ~po3647 & n48396;
  assign n48398 = po3645 & n48397;
  assign n48399 = ~po3646 & ~po3616;
  assign n48400 = po3645 & ~po3647;
  assign n48401 = n48399 & n48400;
  assign n48402 = ~n8209 & n48401;
  assign n48403 = po3645 & po3647;
  assign n48404 = n48399 & n48403;
  assign n48405 = ~n8211 & n48404;
  assign n48406 = ~n48402 & ~n48405;
  assign n48407 = ~n36174 & n48406;
  assign n48408 = ~n48398 & n48407;
  assign n48409 = ~n48395 & n48408;
  assign po2393 = n48392 & n48409;
  assign n48411 = ~pi2083 & ~n46920;
  assign n48412 = ~n48344 & ~n48360;
  assign n48413 = ~n46942 & n48412;
  assign n48414 = pi0408 & ~n48413;
  assign n48415 = ~n48372 & ~n48414;
  assign n48416 = ~pi0425 & n48352;
  assign n48417 = pi0412 & n48416;
  assign n48418 = n48374 & n48417;
  assign n48419 = n48415 & ~n48418;
  assign n48420 = n46920 & ~n48419;
  assign po2394 = n48411 | n48420;
  assign n48422 = ~pi0760 & n35635;
  assign n48423 = ~pi3426 & n48422;
  assign n48424 = ~n13988 & n48423;
  assign n48425 = pi2084 & ~n48423;
  assign po2395 = n48424 | n48425;
  assign n48427 = ~pi0598 & n9365;
  assign n48428 = pi0979 & n48427;
  assign n48429 = ~n47688 & n48428;
  assign n48430 = pi2085 & ~n48428;
  assign po2396 = n48429 | n48430;
  assign n48432 = ~pi2086 & ~n46920;
  assign n48433 = ~n46942 & ~n48360;
  assign n48434 = ~n48359 & n48433;
  assign n48435 = pi0408 & ~n48434;
  assign n48436 = ~n48349 & ~n48435;
  assign n48437 = ~pi0411 & ~pi0425;
  assign n48438 = pi0406 & n48437;
  assign n48439 = n48351 & n48438;
  assign n48440 = n48436 & ~n48439;
  assign n48441 = n46920 & ~n48440;
  assign po2397 = n48432 | n48441;
  assign n48443 = ~n12415 & n48423;
  assign n48444 = pi2087 & ~n48423;
  assign po2398 = n48443 | n48444;
  assign n48446 = ~n15426 & n48277;
  assign n48447 = pi2088 & ~n48277;
  assign po2399 = n48446 | n48447;
  assign n48449 = ~n13701 & n48423;
  assign n48450 = pi2089 & ~n48423;
  assign po2400 = n48449 | n48450;
  assign n48452 = ~pi2090 & ~n47395;
  assign n48453 = ~n12726 & n47395;
  assign po2401 = n48452 | n48453;
  assign n48455 = ~pi2091 & ~n47395;
  assign n48456 = ~n13701 & n47395;
  assign po2402 = n48455 | n48456;
  assign n48458 = ~pi2092 & ~n47395;
  assign n48459 = ~n13398 & n47395;
  assign po2403 = n48458 | n48459;
  assign n48461 = ~pi2093 & ~n47395;
  assign n48462 = ~n12415 & n47395;
  assign po2404 = n48461 | n48462;
  assign n48464 = ~pi2094 & ~n47395;
  assign n48465 = ~n15115 & n47395;
  assign po2405 = n48464 | n48465;
  assign n48467 = ~pi2095 & ~n47395;
  assign n48468 = ~n17368 & n47395;
  assign po2406 = n48467 | n48468;
  assign n48470 = ~pi2096 & ~n47395;
  assign n48471 = ~n10608 & n47395;
  assign po2407 = n48470 | n48471;
  assign n48473 = ~pi2097 & ~n47395;
  assign n48474 = ~n9825 & n47395;
  assign po2408 = n48473 | n48474;
  assign n48476 = ~pi2098 & ~n47395;
  assign n48477 = ~n11181 & n47395;
  assign po2409 = n48476 | n48477;
  assign po2410 = po0493 & ~n31779;
  assign po2411 = ~pi2099 | pi3136;
  assign po2412 = ~n9825 & n44885;
  assign n48482 = pi1749 & ~pi1761;
  assign n48483 = pi3243 & ~pi3317;
  assign n48484 = ~pi3243 & pi3317;
  assign n48485 = ~n48483 & ~n48484;
  assign n48486 = n48482 & ~n48485;
  assign n48487 = ~pi2101 & ~n48486;
  assign n48488 = n38900 & n39500;
  assign n48489 = ~n48487 & ~n48488;
  assign n48490 = ~n9825 & n48488;
  assign po2413 = n48489 | n48490;
  assign n48492 = pi1750 & ~pi1762;
  assign n48493 = pi3219 & ~pi3318;
  assign n48494 = ~pi3219 & pi3318;
  assign n48495 = ~n48493 & ~n48494;
  assign n48496 = n48492 & ~n48495;
  assign n48497 = ~pi2102 & ~n48496;
  assign n48498 = ~n48488 & ~n48497;
  assign n48499 = ~n10608 & n48488;
  assign po2414 = n48498 | n48499;
  assign n48501 = pi1751 & ~pi1857;
  assign n48502 = pi3241 & ~pi3351;
  assign n48503 = ~pi3241 & pi3351;
  assign n48504 = ~n48502 & ~n48503;
  assign n48505 = n48501 & ~n48504;
  assign n48506 = ~pi2103 & ~n48505;
  assign n48507 = ~n48488 & ~n48506;
  assign n48508 = ~n13121 & n48488;
  assign po2415 = n48507 | n48508;
  assign n48510 = pi1752 & ~pi1763;
  assign n48511 = pi3220 & ~pi3349;
  assign n48512 = ~pi3220 & pi3349;
  assign n48513 = ~n48511 & ~n48512;
  assign n48514 = n48510 & ~n48513;
  assign n48515 = ~pi2104 & ~n48514;
  assign n48516 = ~n48488 & ~n48515;
  assign n48517 = ~n13398 & n48488;
  assign po2416 = n48516 | n48517;
  assign n48519 = pi1753 & ~pi1764;
  assign n48520 = pi3242 & ~pi3346;
  assign n48521 = ~pi3242 & pi3346;
  assign n48522 = ~n48520 & ~n48521;
  assign n48523 = n48519 & ~n48522;
  assign n48524 = ~pi2105 & ~n48523;
  assign n48525 = ~n48488 & ~n48524;
  assign n48526 = ~n13988 & n48488;
  assign po2417 = n48525 | n48526;
  assign n48528 = pi1754 & ~pi1765;
  assign n48529 = pi3221 & ~pi3345;
  assign n48530 = ~pi3221 & pi3345;
  assign n48531 = ~n48529 & ~n48530;
  assign n48532 = n48528 & ~n48531;
  assign n48533 = ~pi2106 & ~n48532;
  assign n48534 = ~n48488 & ~n48533;
  assign n48535 = ~n12415 & n48488;
  assign po2418 = n48534 | n48535;
  assign n48537 = pi1755 & ~pi1858;
  assign n48538 = pi3218 & ~pi3348;
  assign n48539 = ~pi3218 & pi3348;
  assign n48540 = ~n48538 & ~n48539;
  assign n48541 = n48537 & ~n48540;
  assign n48542 = ~pi2107 & ~n48541;
  assign n48543 = ~n48488 & ~n48542;
  assign n48544 = ~n14816 & n48488;
  assign po2419 = n48543 | n48544;
  assign n48546 = pi1757 & ~pi1767;
  assign n48547 = pi3223 & ~pi3320;
  assign n48548 = ~pi3223 & pi3320;
  assign n48549 = ~n48547 & ~n48548;
  assign n48550 = n48546 & ~n48549;
  assign n48551 = ~pi2108 & ~n48550;
  assign n48552 = ~n48488 & ~n48551;
  assign n48553 = ~n12061 & n48488;
  assign po2420 = n48552 | n48553;
  assign n48555 = pi1758 & ~pi1768;
  assign n48556 = pi3224 & ~pi3357;
  assign n48557 = ~pi3224 & pi3357;
  assign n48558 = ~n48556 & ~n48557;
  assign n48559 = n48555 & ~n48558;
  assign n48560 = ~pi2109 & ~n48559;
  assign n48561 = ~n48488 & ~n48560;
  assign n48562 = ~n17368 & n48488;
  assign po2421 = n48561 | n48562;
  assign n48564 = pi1760 & ~pi1769;
  assign n48565 = pi3225 & ~pi3321;
  assign n48566 = ~pi3225 & pi3321;
  assign n48567 = ~n48565 & ~n48566;
  assign n48568 = n48564 & ~n48567;
  assign n48569 = ~pi2110 & ~n48568;
  assign n48570 = ~n48488 & ~n48569;
  assign n48571 = ~n11181 & n48488;
  assign po2422 = n48570 | n48571;
  assign n48573 = pi2111 & ~n47510;
  assign n48574 = ~n10608 & n47510;
  assign po2423 = n48573 | n48574;
  assign n48576 = pi2112 & n47561;
  assign po2424 = n47562 | n48576;
  assign n48578 = pi2113 & n48383;
  assign n48579 = pi2799 & pi2825;
  assign n48580 = pi2082 & n48579;
  assign n48581 = pi2600 & n48580;
  assign n48582 = pi2798 & n48581;
  assign n48583 = pi2113 & ~n48582;
  assign n48584 = ~pi2113 & pi2798;
  assign n48585 = n48581 & n48584;
  assign n48586 = ~n48583 & ~n48585;
  assign n48587 = ~n48383 & ~n48586;
  assign n48588 = ~n48578 & ~n48587;
  assign po2425 = n48409 & ~n48588;
  assign n48590 = ~n44983 & n44987;
  assign n48591 = pi2114 & n44983;
  assign n48592 = ~n48590 & n48591;
  assign n48593 = pi2114 & ~n8213;
  assign n48594 = ~n48590 & n48593;
  assign n48595 = ~n8313 & n48594;
  assign n48596 = pi0565 & pi2409;
  assign n48597 = n44991 & n48596;
  assign n48598 = pi3256 & n48597;
  assign n48599 = n48590 & n48598;
  assign n48600 = pi3216 & n48597;
  assign n48601 = n48590 & n48600;
  assign n48602 = ~n48599 & ~n48601;
  assign n48603 = ~n48595 & n48602;
  assign po2426 = n48592 | ~n48603;
  assign n48605 = pi3690 & n47620;
  assign n48606 = pi2115 & ~n47620;
  assign po2427 = n48605 | n48606;
  assign n48608 = pi3689 & n47620;
  assign n48609 = pi2116 & ~n47620;
  assign po2428 = n48608 | n48609;
  assign n48611 = pi3687 & n47620;
  assign n48612 = pi2117 & ~n47620;
  assign po2429 = n48611 | n48612;
  assign n48614 = pi3686 & n47620;
  assign n48615 = pi2118 & ~n47620;
  assign po2430 = n48614 | n48615;
  assign n48617 = pi3685 & n47620;
  assign n48618 = pi2119 & ~n47620;
  assign po2431 = n48617 | n48618;
  assign n48620 = pi3684 & n47620;
  assign n48621 = pi2120 & ~n47620;
  assign po2432 = n48620 | n48621;
  assign n48623 = pi3683 & n47620;
  assign n48624 = pi2121 & ~n47620;
  assign po2433 = n48623 | n48624;
  assign n48626 = ~n10608 & n48277;
  assign n48627 = pi2122 & ~n48277;
  assign po2434 = n48626 | n48627;
  assign n48629 = pi1759 & ~pi1854;
  assign n48630 = pi3240 & ~pi3340;
  assign n48631 = ~pi3240 & pi3340;
  assign n48632 = ~n48630 & ~n48631;
  assign n48633 = n48629 & ~n48632;
  assign n48634 = ~pi2123 & ~n48633;
  assign n48635 = ~n48488 & ~n48634;
  assign n48636 = ~n17199 & n48488;
  assign po2435 = n48635 | n48636;
  assign n48638 = ~pi0711 & n9365;
  assign n48639 = pi0979 & n48638;
  assign n48640 = ~n30267 & n48639;
  assign n48641 = pi2124 & ~n48639;
  assign po2436 = n48640 | n48641;
  assign n48643 = ~n30288 & n48639;
  assign n48644 = pi2125 & ~n48639;
  assign po2437 = n48643 | n48644;
  assign n48646 = ~n24744 & n48639;
  assign n48647 = pi2126 & ~n48639;
  assign po2438 = n48646 | n48647;
  assign n48649 = ~n24769 & n48639;
  assign n48650 = pi2127 & ~n48639;
  assign po2439 = n48649 | n48650;
  assign n48652 = ~n25699 & n48639;
  assign n48653 = pi2128 & ~n48639;
  assign po2440 = n48652 | n48653;
  assign n48655 = ~n25718 & n48639;
  assign n48656 = pi2129 & ~n48639;
  assign po2441 = n48655 | n48656;
  assign n48658 = ~n24256 & n48639;
  assign n48659 = pi2130 & ~n48639;
  assign po2442 = n48658 | n48659;
  assign n48661 = ~n24289 & n48639;
  assign n48662 = pi2131 & ~n48639;
  assign po2443 = n48661 | n48662;
  assign n48664 = ~n24446 & n48639;
  assign n48665 = pi2132 & ~n48639;
  assign po2444 = n48664 | n48665;
  assign n48667 = ~n24265 & n48639;
  assign n48668 = pi2133 & ~n48639;
  assign po2445 = n48667 | n48668;
  assign n48670 = ~n30309 & n48639;
  assign n48671 = pi2134 & ~n48639;
  assign po2446 = n48670 | n48671;
  assign n48673 = ~n30321 & n48639;
  assign n48674 = pi2135 & ~n48639;
  assign po2447 = n48673 | n48674;
  assign n48676 = ~n30333 & n48639;
  assign n48677 = pi2136 & ~n48639;
  assign po2448 = n48676 | n48677;
  assign n48679 = ~n27570 & n48639;
  assign n48680 = pi2137 & ~n48639;
  assign po2449 = n48679 | n48680;
  assign n48682 = ~n25999 & n48639;
  assign n48683 = pi2138 & ~n48639;
  assign po2450 = n48682 | n48683;
  assign n48685 = ~n24488 & n48639;
  assign n48686 = pi2139 & ~n48639;
  assign po2451 = n48685 | n48686;
  assign n48688 = ~n44811 & ~n48105;
  assign n48689 = n36059 & n48688;
  assign n48690 = ~pi2140 & n36128;
  assign po2452 = n48689 | n48690;
  assign n48692 = pi1756 & ~pi1766;
  assign n48693 = pi3222 & ~pi3319;
  assign n48694 = ~pi3222 & pi3319;
  assign n48695 = ~n48693 & ~n48694;
  assign n48696 = n48692 & ~n48695;
  assign n48697 = ~pi2141 & ~n48696;
  assign n48698 = ~n48488 & ~n48697;
  assign n48699 = ~n15115 & n48488;
  assign po2453 = n48698 | n48699;
  assign n48701 = ~pi2142 & n8561;
  assign n48702 = ~n47642 & ~n48701;
  assign po2454 = po3627 & ~n48702;
  assign n48704 = pi2143 & po3853;
  assign po2455 = po0493 & ~n48704;
  assign n48706 = ~n19543 & ~n24340;
  assign po2456 = n19551 | ~n48706;
  assign n48708 = ~n47652 & n48428;
  assign n48709 = pi2144 & ~n48428;
  assign po2457 = n48708 | n48709;
  assign n48711 = ~n47661 & n48428;
  assign n48712 = pi2145 & ~n48428;
  assign po2458 = n48711 | n48712;
  assign n48714 = ~n47670 & n48428;
  assign n48715 = pi2146 & ~n48428;
  assign po2459 = n48714 | n48715;
  assign n48717 = ~n47679 & n48428;
  assign n48718 = pi2147 & ~n48428;
  assign po2460 = n48717 | n48718;
  assign n48720 = ~n47697 & n48428;
  assign n48721 = pi2148 & ~n48428;
  assign po2461 = n48720 | n48721;
  assign n48723 = ~n47706 & n48428;
  assign n48724 = pi2149 & ~n48428;
  assign po2462 = n48723 | n48724;
  assign n48726 = ~n47715 & n48428;
  assign n48727 = pi2150 & ~n48428;
  assign po2463 = n48726 | n48727;
  assign n48729 = ~n46897 & n48428;
  assign n48730 = pi2151 & ~n48428;
  assign po2464 = n48729 | n48730;
  assign n48732 = ~n47724 & n48428;
  assign n48733 = pi2152 & ~n48428;
  assign po2465 = n48732 | n48733;
  assign n48735 = ~n46906 & n48428;
  assign n48736 = pi2153 & ~n48428;
  assign po2466 = n48735 | n48736;
  assign n48738 = ~n47733 & n48428;
  assign n48739 = pi2154 & ~n48428;
  assign po2467 = n48738 | n48739;
  assign n48741 = ~n47742 & n48428;
  assign n48742 = pi2155 & ~n48428;
  assign po2468 = n48741 | n48742;
  assign n48744 = ~n47751 & n48428;
  assign n48745 = pi2156 & ~n48428;
  assign po2469 = n48744 | n48745;
  assign n48747 = ~n47760 & n48428;
  assign n48748 = pi2157 & ~n48428;
  assign po2470 = n48747 | n48748;
  assign n48750 = ~n30540 & n48428;
  assign n48751 = pi2158 & ~n48428;
  assign po2471 = n48750 | n48751;
  assign n48753 = n30709 & ~n46900;
  assign n48754 = pi2159 & ~n30709;
  assign po2472 = n48753 | n48754;
  assign n48756 = n30709 & n46909;
  assign n48757 = pi2160 & ~n30709;
  assign po2473 = n48756 | n48757;
  assign n48759 = ~pi0649 & n9365;
  assign n48760 = pi0979 & n48759;
  assign n48761 = ~n30267 & n48760;
  assign n48762 = pi2161 & ~n48760;
  assign po2474 = n48761 | n48762;
  assign n48764 = ~n30288 & n48760;
  assign n48765 = pi2162 & ~n48760;
  assign po2475 = n48764 | n48765;
  assign n48767 = ~n24744 & n48760;
  assign n48768 = pi2163 & ~n48760;
  assign po2476 = n48767 | n48768;
  assign n48770 = ~n24769 & n48760;
  assign n48771 = pi2164 & ~n48760;
  assign po2477 = n48770 | n48771;
  assign n48773 = ~n25699 & n48760;
  assign n48774 = pi2165 & ~n48760;
  assign po2478 = n48773 | n48774;
  assign n48776 = ~n25718 & n48760;
  assign n48777 = pi2166 & ~n48760;
  assign po2479 = n48776 | n48777;
  assign n48779 = ~n24256 & n48760;
  assign n48780 = pi2167 & ~n48760;
  assign po2480 = n48779 | n48780;
  assign n48782 = ~n24289 & n48760;
  assign n48783 = pi2168 & ~n48760;
  assign po2481 = n48782 | n48783;
  assign n48785 = ~n24446 & n48760;
  assign n48786 = pi2169 & ~n48760;
  assign po2482 = n48785 | n48786;
  assign n48788 = ~n24265 & n48760;
  assign n48789 = pi2170 & ~n48760;
  assign po2483 = n48788 | n48789;
  assign n48791 = ~n30309 & n48760;
  assign n48792 = pi2171 & ~n48760;
  assign po2484 = n48791 | n48792;
  assign n48794 = ~n30321 & n48760;
  assign n48795 = pi2172 & ~n48760;
  assign po2485 = n48794 | n48795;
  assign n48797 = ~n30333 & n48760;
  assign n48798 = pi2173 & ~n48760;
  assign po2486 = n48797 | n48798;
  assign n48800 = ~n27570 & n48760;
  assign n48801 = pi2174 & ~n48760;
  assign po2487 = n48800 | n48801;
  assign n48803 = ~n25999 & n48760;
  assign n48804 = pi2175 & ~n48760;
  assign po2488 = n48803 | n48804;
  assign n48806 = ~n24488 & n48760;
  assign n48807 = pi2176 & ~n48760;
  assign po2489 = n48806 | n48807;
  assign n48809 = ~pi0575 & n9365;
  assign n48810 = pi0979 & n48809;
  assign n48811 = ~n30267 & n48810;
  assign n48812 = pi2177 & ~n48810;
  assign po2490 = n48811 | n48812;
  assign n48814 = ~n30288 & n48810;
  assign n48815 = pi2178 & ~n48810;
  assign po2491 = n48814 | n48815;
  assign n48817 = ~n24744 & n48810;
  assign n48818 = pi2179 & ~n48810;
  assign po2492 = n48817 | n48818;
  assign n48820 = ~n24769 & n48810;
  assign n48821 = pi2180 & ~n48810;
  assign po2493 = n48820 | n48821;
  assign n48823 = ~n25699 & n48810;
  assign n48824 = pi2181 & ~n48810;
  assign po2494 = n48823 | n48824;
  assign n48826 = ~n25718 & n48810;
  assign n48827 = pi2182 & ~n48810;
  assign po2495 = n48826 | n48827;
  assign n48829 = ~n24256 & n48810;
  assign n48830 = pi2183 & ~n48810;
  assign po2496 = n48829 | n48830;
  assign n48832 = ~n24289 & n48810;
  assign n48833 = pi2184 & ~n48810;
  assign po2497 = n48832 | n48833;
  assign n48835 = ~n24446 & n48810;
  assign n48836 = pi2185 & ~n48810;
  assign po2498 = n48835 | n48836;
  assign n48838 = ~n24265 & n48810;
  assign n48839 = pi2186 & ~n48810;
  assign po2499 = n48838 | n48839;
  assign n48841 = ~n30309 & n48810;
  assign n48842 = pi2187 & ~n48810;
  assign po2500 = n48841 | n48842;
  assign n48844 = ~n30321 & n48810;
  assign n48845 = pi2188 & ~n48810;
  assign po2501 = n48844 | n48845;
  assign n48847 = ~n30333 & n48810;
  assign n48848 = pi2189 & ~n48810;
  assign po2502 = n48847 | n48848;
  assign n48850 = ~n27570 & n48810;
  assign n48851 = pi2190 & ~n48810;
  assign po2503 = n48850 | n48851;
  assign n48853 = ~n25999 & n48810;
  assign n48854 = pi2191 & ~n48810;
  assign po2504 = n48853 | n48854;
  assign n48856 = ~n24488 & n48810;
  assign n48857 = pi2192 & ~n48810;
  assign po2505 = n48856 | n48857;
  assign n48859 = po3627 & n33813;
  assign n48860 = pi2193 & n48859;
  assign n48861 = ~n15937 & ~n15992;
  assign n48862 = ~n33813 & ~n48861;
  assign n48863 = po3627 & n48862;
  assign po2506 = n48860 | n48863;
  assign n48865 = ~pi2194 & ~n46920;
  assign n48866 = ~n48372 & ~n48435;
  assign n48867 = n48375 & n48438;
  assign n48868 = n48866 & ~n48867;
  assign n48869 = n46920 & ~n48868;
  assign po2507 = n48865 | n48869;
  assign n48871 = ~pi2195 & ~n46920;
  assign n48872 = ~n46923 & ~n48344;
  assign n48873 = ~n48346 & n48872;
  assign n48874 = pi0408 & ~n48873;
  assign n48875 = ~n48372 & ~n48874;
  assign n48876 = ~pi0406 & pi0425;
  assign n48877 = pi0411 & n48876;
  assign n48878 = n48375 & n48877;
  assign n48879 = n48875 & ~n48878;
  assign n48880 = n46920 & ~n48879;
  assign po2508 = n48871 | n48880;
  assign n48882 = ~pi2196 & ~n46920;
  assign n48883 = ~n48349 & ~n48874;
  assign n48884 = n48351 & n48877;
  assign n48885 = n48883 & ~n48884;
  assign n48886 = n46920 & ~n48885;
  assign po2509 = n48882 | n48886;
  assign n48888 = ~pi2197 & ~n46920;
  assign n48889 = ~n48348 & ~n48372;
  assign n48890 = n48353 & n48375;
  assign n48891 = n48889 & ~n48890;
  assign n48892 = n46920 & ~n48891;
  assign po2510 = n48888 | n48892;
  assign n48894 = ~pi2198 & ~n46920;
  assign n48895 = ~n46923 & n48412;
  assign n48896 = pi0408 & ~n48895;
  assign n48897 = ~n48349 & ~n48896;
  assign n48898 = ~pi0406 & ~pi0425;
  assign n48899 = pi0411 & n48898;
  assign n48900 = n48351 & n48899;
  assign n48901 = n48897 & ~n48900;
  assign n48902 = n46920 & ~n48901;
  assign po2511 = n48894 | n48902;
  assign n48904 = ~pi2199 & ~n46920;
  assign n48905 = ~n48372 & ~n48896;
  assign n48906 = n48375 & n48899;
  assign n48907 = n48905 & ~n48906;
  assign n48908 = n46920 & ~n48907;
  assign po2512 = n48904 | n48908;
  assign n48910 = ~pi2200 & ~n46920;
  assign n48911 = ~n48349 & ~n48414;
  assign n48912 = pi0408 & n48416;
  assign n48913 = n46934 & n48912;
  assign n48914 = n48911 & ~n48913;
  assign n48915 = n46920 & ~n48914;
  assign po2513 = n48910 | n48915;
  assign n48917 = ~pi1050 & n35504;
  assign n48918 = ~pi3426 & n48917;
  assign n48919 = ~n12726 & n48918;
  assign n48920 = pi2201 & ~n48918;
  assign po2514 = n48919 | n48920;
  assign n48922 = ~n13701 & n48918;
  assign n48923 = pi2202 & ~n48918;
  assign po2515 = n48922 | n48923;
  assign n48925 = ~n13121 & n48918;
  assign n48926 = pi2203 & ~n48918;
  assign po2516 = n48925 | n48926;
  assign n48928 = ~n13398 & n48918;
  assign n48929 = pi2204 & ~n48918;
  assign po2517 = n48928 | n48929;
  assign n48931 = ~n13988 & n48918;
  assign n48932 = pi2205 & ~n48918;
  assign po2518 = n48931 | n48932;
  assign n48934 = ~n12415 & n48918;
  assign n48935 = pi2206 & ~n48918;
  assign po2519 = n48934 | n48935;
  assign n48937 = ~n14816 & n48918;
  assign n48938 = pi2207 & ~n48918;
  assign po2520 = n48937 | n48938;
  assign n48940 = ~n15115 & n48918;
  assign n48941 = pi2208 & ~n48918;
  assign po2521 = n48940 | n48941;
  assign n48943 = ~n12061 & n48918;
  assign n48944 = pi2209 & ~n48918;
  assign po2522 = n48943 | n48944;
  assign n48946 = ~n9825 & n48918;
  assign n48947 = pi2210 & ~n48918;
  assign po2523 = n48946 | n48947;
  assign n48949 = ~n10608 & n48918;
  assign n48950 = pi2211 & ~n48918;
  assign po2524 = n48949 | n48950;
  assign n48952 = ~n15426 & n48918;
  assign n48953 = pi2212 & ~n48918;
  assign po2525 = n48952 | n48953;
  assign n48955 = ~n14403 & n48918;
  assign n48956 = pi2213 & ~n48918;
  assign po2526 = n48955 | n48956;
  assign n48958 = ~n11181 & n48918;
  assign n48959 = pi2214 & ~n48918;
  assign po2527 = n48958 | n48959;
  assign n48961 = ~pi0983 & n35499;
  assign n48962 = ~pi3426 & n48961;
  assign n48963 = ~n12726 & n48962;
  assign n48964 = pi2215 & ~n48962;
  assign po2528 = n48963 | n48964;
  assign n48966 = ~n13701 & n48962;
  assign n48967 = pi2216 & ~n48962;
  assign po2529 = n48966 | n48967;
  assign n48969 = ~n13121 & n48962;
  assign n48970 = pi2217 & ~n48962;
  assign po2530 = n48969 | n48970;
  assign n48972 = ~n13398 & n48962;
  assign n48973 = pi2218 & ~n48962;
  assign po2531 = n48972 | n48973;
  assign n48975 = ~n13988 & n48962;
  assign n48976 = pi2219 & ~n48962;
  assign po2532 = n48975 | n48976;
  assign n48978 = ~n12415 & n48962;
  assign n48979 = pi2220 & ~n48962;
  assign po2533 = n48978 | n48979;
  assign n48981 = ~n14816 & n48962;
  assign n48982 = pi2221 & ~n48962;
  assign po2534 = n48981 | n48982;
  assign n48984 = ~n15115 & n48962;
  assign n48985 = pi2222 & ~n48962;
  assign po2535 = n48984 | n48985;
  assign n48987 = ~n12061 & n48962;
  assign n48988 = pi2223 & ~n48962;
  assign po2536 = n48987 | n48988;
  assign n48990 = ~n9825 & n48962;
  assign n48991 = pi2224 & ~n48962;
  assign po2537 = n48990 | n48991;
  assign n48993 = ~n10608 & n48962;
  assign n48994 = pi2225 & ~n48962;
  assign po2538 = n48993 | n48994;
  assign n48996 = ~n15426 & n48962;
  assign n48997 = pi2226 & ~n48962;
  assign po2539 = n48996 | n48997;
  assign n48999 = ~n14403 & n48962;
  assign n49000 = pi2227 & ~n48962;
  assign po2540 = n48999 | n49000;
  assign n49002 = ~n11181 & n48962;
  assign n49003 = pi2228 & ~n48962;
  assign po2541 = n49002 | n49003;
  assign n49005 = ~pi1011 & n35463;
  assign n49006 = ~pi3426 & n49005;
  assign n49007 = ~n12726 & n49006;
  assign n49008 = pi2229 & ~n49006;
  assign po2542 = n49007 | n49008;
  assign n49010 = ~n13701 & n49006;
  assign n49011 = pi2230 & ~n49006;
  assign po2543 = n49010 | n49011;
  assign n49013 = ~n13121 & n49006;
  assign n49014 = pi2231 & ~n49006;
  assign po2544 = n49013 | n49014;
  assign n49016 = ~n13398 & n49006;
  assign n49017 = pi2232 & ~n49006;
  assign po2545 = n49016 | n49017;
  assign n49019 = ~n13988 & n49006;
  assign n49020 = pi2233 & ~n49006;
  assign po2546 = n49019 | n49020;
  assign n49022 = ~n12415 & n49006;
  assign n49023 = pi2234 & ~n49006;
  assign po2547 = n49022 | n49023;
  assign n49025 = ~n14816 & n49006;
  assign n49026 = pi2235 & ~n49006;
  assign po2548 = n49025 | n49026;
  assign n49028 = ~n15115 & n49006;
  assign n49029 = pi2236 & ~n49006;
  assign po2549 = n49028 | n49029;
  assign n49031 = ~n12061 & n49006;
  assign n49032 = pi2237 & ~n49006;
  assign po2550 = n49031 | n49032;
  assign n49034 = ~n9825 & n49006;
  assign n49035 = pi2238 & ~n49006;
  assign po2551 = n49034 | n49035;
  assign n49037 = ~n10608 & n49006;
  assign n49038 = pi2239 & ~n49006;
  assign po2552 = n49037 | n49038;
  assign n49040 = ~n15426 & n49006;
  assign n49041 = pi2240 & ~n49006;
  assign po2553 = n49040 | n49041;
  assign n49043 = ~n14403 & n49006;
  assign n49044 = pi2241 & ~n49006;
  assign po2554 = n49043 | n49044;
  assign n49046 = ~n11181 & n49006;
  assign n49047 = pi2242 & ~n49006;
  assign po2555 = n49046 | n49047;
  assign n49049 = ~pi0984 & n35514;
  assign n49050 = ~pi3426 & n49049;
  assign n49051 = ~n12726 & n49050;
  assign n49052 = pi2243 & ~n49050;
  assign po2556 = n49051 | n49052;
  assign n49054 = ~n13701 & n49050;
  assign n49055 = pi2244 & ~n49050;
  assign po2557 = n49054 | n49055;
  assign n49057 = ~n13121 & n49050;
  assign n49058 = pi2245 & ~n49050;
  assign po2558 = n49057 | n49058;
  assign n49060 = ~n13398 & n49050;
  assign n49061 = pi2246 & ~n49050;
  assign po2559 = n49060 | n49061;
  assign n49063 = ~n13988 & n49050;
  assign n49064 = pi2247 & ~n49050;
  assign po2560 = n49063 | n49064;
  assign n49066 = ~n12415 & n49050;
  assign n49067 = pi2248 & ~n49050;
  assign po2561 = n49066 | n49067;
  assign n49069 = ~n14816 & n49050;
  assign n49070 = pi2249 & ~n49050;
  assign po2562 = n49069 | n49070;
  assign n49072 = ~n15115 & n49050;
  assign n49073 = pi2250 & ~n49050;
  assign po2563 = n49072 | n49073;
  assign n49075 = ~n12061 & n49050;
  assign n49076 = pi2251 & ~n49050;
  assign po2564 = n49075 | n49076;
  assign n49078 = ~n9825 & n49050;
  assign n49079 = pi2252 & ~n49050;
  assign po2565 = n49078 | n49079;
  assign n49081 = ~n10608 & n49050;
  assign n49082 = pi2253 & ~n49050;
  assign po2566 = n49081 | n49082;
  assign n49084 = ~n15426 & n49050;
  assign n49085 = pi2254 & ~n49050;
  assign po2567 = n49084 | n49085;
  assign n49087 = ~n14403 & n49050;
  assign n49088 = pi2255 & ~n49050;
  assign po2568 = n49087 | n49088;
  assign n49090 = ~n11181 & n49050;
  assign n49091 = pi2256 & ~n49050;
  assign po2569 = n49090 | n49091;
  assign n49093 = pi0992 & ~pi3426;
  assign n49094 = ~n9391 & ~n49093;
  assign n49095 = ~n9388 & n49094;
  assign n49096 = ~n9394 & ~n49095;
  assign n49097 = ~n37833 & n49096;
  assign n49098 = pi2257 & ~n49096;
  assign po2570 = n49097 | n49098;
  assign n49100 = ~n37586 & n49096;
  assign n49101 = pi2258 & ~n49096;
  assign po2571 = n49100 | n49101;
  assign n49103 = ~n37867 & n49096;
  assign n49104 = pi2259 & ~n49096;
  assign po2572 = n49103 | n49104;
  assign n49106 = ~n37884 & n49096;
  assign n49107 = pi2260 & ~n49096;
  assign po2573 = n49106 | n49107;
  assign n49109 = ~n9407 & ~n9408;
  assign n49110 = pi0993 & ~pi3426;
  assign n49111 = n49109 & ~n49110;
  assign n49112 = ~n9411 & ~n49111;
  assign n49113 = ~n37833 & n49112;
  assign n49114 = pi2261 & ~n49112;
  assign po2574 = n49113 | n49114;
  assign n49116 = ~n37586 & n49112;
  assign n49117 = pi2262 & ~n49112;
  assign po2575 = n49116 | n49117;
  assign n49119 = ~n37850 & n49112;
  assign n49120 = pi2263 & ~n49112;
  assign po2576 = n49119 | n49120;
  assign n49122 = ~n37867 & n49112;
  assign n49123 = pi2264 & ~n49112;
  assign po2577 = n49122 | n49123;
  assign n49125 = ~n37884 & n49112;
  assign n49126 = pi2265 & ~n49112;
  assign po2578 = n49125 | n49126;
  assign n49128 = ~n37901 & n49112;
  assign n49129 = pi2266 & ~n49112;
  assign po2579 = n49128 | n49129;
  assign n49131 = ~n37918 & n49112;
  assign n49132 = pi2267 & ~n49112;
  assign po2580 = n49131 | n49132;
  assign n49134 = ~n37935 & n49112;
  assign n49135 = pi2268 & ~n49112;
  assign po2581 = n49134 | n49135;
  assign n49137 = ~n37613 & n49112;
  assign n49138 = pi2269 & ~n49112;
  assign po2582 = n49137 | n49138;
  assign n49140 = ~n37952 & n49112;
  assign n49141 = pi2270 & ~n49112;
  assign po2583 = n49140 | n49141;
  assign n49143 = pi0994 & ~pi3426;
  assign n49144 = ~n9369 & ~n49143;
  assign n49145 = ~n9364 & n49144;
  assign n49146 = ~n9372 & ~n49145;
  assign n49147 = ~n37833 & n49146;
  assign n49148 = pi2271 & ~n49146;
  assign po2584 = n49147 | n49148;
  assign n49150 = ~n37586 & n49146;
  assign n49151 = pi2272 & ~n49146;
  assign po2585 = n49150 | n49151;
  assign n49153 = ~n37867 & n49146;
  assign n49154 = pi2273 & ~n49146;
  assign po2586 = n49153 | n49154;
  assign n49156 = ~n37901 & n49146;
  assign n49157 = pi2274 & ~n49146;
  assign po2587 = n49156 | n49157;
  assign n49159 = ~n39032 & n47806;
  assign n49160 = pi2275 & ~n47806;
  assign po2588 = n49159 | n49160;
  assign n49162 = ~n39047 & n47806;
  assign n49163 = pi2276 & ~n47806;
  assign po2589 = n49162 | n49163;
  assign n49165 = ~n39062 & n47806;
  assign n49166 = pi2277 & ~n47806;
  assign po2590 = n49165 | n49166;
  assign n49168 = ~n39077 & n47806;
  assign n49169 = pi2278 & ~n47806;
  assign po2591 = n49168 | n49169;
  assign n49171 = ~n12726 & n48282;
  assign n49172 = pi2279 & ~n48282;
  assign po2592 = n49171 | n49172;
  assign n49174 = ~n13701 & n48282;
  assign n49175 = pi2280 & ~n48282;
  assign po2593 = n49174 | n49175;
  assign n49177 = ~n13121 & n48282;
  assign n49178 = pi2281 & ~n48282;
  assign po2594 = n49177 | n49178;
  assign n49180 = ~n13398 & n48282;
  assign n49181 = pi2282 & ~n48282;
  assign po2595 = n49180 | n49181;
  assign n49183 = ~n13988 & n48282;
  assign n49184 = pi2283 & ~n48282;
  assign po2596 = n49183 | n49184;
  assign n49186 = ~n12415 & n48282;
  assign n49187 = pi2284 & ~n48282;
  assign po2597 = n49186 | n49187;
  assign n49189 = ~n14816 & n48282;
  assign n49190 = pi2285 & ~n48282;
  assign po2598 = n49189 | n49190;
  assign n49192 = ~n15115 & n48282;
  assign n49193 = pi2286 & ~n48282;
  assign po2599 = n49192 | n49193;
  assign n49195 = ~n9825 & n48282;
  assign n49196 = pi2287 & ~n48282;
  assign po2600 = n49195 | n49196;
  assign n49198 = ~n10608 & n48282;
  assign n49199 = pi2288 & ~n48282;
  assign po2601 = n49198 | n49199;
  assign n49201 = ~n15426 & n48282;
  assign n49202 = pi2289 & ~n48282;
  assign po2602 = n49201 | n49202;
  assign n49204 = ~n14403 & n48282;
  assign n49205 = pi2290 & ~n48282;
  assign po2603 = n49204 | n49205;
  assign n49207 = ~n11181 & n48282;
  assign n49208 = pi2291 & ~n48282;
  assign po2604 = n49207 | n49208;
  assign n49210 = ~n12726 & n48277;
  assign n49211 = pi2292 & ~n48277;
  assign po2605 = n49210 | n49211;
  assign n49213 = ~n13121 & n48277;
  assign n49214 = pi2293 & ~n48277;
  assign po2606 = n49213 | n49214;
  assign n49216 = ~n13398 & n48277;
  assign n49217 = pi2294 & ~n48277;
  assign po2607 = n49216 | n49217;
  assign n49219 = ~n13988 & n48277;
  assign n49220 = pi2295 & ~n48277;
  assign po2608 = n49219 | n49220;
  assign n49222 = ~n12415 & n48277;
  assign n49223 = pi2296 & ~n48277;
  assign po2609 = n49222 | n49223;
  assign n49225 = ~n14816 & n48277;
  assign n49226 = pi2297 & ~n48277;
  assign po2610 = n49225 | n49226;
  assign n49228 = ~n15115 & n48277;
  assign n49229 = pi2298 & ~n48277;
  assign po2611 = n49228 | n49229;
  assign n49231 = ~n12061 & n48277;
  assign n49232 = pi2299 & ~n48277;
  assign po2612 = n49231 | n49232;
  assign n49234 = ~n9825 & n48277;
  assign n49235 = pi2300 & ~n48277;
  assign po2613 = n49234 | n49235;
  assign n49237 = ~n14403 & n48277;
  assign n49238 = pi2301 & ~n48277;
  assign po2614 = n49237 | n49238;
  assign n49240 = ~n11181 & n48277;
  assign n49241 = pi2302 & ~n48277;
  assign po2615 = n49240 | n49241;
  assign n49243 = ~n12726 & n48423;
  assign n49244 = pi2303 & ~n48423;
  assign po2616 = n49243 | n49244;
  assign n49246 = ~n13121 & n48423;
  assign n49247 = pi2304 & ~n48423;
  assign po2617 = n49246 | n49247;
  assign n49249 = ~n13398 & n48423;
  assign n49250 = pi2305 & ~n48423;
  assign po2618 = n49249 | n49250;
  assign n49252 = ~n14816 & n48423;
  assign n49253 = pi2306 & ~n48423;
  assign po2619 = n49252 | n49253;
  assign n49255 = ~n15115 & n48423;
  assign n49256 = pi2307 & ~n48423;
  assign po2620 = n49255 | n49256;
  assign n49258 = ~n12061 & n48423;
  assign n49259 = pi2308 & ~n48423;
  assign po2621 = n49258 | n49259;
  assign n49261 = ~n9825 & n48423;
  assign n49262 = pi2309 & ~n48423;
  assign po2622 = n49261 | n49262;
  assign n49264 = ~n10608 & n48423;
  assign n49265 = pi2310 & ~n48423;
  assign po2623 = n49264 | n49265;
  assign n49267 = ~n15426 & n48423;
  assign n49268 = pi2311 & ~n48423;
  assign po2624 = n49267 | n49268;
  assign n49270 = ~n14403 & n48423;
  assign n49271 = pi2312 & ~n48423;
  assign po2625 = n49270 | n49271;
  assign n49273 = ~n11181 & n48423;
  assign n49274 = pi2313 & ~n48423;
  assign po2626 = n49273 | n49274;
  assign n49276 = ~pi0945 & n35630;
  assign n49277 = ~pi3426 & n49276;
  assign n49278 = ~n12726 & n49277;
  assign n49279 = pi2314 & ~n49277;
  assign po2627 = n49278 | n49279;
  assign n49281 = ~n13701 & n49277;
  assign n49282 = pi2315 & ~n49277;
  assign po2628 = n49281 | n49282;
  assign n49284 = ~n13121 & n49277;
  assign n49285 = pi2316 & ~n49277;
  assign po2629 = n49284 | n49285;
  assign n49287 = ~n13398 & n49277;
  assign n49288 = pi2317 & ~n49277;
  assign po2630 = n49287 | n49288;
  assign n49290 = ~n13988 & n49277;
  assign n49291 = pi2318 & ~n49277;
  assign po2631 = n49290 | n49291;
  assign n49293 = ~n12415 & n49277;
  assign n49294 = pi2319 & ~n49277;
  assign po2632 = n49293 | n49294;
  assign n49296 = ~n14816 & n49277;
  assign n49297 = pi2320 & ~n49277;
  assign po2633 = n49296 | n49297;
  assign n49299 = ~n15115 & n49277;
  assign n49300 = pi2321 & ~n49277;
  assign po2634 = n49299 | n49300;
  assign n49302 = ~n12061 & n49277;
  assign n49303 = pi2322 & ~n49277;
  assign po2635 = n49302 | n49303;
  assign n49305 = ~n9825 & n49277;
  assign n49306 = pi2323 & ~n49277;
  assign po2636 = n49305 | n49306;
  assign n49308 = ~n10608 & n49277;
  assign n49309 = pi2324 & ~n49277;
  assign po2637 = n49308 | n49309;
  assign n49311 = ~n15426 & n49277;
  assign n49312 = pi2325 & ~n49277;
  assign po2638 = n49311 | n49312;
  assign n49314 = ~n14403 & n49277;
  assign n49315 = pi2326 & ~n49277;
  assign po2639 = n49314 | n49315;
  assign n49317 = ~n11181 & n49277;
  assign n49318 = pi2327 & ~n49277;
  assign po2640 = n49317 | n49318;
  assign n49320 = ~pi2328 & ~n46586;
  assign n49321 = pi2472 & n46972;
  assign n49322 = ~pi2328 & ~n46972;
  assign n49323 = ~n49321 & ~n49322;
  assign n49324 = n46586 & ~n49323;
  assign po2641 = n49320 | n49324;
  assign n49326 = ~pi2329 & ~n46586;
  assign n49327 = pi2400 & n46972;
  assign n49328 = ~pi2329 & ~n46972;
  assign n49329 = ~n49327 & ~n49328;
  assign n49330 = n46586 & ~n49329;
  assign po2642 = n49326 | n49330;
  assign n49332 = pi3517 & n46972;
  assign n49333 = pi2330 & ~n46972;
  assign n49334 = ~n49332 & ~n49333;
  assign n49335 = n46586 & ~n49334;
  assign n49336 = pi2330 & ~n46586;
  assign po2643 = n49335 | n49336;
  assign n49338 = pi3508 & n46972;
  assign n49339 = pi2331 & ~n46972;
  assign n49340 = ~n49338 & ~n49339;
  assign n49341 = n46586 & ~n49340;
  assign n49342 = pi2331 & ~n46586;
  assign po2644 = n49341 | n49342;
  assign n49344 = pi3509 & n46972;
  assign n49345 = pi2332 & ~n46972;
  assign n49346 = ~n49344 & ~n49345;
  assign n49347 = n46586 & ~n49346;
  assign n49348 = pi2332 & ~n46586;
  assign po2645 = n49347 | n49348;
  assign n49350 = pi3521 & n46972;
  assign n49351 = pi2333 & ~n46972;
  assign n49352 = ~n49350 & ~n49351;
  assign n49353 = n46586 & ~n49352;
  assign n49354 = pi2333 & ~n46586;
  assign po2646 = n49353 | n49354;
  assign n49356 = pi3510 & n46972;
  assign n49357 = pi2334 & ~n46972;
  assign n49358 = ~n49356 & ~n49357;
  assign n49359 = n46586 & ~n49358;
  assign n49360 = pi2334 & ~n46586;
  assign po2647 = n49359 | n49360;
  assign n49362 = ~pi2335 & ~n46586;
  assign n49363 = pi2408 & n46972;
  assign n49364 = ~pi2335 & ~n46972;
  assign n49365 = ~n49363 & ~n49364;
  assign n49366 = n46586 & ~n49365;
  assign po2648 = n49362 | n49366;
  assign n49368 = pi3520 & n47897;
  assign n49369 = pi2336 & ~n47897;
  assign n49370 = ~n49368 & ~n49369;
  assign n49371 = n46586 & ~n49370;
  assign n49372 = pi2336 & ~n46586;
  assign po2649 = n49371 | n49372;
  assign n49374 = pi3398 & n47897;
  assign n49375 = pi2337 & ~n47897;
  assign n49376 = ~n49374 & ~n49375;
  assign n49377 = n46586 & ~n49376;
  assign n49378 = pi2337 & ~n46586;
  assign po2650 = n49377 | n49378;
  assign n49380 = ~pi2338 & ~n46586;
  assign n49381 = pi2514 & n47897;
  assign n49382 = ~pi2338 & ~n47897;
  assign n49383 = ~n49381 & ~n49382;
  assign n49384 = n46586 & ~n49383;
  assign po2651 = n49380 | n49384;
  assign n49386 = pi3512 & n47897;
  assign n49387 = pi2339 & ~n47897;
  assign n49388 = ~n49386 & ~n49387;
  assign n49389 = n46586 & ~n49388;
  assign n49390 = pi2339 & ~n46586;
  assign po2652 = n49389 | n49390;
  assign n49392 = ~pi2340 & ~n46586;
  assign n49393 = pi2400 & n47897;
  assign n49394 = ~pi2340 & ~n47897;
  assign n49395 = ~n49393 & ~n49394;
  assign n49396 = n46586 & ~n49395;
  assign po2653 = n49392 | n49396;
  assign n49398 = pi3513 & n47897;
  assign n49399 = pi2341 & ~n47897;
  assign n49400 = ~n49398 & ~n49399;
  assign n49401 = n46586 & ~n49400;
  assign n49402 = pi2341 & ~n46586;
  assign po2654 = n49401 | n49402;
  assign n49404 = pi3504 & n47897;
  assign n49405 = pi2342 & ~n47897;
  assign n49406 = ~n49404 & ~n49405;
  assign n49407 = n46586 & ~n49406;
  assign n49408 = pi2342 & ~n46586;
  assign po2655 = n49407 | n49408;
  assign n49410 = pi3514 & n47897;
  assign n49411 = pi2343 & ~n47897;
  assign n49412 = ~n49410 & ~n49411;
  assign n49413 = n46586 & ~n49412;
  assign n49414 = pi2343 & ~n46586;
  assign po2656 = n49413 | n49414;
  assign n49416 = pi3518 & n47897;
  assign n49417 = pi2344 & ~n47897;
  assign n49418 = ~n49416 & ~n49417;
  assign n49419 = n46586 & ~n49418;
  assign n49420 = pi2344 & ~n46586;
  assign po2657 = n49419 | n49420;
  assign n49422 = pi3516 & n47897;
  assign n49423 = pi2345 & ~n47897;
  assign n49424 = ~n49422 & ~n49423;
  assign n49425 = n46586 & ~n49424;
  assign n49426 = pi2345 & ~n46586;
  assign po2658 = n49425 | n49426;
  assign n49428 = pi3517 & n47897;
  assign n49429 = pi2346 & ~n47897;
  assign n49430 = ~n49428 & ~n49429;
  assign n49431 = n46586 & ~n49430;
  assign n49432 = pi2346 & ~n46586;
  assign po2659 = n49431 | n49432;
  assign n49434 = pi3508 & n47897;
  assign n49435 = pi2347 & ~n47897;
  assign n49436 = ~n49434 & ~n49435;
  assign n49437 = n46586 & ~n49436;
  assign n49438 = pi2347 & ~n46586;
  assign po2660 = n49437 | n49438;
  assign n49440 = pi3509 & n47897;
  assign n49441 = pi2348 & ~n47897;
  assign n49442 = ~n49440 & ~n49441;
  assign n49443 = n46586 & ~n49442;
  assign n49444 = pi2348 & ~n46586;
  assign po2661 = n49443 | n49444;
  assign n49446 = pi3521 & n47897;
  assign n49447 = pi2349 & ~n47897;
  assign n49448 = ~n49446 & ~n49447;
  assign n49449 = n46586 & ~n49448;
  assign n49450 = pi2349 & ~n46586;
  assign po2662 = n49449 | n49450;
  assign n49452 = pi3510 & n47897;
  assign n49453 = pi2350 & ~n47897;
  assign n49454 = ~n49452 & ~n49453;
  assign n49455 = n46586 & ~n49454;
  assign n49456 = pi2350 & ~n46586;
  assign po2663 = n49455 | n49456;
  assign n49458 = pi3520 & n46979;
  assign n49459 = pi2351 & ~n46979;
  assign n49460 = ~n49458 & ~n49459;
  assign n49461 = n46586 & ~n49460;
  assign n49462 = pi2351 & ~n46586;
  assign po2664 = n49461 | n49462;
  assign n49464 = pi3398 & n46979;
  assign n49465 = pi2352 & ~n46979;
  assign n49466 = ~n49464 & ~n49465;
  assign n49467 = n46586 & ~n49466;
  assign n49468 = pi2352 & ~n46586;
  assign po2665 = n49467 | n49468;
  assign n49470 = ~pi2353 & ~n46586;
  assign n49471 = pi2472 & n46979;
  assign n49472 = ~pi2353 & ~n46979;
  assign n49473 = ~n49471 & ~n49472;
  assign n49474 = n46586 & ~n49473;
  assign po2666 = n49470 | n49474;
  assign n49476 = ~pi2354 & ~n46586;
  assign n49477 = pi2400 & n46979;
  assign n49478 = ~pi2354 & ~n46979;
  assign n49479 = ~n49477 & ~n49478;
  assign n49480 = n46586 & ~n49479;
  assign po2667 = n49476 | n49480;
  assign n49482 = pi3504 & n46979;
  assign n49483 = pi2355 & ~n46979;
  assign n49484 = ~n49482 & ~n49483;
  assign n49485 = n46586 & ~n49484;
  assign n49486 = pi2355 & ~n46586;
  assign po2668 = n49485 | n49486;
  assign n49488 = pi3518 & n46979;
  assign n49489 = pi2356 & ~n46979;
  assign n49490 = ~n49488 & ~n49489;
  assign n49491 = n46586 & ~n49490;
  assign n49492 = pi2356 & ~n46586;
  assign po2669 = n49491 | n49492;
  assign n49494 = pi3508 & n46979;
  assign n49495 = pi2357 & ~n46979;
  assign n49496 = ~n49494 & ~n49495;
  assign n49497 = n46586 & ~n49496;
  assign n49498 = pi2357 & ~n46586;
  assign po2670 = n49497 | n49498;
  assign n49500 = ~pi2358 & ~n46586;
  assign n49501 = pi2408 & n46979;
  assign n49502 = ~pi2358 & ~n46979;
  assign n49503 = ~n49501 & ~n49502;
  assign n49504 = n46586 & ~n49503;
  assign po2671 = n49500 | n49504;
  assign n49506 = pi3520 & n47970;
  assign n49507 = pi2359 & ~n47970;
  assign n49508 = ~n49506 & ~n49507;
  assign n49509 = n46586 & ~n49508;
  assign n49510 = pi2359 & ~n46586;
  assign po2672 = n49509 | n49510;
  assign n49512 = pi3398 & n47970;
  assign n49513 = pi2360 & ~n47970;
  assign n49514 = ~n49512 & ~n49513;
  assign n49515 = n46586 & ~n49514;
  assign n49516 = pi2360 & ~n46586;
  assign po2673 = n49515 | n49516;
  assign n49518 = pi3392 & n47970;
  assign n49519 = pi2361 & ~n47970;
  assign n49520 = ~n49518 & ~n49519;
  assign n49521 = n46586 & ~n49520;
  assign n49522 = pi2361 & ~n46586;
  assign po2674 = n49521 | n49522;
  assign n49524 = ~pi2362 & ~n46586;
  assign n49525 = pi2514 & n47970;
  assign n49526 = ~pi2362 & ~n47970;
  assign n49527 = ~n49525 & ~n49526;
  assign n49528 = n46586 & ~n49527;
  assign po2675 = n49524 | n49528;
  assign n49530 = pi2363 & ~n47970;
  assign n49531 = pi3512 & n47970;
  assign n49532 = ~n49530 & ~n49531;
  assign n49533 = n46586 & ~n49532;
  assign n49534 = pi2363 & ~n46586;
  assign po2676 = n49533 | n49534;
  assign n49536 = ~pi2364 & ~n46586;
  assign n49537 = pi2400 & n47970;
  assign n49538 = ~pi2364 & ~n47970;
  assign n49539 = ~n49537 & ~n49538;
  assign n49540 = n46586 & ~n49539;
  assign po2677 = n49536 | n49540;
  assign n49542 = pi3513 & n47970;
  assign n49543 = pi2365 & ~n47970;
  assign n49544 = ~n49542 & ~n49543;
  assign n49545 = n46586 & ~n49544;
  assign n49546 = pi2365 & ~n46586;
  assign po2678 = n49545 | n49546;
  assign n49548 = pi3514 & n47970;
  assign n49549 = pi2366 & ~n47970;
  assign n49550 = ~n49548 & ~n49549;
  assign n49551 = n46586 & ~n49550;
  assign n49552 = pi2366 & ~n46586;
  assign po2679 = n49551 | n49552;
  assign n49554 = pi3518 & n47970;
  assign n49555 = pi2367 & ~n47970;
  assign n49556 = ~n49554 & ~n49555;
  assign n49557 = n46586 & ~n49556;
  assign n49558 = pi2367 & ~n46586;
  assign po2680 = n49557 | n49558;
  assign n49560 = pi3517 & n47970;
  assign n49561 = pi2368 & ~n47970;
  assign n49562 = ~n49560 & ~n49561;
  assign n49563 = n46586 & ~n49562;
  assign n49564 = pi2368 & ~n46586;
  assign po2681 = n49563 | n49564;
  assign n49566 = pi3508 & n47970;
  assign n49567 = pi2369 & ~n47970;
  assign n49568 = ~n49566 & ~n49567;
  assign n49569 = n46586 & ~n49568;
  assign n49570 = pi2369 & ~n46586;
  assign po2682 = n49569 | n49570;
  assign n49572 = pi3509 & n47970;
  assign n49573 = pi2370 & ~n47970;
  assign n49574 = ~n49572 & ~n49573;
  assign n49575 = n46586 & ~n49574;
  assign n49576 = pi2370 & ~n46586;
  assign po2683 = n49575 | n49576;
  assign n49578 = pi3521 & n47970;
  assign n49579 = pi2371 & ~n47970;
  assign n49580 = ~n49578 & ~n49579;
  assign n49581 = n46586 & ~n49580;
  assign n49582 = pi2371 & ~n46586;
  assign po2684 = n49581 | n49582;
  assign n49584 = pi3510 & n47970;
  assign n49585 = pi2372 & ~n47970;
  assign n49586 = ~n49584 & ~n49585;
  assign n49587 = n46586 & ~n49586;
  assign n49588 = pi2372 & ~n46586;
  assign po2685 = n49587 | n49588;
  assign n49590 = n9415 & ~n14152;
  assign n49591 = ~n9415 & ~n13701;
  assign n49592 = ~n49590 & ~n49591;
  assign n49593 = n9361 & n49592;
  assign n49594 = ~n9415 & ~n14134;
  assign n49595 = ~n49590 & ~n49594;
  assign n49596 = ~n9361 & n49595;
  assign n49597 = ~n49593 & ~n49596;
  assign n49598 = n9377 & n49597;
  assign n49599 = pi0406 & n47131;
  assign n49600 = ~n49598 & ~n49599;
  assign n49601 = po3831 & ~n49600;
  assign n49602 = pi2373 & ~po3831;
  assign po2686 = n49601 | n49602;
  assign n49604 = n9415 & ~n13424;
  assign n49605 = ~n9415 & ~n13398;
  assign n49606 = ~n49604 & ~n49605;
  assign n49607 = n9361 & n49606;
  assign n49608 = ~n9415 & ~n13451;
  assign n49609 = ~n49604 & ~n49608;
  assign n49610 = ~n9361 & n49609;
  assign n49611 = ~n49607 & ~n49610;
  assign n49612 = n9377 & n49611;
  assign n49613 = pi0426 & n47131;
  assign n49614 = ~n49612 & ~n49613;
  assign n49615 = po3831 & ~n49614;
  assign n49616 = pi2374 & ~po3831;
  assign po2687 = n49615 | n49616;
  assign n49618 = n9377 & n36443;
  assign n49619 = pi0421 & n47131;
  assign n49620 = ~n49618 & ~n49619;
  assign n49621 = po3831 & ~n49620;
  assign n49622 = pi2375 & ~po3831;
  assign po2688 = n49621 | n49622;
  assign n49624 = n9377 & n36451;
  assign n49625 = pi0405 & n47131;
  assign n49626 = ~n49624 & ~n49625;
  assign n49627 = po3831 & ~n49626;
  assign n49628 = pi2376 & ~po3831;
  assign po2689 = n49627 | n49628;
  assign n49630 = n9415 & ~n14857;
  assign n49631 = ~n9415 & ~n15426;
  assign n49632 = ~n49630 & ~n49631;
  assign n49633 = n9361 & n49632;
  assign n49634 = ~n9415 & ~n15146;
  assign n49635 = ~n49630 & ~n49634;
  assign n49636 = ~n9361 & n49635;
  assign n49637 = ~n49633 & ~n49636;
  assign n49638 = n9377 & n49637;
  assign n49639 = pi0422 & n47131;
  assign n49640 = ~n49638 & ~n49639;
  assign n49641 = po3831 & ~n49640;
  assign n49642 = pi2377 & ~po3831;
  assign po2690 = n49641 | n49642;
  assign n49644 = n9415 & ~n14502;
  assign n49645 = ~n9415 & ~n14403;
  assign n49646 = ~n49644 & ~n49645;
  assign n49647 = n9361 & n49646;
  assign n49648 = ~n9415 & ~n14458;
  assign n49649 = ~n49644 & ~n49648;
  assign n49650 = ~n9361 & n49649;
  assign n49651 = ~n49647 & ~n49650;
  assign n49652 = n9377 & n49651;
  assign n49653 = pi0423 & n47131;
  assign n49654 = ~n49652 & ~n49653;
  assign n49655 = po3831 & ~n49654;
  assign n49656 = pi2378 & ~po3831;
  assign po2691 = n49655 | n49656;
  assign n49658 = ~pi2379 & ~n42183;
  assign n49659 = n20363 & n49658;
  assign n49660 = pi2379 & ~n49658;
  assign po2692 = n49659 | n49660;
  assign n49662 = pi1093 & n20355;
  assign n49663 = ~n19549 & ~n49662;
  assign n49664 = ~n19544 & ~n19546;
  assign n49665 = ~n9352 & ~n49664;
  assign n49666 = ~n41535 & ~n49665;
  assign n49667 = ~n9352 & ~n19547;
  assign n49668 = ~n49666 & n49667;
  assign n49669 = ~n49663 & n49668;
  assign n49670 = pi2380 & n49666;
  assign po2693 = n49669 | n49670;
  assign n49672 = pi3328 & pi3541;
  assign n49673 = ~pi3213 & ~n49672;
  assign n49674 = ~pi3328 & n49673;
  assign n49675 = pi2777 & ~po3627;
  assign n49676 = ~pi2974 & pi3328;
  assign n49677 = ~n49675 & ~n49676;
  assign n49678 = ~pi2381 & pi3328;
  assign n49679 = n49677 & n49678;
  assign n49680 = ~n49674 & ~n49679;
  assign n49681 = ~pi3375 & ~n49673;
  assign n49682 = n49677 & ~n49681;
  assign n49683 = pi3328 & n49682;
  assign po2694 = ~n49680 | n49683;
  assign n49685 = pi2382 & n8561;
  assign n49686 = ~n10808 & ~n10811;
  assign n49687 = n35527 & ~n35534;
  assign n49688 = n49686 & n49687;
  assign n49689 = n35528 & n49688;
  assign n49690 = ~n8561 & ~n49689;
  assign n49691 = ~n49685 & ~n49690;
  assign po2695 = po3627 & ~n49691;
  assign n49693 = ~n8561 & n9345;
  assign n49694 = n36116 & n49693;
  assign n49695 = pi0414 & n49694;
  assign n49696 = ~pi2383 & n8561;
  assign n49697 = ~n49695 & ~n49696;
  assign po2696 = po3627 & ~n49697;
  assign n49699 = pi2384 & n8561;
  assign n49700 = ~n25623 & ~n49699;
  assign po2697 = po3627 & ~n49700;
  assign n49702 = n38725 & n38736;
  assign n49703 = pi3502 & n38740;
  assign n49704 = n38732 & n49703;
  assign n49705 = n38723 & n49704;
  assign n49706 = n49702 & n49705;
  assign po3574 = n38738 & n49706;
  assign n49708 = n38781 & po3574;
  assign n49709 = pi0853 & n49708;
  assign n49710 = pi2385 & ~n49708;
  assign po2698 = n49709 | n49710;
  assign po2699 = pi1835 | ~po3853;
  assign n49713 = pi1838 & pi2760;
  assign n49714 = ~pi1838 & ~pi2760;
  assign n49715 = ~n49713 & ~n49714;
  assign n49716 = pi1705 & pi2506;
  assign n49717 = ~pi1705 & ~pi2506;
  assign n49718 = ~n49716 & ~n49717;
  assign n49719 = n49715 & n49718;
  assign n49720 = pi1828 & pi2771;
  assign n49721 = ~pi1828 & ~pi2771;
  assign n49722 = ~n49720 & ~n49721;
  assign n49723 = pi1829 & pi2523;
  assign n49724 = ~pi1829 & ~pi2523;
  assign n49725 = ~n49723 & ~n49724;
  assign n49726 = n49722 & n49725;
  assign n49727 = pi1836 & pi2507;
  assign n49728 = ~pi1836 & ~pi2507;
  assign n49729 = ~n49727 & ~n49728;
  assign n49730 = pi1837 & pi2772;
  assign n49731 = ~pi1837 & ~pi2772;
  assign n49732 = ~n49730 & ~n49731;
  assign n49733 = n49729 & n49732;
  assign n49734 = ~pi1792 & pi2770;
  assign n49735 = pi1792 & ~pi2770;
  assign n49736 = ~n49734 & ~n49735;
  assign n49737 = n49733 & ~n49736;
  assign n49738 = n49726 & n49737;
  assign n49739 = n49719 & n49738;
  assign n49740 = pi2386 & ~n49739;
  assign n49741 = ~pi2386 & n49739;
  assign po2700 = n49740 | n49741;
  assign n49743 = pi3510 & n46979;
  assign n49744 = pi2388 & ~n46979;
  assign n49745 = ~n49743 & ~n49744;
  assign n49746 = n46586 & ~n49745;
  assign n49747 = pi2388 & ~n46586;
  assign po2702 = n49746 | n49747;
  assign n49749 = pi3511 & n47970;
  assign n49750 = pi2389 & ~n47970;
  assign n49751 = ~n49749 & ~n49750;
  assign n49752 = n46586 & ~n49751;
  assign n49753 = pi2389 & ~n46586;
  assign po2703 = n49752 | n49753;
  assign n49755 = pi3519 & n46979;
  assign n49756 = pi2390 & ~n46979;
  assign n49757 = ~n49755 & ~n49756;
  assign n49758 = n46586 & ~n49757;
  assign n49759 = pi2390 & ~n46586;
  assign po2704 = n49758 | n49759;
  assign n49761 = pi3513 & n46979;
  assign n49762 = pi2391 & ~n46979;
  assign n49763 = ~n49761 & ~n49762;
  assign n49764 = n46586 & ~n49763;
  assign n49765 = pi2391 & ~n46586;
  assign po2705 = n49764 | n49765;
  assign n49767 = n9415 & ~n12163;
  assign n49768 = ~n9415 & ~n12726;
  assign n49769 = ~n49767 & ~n49768;
  assign n49770 = n9361 & n49769;
  assign n49771 = ~n9415 & ~n12445;
  assign n49772 = ~n49767 & ~n49771;
  assign n49773 = ~n9361 & n49772;
  assign n49774 = ~n49770 & ~n49773;
  assign n49775 = n9377 & n49774;
  assign n49776 = pi0424 & n47131;
  assign n49777 = ~n49775 & ~n49776;
  assign n49778 = po3831 & ~n49777;
  assign n49779 = pi2392 & ~po3831;
  assign po2706 = n49778 | n49779;
  assign n49781 = ~pi2393 & ~n47395;
  assign n49782 = ~n13988 & n47395;
  assign po2707 = n49781 | n49782;
  assign n49784 = ~pi2394 & ~n47395;
  assign n49785 = ~n17199 & n47395;
  assign po2708 = n49784 | n49785;
  assign n49787 = ~pi2395 & ~n47395;
  assign n49788 = ~n14403 & n47395;
  assign po2709 = n49787 | n49788;
  assign n49790 = ~pi2396 & ~n47395;
  assign n49791 = ~n12061 & n47395;
  assign po2710 = n49790 | n49791;
  assign n49793 = ~pi2397 & ~n47395;
  assign n49794 = ~n14816 & n47395;
  assign po2711 = n49793 | n49794;
  assign n49796 = ~pi2398 & ~n47395;
  assign n49797 = ~n13121 & n47395;
  assign po2712 = n49796 | n49797;
  assign n49799 = ~n14816 & ~n15115;
  assign n49800 = ~n11181 & n49799;
  assign n49801 = ~n12061 & n49800;
  assign n49802 = ~pi0944 & n9365;
  assign n49803 = ~n49801 & n49802;
  assign n49804 = ~n12061 & n49803;
  assign n49805 = pi2400 & ~n49803;
  assign po2714 = n49804 | n49805;
  assign n49807 = ~pi2976 & pi3361;
  assign n49808 = ~n36205 & ~n49807;
  assign n49809 = pi3361 & n49808;
  assign n49810 = ~pi2401 & n49809;
  assign n49811 = ~pi1931 & pi3361;
  assign n49812 = pi3361 & pi3543;
  assign n49813 = ~pi3212 & ~n49812;
  assign n49814 = pi3189 & ~n49813;
  assign n49815 = n49811 & ~n49814;
  assign n49816 = n49808 & n49815;
  assign n49817 = ~pi3361 & n49813;
  assign n49818 = ~n49816 & ~n49817;
  assign po2715 = n49810 | ~n49818;
  assign n49820 = ~pi3442 & ~pi3537;
  assign n49821 = ~pi2100 & ~n49820;
  assign n49822 = pi2402 & n49821;
  assign n49823 = pi3269 & ~po3627;
  assign po2716 = ~n49822 & ~n49823;
  assign n49825 = ~pi3239 & pi3360;
  assign n49826 = ~n36512 & ~n49825;
  assign n49827 = pi3360 & n49826;
  assign n49828 = ~pi2403 & n49827;
  assign n49829 = ~pi1931 & pi3360;
  assign n49830 = pi3360 & pi3542;
  assign n49831 = ~pi3232 & ~n49830;
  assign n49832 = pi3226 & ~n49831;
  assign n49833 = n49829 & ~n49832;
  assign n49834 = n49826 & n49833;
  assign n49835 = ~pi3360 & n49831;
  assign n49836 = ~n49834 & ~n49835;
  assign po2717 = n49828 | ~n49836;
  assign n49838 = ~n13121 & ~n13988;
  assign n49839 = ~n12415 & n49838;
  assign n49840 = ~n13398 & n49839;
  assign n49841 = n49802 & ~n49840;
  assign n49842 = ~n13988 & n49841;
  assign n49843 = pi2404 & ~n49841;
  assign po2718 = n49842 | n49843;
  assign n49845 = ~n12415 & n49841;
  assign n49846 = pi2405 & ~n49841;
  assign po2719 = n49845 | n49846;
  assign n49848 = ~pi2406 & ~n46586;
  assign n49849 = pi2472 & n47897;
  assign n49850 = ~pi2406 & ~n47897;
  assign n49851 = ~n49849 & ~n49850;
  assign n49852 = n46586 & ~n49851;
  assign po2720 = n49848 | n49852;
  assign n49854 = ~pi2407 & ~n46586;
  assign n49855 = pi2472 & n47970;
  assign n49856 = ~pi2407 & ~n47970;
  assign n49857 = ~n49855 & ~n49856;
  assign n49858 = n46586 & ~n49857;
  assign po2721 = n49854 | n49858;
  assign n49860 = ~n11181 & n49803;
  assign n49861 = pi2408 & ~n49803;
  assign po2722 = n49860 | n49861;
  assign n49863 = ~n13121 & n49841;
  assign n49864 = pi2409 & ~n49841;
  assign po2723 = n49863 | n49864;
  assign n49866 = pi0999 & ~pi3426;
  assign n49867 = ~n10830 & ~n49866;
  assign n49868 = ~n10834 & n49867;
  assign n49869 = ~n10835 & ~n49868;
  assign n49870 = n38156 & n49869;
  assign n49871 = pi2410 & ~n49869;
  assign po2724 = n49870 | n49871;
  assign n49873 = ~n38488 & n49869;
  assign n49874 = pi2411 & ~n49869;
  assign po2725 = n49873 | n49874;
  assign n49876 = n38095 & n49869;
  assign n49877 = pi2412 & ~n49869;
  assign po2726 = n49876 | n49877;
  assign n49879 = ~n38413 & n49869;
  assign n49880 = pi2413 & ~n49869;
  assign po2727 = n49879 | n49880;
  assign n49882 = pi3691 & n47620;
  assign n49883 = pi2414 & ~n47620;
  assign po2728 = n49882 | n49883;
  assign n49885 = ~n8589 & n9424;
  assign n49886 = ~n8577 & n49885;
  assign n49887 = ~n8567 & ~n49886;
  assign n49888 = ~n9352 & n49887;
  assign n49889 = pi2796 & pi3245;
  assign n49890 = pi1029 & ~pi3245;
  assign n49891 = ~n49889 & ~n49890;
  assign n49892 = n49888 & ~n49891;
  assign n49893 = pi2415 & ~n49888;
  assign po2729 = n49892 | n49893;
  assign n49895 = ~pi2416 & ~n42536;
  assign n49896 = ~pi3290 & n46883;
  assign n49897 = pi2416 & n49896;
  assign n49898 = ~pi2416 & ~n49896;
  assign n49899 = ~n49897 & ~n49898;
  assign n49900 = n42536 & ~n49899;
  assign po2730 = n49895 | n49900;
  assign n49902 = ~n8561 & ~n36385;
  assign n49903 = ~pi2417 & n8561;
  assign po2731 = n49902 | n49903;
  assign n49905 = pi3692 & n47620;
  assign n49906 = pi2418 & ~n47620;
  assign po2732 = n49905 | n49906;
  assign n49908 = pi2419 & ~n46873;
  assign n49909 = ~n48590 & n49908;
  assign po2733 = n48599 | n49909;
  assign n49911 = n30709 & n47655;
  assign n49912 = pi2420 & ~n30709;
  assign po2734 = n49911 | n49912;
  assign n49914 = n30709 & n47664;
  assign n49915 = pi2421 & ~n30709;
  assign po2735 = n49914 | n49915;
  assign n49917 = n30709 & n47673;
  assign n49918 = pi2422 & ~n30709;
  assign po2736 = n49917 | n49918;
  assign n49920 = n30709 & n47682;
  assign n49921 = pi2423 & ~n30709;
  assign po2737 = n49920 | n49921;
  assign n49923 = n30709 & n47691;
  assign n49924 = pi2424 & ~n30709;
  assign po2738 = n49923 | n49924;
  assign n49926 = n30709 & n47700;
  assign n49927 = pi2425 & ~n30709;
  assign po2739 = n49926 | n49927;
  assign n49929 = n30709 & n47709;
  assign n49930 = pi2426 & ~n30709;
  assign po2740 = n49929 | n49930;
  assign n49932 = n30709 & n47718;
  assign n49933 = pi2427 & ~n30709;
  assign po2741 = n49932 | n49933;
  assign n49935 = n30709 & n47727;
  assign n49936 = pi2428 & ~n30709;
  assign po2742 = n49935 | n49936;
  assign n49938 = n30709 & n47736;
  assign n49939 = pi2429 & ~n30709;
  assign po2743 = n49938 | n49939;
  assign n49941 = n30709 & n47745;
  assign n49942 = pi2430 & ~n30709;
  assign po2744 = n49941 | n49942;
  assign n49944 = n30709 & n47763;
  assign n49945 = pi2431 & ~n30709;
  assign po2745 = n49944 | n49945;
  assign n49947 = ~n37850 & n49096;
  assign n49948 = pi2432 & ~n49096;
  assign po2746 = n49947 | n49948;
  assign n49950 = ~n37901 & n49096;
  assign n49951 = pi2433 & ~n49096;
  assign po2747 = n49950 | n49951;
  assign n49953 = ~n37918 & n49096;
  assign n49954 = pi2434 & ~n49096;
  assign po2748 = n49953 | n49954;
  assign n49956 = ~n37935 & n49096;
  assign n49957 = pi2435 & ~n49096;
  assign po2749 = n49956 | n49957;
  assign n49959 = ~n37613 & n49096;
  assign n49960 = pi2436 & ~n49096;
  assign po2750 = n49959 | n49960;
  assign n49962 = ~n37952 & n49096;
  assign n49963 = pi2437 & ~n49096;
  assign po2751 = n49962 | n49963;
  assign n49965 = ~n39032 & n49112;
  assign n49966 = pi2438 & ~n49112;
  assign po2752 = n49965 | n49966;
  assign n49968 = ~n39047 & n49112;
  assign n49969 = pi2439 & ~n49112;
  assign po2753 = n49968 | n49969;
  assign n49971 = ~n39062 & n49112;
  assign n49972 = pi2440 & ~n49112;
  assign po2754 = n49971 | n49972;
  assign n49974 = ~n39077 & n49112;
  assign n49975 = pi2441 & ~n49112;
  assign po2755 = n49974 | n49975;
  assign n49977 = ~n37850 & n49146;
  assign n49978 = pi2442 & ~n49146;
  assign po2756 = n49977 | n49978;
  assign n49980 = ~n37884 & n49146;
  assign n49981 = pi2443 & ~n49146;
  assign po2757 = n49980 | n49981;
  assign n49983 = ~n37918 & n49146;
  assign n49984 = pi2444 & ~n49146;
  assign po2758 = n49983 | n49984;
  assign n49986 = ~n37935 & n49146;
  assign n49987 = pi2445 & ~n49146;
  assign po2759 = n49986 | n49987;
  assign n49989 = ~n37613 & n49146;
  assign n49990 = pi2446 & ~n49146;
  assign po2760 = n49989 | n49990;
  assign n49992 = ~n37952 & n49146;
  assign n49993 = pi2447 & ~n49146;
  assign po2761 = n49992 | n49993;
  assign n49995 = pi2794 & pi3245;
  assign n49996 = pi1028 & ~pi3245;
  assign n49997 = ~n49995 & ~n49996;
  assign n49998 = n49888 & ~n49997;
  assign n49999 = pi2448 & ~n49888;
  assign po2762 = n49998 | n49999;
  assign n50001 = pi2644 & pi3245;
  assign n50002 = pi1030 & ~pi3245;
  assign n50003 = ~n50001 & ~n50002;
  assign n50004 = n49888 & ~n50003;
  assign n50005 = pi2449 & ~n49888;
  assign po2763 = n50004 | n50005;
  assign n50007 = pi2797 & pi3245;
  assign n50008 = pi1031 & ~pi3245;
  assign n50009 = ~n50007 & ~n50008;
  assign n50010 = n49888 & ~n50009;
  assign n50011 = pi2450 & ~n49888;
  assign po2764 = n50010 | n50011;
  assign n50013 = pi2645 & pi3245;
  assign n50014 = pi1013 & ~pi3245;
  assign n50015 = ~n50013 & ~n50014;
  assign n50016 = n49888 & ~n50015;
  assign n50017 = pi2451 & ~n49888;
  assign po2765 = n50016 | n50017;
  assign n50019 = pi0997 & ~pi3426;
  assign n50020 = ~n10847 & ~n50019;
  assign n50021 = ~n10846 & n50020;
  assign n50022 = ~n10850 & ~n50021;
  assign n50023 = ~n38413 & n50022;
  assign n50024 = pi2452 & ~n50022;
  assign po2766 = n50023 | n50024;
  assign n50026 = ~n38428 & n50022;
  assign n50027 = pi2453 & ~n50022;
  assign po2767 = n50026 | n50027;
  assign n50029 = ~n38443 & n50022;
  assign n50030 = pi2454 & ~n50022;
  assign po2768 = n50029 | n50030;
  assign n50032 = ~n38458 & n50022;
  assign n50033 = pi2455 & ~n50022;
  assign po2769 = n50032 | n50033;
  assign n50035 = ~n38473 & n50022;
  assign n50036 = pi2456 & ~n50022;
  assign po2770 = n50035 | n50036;
  assign n50038 = n38139 & n50022;
  assign n50039 = pi2457 & ~n50022;
  assign po2771 = n50038 | n50039;
  assign n50041 = n38156 & n50022;
  assign n50042 = pi2458 & ~n50022;
  assign po2772 = n50041 | n50042;
  assign n50044 = n38190 & n50022;
  assign n50045 = pi2459 & ~n50022;
  assign po2773 = n50044 | n50045;
  assign n50047 = n38207 & n50022;
  assign n50048 = pi2460 & ~n50022;
  assign po2774 = n50047 | n50048;
  assign n50050 = ~n38428 & n49869;
  assign n50051 = pi2461 & ~n49869;
  assign po2775 = n50050 | n50051;
  assign n50053 = ~n38443 & n49869;
  assign n50054 = pi2462 & ~n49869;
  assign po2776 = n50053 | n50054;
  assign n50056 = n38122 & n49869;
  assign n50057 = pi2463 & ~n49869;
  assign po2777 = n50056 | n50057;
  assign n50059 = ~n38458 & n49869;
  assign n50060 = pi2464 & ~n49869;
  assign po2778 = n50059 | n50060;
  assign n50062 = ~n38473 & n49869;
  assign n50063 = pi2465 & ~n49869;
  assign po2779 = n50062 | n50063;
  assign n50065 = n38139 & n49869;
  assign n50066 = pi2466 & ~n49869;
  assign po2780 = n50065 | n50066;
  assign n50068 = n38173 & n49869;
  assign n50069 = pi2467 & ~n49869;
  assign po2781 = n50068 | n50069;
  assign n50071 = n38190 & n49869;
  assign n50072 = pi2468 & ~n49869;
  assign po2782 = n50071 | n50072;
  assign n50074 = n38207 & n49869;
  assign n50075 = pi2469 & ~n49869;
  assign po2783 = n50074 | n50075;
  assign n50077 = ~n38503 & n49869;
  assign n50078 = pi2470 & ~n49869;
  assign po2784 = n50077 | n50078;
  assign n50080 = ~pi2471 & ~n46586;
  assign n50081 = pi2408 & n47970;
  assign n50082 = ~pi2471 & ~n47970;
  assign n50083 = ~n50081 & ~n50082;
  assign n50084 = n46586 & ~n50083;
  assign po2785 = n50080 | n50084;
  assign n50086 = ~n14816 & n49803;
  assign n50087 = pi2472 & ~n49803;
  assign po2786 = n50086 | n50087;
  assign n50089 = ~n13398 & n49841;
  assign n50090 = pi2473 & ~n49841;
  assign po2787 = n50089 | n50090;
  assign n50092 = n38250 & n48086;
  assign n50093 = pi2474 & ~n38262;
  assign po2788 = n50092 | n50093;
  assign n50095 = pi2475 & n33813;
  assign n50096 = pi3432 & ~n33813;
  assign po2789 = n50095 | n50096;
  assign n50098 = pi2476 & n33813;
  assign n50099 = pi3453 & ~n33813;
  assign po2790 = n50098 | n50099;
  assign n50101 = pi2477 & n33813;
  assign n50102 = pi3454 & ~n33813;
  assign po2791 = n50101 | n50102;
  assign n50104 = pi2478 & n33813;
  assign n50105 = pi3455 & ~n33813;
  assign po2792 = n50104 | n50105;
  assign n50107 = pi2479 & n33813;
  assign n50108 = pi3434 & ~n33813;
  assign po2793 = n50107 | n50108;
  assign n50110 = pi2480 & n33813;
  assign n50111 = pi3456 & ~n33813;
  assign po2794 = n50110 | n50111;
  assign n50113 = pi2481 & n33813;
  assign n50114 = pi3457 & ~n33813;
  assign po2795 = n50113 | n50114;
  assign n50116 = pi2482 & n33813;
  assign n50117 = pi3433 & ~n33813;
  assign po2796 = n50116 | n50117;
  assign n50119 = pi2483 & n33813;
  assign n50120 = pi3437 & ~n33813;
  assign po2797 = n50119 | n50120;
  assign n50122 = pi2484 & n33813;
  assign n50123 = pi3458 & ~n33813;
  assign po2798 = n50122 | n50123;
  assign n50125 = pi2485 & n33813;
  assign n50126 = pi3450 & ~n33813;
  assign po2799 = n50125 | n50126;
  assign n50128 = ~n8561 & ~n48102;
  assign n50129 = pi2486 & n8561;
  assign n50130 = ~n50128 & ~n50129;
  assign po2800 = po3627 & n50130;
  assign n50132 = ~pi2487 & n8561;
  assign n50133 = ~n49694 & ~n50132;
  assign po2801 = po3627 & ~n50133;
  assign n50135 = n10805 & ~n35655;
  assign n50136 = n36059 & ~n50135;
  assign n50137 = pi2488 & n36128;
  assign po2802 = n50136 | n50137;
  assign n50139 = ~n9377 & ~n47131;
  assign n50140 = n49693 & ~n50139;
  assign n50141 = pi2489 & n8561;
  assign n50142 = ~n50140 & ~n50141;
  assign n50143 = n9345 & n15589;
  assign n50144 = ~n8561 & n50143;
  assign n50145 = n50142 & ~n50144;
  assign po2803 = po3627 & ~n50145;
  assign n50147 = pi2490 & n8561;
  assign n50148 = ~n50140 & ~n50147;
  assign n50149 = ~pi0408 & n15589;
  assign n50150 = n9345 & n50149;
  assign n50151 = ~n8561 & n50150;
  assign n50152 = n50148 & ~n50151;
  assign po2804 = po3627 & ~n50152;
  assign n50154 = pi0420 & n47131;
  assign n50155 = pi0408 & n9377;
  assign n50156 = ~n50154 & ~n50155;
  assign n50157 = n49693 & ~n50156;
  assign n50158 = ~pi2491 & n8561;
  assign n50159 = ~n50157 & ~n50158;
  assign po2805 = po3627 & ~n50159;
  assign n50161 = ~pi3417 & po3745;
  assign n50162 = po0493 & ~n50161;
  assign n50163 = ~pi3337 & ~pi3389;
  assign po3743 = pi3568 & n50163;
  assign po2806 = n50162 & po3743;
  assign n50166 = pi3398 & po3850;
  assign n50167 = ~pi3481 & n50166;
  assign n50168 = pi2492 & pi3481;
  assign po2807 = n50167 | n50168;
  assign n50170 = n11157 & n38277;
  assign n50171 = pi2493 & ~n50170;
  assign n50172 = ~n12726 & n50170;
  assign po2808 = n50171 | n50172;
  assign n50174 = pi2494 & ~n50170;
  assign n50175 = ~n13701 & n50170;
  assign po2809 = n50174 | n50175;
  assign n50177 = pi2495 & ~n50170;
  assign n50178 = ~n13121 & n50170;
  assign po2810 = n50177 | n50178;
  assign n50180 = pi2496 & ~n50170;
  assign n50181 = ~n13398 & n50170;
  assign po2811 = n50180 | n50181;
  assign n50183 = pi2497 & ~n50170;
  assign n50184 = ~n13988 & n50170;
  assign po2812 = n50183 | n50184;
  assign n50186 = pi2498 & ~n50170;
  assign n50187 = ~n14816 & n50170;
  assign po2813 = n50186 | n50187;
  assign n50189 = pi2499 & ~n50170;
  assign n50190 = ~n12061 & n50170;
  assign po2814 = n50189 | n50190;
  assign n50192 = pi2500 & ~n50170;
  assign n50193 = ~n15426 & n50170;
  assign po2815 = n50192 | n50193;
  assign n50195 = pi2501 & ~n50170;
  assign n50196 = ~n14403 & n50170;
  assign po2816 = n50195 | n50196;
  assign n50198 = pi2502 & ~n50170;
  assign n50199 = ~n11181 & n50170;
  assign po2817 = n50198 | n50199;
  assign n50201 = n9646 & n38277;
  assign n50202 = pi2503 & ~n50201;
  assign n50203 = ~n13121 & n50201;
  assign n50204 = ~n50202 & ~n50203;
  assign n50205 = n13121 & n13988;
  assign n50206 = n13398 & n50205;
  assign n50207 = n50201 & n50206;
  assign n50208 = n12415 & n50207;
  assign po2818 = ~n50204 | n50208;
  assign n50210 = pi2504 & ~n50201;
  assign n50211 = ~n13398 & n50201;
  assign n50212 = ~n50210 & ~n50211;
  assign po2819 = n50208 | ~n50212;
  assign n50214 = pi2505 & ~n50201;
  assign n50215 = ~n12415 & n50201;
  assign n50216 = ~n50214 & ~n50215;
  assign po2820 = n50208 | ~n50216;
  assign n50218 = ~pi2523 & ~pi2771;
  assign n50219 = ~pi2506 & n50218;
  assign n50220 = pi2506 & ~n50218;
  assign n50221 = ~n50219 & ~n50220;
  assign po2821 = ~n49739 & n50221;
  assign n50223 = ~pi2506 & ~pi2760;
  assign n50224 = n50218 & n50223;
  assign n50225 = ~pi2772 & n50224;
  assign n50226 = ~pi2507 & n50225;
  assign n50227 = pi2507 & ~n50225;
  assign n50228 = ~n50226 & ~n50227;
  assign po2822 = ~n49739 & n50228;
  assign n50230 = ~pi2510 & ~n42536;
  assign n50231 = pi2510 & n41247;
  assign n50232 = ~pi2510 & ~n41247;
  assign n50233 = ~n50231 & ~n50232;
  assign n50234 = n42536 & ~n50233;
  assign po2825 = n50230 | n50234;
  assign n50236 = n30709 & n47754;
  assign n50237 = pi2511 & ~n30709;
  assign po2826 = n50236 | n50237;
  assign n50239 = pi2512 & ~n50170;
  assign n50240 = ~n15115 & n50170;
  assign po2827 = n50239 | n50240;
  assign n50242 = pi2513 & ~n50170;
  assign n50243 = ~n12415 & n50170;
  assign po2828 = n50242 | n50243;
  assign n50245 = ~n15115 & n49803;
  assign n50246 = pi2514 & ~n49803;
  assign po2829 = n50245 | n50246;
  assign n50248 = pi2515 & n32787;
  assign po2830 = n46808 | n50248;
  assign n50250 = pi2516 & n33813;
  assign n50251 = pi3460 & ~n33813;
  assign po2831 = n50250 | n50251;
  assign n50253 = pi2517 & n33813;
  assign n50254 = pi3459 & ~n33813;
  assign po2832 = n50253 | n50254;
  assign n50256 = pi2518 & n33813;
  assign n50257 = pi3478 & ~n33813;
  assign po2833 = n50256 | n50257;
  assign n50259 = ~pi2519 & ~n46586;
  assign n50260 = pi2408 & n47897;
  assign n50261 = ~pi2519 & ~n47897;
  assign n50262 = ~n50260 & ~n50261;
  assign n50263 = n46586 & ~n50262;
  assign po2834 = n50259 | n50263;
  assign n50265 = n38095 & n50022;
  assign n50266 = pi2520 & ~n50022;
  assign po2835 = n50265 | n50266;
  assign n50268 = pi2522 & ~n50201;
  assign n50269 = ~n13988 & n50201;
  assign n50270 = ~n50268 & ~n50269;
  assign po2837 = n50208 | ~n50270;
  assign po2838 = pi2523 & ~n49739;
  assign n50273 = ~n38503 & n50022;
  assign n50274 = pi2524 & ~n50022;
  assign po2839 = n50273 | n50274;
  assign n50276 = n38173 & n50022;
  assign n50277 = pi2525 & ~n50022;
  assign po2840 = n50276 | n50277;
  assign n50279 = ~n38488 & n50022;
  assign n50280 = pi2526 & ~n50022;
  assign po2841 = n50279 | n50280;
  assign n50282 = n38122 & n50022;
  assign n50283 = pi2527 & ~n50022;
  assign po2842 = n50282 | n50283;
  assign n50285 = ~pi0990 & n37646;
  assign n50286 = ~pi3426 & n50285;
  assign n50287 = ~n13398 & n50286;
  assign n50288 = pi2528 & ~n50286;
  assign po2843 = n50287 | n50288;
  assign n50290 = ~n8612 & n35527;
  assign n50291 = ~n8561 & ~n50290;
  assign n50292 = n36451 & n50291;
  assign n50293 = pi2529 & ~n50291;
  assign po2844 = n50292 | n50293;
  assign n50295 = pi0998 & ~pi3426;
  assign n50296 = ~n10839 & ~n50295;
  assign n50297 = ~n10842 & n50296;
  assign n50298 = ~n10843 & ~n50297;
  assign n50299 = pi2530 & ~n50298;
  assign n50300 = n38156 & n50298;
  assign po2845 = n50299 | n50300;
  assign n50302 = ~n13121 & n50286;
  assign n50303 = pi2531 & ~n50286;
  assign po2846 = n50302 | n50303;
  assign n50305 = ~pi1051 & n37651;
  assign n50306 = ~pi3426 & n50305;
  assign n50307 = ~n11181 & n50306;
  assign n50308 = pi2532 & ~n50306;
  assign po2847 = n50307 | n50308;
  assign n50310 = pi0996 & ~pi3426;
  assign n50311 = ~n10822 & ~n50310;
  assign n50312 = ~n10818 & n50311;
  assign n50313 = ~n10825 & ~n50312;
  assign n50314 = pi2533 & ~n50313;
  assign n50315 = n38173 & n50313;
  assign po2848 = n50314 | n50315;
  assign n50317 = ~n15426 & n50306;
  assign n50318 = pi2534 & ~n50306;
  assign po2849 = n50317 | n50318;
  assign n50320 = pi2535 & ~n50313;
  assign n50321 = n38095 & n50313;
  assign po2850 = n50320 | n50321;
  assign n50323 = ~n13988 & n50306;
  assign n50324 = pi2536 & ~n50306;
  assign po2851 = n50323 | n50324;
  assign n50326 = n24309 & n25551;
  assign n50327 = ~n24488 & n50326;
  assign n50328 = pi2537 & ~n50326;
  assign po2852 = n50327 | n50328;
  assign n50330 = ~n27570 & n50326;
  assign n50331 = pi2538 & ~n50326;
  assign po2853 = n50330 | n50331;
  assign n50333 = pi2539 & ~n49096;
  assign n50334 = ~n39062 & n49096;
  assign po2854 = n50333 | n50334;
  assign n50336 = pi2540 & ~n50291;
  assign n50337 = n48074 & n50291;
  assign po2855 = n50336 | n50337;
  assign n50339 = ~n24256 & n50326;
  assign n50340 = pi2541 & ~n50326;
  assign po2856 = n50339 | n50340;
  assign n50342 = ~pi0991 & n37641;
  assign n50343 = ~pi3426 & n50342;
  assign n50344 = ~n11181 & n50343;
  assign n50345 = pi2542 & ~n50343;
  assign po2857 = n50344 | n50345;
  assign n50347 = ~n10608 & n50343;
  assign n50348 = pi2543 & ~n50343;
  assign po2858 = n50347 | n50348;
  assign n50350 = pi2544 & ~n50298;
  assign n50351 = n38190 & n50298;
  assign po2859 = n50350 | n50351;
  assign n50353 = ~n15426 & n50343;
  assign n50354 = pi2545 & ~n50343;
  assign po2860 = n50353 | n50354;
  assign n50356 = ~n12415 & n50343;
  assign n50357 = pi2546 & ~n50343;
  assign po2861 = n50356 | n50357;
  assign n50359 = ~n15115 & n50343;
  assign n50360 = pi2547 & ~n50343;
  assign po2862 = n50359 | n50360;
  assign n50362 = ~n13121 & n50343;
  assign n50363 = pi2548 & ~n50343;
  assign po2863 = n50362 | n50363;
  assign n50365 = pi2549 & ~n50291;
  assign n50366 = n48060 & n50291;
  assign po2864 = n50365 | n50366;
  assign n50368 = ~pi0987 & n37277;
  assign n50369 = ~pi3426 & n50368;
  assign n50370 = ~n12726 & n50369;
  assign n50371 = pi2550 & ~n50369;
  assign po2865 = n50370 | n50371;
  assign n50373 = pi2551 & ~n50291;
  assign n50374 = n48032 & n50291;
  assign po2866 = n50373 | n50374;
  assign n50376 = ~pi0920 & n37628;
  assign n50377 = ~pi3426 & n50376;
  assign n50378 = ~n11181 & n50377;
  assign n50379 = pi2552 & ~n50377;
  assign po2867 = n50378 | n50379;
  assign n50381 = pi2553 & ~n50291;
  assign n50382 = n48018 & n50291;
  assign po2868 = n50381 | n50382;
  assign n50384 = pi2554 & ~n49888;
  assign n50385 = pi2540 & pi3245;
  assign n50386 = pi1039 & ~pi3245;
  assign n50387 = ~n50385 & ~n50386;
  assign n50388 = n49888 & ~n50387;
  assign po2869 = n50384 | n50388;
  assign po2870 = pi0955 & ~pi3250;
  assign n50391 = pi2556 & ~n49888;
  assign n50392 = pi2551 & pi3245;
  assign n50393 = pi1033 & ~pi3245;
  assign n50394 = ~n50392 & ~n50393;
  assign n50395 = n49888 & ~n50394;
  assign po2871 = n50391 | n50395;
  assign n50397 = ~pi2529 & pi3245;
  assign n50398 = ~pi1036 & ~pi3245;
  assign n50399 = ~n50397 & ~n50398;
  assign n50400 = n49888 & n50399;
  assign n50401 = pi2557 & ~n49888;
  assign po2872 = n50400 | n50401;
  assign n50403 = ~pi2647 & pi3245;
  assign n50404 = ~pi1035 & ~pi3245;
  assign n50405 = ~n50403 & ~n50404;
  assign n50406 = n49888 & n50405;
  assign n50407 = pi2558 & ~n49888;
  assign po2873 = n50406 | n50407;
  assign n50409 = pi2559 & ~n49888;
  assign n50410 = pi2549 & pi3245;
  assign n50411 = pi1012 & ~pi3245;
  assign n50412 = ~n50410 & ~n50411;
  assign n50413 = n49888 & ~n50412;
  assign po2874 = n50409 | n50413;
  assign n50415 = ~n15115 & n50377;
  assign n50416 = pi2560 & ~n50377;
  assign po2875 = n50415 | n50416;
  assign n50418 = ~n9825 & n50377;
  assign n50419 = pi2561 & ~n50377;
  assign po2876 = n50418 | n50419;
  assign n50421 = ~pi1010 & n37267;
  assign n50422 = ~pi3426 & n50421;
  assign n50423 = ~n11181 & n50422;
  assign n50424 = pi2562 & ~n50422;
  assign po2877 = n50423 | n50424;
  assign n50426 = ~n13398 & n50422;
  assign n50427 = pi2563 & ~n50422;
  assign po2878 = n50426 | n50427;
  assign n50429 = ~n15426 & n50286;
  assign n50430 = pi2565 & ~n50286;
  assign po2880 = n50429 | n50430;
  assign n50432 = ~n13701 & n50377;
  assign n50433 = pi2566 & ~n50377;
  assign po2881 = n50432 | n50433;
  assign n50435 = ~pi0758 & n9365;
  assign n50436 = ~pi3424 & ~n50435;
  assign n50437 = ~n13701 & ~n50436;
  assign n50438 = pi2568 & n50436;
  assign po2883 = n50437 | n50438;
  assign n50440 = ~n13121 & ~n50436;
  assign n50441 = pi2569 & n50436;
  assign po2884 = n50440 | n50441;
  assign n50443 = ~n13398 & ~n50436;
  assign n50444 = pi2570 & n50436;
  assign po2885 = n50443 | n50444;
  assign n50446 = ~n13988 & ~n50436;
  assign n50447 = pi2571 & n50436;
  assign po2886 = n50446 | n50447;
  assign n50449 = ~n12415 & ~n50436;
  assign n50450 = pi2572 & n50436;
  assign po2887 = n50449 | n50450;
  assign n50452 = ~n14816 & ~n50436;
  assign n50453 = pi2573 & n50436;
  assign po2888 = n50452 | n50453;
  assign n50455 = ~n15115 & ~n50436;
  assign n50456 = pi2574 & n50436;
  assign po2889 = n50455 | n50456;
  assign n50458 = ~n12061 & ~n50436;
  assign n50459 = pi2575 & n50436;
  assign po2890 = n50458 | n50459;
  assign n50461 = ~n17368 & ~n50436;
  assign n50462 = pi2576 & n50436;
  assign po2891 = n50461 | n50462;
  assign n50464 = ~n17199 & ~n50436;
  assign n50465 = pi2577 & n50436;
  assign po2892 = n50464 | n50465;
  assign n50467 = ~n9825 & ~n50436;
  assign n50468 = pi2578 & n50436;
  assign po2893 = n50467 | n50468;
  assign n50470 = ~n10608 & ~n50436;
  assign n50471 = pi2579 & n50436;
  assign po2894 = n50470 | n50471;
  assign n50473 = ~n15426 & ~n50436;
  assign n50474 = pi2580 & n50436;
  assign po2895 = n50473 | n50474;
  assign n50476 = ~n14403 & ~n50436;
  assign n50477 = pi2581 & n50436;
  assign po2896 = n50476 | n50477;
  assign n50479 = ~n11181 & ~n50436;
  assign n50480 = pi2582 & n50436;
  assign po2897 = n50479 | n50480;
  assign n50482 = ~pi0581 & pi3535;
  assign n50483 = pi0478 & n50482;
  assign n50484 = n12726 & ~n50482;
  assign n50485 = ~n50483 & ~n50484;
  assign n50486 = ~pi0982 & n9365;
  assign n50487 = ~n50482 & ~n50486;
  assign n50488 = n50485 & ~n50487;
  assign n50489 = pi2583 & n50487;
  assign po2898 = n50488 | n50489;
  assign n50491 = pi0477 & n50482;
  assign n50492 = n13701 & ~n50482;
  assign n50493 = ~n50491 & ~n50492;
  assign n50494 = ~n50487 & n50493;
  assign n50495 = pi2584 & n50487;
  assign po2899 = n50494 | n50495;
  assign n50497 = pi0476 & n50482;
  assign n50498 = n13121 & ~n50482;
  assign n50499 = ~n50497 & ~n50498;
  assign n50500 = ~n50487 & n50499;
  assign n50501 = pi2585 & n50487;
  assign po2900 = n50500 | n50501;
  assign n50503 = pi0475 & n50482;
  assign n50504 = n13398 & ~n50482;
  assign n50505 = ~n50503 & ~n50504;
  assign n50506 = ~n50487 & n50505;
  assign n50507 = pi2586 & n50487;
  assign po2901 = n50506 | n50507;
  assign n50509 = pi0474 & n50482;
  assign n50510 = n12415 & ~n50482;
  assign n50511 = ~n50509 & ~n50510;
  assign n50512 = ~n50487 & n50511;
  assign n50513 = pi2587 & n50487;
  assign po2902 = n50512 | n50513;
  assign n50515 = pi0473 & n50482;
  assign n50516 = n14816 & ~n50482;
  assign n50517 = ~n50515 & ~n50516;
  assign n50518 = ~n50487 & n50517;
  assign n50519 = pi2588 & n50487;
  assign po2903 = n50518 | n50519;
  assign n50521 = pi0472 & n50482;
  assign n50522 = n15115 & ~n50482;
  assign n50523 = ~n50521 & ~n50522;
  assign n50524 = ~n50487 & n50523;
  assign n50525 = pi2589 & n50487;
  assign po2904 = n50524 | n50525;
  assign n50527 = pi0697 & n50482;
  assign n50528 = n12061 & ~n50482;
  assign n50529 = ~n50527 & ~n50528;
  assign n50530 = ~n50487 & n50529;
  assign n50531 = pi2590 & n50487;
  assign po2905 = n50530 | n50531;
  assign n50533 = pi0471 & n50482;
  assign n50534 = n17368 & ~n50482;
  assign n50535 = ~n50533 & ~n50534;
  assign n50536 = ~n50487 & n50535;
  assign n50537 = pi2591 & n50487;
  assign po2906 = n50536 | n50537;
  assign n50539 = pi0470 & n50482;
  assign n50540 = n17199 & ~n50482;
  assign n50541 = ~n50539 & ~n50540;
  assign n50542 = ~n50487 & n50541;
  assign n50543 = pi2592 & n50487;
  assign po2907 = n50542 | n50543;
  assign n50545 = pi0469 & n50482;
  assign n50546 = n9825 & ~n50482;
  assign n50547 = ~n50545 & ~n50546;
  assign n50548 = ~n50487 & n50547;
  assign n50549 = pi2593 & n50487;
  assign po2908 = n50548 | n50549;
  assign n50551 = pi0468 & n50482;
  assign n50552 = n10608 & ~n50482;
  assign n50553 = ~n50551 & ~n50552;
  assign n50554 = ~n50487 & n50553;
  assign n50555 = pi2594 & n50487;
  assign po2909 = n50554 | n50555;
  assign n50557 = pi0467 & n50482;
  assign n50558 = n15426 & ~n50482;
  assign n50559 = ~n50557 & ~n50558;
  assign n50560 = ~n50487 & n50559;
  assign n50561 = pi2595 & n50487;
  assign po2910 = n50560 | n50561;
  assign n50563 = pi0466 & n50482;
  assign n50564 = n14403 & ~n50482;
  assign n50565 = ~n50563 & ~n50564;
  assign n50566 = ~n50487 & n50565;
  assign n50567 = pi2596 & n50487;
  assign po2911 = n50566 | n50567;
  assign n50569 = pi0696 & n50482;
  assign n50570 = n11181 & ~n50482;
  assign n50571 = ~n50569 & ~n50570;
  assign n50572 = ~n50487 & n50571;
  assign n50573 = pi2597 & n50487;
  assign po2912 = n50572 | n50573;
  assign po2913 = ~pi3429 & ~pi3639;
  assign n50576 = pi1738 & pi3647;
  assign n50577 = ~n50487 & n50576;
  assign po2914 = pi2598 | n50577;
  assign n50579 = pi2600 & n48383;
  assign n50580 = ~pi2600 & n48385;
  assign n50581 = pi2799 & n50580;
  assign n50582 = pi2600 & ~n48386;
  assign n50583 = ~n50581 & ~n50582;
  assign n50584 = ~n48383 & ~n50583;
  assign n50585 = ~n50579 & ~n50584;
  assign po2916 = n48409 & ~n50585;
  assign po2917 = pi3428 & ~pi3556;
  assign n50588 = ~pi1422 & ~n39524;
  assign n50589 = n46808 & ~n50588;
  assign n50590 = n10782 & n39526;
  assign n50591 = ~n50589 & ~n50590;
  assign n50592 = n8601 & n39526;
  assign n50593 = pi0975 & n50592;
  assign n50594 = ~pi2601 & ~n50593;
  assign po2918 = ~n50591 | ~n50594;
  assign n50596 = ~n12726 & n50422;
  assign n50597 = pi2602 & ~n50422;
  assign po2919 = n50596 | n50597;
  assign n50599 = ~pi0989 & n37252;
  assign n50600 = ~pi3426 & n50599;
  assign n50601 = ~n11181 & n50600;
  assign n50602 = pi2603 & ~n50600;
  assign po2920 = n50601 | n50602;
  assign po2921 = po0767 & ~n50161;
  assign n50605 = pi2492 & pi3441;
  assign n50606 = ~pi2604 & n50605;
  assign po2922 = pi2604 | n50606;
  assign n50608 = n24251 & n25522;
  assign n50609 = ~n47652 & n50608;
  assign n50610 = pi2605 & ~n50608;
  assign po2923 = n50609 | n50610;
  assign n50612 = ~n47661 & n50608;
  assign n50613 = pi2606 & ~n50608;
  assign po2924 = n50612 | n50613;
  assign n50615 = ~n47733 & n50608;
  assign n50616 = pi2607 & ~n50608;
  assign po2925 = n50615 | n50616;
  assign n50618 = ~n47742 & n50608;
  assign n50619 = pi2608 & ~n50608;
  assign po2926 = n50618 | n50619;
  assign n50621 = ~n47751 & n50608;
  assign n50622 = pi2609 & ~n50608;
  assign po2927 = n50621 | n50622;
  assign n50624 = ~n47760 & n50608;
  assign n50625 = pi2610 & ~n50608;
  assign po2928 = n50624 | n50625;
  assign n50627 = n24309 & n25522;
  assign n50628 = ~n47652 & n50627;
  assign n50629 = pi2611 & ~n50627;
  assign po2929 = n50628 | n50629;
  assign n50631 = ~n47661 & n50627;
  assign n50632 = pi2612 & ~n50627;
  assign po2930 = n50631 | n50632;
  assign n50634 = ~n47733 & n50627;
  assign n50635 = pi2613 & ~n50627;
  assign po2931 = n50634 | n50635;
  assign n50637 = ~n47742 & n50627;
  assign n50638 = pi2614 & ~n50627;
  assign po2932 = n50637 | n50638;
  assign n50640 = ~n15426 & n50600;
  assign n50641 = pi2615 & ~n50600;
  assign po2933 = n50640 | n50641;
  assign n50643 = ~n47751 & n50627;
  assign n50644 = pi2616 & ~n50627;
  assign po2934 = n50643 | n50644;
  assign n50646 = ~n47760 & n50627;
  assign n50647 = pi2617 & ~n50627;
  assign po2935 = n50646 | n50647;
  assign n50649 = n24251 & n25520;
  assign n50650 = ~n47652 & n50649;
  assign n50651 = pi2618 & ~n50649;
  assign po2936 = n50650 | n50651;
  assign n50653 = ~n47661 & n50649;
  assign n50654 = pi2619 & ~n50649;
  assign po2937 = n50653 | n50654;
  assign n50656 = ~n47733 & n50649;
  assign n50657 = pi2620 & ~n50649;
  assign po2938 = n50656 | n50657;
  assign n50659 = ~n47742 & n50649;
  assign n50660 = pi2621 & ~n50649;
  assign po2939 = n50659 | n50660;
  assign n50662 = ~n47751 & n50649;
  assign n50663 = pi2622 & ~n50649;
  assign po2940 = n50662 | n50663;
  assign n50665 = ~n47760 & n50649;
  assign n50666 = pi2623 & ~n50649;
  assign po2941 = n50665 | n50666;
  assign n50668 = n24309 & n25520;
  assign n50669 = ~n47652 & n50668;
  assign n50670 = pi2624 & ~n50668;
  assign po2942 = n50669 | n50670;
  assign n50672 = ~n47661 & n50668;
  assign n50673 = pi2625 & ~n50668;
  assign po2943 = n50672 | n50673;
  assign n50675 = ~n47733 & n50668;
  assign n50676 = pi2626 & ~n50668;
  assign po2944 = n50675 | n50676;
  assign n50678 = ~n47742 & n50668;
  assign n50679 = pi2627 & ~n50668;
  assign po2945 = n50678 | n50679;
  assign n50681 = ~n47751 & n50668;
  assign n50682 = pi2628 & ~n50668;
  assign po2946 = n50681 | n50682;
  assign n50684 = ~n47760 & n50668;
  assign n50685 = pi2629 & ~n50668;
  assign po2947 = n50684 | n50685;
  assign n50687 = ~n30267 & n50326;
  assign n50688 = pi2630 & ~n50326;
  assign po2948 = n50687 | n50688;
  assign n50690 = ~n30288 & n50326;
  assign n50691 = pi2631 & ~n50326;
  assign po2949 = n50690 | n50691;
  assign n50693 = ~n24744 & n50326;
  assign n50694 = pi2632 & ~n50326;
  assign po2950 = n50693 | n50694;
  assign n50696 = ~n24769 & n50326;
  assign n50697 = pi2633 & ~n50326;
  assign po2951 = n50696 | n50697;
  assign n50699 = ~n25699 & n50326;
  assign n50700 = pi2634 & ~n50326;
  assign po2952 = n50699 | n50700;
  assign n50702 = ~n25718 & n50326;
  assign n50703 = pi2635 & ~n50326;
  assign po2953 = n50702 | n50703;
  assign n50705 = ~n24289 & n50326;
  assign n50706 = pi2636 & ~n50326;
  assign po2954 = n50705 | n50706;
  assign n50708 = ~n24446 & n50326;
  assign n50709 = pi2637 & ~n50326;
  assign po2955 = n50708 | n50709;
  assign n50711 = ~n24265 & n50326;
  assign n50712 = pi2638 & ~n50326;
  assign po2956 = n50711 | n50712;
  assign n50714 = ~n30309 & n50326;
  assign n50715 = pi2639 & ~n50326;
  assign po2957 = n50714 | n50715;
  assign n50717 = ~n30321 & n50326;
  assign n50718 = pi2640 & ~n50326;
  assign po2958 = n50717 | n50718;
  assign n50720 = ~n30333 & n50326;
  assign n50721 = pi2641 & ~n50326;
  assign po2959 = n50720 | n50721;
  assign n50723 = ~n25999 & n50326;
  assign n50724 = pi2642 & ~n50326;
  assign po2960 = n50723 | n50724;
  assign n50726 = n38764 & po3574;
  assign n50727 = ~pi2643 & ~n50726;
  assign n50728 = pi0731 & n50726;
  assign po2961 = n50727 | n50728;
  assign n50730 = pi2644 & ~n50291;
  assign n50731 = n47990 & n50291;
  assign po2962 = n50730 | n50731;
  assign n50733 = pi2645 & ~n50291;
  assign n50734 = n48004 & n50291;
  assign po2963 = n50733 | n50734;
  assign n50736 = pi2646 & ~n50291;
  assign n50737 = n48046 & n50291;
  assign po2964 = n50736 | n50737;
  assign n50739 = n36443 & n50291;
  assign n50740 = pi2647 & ~n50291;
  assign po2965 = n50739 | n50740;
  assign n50742 = ~n13701 & n50369;
  assign n50743 = pi2648 & ~n50369;
  assign po2966 = n50742 | n50743;
  assign n50745 = ~n13121 & n50369;
  assign n50746 = pi2649 & ~n50369;
  assign po2967 = n50745 | n50746;
  assign n50748 = ~n13398 & n50369;
  assign n50749 = pi2650 & ~n50369;
  assign po2968 = n50748 | n50749;
  assign n50751 = ~n13988 & n50369;
  assign n50752 = pi2651 & ~n50369;
  assign po2969 = n50751 | n50752;
  assign n50754 = ~n12415 & n50369;
  assign n50755 = pi2652 & ~n50369;
  assign po2970 = n50754 | n50755;
  assign n50757 = ~n14816 & n50369;
  assign n50758 = pi2653 & ~n50369;
  assign po2971 = n50757 | n50758;
  assign n50760 = ~n15115 & n50369;
  assign n50761 = pi2654 & ~n50369;
  assign po2972 = n50760 | n50761;
  assign n50763 = ~n12061 & n50369;
  assign n50764 = pi2655 & ~n50369;
  assign po2973 = n50763 | n50764;
  assign n50766 = ~n9825 & n50369;
  assign n50767 = pi2656 & ~n50369;
  assign po2974 = n50766 | n50767;
  assign n50769 = ~n10608 & n50369;
  assign n50770 = pi2657 & ~n50369;
  assign po2975 = n50769 | n50770;
  assign n50772 = ~n15426 & n50369;
  assign n50773 = pi2658 & ~n50369;
  assign po2976 = n50772 | n50773;
  assign n50775 = ~n14403 & n50369;
  assign n50776 = pi2659 & ~n50369;
  assign po2977 = n50775 | n50776;
  assign n50778 = ~n11181 & n50369;
  assign n50779 = pi2660 & ~n50369;
  assign po2978 = n50778 | n50779;
  assign n50781 = ~pi0988 & n37272;
  assign n50782 = ~pi3426 & n50781;
  assign n50783 = ~n12726 & n50782;
  assign n50784 = pi2661 & ~n50782;
  assign po2979 = n50783 | n50784;
  assign n50786 = ~n13701 & n50782;
  assign n50787 = pi2662 & ~n50782;
  assign po2980 = n50786 | n50787;
  assign n50789 = ~n13121 & n50782;
  assign n50790 = pi2663 & ~n50782;
  assign po2981 = n50789 | n50790;
  assign n50792 = ~n13398 & n50782;
  assign n50793 = pi2664 & ~n50782;
  assign po2982 = n50792 | n50793;
  assign n50795 = ~n13988 & n50782;
  assign n50796 = pi2665 & ~n50782;
  assign po2983 = n50795 | n50796;
  assign n50798 = ~n12415 & n50782;
  assign n50799 = pi2666 & ~n50782;
  assign po2984 = n50798 | n50799;
  assign n50801 = ~n14816 & n50782;
  assign n50802 = pi2667 & ~n50782;
  assign po2985 = n50801 | n50802;
  assign n50804 = ~n15115 & n50782;
  assign n50805 = pi2668 & ~n50782;
  assign po2986 = n50804 | n50805;
  assign n50807 = ~n12061 & n50782;
  assign n50808 = pi2669 & ~n50782;
  assign po2987 = n50807 | n50808;
  assign n50810 = ~n9825 & n50782;
  assign n50811 = pi2670 & ~n50782;
  assign po2988 = n50810 | n50811;
  assign n50813 = ~n10608 & n50782;
  assign n50814 = pi2671 & ~n50782;
  assign po2989 = n50813 | n50814;
  assign n50816 = ~n15426 & n50782;
  assign n50817 = pi2672 & ~n50782;
  assign po2990 = n50816 | n50817;
  assign n50819 = ~n14403 & n50782;
  assign n50820 = pi2673 & ~n50782;
  assign po2991 = n50819 | n50820;
  assign n50822 = ~n11181 & n50782;
  assign n50823 = pi2674 & ~n50782;
  assign po2992 = n50822 | n50823;
  assign n50825 = ~n12726 & n50600;
  assign n50826 = pi2675 & ~n50600;
  assign po2993 = n50825 | n50826;
  assign n50828 = ~n13701 & n50600;
  assign n50829 = pi2676 & ~n50600;
  assign po2994 = n50828 | n50829;
  assign n50831 = ~n13121 & n50600;
  assign n50832 = pi2677 & ~n50600;
  assign po2995 = n50831 | n50832;
  assign n50834 = ~n13398 & n50600;
  assign n50835 = pi2678 & ~n50600;
  assign po2996 = n50834 | n50835;
  assign n50837 = ~n13988 & n50600;
  assign n50838 = pi2679 & ~n50600;
  assign po2997 = n50837 | n50838;
  assign n50840 = ~n12415 & n50600;
  assign n50841 = pi2680 & ~n50600;
  assign po2998 = n50840 | n50841;
  assign n50843 = ~n14816 & n50600;
  assign n50844 = pi2681 & ~n50600;
  assign po2999 = n50843 | n50844;
  assign n50846 = ~n15115 & n50600;
  assign n50847 = pi2682 & ~n50600;
  assign po3000 = n50846 | n50847;
  assign n50849 = ~n12061 & n50600;
  assign n50850 = pi2683 & ~n50600;
  assign po3001 = n50849 | n50850;
  assign n50852 = ~n9825 & n50600;
  assign n50853 = pi2684 & ~n50600;
  assign po3002 = n50852 | n50853;
  assign n50855 = ~n10608 & n50600;
  assign n50856 = pi2685 & ~n50600;
  assign po3003 = n50855 | n50856;
  assign n50858 = ~n14403 & n50600;
  assign n50859 = pi2686 & ~n50600;
  assign po3004 = n50858 | n50859;
  assign n50861 = ~n13701 & n50422;
  assign n50862 = pi2687 & ~n50422;
  assign po3005 = n50861 | n50862;
  assign n50864 = ~n13121 & n50422;
  assign n50865 = pi2688 & ~n50422;
  assign po3006 = n50864 | n50865;
  assign n50867 = ~n13988 & n50422;
  assign n50868 = pi2689 & ~n50422;
  assign po3007 = n50867 | n50868;
  assign n50870 = ~n12415 & n50422;
  assign n50871 = pi2690 & ~n50422;
  assign po3008 = n50870 | n50871;
  assign n50873 = ~n14816 & n50422;
  assign n50874 = pi2691 & ~n50422;
  assign po3009 = n50873 | n50874;
  assign n50876 = ~n15115 & n50422;
  assign n50877 = pi2692 & ~n50422;
  assign po3010 = n50876 | n50877;
  assign n50879 = ~n12061 & n50422;
  assign n50880 = pi2693 & ~n50422;
  assign po3011 = n50879 | n50880;
  assign n50882 = ~n9825 & n50422;
  assign n50883 = pi2694 & ~n50422;
  assign po3012 = n50882 | n50883;
  assign n50885 = ~n10608 & n50422;
  assign n50886 = pi2695 & ~n50422;
  assign po3013 = n50885 | n50886;
  assign n50888 = ~n15426 & n50422;
  assign n50889 = pi2696 & ~n50422;
  assign po3014 = n50888 | n50889;
  assign n50891 = ~n14403 & n50422;
  assign n50892 = pi2697 & ~n50422;
  assign po3015 = n50891 | n50892;
  assign n50894 = pi2698 & ~n49096;
  assign n50895 = ~n39032 & n49096;
  assign po3016 = n50894 | n50895;
  assign n50897 = pi2699 & ~n49096;
  assign n50898 = ~n39047 & n49096;
  assign po3017 = n50897 | n50898;
  assign n50900 = pi2700 & ~n49096;
  assign n50901 = ~n39077 & n49096;
  assign po3018 = n50900 | n50901;
  assign n50903 = pi2701 & ~n49146;
  assign n50904 = ~n39032 & n49146;
  assign po3019 = n50903 | n50904;
  assign n50906 = pi2702 & ~n49146;
  assign n50907 = ~n39047 & n49146;
  assign po3020 = n50906 | n50907;
  assign n50909 = pi2703 & ~n49146;
  assign n50910 = ~n39062 & n49146;
  assign po3021 = n50909 | n50910;
  assign n50912 = pi2704 & ~n49888;
  assign n50913 = pi2553 & pi3245;
  assign n50914 = pi1032 & ~pi3245;
  assign n50915 = ~n50913 & ~n50914;
  assign n50916 = n49888 & ~n50915;
  assign po3022 = n50912 | n50916;
  assign n50918 = pi2705 & ~n49888;
  assign n50919 = pi2646 & pi3245;
  assign n50920 = pi1034 & ~pi3245;
  assign n50921 = ~n50919 & ~n50920;
  assign n50922 = n49888 & ~n50921;
  assign po3023 = n50918 | n50922;
  assign n50924 = pi1037 & ~pi3245;
  assign n50925 = pi2953 & pi3245;
  assign n50926 = ~n50924 & ~n50925;
  assign n50927 = n49888 & ~n50926;
  assign n50928 = pi2706 & ~n49888;
  assign po3024 = n50927 | n50928;
  assign n50930 = pi1038 & ~pi3245;
  assign n50931 = pi2788 & pi3245;
  assign n50932 = ~n50930 & ~n50931;
  assign n50933 = n49888 & ~n50932;
  assign n50934 = pi2707 & ~n49888;
  assign po3025 = n50933 | n50934;
  assign n50936 = ~n12726 & n50306;
  assign n50937 = pi2708 & ~n50306;
  assign po3026 = n50936 | n50937;
  assign n50939 = ~n13701 & n50306;
  assign n50940 = pi2709 & ~n50306;
  assign po3027 = n50939 | n50940;
  assign n50942 = ~n13121 & n50306;
  assign n50943 = pi2710 & ~n50306;
  assign po3028 = n50942 | n50943;
  assign n50945 = ~n13398 & n50306;
  assign n50946 = pi2711 & ~n50306;
  assign po3029 = n50945 | n50946;
  assign n50948 = ~n12415 & n50306;
  assign n50949 = pi2712 & ~n50306;
  assign po3030 = n50948 | n50949;
  assign n50951 = ~n14816 & n50306;
  assign n50952 = pi2713 & ~n50306;
  assign po3031 = n50951 | n50952;
  assign n50954 = ~n15115 & n50306;
  assign n50955 = pi2714 & ~n50306;
  assign po3032 = n50954 | n50955;
  assign n50957 = ~n12061 & n50306;
  assign n50958 = pi2715 & ~n50306;
  assign po3033 = n50957 | n50958;
  assign n50960 = ~n9825 & n50306;
  assign n50961 = pi2716 & ~n50306;
  assign po3034 = n50960 | n50961;
  assign n50963 = ~n10608 & n50306;
  assign n50964 = pi2717 & ~n50306;
  assign po3035 = n50963 | n50964;
  assign n50966 = ~n14403 & n50306;
  assign n50967 = pi2718 & ~n50306;
  assign po3036 = n50966 | n50967;
  assign n50969 = ~n12726 & n50286;
  assign n50970 = pi2719 & ~n50286;
  assign po3037 = n50969 | n50970;
  assign n50972 = ~n13701 & n50286;
  assign n50973 = pi2720 & ~n50286;
  assign po3038 = n50972 | n50973;
  assign n50975 = ~n13988 & n50286;
  assign n50976 = pi2721 & ~n50286;
  assign po3039 = n50975 | n50976;
  assign n50978 = ~n12415 & n50286;
  assign n50979 = pi2722 & ~n50286;
  assign po3040 = n50978 | n50979;
  assign n50981 = ~n14816 & n50286;
  assign n50982 = pi2723 & ~n50286;
  assign po3041 = n50981 | n50982;
  assign n50984 = ~n15115 & n50286;
  assign n50985 = pi2724 & ~n50286;
  assign po3042 = n50984 | n50985;
  assign n50987 = ~n10608 & n50286;
  assign n50988 = pi2725 & ~n50286;
  assign po3043 = n50987 | n50988;
  assign n50990 = ~n14403 & n50286;
  assign n50991 = pi2726 & ~n50286;
  assign po3044 = n50990 | n50991;
  assign n50993 = ~n11181 & n50286;
  assign n50994 = pi2727 & ~n50286;
  assign po3045 = n50993 | n50994;
  assign n50996 = ~n12726 & n50377;
  assign n50997 = pi2728 & ~n50377;
  assign po3046 = n50996 | n50997;
  assign n50999 = ~n13121 & n50377;
  assign n51000 = pi2729 & ~n50377;
  assign po3047 = n50999 | n51000;
  assign n51002 = ~n13398 & n50377;
  assign n51003 = pi2730 & ~n50377;
  assign po3048 = n51002 | n51003;
  assign n51005 = ~n13988 & n50377;
  assign n51006 = pi2731 & ~n50377;
  assign po3049 = n51005 | n51006;
  assign n51008 = ~n12415 & n50377;
  assign n51009 = pi2732 & ~n50377;
  assign po3050 = n51008 | n51009;
  assign n51011 = ~n14816 & n50377;
  assign n51012 = pi2733 & ~n50377;
  assign po3051 = n51011 | n51012;
  assign n51014 = ~n12061 & n50377;
  assign n51015 = pi2734 & ~n50377;
  assign po3052 = n51014 | n51015;
  assign n51017 = ~n10608 & n50377;
  assign n51018 = pi2735 & ~n50377;
  assign po3053 = n51017 | n51018;
  assign n51020 = ~n15426 & n50377;
  assign n51021 = pi2736 & ~n50377;
  assign po3054 = n51020 | n51021;
  assign n51023 = ~n14403 & n50377;
  assign n51024 = pi2737 & ~n50377;
  assign po3055 = n51023 | n51024;
  assign n51026 = ~n12726 & n50343;
  assign n51027 = pi2738 & ~n50343;
  assign po3056 = n51026 | n51027;
  assign n51029 = ~n13701 & n50343;
  assign n51030 = pi2739 & ~n50343;
  assign po3057 = n51029 | n51030;
  assign n51032 = ~n13398 & n50343;
  assign n51033 = pi2740 & ~n50343;
  assign po3058 = n51032 | n51033;
  assign n51035 = ~n13988 & n50343;
  assign n51036 = pi2741 & ~n50343;
  assign po3059 = n51035 | n51036;
  assign n51038 = ~n14816 & n50343;
  assign n51039 = pi2742 & ~n50343;
  assign po3060 = n51038 | n51039;
  assign n51041 = ~n12061 & n50343;
  assign n51042 = pi2743 & ~n50343;
  assign po3061 = n51041 | n51042;
  assign n51044 = ~n9825 & n50343;
  assign n51045 = pi2744 & ~n50343;
  assign po3062 = n51044 | n51045;
  assign n51047 = ~n14403 & n50343;
  assign n51048 = pi2745 & ~n50343;
  assign po3063 = n51047 | n51048;
  assign n51050 = pi2746 & ~n50313;
  assign n51051 = n38122 & n50313;
  assign po3064 = n51050 | n51051;
  assign n51053 = pi2747 & ~n50313;
  assign n51054 = n38139 & n50313;
  assign po3065 = n51053 | n51054;
  assign n51056 = pi2748 & ~n50313;
  assign n51057 = n38156 & n50313;
  assign po3066 = n51056 | n51057;
  assign n51059 = pi2749 & ~n50313;
  assign n51060 = n38190 & n50313;
  assign po3067 = n51059 | n51060;
  assign n51062 = pi2750 & ~n50313;
  assign n51063 = n38207 & n50313;
  assign po3068 = n51062 | n51063;
  assign n51065 = pi2751 & ~n49146;
  assign n51066 = ~n39077 & n49146;
  assign po3069 = n51065 | n51066;
  assign n51068 = pi2752 & ~n50298;
  assign n51069 = n38095 & n50298;
  assign po3070 = n51068 | n51069;
  assign n51071 = pi2753 & ~n50298;
  assign n51072 = n38122 & n50298;
  assign po3071 = n51071 | n51072;
  assign n51074 = pi2754 & ~n50298;
  assign n51075 = n38139 & n50298;
  assign po3072 = n51074 | n51075;
  assign n51077 = pi2755 & ~n50298;
  assign n51078 = n38173 & n50298;
  assign po3073 = n51077 | n51078;
  assign n51080 = pi2756 & ~n50298;
  assign n51081 = n38207 & n50298;
  assign po3074 = n51080 | n51081;
  assign n51083 = ~pi2757 & n8561;
  assign n51084 = ~pi0405 & n47782;
  assign n51085 = pi0420 & n51084;
  assign n51086 = pi0421 & n51085;
  assign n51087 = ~n51083 & ~n51086;
  assign po3075 = po3627 & ~n51087;
  assign n51089 = ~pi2758 & n8561;
  assign n51090 = ~n47785 & ~n51089;
  assign po3076 = po3627 & ~n51090;
  assign n51092 = ~pi2759 & ~n48192;
  assign n51093 = ~pi2759 & pi3199;
  assign n51094 = n48194 & n51093;
  assign n51095 = pi2759 & ~n48195;
  assign n51096 = ~n51094 & ~n51095;
  assign n51097 = n48192 & n51096;
  assign n51098 = ~n51092 & ~n51097;
  assign po3077 = ~n36174 & n51098;
  assign n51100 = ~pi2760 & ~n50219;
  assign n51101 = pi2760 & n50219;
  assign n51102 = ~n51100 & ~n51101;
  assign po3078 = ~n49739 & ~n51102;
  assign n51104 = ~pi2761 & ~n50726;
  assign n51105 = pi0730 & n50726;
  assign po3079 = n51104 | n51105;
  assign n51107 = ~pi2762 & ~n50726;
  assign n51108 = pi0938 & n50726;
  assign po3080 = n51107 | n51108;
  assign n51110 = pi2763 & n8561;
  assign n51111 = ~n50140 & ~n51110;
  assign po3081 = po3627 & ~n51111;
  assign n51113 = pi0465 & n50482;
  assign n51114 = n13988 & ~n50482;
  assign n51115 = ~n51113 & ~n51114;
  assign n51116 = ~n50487 & n51115;
  assign n51117 = pi2764 & n50487;
  assign po3082 = n51116 | n51117;
  assign n51119 = ~n41540 & n41542;
  assign po3084 = pi2766 | n51119;
  assign n51121 = ~n46577 & ~n46588;
  assign n51122 = n46588 & ~n51121;
  assign n51123 = ~n46960 & n51122;
  assign n51124 = pi2767 & n51121;
  assign po3085 = n51123 | n51124;
  assign n51126 = ~n12726 & ~n50436;
  assign n51127 = pi2768 & n50436;
  assign po3086 = n51126 | n51127;
  assign n51129 = pi2769 & n39529;
  assign po3087 = n46822 | n51129;
  assign n51131 = ~pi2772 & n50218;
  assign n51132 = ~pi2507 & n51131;
  assign n51133 = n50223 & n51132;
  assign n51134 = ~pi2770 & ~n51133;
  assign n51135 = pi2770 & n51133;
  assign n51136 = ~n51134 & ~n51135;
  assign po3088 = ~n49739 & ~n51136;
  assign n51138 = pi2523 & ~pi2771;
  assign n51139 = ~pi2523 & pi2771;
  assign n51140 = ~n51138 & ~n51139;
  assign po3089 = ~n49739 & ~n51140;
  assign n51142 = ~pi2760 & n50219;
  assign n51143 = pi2772 & n51142;
  assign n51144 = ~pi2772 & ~n51142;
  assign n51145 = ~n51143 & ~n51144;
  assign po3090 = ~n49739 & ~n51145;
  assign n51147 = ~n12061 & n50286;
  assign n51148 = pi2773 & ~n50286;
  assign po3091 = n51147 | n51148;
  assign n51150 = ~n9825 & n50286;
  assign n51151 = pi2774 & ~n50286;
  assign po3092 = n51150 | n51151;
  assign n51153 = n38752 & po3574;
  assign n51154 = ~pi2775 & ~n51153;
  assign n51155 = pi0824 & n51153;
  assign po3093 = n51154 | n51155;
  assign n51157 = ~n38488 & n50313;
  assign n51158 = pi2776 & ~n50313;
  assign po3094 = n51157 | n51158;
  assign n51160 = n38252 & n38262;
  assign n51161 = ~n38253 & n51160;
  assign n51162 = pi2777 & ~n38262;
  assign po3095 = n51161 | n51162;
  assign n51164 = ~pi0598 & n30707;
  assign n51165 = ~n9352 & n51164;
  assign n51166 = ~n47751 & n51165;
  assign n51167 = pi2778 & ~n51165;
  assign po3096 = n51166 | n51167;
  assign n51169 = n9345 & n35827;
  assign n51170 = ~n8561 & n51169;
  assign n51171 = ~pi0422 & n51170;
  assign n51172 = pi2779 & n8561;
  assign po3097 = n51171 | n51172;
  assign n51174 = ~n38473 & n50313;
  assign n51175 = pi2780 & ~n50313;
  assign po3098 = n51174 | n51175;
  assign n51177 = ~n46897 & n50627;
  assign n51178 = pi2781 & ~n50627;
  assign po3099 = n51177 | n51178;
  assign n51180 = ~n47697 & n50627;
  assign n51181 = pi2782 & ~n50627;
  assign po3100 = n51180 | n51181;
  assign n51183 = ~pi0575 & n30707;
  assign n51184 = ~n9352 & n51183;
  assign n51185 = ~n24446 & n51184;
  assign n51186 = pi2783 & ~n51184;
  assign po3101 = n51185 | n51186;
  assign n51188 = ~n24744 & n51184;
  assign n51189 = pi2784 & ~n51184;
  assign po3102 = n51188 | n51189;
  assign n51191 = pi2785 & ~n45004;
  assign n51192 = ~n48590 & n51191;
  assign n51193 = pi0565 & ~pi3146;
  assign n51194 = n48590 & n51193;
  assign po3103 = n51192 | n51194;
  assign n51196 = n38766 & po3574;
  assign n51197 = ~pi2786 & ~n51196;
  assign n51198 = pi0858 & n51196;
  assign po3104 = n51197 | n51198;
  assign n51200 = ~n47688 & n51165;
  assign n51201 = pi2787 & ~n51165;
  assign po3105 = n51200 | n51201;
  assign n51203 = pi2788 & ~n50291;
  assign n51204 = n49651 & n50291;
  assign po3106 = n51203 | n51204;
  assign n51206 = ~n36384 & n49693;
  assign n51207 = pi2789 & n8561;
  assign po3107 = n51206 | n51207;
  assign n51209 = n38760 & po3574;
  assign n51210 = ~pi2790 & ~n51209;
  assign n51211 = pi0851 & n51209;
  assign po3108 = n51210 | n51211;
  assign n51213 = n38770 & po3574;
  assign n51214 = ~pi2791 & ~n51213;
  assign n51215 = pi0938 & n51213;
  assign po3109 = n51214 | n51215;
  assign n51217 = n38749 & po3574;
  assign n51218 = ~pi0823 & n51217;
  assign n51219 = pi2792 & ~n51217;
  assign po3110 = ~n51218 & ~n51219;
  assign n51221 = ~pi0649 & n30707;
  assign n51222 = ~n9352 & n51221;
  assign n51223 = ~n24256 & n51222;
  assign n51224 = pi2793 & ~n51222;
  assign po3111 = n51223 | n51224;
  assign n51226 = pi2794 & ~n50291;
  assign n51227 = n49774 & n50291;
  assign po3112 = n51226 | n51227;
  assign n51229 = pi0422 & n51170;
  assign n51230 = pi2795 & n8561;
  assign po3113 = n51229 | n51230;
  assign n51232 = pi2796 & ~n50291;
  assign n51233 = n49597 & n50291;
  assign po3114 = n51232 | n51233;
  assign n51235 = pi2797 & ~n50291;
  assign n51236 = n49611 & n50291;
  assign po3115 = n51235 | n51236;
  assign n51238 = ~pi2798 & n48383;
  assign n51239 = pi2798 & ~n48383;
  assign n51240 = ~n51238 & ~n51239;
  assign po3116 = n48409 & n51240;
  assign n51242 = ~pi2799 & n48383;
  assign n51243 = ~pi2799 & ~n48385;
  assign n51244 = ~n48386 & ~n51243;
  assign n51245 = ~n48383 & ~n51244;
  assign n51246 = ~n51242 & ~n51245;
  assign po3117 = n48409 & n51246;
  assign n51248 = po3745 & n42233;
  assign po3118 = n33823 & n51248;
  assign n51250 = ~n27570 & n51222;
  assign n51251 = pi2801 & ~n51222;
  assign po3119 = n51250 | n51251;
  assign n51253 = ~n8561 & ~n36434;
  assign n51254 = ~pi2802 & n8561;
  assign po3120 = n51253 | n51254;
  assign n51256 = ~n30333 & n51222;
  assign n51257 = pi2803 & ~n51222;
  assign po3121 = n51256 | n51257;
  assign n51259 = ~n30309 & n51222;
  assign n51260 = pi2804 & ~n51222;
  assign po3122 = n51259 | n51260;
  assign n51262 = ~n24265 & n51222;
  assign n51263 = pi2805 & ~n51222;
  assign po3123 = n51262 | n51263;
  assign n51265 = ~pi2806 & ~n51213;
  assign n51266 = pi0785 & n51213;
  assign po3124 = n51265 | n51266;
  assign n51268 = ~n25699 & n51222;
  assign n51269 = pi2807 & ~n51222;
  assign po3125 = n51268 | n51269;
  assign n51271 = ~n24769 & n51222;
  assign n51272 = pi2808 & ~n51222;
  assign po3126 = n51271 | n51272;
  assign n51274 = ~n30288 & n51222;
  assign n51275 = pi2809 & ~n51222;
  assign po3127 = n51274 | n51275;
  assign n51277 = ~n38473 & n50298;
  assign n51278 = pi2810 & ~n50298;
  assign po3128 = n51277 | n51278;
  assign n51280 = ~pi2811 & ~n51213;
  assign n51281 = pi0852 & n51213;
  assign po3129 = n51280 | n51281;
  assign n51283 = ~n8561 & ~n24376;
  assign n51284 = pi2812 & n8561;
  assign n51285 = ~n51283 & ~n51284;
  assign po3130 = ~po3897 & ~n51285;
  assign n51287 = pi2813 & n15547;
  assign n51288 = ~pi2813 & n48394;
  assign n51289 = ~pi3682 & ~po3616;
  assign n51290 = n51288 & n51289;
  assign n51291 = ~n51287 & ~n51290;
  assign n51292 = ~pi2813 & po3616;
  assign n51293 = pi3682 & n51292;
  assign n51294 = po3645 & n51293;
  assign n51295 = ~po3646 & n51294;
  assign n51296 = po3647 & n51295;
  assign po3131 = ~n51291 | n51296;
  assign n51298 = ~pi2815 & ~n51209;
  assign n51299 = pi0824 & n51209;
  assign po3133 = n51298 | n51299;
  assign n51301 = ~pi2779 & ~pi3257;
  assign n51302 = ~n8307 & ~n51301;
  assign n51303 = ~n16460 & ~n44983;
  assign n51304 = n8196 & n51303;
  assign n51305 = n51302 & n51304;
  assign n51306 = pi3698 & n51305;
  assign n51307 = pi2816 & ~n51305;
  assign po3134 = n51306 | n51307;
  assign n51309 = pi3696 & n51305;
  assign n51310 = pi2817 & ~n51305;
  assign po3135 = n51309 | n51310;
  assign n51312 = ~pi2818 & ~n51153;
  assign n51313 = pi0821 & n51153;
  assign po3136 = n51312 | n51313;
  assign n51315 = pi3689 & n51305;
  assign n51316 = pi2819 & ~n51305;
  assign po3137 = n51315 | n51316;
  assign n51318 = ~pi0955 & n31013;
  assign n51319 = ~n31887 & ~n51318;
  assign po3138 = pi3635 & ~n51319;
  assign n51321 = n38772 & po3574;
  assign n51322 = ~pi2821 & ~n51321;
  assign n51323 = pi0938 & n51321;
  assign po3139 = n51322 | n51323;
  assign n51325 = ~pi2822 & ~n51321;
  assign n51326 = pi0851 & n51321;
  assign po3140 = n51325 | n51326;
  assign n51328 = ~pi2823 & ~n51217;
  assign n51329 = pi0857 & n51217;
  assign po3141 = n51328 | n51329;
  assign n51331 = ~pi2824 & ~n42536;
  assign n51332 = pi2824 & n41246;
  assign n51333 = ~pi2824 & ~n41246;
  assign n51334 = ~n51332 & ~n51333;
  assign n51335 = n42536 & ~n51334;
  assign po3142 = n51331 | n51335;
  assign n51337 = pi2825 & n48383;
  assign n51338 = ~pi2798 & pi2825;
  assign n51339 = pi2798 & ~pi2825;
  assign n51340 = ~n51338 & ~n51339;
  assign n51341 = ~n48383 & ~n51340;
  assign n51342 = ~n51337 & ~n51341;
  assign po3143 = n48409 & ~n51342;
  assign n51344 = pi3690 & n51305;
  assign n51345 = pi2826 & ~n51305;
  assign po3144 = n51344 | n51345;
  assign n51347 = pi3688 & n51305;
  assign n51348 = pi2827 & ~n51305;
  assign po3145 = n51347 | n51348;
  assign n51350 = pi3687 & n51305;
  assign n51351 = pi2828 & ~n51305;
  assign po3146 = n51350 | n51351;
  assign n51353 = pi3686 & n51305;
  assign n51354 = pi2829 & ~n51305;
  assign po3147 = n51353 | n51354;
  assign n51356 = pi3685 & n51305;
  assign n51357 = pi2830 & ~n51305;
  assign po3148 = n51356 | n51357;
  assign n51359 = pi3684 & n51305;
  assign n51360 = pi2831 & ~n51305;
  assign po3149 = n51359 | n51360;
  assign n51362 = pi3697 & n51305;
  assign n51363 = pi2832 & ~n51305;
  assign po3150 = n51362 | n51363;
  assign n51365 = pi3695 & n51305;
  assign n51366 = pi2833 & ~n51305;
  assign po3151 = n51365 | n51366;
  assign n51368 = pi3694 & n51305;
  assign n51369 = pi2834 & ~n51305;
  assign po3152 = n51368 | n51369;
  assign n51371 = pi3693 & n51305;
  assign n51372 = pi2835 & ~n51305;
  assign po3153 = n51371 | n51372;
  assign n51374 = pi3683 & n51305;
  assign n51375 = pi2836 & ~n51305;
  assign po3154 = n51374 | n51375;
  assign n51377 = ~pi2837 & ~n51209;
  assign n51378 = pi0785 & n51209;
  assign po3155 = n51377 | n51378;
  assign n51380 = ~pi2838 & ~n51321;
  assign n51381 = pi0852 & n51321;
  assign po3156 = n51380 | n51381;
  assign n51383 = ~pi2839 & ~n51321;
  assign n51384 = pi0860 & n51321;
  assign po3157 = n51383 | n51384;
  assign n51386 = n24309 & n25554;
  assign n51387 = ~n25999 & n51386;
  assign n51388 = pi2840 & ~n51386;
  assign po3158 = n51387 | n51388;
  assign n51390 = ~pi0711 & n30707;
  assign n51391 = ~n9352 & n51390;
  assign n51392 = ~n30267 & n51391;
  assign n51393 = pi2841 & ~n51391;
  assign po3159 = n51392 | n51393;
  assign n51395 = ~n30288 & n51391;
  assign n51396 = pi2842 & ~n51391;
  assign po3160 = n51395 | n51396;
  assign n51398 = ~n24744 & n51391;
  assign n51399 = pi2843 & ~n51391;
  assign po3161 = n51398 | n51399;
  assign n51401 = ~n24769 & n51391;
  assign n51402 = pi2844 & ~n51391;
  assign po3162 = n51401 | n51402;
  assign n51404 = ~n25699 & n51391;
  assign n51405 = pi2845 & ~n51391;
  assign po3163 = n51404 | n51405;
  assign n51407 = ~n25718 & n51391;
  assign n51408 = pi2846 & ~n51391;
  assign po3164 = n51407 | n51408;
  assign n51410 = ~n24256 & n51391;
  assign n51411 = pi2847 & ~n51391;
  assign po3165 = n51410 | n51411;
  assign n51413 = ~n24289 & n51391;
  assign n51414 = pi2848 & ~n51391;
  assign po3166 = n51413 | n51414;
  assign n51416 = ~n24446 & n51391;
  assign n51417 = pi2849 & ~n51391;
  assign po3167 = n51416 | n51417;
  assign n51419 = ~n24265 & n51391;
  assign n51420 = pi2850 & ~n51391;
  assign po3168 = n51419 | n51420;
  assign n51422 = ~n30309 & n51391;
  assign n51423 = pi2851 & ~n51391;
  assign po3169 = n51422 | n51423;
  assign n51425 = ~n30321 & n51391;
  assign n51426 = pi2852 & ~n51391;
  assign po3170 = n51425 | n51426;
  assign n51428 = ~n30333 & n51391;
  assign n51429 = pi2853 & ~n51391;
  assign po3171 = n51428 | n51429;
  assign n51431 = ~n27570 & n51391;
  assign n51432 = pi2854 & ~n51391;
  assign po3172 = n51431 | n51432;
  assign n51434 = ~n25999 & n51391;
  assign n51435 = pi2855 & ~n51391;
  assign po3173 = n51434 | n51435;
  assign n51437 = ~n24488 & n51391;
  assign n51438 = pi2856 & ~n51391;
  assign po3174 = n51437 | n51438;
  assign n51440 = ~pi2857 & ~n51321;
  assign n51441 = pi0825 & n51321;
  assign po3175 = n51440 | n51441;
  assign n51443 = ~pi2858 & ~n51321;
  assign n51444 = pi0854 & n51321;
  assign po3176 = n51443 | n51444;
  assign n51446 = n38775 & po3574;
  assign n51447 = ~pi2859 & ~n51446;
  assign n51448 = pi0860 & n51446;
  assign po3177 = n51447 | n51448;
  assign n51450 = pi3246 & po3574;
  assign n51451 = n33319 & n51450;
  assign n51452 = ~pi3266 & n51451;
  assign n51453 = pi0855 & n51452;
  assign n51454 = ~pi2860 & ~n51452;
  assign po3178 = n51453 | n51454;
  assign n51456 = ~n46906 & n50608;
  assign n51457 = pi2861 & ~n50608;
  assign po3179 = n51456 | n51457;
  assign n51459 = ~n47670 & n50627;
  assign n51460 = pi2862 & ~n50627;
  assign po3180 = n51459 | n51460;
  assign n51462 = ~n47679 & n50627;
  assign n51463 = pi2863 & ~n50627;
  assign po3181 = n51462 | n51463;
  assign n51465 = ~n47688 & n50627;
  assign n51466 = pi2864 & ~n50627;
  assign po3182 = n51465 | n51466;
  assign n51468 = ~n47706 & n50627;
  assign n51469 = pi2865 & ~n50627;
  assign po3183 = n51468 | n51469;
  assign n51471 = ~n47715 & n50627;
  assign n51472 = pi2866 & ~n50627;
  assign po3184 = n51471 | n51472;
  assign n51474 = ~n47724 & n50627;
  assign n51475 = pi2867 & ~n50627;
  assign po3185 = n51474 | n51475;
  assign n51477 = ~n46906 & n50627;
  assign n51478 = pi2868 & ~n50627;
  assign po3186 = n51477 | n51478;
  assign n51480 = ~n46906 & n50649;
  assign n51481 = pi2869 & ~n50649;
  assign po3187 = n51480 | n51481;
  assign n51483 = ~n47670 & n50668;
  assign n51484 = pi2870 & ~n50668;
  assign po3188 = n51483 | n51484;
  assign n51486 = ~n47679 & n50668;
  assign n51487 = pi2871 & ~n50668;
  assign po3189 = n51486 | n51487;
  assign n51489 = ~n47688 & n50668;
  assign n51490 = pi2872 & ~n50668;
  assign po3190 = n51489 | n51490;
  assign n51492 = ~n47697 & n50668;
  assign n51493 = pi2873 & ~n50668;
  assign po3191 = n51492 | n51493;
  assign n51495 = ~n47706 & n50668;
  assign n51496 = pi2874 & ~n50668;
  assign po3192 = n51495 | n51496;
  assign n51498 = ~n47715 & n50668;
  assign n51499 = pi2875 & ~n50668;
  assign po3193 = n51498 | n51499;
  assign n51501 = ~n46897 & n50668;
  assign n51502 = pi2876 & ~n50668;
  assign po3194 = n51501 | n51502;
  assign n51504 = ~n47724 & n50668;
  assign n51505 = pi2877 & ~n50668;
  assign po3195 = n51504 | n51505;
  assign n51507 = ~n46906 & n50668;
  assign n51508 = pi2878 & ~n50668;
  assign po3196 = n51507 | n51508;
  assign n51510 = ~n30540 & n50668;
  assign n51511 = pi2879 & ~n50668;
  assign po3197 = n51510 | n51511;
  assign n51513 = ~pi2880 & ~n51321;
  assign n51514 = pi0824 & n51321;
  assign po3198 = n51513 | n51514;
  assign n51516 = ~pi2881 & ~n51217;
  assign n51517 = pi0730 & n51217;
  assign po3199 = n51516 | n51517;
  assign n51519 = ~pi2882 & ~n51153;
  assign n51520 = ~pi0937 & n51153;
  assign po3200 = n51519 | n51520;
  assign n51522 = ~pi2883 & ~n51217;
  assign n51523 = pi0858 & n51217;
  assign po3201 = n51522 | n51523;
  assign n51525 = ~pi2884 & ~n51321;
  assign n51526 = pi0731 & n51321;
  assign po3202 = n51525 | n51526;
  assign n51528 = ~pi2885 & ~n51209;
  assign n51529 = pi0856 & n51209;
  assign po3203 = n51528 | n51529;
  assign n51531 = ~pi2886 & ~n51196;
  assign n51532 = pi0856 & n51196;
  assign po3204 = n51531 | n51532;
  assign n51534 = n38757 & po3574;
  assign n51535 = ~pi2887 & ~n51534;
  assign n51536 = pi0825 & n51534;
  assign po3205 = n51535 | n51536;
  assign n51538 = ~n30267 & n51386;
  assign n51539 = pi2888 & ~n51386;
  assign po3206 = n51538 | n51539;
  assign n51541 = ~n30288 & n51386;
  assign n51542 = pi2889 & ~n51386;
  assign po3207 = n51541 | n51542;
  assign n51544 = ~n24769 & n51386;
  assign n51545 = pi2890 & ~n51386;
  assign po3208 = n51544 | n51545;
  assign n51547 = ~n24256 & n51386;
  assign n51548 = pi2891 & ~n51386;
  assign po3209 = n51547 | n51548;
  assign n51550 = ~n24289 & n51386;
  assign n51551 = pi2892 & ~n51386;
  assign po3210 = n51550 | n51551;
  assign n51553 = ~n24446 & n51386;
  assign n51554 = pi2893 & ~n51386;
  assign po3211 = n51553 | n51554;
  assign n51556 = ~n24265 & n51386;
  assign n51557 = pi2894 & ~n51386;
  assign po3212 = n51556 | n51557;
  assign n51559 = ~n30333 & n51386;
  assign n51560 = pi2895 & ~n51386;
  assign po3213 = n51559 | n51560;
  assign n51562 = ~n27570 & n51386;
  assign n51563 = pi2896 & ~n51386;
  assign po3214 = n51562 | n51563;
  assign n51565 = ~n24488 & n51386;
  assign n51566 = pi2897 & ~n51386;
  assign po3215 = n51565 | n51566;
  assign n51568 = ~pi2898 & ~n51213;
  assign n51569 = pi0730 & n51213;
  assign po3216 = n51568 | n51569;
  assign n51571 = ~pi2899 & ~n51153;
  assign n51572 = pi0823 & n51153;
  assign po3217 = n51571 | n51572;
  assign n51574 = ~pi2900 & ~n51534;
  assign n51575 = pi0731 & n51534;
  assign po3218 = n51574 | n51575;
  assign n51577 = ~pi2901 & ~n51534;
  assign n51578 = pi0856 & n51534;
  assign po3219 = n51577 | n51578;
  assign n51580 = ~pi2902 & ~n51213;
  assign n51581 = pi0853 & n51213;
  assign po3220 = n51580 | n51581;
  assign n51583 = ~pi2903 & ~n51217;
  assign n51584 = pi0938 & n51217;
  assign po3221 = n51583 | n51584;
  assign n51586 = ~pi2904 & ~n51213;
  assign n51587 = pi0855 & n51213;
  assign po3222 = n51586 | n51587;
  assign n51589 = ~pi2905 & ~n51217;
  assign n51590 = pi0860 & n51217;
  assign po3223 = n51589 | n51590;
  assign n51592 = ~pi2906 & ~n51209;
  assign n51593 = pi0855 & n51209;
  assign po3224 = n51592 | n51593;
  assign n51595 = ~pi2907 & ~n51534;
  assign n51596 = pi0852 & n51534;
  assign po3225 = n51595 | n51596;
  assign n51598 = ~pi2908 & ~n51534;
  assign n51599 = pi0854 & n51534;
  assign po3226 = n51598 | n51599;
  assign n51601 = ~pi2909 & ~n51209;
  assign n51602 = pi0854 & n51209;
  assign po3227 = n51601 | n51602;
  assign n51604 = ~pi2910 & ~n51209;
  assign n51605 = pi0825 & n51209;
  assign po3228 = n51604 | n51605;
  assign n51607 = ~n8561 & ~n24361;
  assign n51608 = pi2911 & n8561;
  assign n51609 = ~n51607 & ~n51608;
  assign po3229 = ~po3897 & ~n51609;
  assign n51611 = pi2912 & n8561;
  assign n51612 = ~n8561 & ~n24369;
  assign n51613 = ~n51611 & ~n51612;
  assign po3230 = ~po3897 & ~n51613;
  assign n51615 = pi2913 & n8561;
  assign n51616 = ~n8561 & ~n24354;
  assign n51617 = ~n51615 & ~n51616;
  assign po3231 = ~po3897 & ~n51617;
  assign n51619 = ~n30309 & n51386;
  assign n51620 = pi2914 & ~n51386;
  assign po3232 = n51619 | n51620;
  assign n51622 = ~pi2915 & ~n51153;
  assign n51623 = pi0857 & n51153;
  assign po3233 = n51622 | n51623;
  assign n51625 = ~n47652 & n51165;
  assign n51626 = pi2916 & ~n51165;
  assign po3234 = n51625 | n51626;
  assign n51628 = ~n47661 & n51165;
  assign n51629 = pi2917 & ~n51165;
  assign po3235 = n51628 | n51629;
  assign n51631 = ~n47670 & n51165;
  assign n51632 = pi2918 & ~n51165;
  assign po3236 = n51631 | n51632;
  assign n51634 = ~n47679 & n51165;
  assign n51635 = pi2919 & ~n51165;
  assign po3237 = n51634 | n51635;
  assign n51637 = ~n47697 & n51165;
  assign n51638 = pi2920 & ~n51165;
  assign po3238 = n51637 | n51638;
  assign n51640 = ~n47706 & n51165;
  assign n51641 = pi2921 & ~n51165;
  assign po3239 = n51640 | n51641;
  assign n51643 = ~n47715 & n51165;
  assign n51644 = pi2922 & ~n51165;
  assign po3240 = n51643 | n51644;
  assign n51646 = ~n46897 & n51165;
  assign n51647 = pi2923 & ~n51165;
  assign po3241 = n51646 | n51647;
  assign n51649 = ~n47724 & n51165;
  assign n51650 = pi2924 & ~n51165;
  assign po3242 = n51649 | n51650;
  assign n51652 = ~n46906 & n51165;
  assign n51653 = pi2925 & ~n51165;
  assign po3243 = n51652 | n51653;
  assign n51655 = ~n47733 & n51165;
  assign n51656 = pi2926 & ~n51165;
  assign po3244 = n51655 | n51656;
  assign n51658 = ~n47742 & n51165;
  assign n51659 = pi2927 & ~n51165;
  assign po3245 = n51658 | n51659;
  assign n51661 = ~n47760 & n51165;
  assign n51662 = pi2928 & ~n51165;
  assign po3246 = n51661 | n51662;
  assign n51664 = ~n30540 & n51165;
  assign n51665 = pi2929 & ~n51165;
  assign po3247 = n51664 | n51665;
  assign n51667 = ~pi2930 & ~n51153;
  assign n51668 = pi0825 & n51153;
  assign po3248 = n51667 | n51668;
  assign n51670 = ~n30267 & n51222;
  assign n51671 = pi2931 & ~n51222;
  assign po3249 = n51670 | n51671;
  assign n51673 = ~n24744 & n51222;
  assign n51674 = pi2932 & ~n51222;
  assign po3250 = n51673 | n51674;
  assign n51676 = ~n25718 & n51222;
  assign n51677 = pi2933 & ~n51222;
  assign po3251 = n51676 | n51677;
  assign n51679 = ~n24289 & n51222;
  assign n51680 = pi2934 & ~n51222;
  assign po3252 = n51679 | n51680;
  assign n51682 = ~n24446 & n51222;
  assign n51683 = pi2935 & ~n51222;
  assign po3253 = n51682 | n51683;
  assign n51685 = ~n30321 & n51222;
  assign n51686 = pi2936 & ~n51222;
  assign po3254 = n51685 | n51686;
  assign n51688 = ~n25999 & n51222;
  assign n51689 = pi2937 & ~n51222;
  assign po3255 = n51688 | n51689;
  assign n51691 = ~n24488 & n51222;
  assign n51692 = pi2938 & ~n51222;
  assign po3256 = n51691 | n51692;
  assign n51694 = ~n30267 & n51184;
  assign n51695 = pi2939 & ~n51184;
  assign po3257 = n51694 | n51695;
  assign n51697 = ~n30288 & n51184;
  assign n51698 = pi2940 & ~n51184;
  assign po3258 = n51697 | n51698;
  assign n51700 = ~n24769 & n51184;
  assign n51701 = pi2941 & ~n51184;
  assign po3259 = n51700 | n51701;
  assign n51703 = ~n25699 & n51184;
  assign n51704 = pi2942 & ~n51184;
  assign po3260 = n51703 | n51704;
  assign n51706 = ~n25718 & n51184;
  assign n51707 = pi2943 & ~n51184;
  assign po3261 = n51706 | n51707;
  assign n51709 = ~n24256 & n51184;
  assign n51710 = pi2944 & ~n51184;
  assign po3262 = n51709 | n51710;
  assign n51712 = ~n24289 & n51184;
  assign n51713 = pi2945 & ~n51184;
  assign po3263 = n51712 | n51713;
  assign n51715 = ~n24265 & n51184;
  assign n51716 = pi2946 & ~n51184;
  assign po3264 = n51715 | n51716;
  assign n51718 = ~n30309 & n51184;
  assign n51719 = pi2947 & ~n51184;
  assign po3265 = n51718 | n51719;
  assign n51721 = ~n30321 & n51184;
  assign n51722 = pi2948 & ~n51184;
  assign po3266 = n51721 | n51722;
  assign n51724 = ~n30333 & n51184;
  assign n51725 = pi2949 & ~n51184;
  assign po3267 = n51724 | n51725;
  assign n51727 = ~n24488 & n51184;
  assign n51728 = pi2950 & ~n51184;
  assign po3268 = n51727 | n51728;
  assign n51730 = pi1930 & ~n8561;
  assign n51731 = pi2951 & ~n51730;
  assign n51732 = ~pi1826 & n51730;
  assign n51733 = ~n51731 & ~n51732;
  assign po3269 = po3627 & ~n51733;
  assign n51735 = pi2952 & ~n51730;
  assign n51736 = ~pi1825 & n51730;
  assign n51737 = ~n51735 & ~n51736;
  assign po3270 = po3627 & ~n51737;
  assign n51739 = pi2953 & ~n50291;
  assign n51740 = n49637 & n50291;
  assign po3271 = n51739 | n51740;
  assign n51742 = ~pi2954 & ~n51534;
  assign n51743 = pi0824 & n51534;
  assign po3272 = n51742 | n51743;
  assign n51745 = ~pi2955 & ~n51534;
  assign n51746 = pi0859 & n51534;
  assign po3273 = n51745 | n51746;
  assign n51748 = ~pi2956 & ~n51209;
  assign n51749 = pi0731 & n51209;
  assign po3274 = n51748 | n51749;
  assign n51751 = ~pi2957 & ~n51153;
  assign n51752 = pi0860 & n51153;
  assign po3275 = n51751 | n51752;
  assign n51754 = ~pi2958 & ~n51153;
  assign n51755 = pi0852 & n51153;
  assign po3276 = n51754 | n51755;
  assign n51757 = ~pi2959 & ~n51196;
  assign n51758 = pi0857 & n51196;
  assign po3277 = n51757 | n51758;
  assign n51760 = ~n38413 & n50313;
  assign n51761 = pi2960 & ~n50313;
  assign po3278 = n51760 | n51761;
  assign n51763 = ~n38428 & n50313;
  assign n51764 = pi2961 & ~n50313;
  assign po3279 = n51763 | n51764;
  assign n51766 = ~n38443 & n50313;
  assign n51767 = pi2962 & ~n50313;
  assign po3280 = n51766 | n51767;
  assign n51769 = ~n38458 & n50313;
  assign n51770 = pi2963 & ~n50313;
  assign po3281 = n51769 | n51770;
  assign n51772 = ~n38503 & n50313;
  assign n51773 = pi2964 & ~n50313;
  assign po3282 = n51772 | n51773;
  assign n51775 = ~n38413 & n50298;
  assign n51776 = pi2965 & ~n50298;
  assign po3283 = n51775 | n51776;
  assign n51778 = ~n38458 & n50298;
  assign n51779 = pi2966 & ~n50298;
  assign po3284 = n51778 | n51779;
  assign n51781 = ~n38488 & n50298;
  assign n51782 = pi2967 & ~n50298;
  assign po3285 = n51781 | n51782;
  assign n51784 = ~n38503 & n50298;
  assign n51785 = pi2968 & ~n50298;
  assign po3286 = n51784 | n51785;
  assign n51787 = ~n30321 & n51386;
  assign n51788 = pi2969 & ~n51386;
  assign po3287 = n51787 | n51788;
  assign n51790 = ~pi2970 & ~n51213;
  assign n51791 = pi0851 & n51213;
  assign po3288 = n51790 | n51791;
  assign n51793 = ~pi2971 & ~n51153;
  assign n51794 = pi0851 & n51153;
  assign po3289 = n51793 | n51794;
  assign n51796 = ~pi2972 & ~n51196;
  assign n51797 = pi0825 & n51196;
  assign po3290 = n51796 | n51797;
  assign n51799 = ~pi2973 & ~n51217;
  assign n51800 = pi0821 & n51217;
  assign po3291 = n51799 | n51800;
  assign n51802 = ~pi0833 & ~n9352;
  assign n51803 = pi3237 & ~n51802;
  assign n51804 = ~pi2974 & n51803;
  assign n51805 = ~n13398 & n51802;
  assign po3292 = n51804 | n51805;
  assign n51807 = pi3239 & ~n51802;
  assign n51808 = ~pi2975 & n51807;
  assign n51809 = ~n15115 & n51802;
  assign po3293 = n51808 | n51809;
  assign n51811 = pi3227 & ~n51802;
  assign n51812 = ~pi2976 & n51811;
  assign n51813 = ~n11181 & n51802;
  assign po3294 = n51812 | n51813;
  assign n51815 = ~pi2977 & ~n51196;
  assign n51816 = pi0852 & n51196;
  assign po3295 = n51815 | n51816;
  assign n51818 = ~pi1000 & n9365;
  assign n51819 = ~n14816 & n51818;
  assign n51820 = pi2978 & ~n51818;
  assign po3296 = n51819 | n51820;
  assign n51822 = ~n15115 & n51818;
  assign n51823 = pi2979 & ~n51818;
  assign po3297 = n51822 | n51823;
  assign n51825 = ~n12061 & n51818;
  assign n51826 = pi2980 & ~n51818;
  assign po3298 = n51825 | n51826;
  assign n51828 = ~n11181 & n51818;
  assign n51829 = pi2981 & ~n51818;
  assign po3299 = n51828 | n51829;
  assign n51831 = ~n8561 & n24813;
  assign n51832 = ~pi2982 & n8561;
  assign n51833 = ~n51831 & ~n51832;
  assign po3300 = po3627 & ~n51833;
  assign n51835 = ~n8561 & n34038;
  assign n51836 = pi0421 & n45053;
  assign n51837 = n51835 & n51836;
  assign n51838 = ~pi2983 & n8561;
  assign n51839 = ~n51837 & ~n51838;
  assign po3301 = po3627 & ~n51839;
  assign n51841 = ~pi2984 & ~n51196;
  assign n51842 = pi0854 & n51196;
  assign po3302 = n51841 | n51842;
  assign n51844 = pi2985 & ~n39893;
  assign n51845 = pi3686 & n39893;
  assign po3303 = n51844 | n51845;
  assign n51847 = ~n12061 & n50201;
  assign n51848 = pi2986 & ~n50201;
  assign po3304 = n51847 | n51848;
  assign n51850 = ~n17199 & n50201;
  assign n51851 = pi2987 & ~n50201;
  assign po3305 = n51850 | n51851;
  assign n51853 = ~n9825 & n50201;
  assign n51854 = pi2988 & ~n50201;
  assign po3306 = n51853 | n51854;
  assign n51856 = ~n10608 & n50201;
  assign n51857 = pi2989 & ~n50201;
  assign po3307 = n51856 | n51857;
  assign n51859 = ~n11181 & n50201;
  assign n51860 = pi2990 & ~n50201;
  assign po3308 = n51859 | n51860;
  assign n51862 = ~pi2991 & ~n51196;
  assign n51863 = pi0851 & n51196;
  assign po3309 = n51862 | n51863;
  assign n51865 = ~pi2994 & ~n51534;
  assign n51866 = pi0823 & n51534;
  assign po3312 = n51865 | n51866;
  assign n51868 = ~pi2995 & ~n51534;
  assign n51869 = pi0730 & n51534;
  assign po3313 = n51868 | n51869;
  assign n51871 = ~pi2996 & ~n51534;
  assign n51872 = pi0853 & n51534;
  assign po3314 = n51871 | n51872;
  assign n51874 = ~pi2997 & ~n51534;
  assign n51875 = pi0785 & n51534;
  assign po3315 = n51874 | n51875;
  assign n51877 = ~pi2998 & ~n51534;
  assign n51878 = pi0855 & n51534;
  assign po3316 = n51877 | n51878;
  assign n51880 = ~pi2999 & ~n51534;
  assign n51881 = pi0857 & n51534;
  assign po3317 = n51880 | n51881;
  assign n51883 = ~pi3000 & ~n51534;
  assign n51884 = pi0858 & n51534;
  assign po3318 = n51883 | n51884;
  assign n51886 = ~pi3001 & ~n51534;
  assign n51887 = pi0821 & n51534;
  assign po3319 = n51886 | n51887;
  assign n51889 = ~pi3002 & ~n51321;
  assign n51890 = pi0823 & n51321;
  assign po3320 = n51889 | n51890;
  assign n51892 = ~pi3003 & ~n51321;
  assign n51893 = pi0859 & n51321;
  assign po3321 = n51892 | n51893;
  assign n51895 = ~pi3004 & ~n51321;
  assign n51896 = pi0730 & n51321;
  assign po3322 = n51895 | n51896;
  assign n51898 = ~pi3005 & ~n51321;
  assign n51899 = pi0853 & n51321;
  assign po3323 = n51898 | n51899;
  assign n51901 = ~pi3006 & ~n51321;
  assign n51902 = pi0785 & n51321;
  assign po3324 = n51901 | n51902;
  assign n51904 = ~pi3007 & ~n51321;
  assign n51905 = pi0855 & n51321;
  assign po3325 = n51904 | n51905;
  assign n51907 = ~pi3008 & ~n51321;
  assign n51908 = pi0821 & n51321;
  assign po3326 = n51907 | n51908;
  assign n51910 = ~pi3009 & ~n51196;
  assign n51911 = pi0824 & n51196;
  assign po3327 = n51910 | n51911;
  assign n51913 = ~pi3010 & ~n51196;
  assign n51914 = pi0823 & n51196;
  assign po3328 = n51913 | n51914;
  assign n51916 = ~pi3011 & ~n51196;
  assign n51917 = pi0730 & n51196;
  assign po3329 = n51916 | n51917;
  assign n51919 = ~pi3012 & ~n51196;
  assign n51920 = pi0860 & n51196;
  assign po3330 = n51919 | n51920;
  assign n51922 = ~pi3013 & ~n51196;
  assign n51923 = pi0853 & n51196;
  assign po3331 = n51922 | n51923;
  assign n51925 = ~pi3014 & ~n51196;
  assign n51926 = pi0785 & n51196;
  assign po3332 = n51925 | n51926;
  assign n51928 = ~pi3015 & ~n51196;
  assign n51929 = pi0855 & n51196;
  assign po3333 = n51928 | n51929;
  assign n51931 = ~pi3016 & ~n51196;
  assign n51932 = pi0821 & n51196;
  assign po3334 = n51931 | n51932;
  assign n51934 = ~pi3017 & ~n51209;
  assign n51935 = pi0823 & n51209;
  assign po3335 = n51934 | n51935;
  assign n51937 = ~pi3018 & ~n51209;
  assign n51938 = pi0730 & n51209;
  assign po3336 = n51937 | n51938;
  assign n51940 = ~pi3019 & ~n51209;
  assign n51941 = pi0938 & n51209;
  assign po3337 = n51940 | n51941;
  assign n51943 = ~pi3020 & ~n51209;
  assign n51944 = pi0860 & n51209;
  assign po3338 = n51943 | n51944;
  assign n51946 = ~pi3021 & ~n51209;
  assign n51947 = pi0852 & n51209;
  assign po3339 = n51946 | n51947;
  assign n51949 = ~pi3022 & ~n51209;
  assign n51950 = pi0853 & n51209;
  assign po3340 = n51949 | n51950;
  assign n51952 = ~pi3023 & ~n51209;
  assign n51953 = pi0857 & n51209;
  assign po3341 = n51952 | n51953;
  assign n51955 = ~pi3024 & ~n51209;
  assign n51956 = pi0858 & n51209;
  assign po3342 = n51955 | n51956;
  assign n51958 = ~pi3025 & ~n51209;
  assign n51959 = pi0821 & n51209;
  assign po3343 = n51958 | n51959;
  assign n51961 = ~pi3026 & ~n51446;
  assign n51962 = pi0824 & n51446;
  assign po3344 = n51961 | n51962;
  assign n51964 = ~pi3027 & ~n51446;
  assign n51965 = pi0731 & n51446;
  assign po3345 = n51964 | n51965;
  assign n51967 = ~pi3028 & ~n51446;
  assign n51968 = pi0852 & n51446;
  assign po3346 = n51967 | n51968;
  assign n51970 = ~pi3029 & ~n51446;
  assign n51971 = pi0854 & n51446;
  assign po3347 = n51970 | n51971;
  assign n51973 = ~pi3030 & ~n51446;
  assign n51974 = pi0856 & n51446;
  assign po3348 = n51973 | n51974;
  assign n51976 = ~pi3031 & ~n51446;
  assign n51977 = pi0858 & n51446;
  assign po3349 = n51976 | n51977;
  assign n51979 = ~pi3032 & ~n51446;
  assign n51980 = pi0821 & n51446;
  assign po3350 = n51979 | n51980;
  assign n51982 = ~pi3033 & ~n51217;
  assign n51983 = pi0824 & n51217;
  assign po3351 = n51982 | n51983;
  assign n51985 = ~pi3034 & ~n51217;
  assign n51986 = pi0859 & n51217;
  assign po3352 = n51985 | n51986;
  assign n51988 = ~pi3035 & ~n51217;
  assign n51989 = pi0731 & n51217;
  assign po3353 = n51988 | n51989;
  assign n51991 = ~pi3036 & ~n51217;
  assign n51992 = pi0851 & n51217;
  assign po3354 = n51991 | n51992;
  assign n51994 = ~pi3037 & ~n51217;
  assign n51995 = pi0852 & n51217;
  assign po3355 = n51994 | n51995;
  assign n51997 = ~pi3038 & ~n51217;
  assign n51998 = pi0854 & n51217;
  assign po3356 = n51997 | n51998;
  assign n52000 = ~pi3039 & ~n51217;
  assign n52001 = pi0825 & n51217;
  assign po3357 = n52000 | n52001;
  assign n52003 = ~pi3040 & ~n51213;
  assign n52004 = pi0823 & n51213;
  assign po3358 = n52003 | n52004;
  assign n52006 = ~pi3041 & ~n51213;
  assign n52007 = pi0860 & n51213;
  assign po3359 = n52006 | n52007;
  assign n52009 = ~pi3042 & ~n51213;
  assign n52010 = pi0821 & n51213;
  assign po3360 = n52009 | n52010;
  assign n52012 = ~pi3043 & ~n51213;
  assign n52013 = pi0854 & n51213;
  assign po3361 = n52012 | n52013;
  assign n52015 = ~pi3044 & ~n51213;
  assign n52016 = pi0825 & n51213;
  assign po3362 = n52015 | n52016;
  assign n52018 = ~pi3045 & ~n51213;
  assign n52019 = pi0856 & n51213;
  assign po3363 = n52018 | n52019;
  assign n52021 = ~pi3046 & ~n51213;
  assign n52022 = pi0858 & n51213;
  assign po3364 = n52021 | n52022;
  assign n52024 = ~pi3047 & ~n51213;
  assign n52025 = ~pi0937 & n51213;
  assign po3365 = n52024 | n52025;
  assign n52027 = ~pi3048 & ~n51153;
  assign n52028 = pi0859 & n51153;
  assign po3366 = n52027 | n52028;
  assign n52030 = ~pi3049 & ~n51153;
  assign n52031 = pi0730 & n51153;
  assign po3367 = n52030 | n52031;
  assign n52033 = ~pi3050 & ~n51153;
  assign n52034 = pi0731 & n51153;
  assign po3368 = n52033 | n52034;
  assign n52036 = ~pi3051 & ~n51153;
  assign n52037 = pi0853 & n51153;
  assign po3369 = n52036 | n52037;
  assign n52039 = ~pi3052 & ~n51153;
  assign n52040 = pi0854 & n51153;
  assign po3370 = n52039 | n52040;
  assign n52042 = ~pi3053 & ~n51153;
  assign n52043 = pi0785 & n51153;
  assign po3371 = n52042 | n52043;
  assign n52045 = ~pi3054 & ~n51153;
  assign n52046 = pi0855 & n51153;
  assign po3372 = n52045 | n52046;
  assign n52048 = pi0853 & n51452;
  assign n52049 = pi3055 & ~n51452;
  assign po3373 = n52048 | n52049;
  assign n52051 = ~pi3056 & ~n51196;
  assign n52052 = pi0731 & n51196;
  assign po3374 = n52051 | n52052;
  assign n52054 = ~pi3057 & ~n51446;
  assign n52055 = pi0785 & n51446;
  assign po3375 = n52054 | n52055;
  assign n52057 = ~pi3058 & ~n51446;
  assign n52058 = pi0825 & n51446;
  assign po3376 = n52057 | n52058;
  assign n52060 = ~n25718 & n51386;
  assign n52061 = pi3059 & ~n51386;
  assign po3377 = n52060 | n52061;
  assign n52063 = ~pi3060 & ~n51446;
  assign n52064 = pi0851 & n51446;
  assign po3378 = n52063 | n52064;
  assign n52066 = ~pi3061 & ~n51213;
  assign n52067 = pi0824 & n51213;
  assign po3379 = n52066 | n52067;
  assign n52069 = ~pi3062 & ~n51446;
  assign n52070 = pi0938 & n51446;
  assign po3380 = n52069 | n52070;
  assign n52072 = ~n14403 & n50201;
  assign n52073 = pi3063 & ~n50201;
  assign po3381 = n52072 | n52073;
  assign n52075 = ~pi3064 & ~n51217;
  assign n52076 = pi0855 & n51217;
  assign po3382 = n52075 | n52076;
  assign n52078 = ~pi3065 & n8561;
  assign n52079 = ~n47780 & ~n52078;
  assign po3383 = po3627 & ~n52079;
  assign n52081 = ~pi3066 & ~n51209;
  assign n52082 = pi0859 & n51209;
  assign po3384 = n52081 | n52082;
  assign n52084 = ~pi3067 & ~n51534;
  assign n52085 = pi0851 & n51534;
  assign po3385 = n52084 | n52085;
  assign n52087 = pi3217 & ~n51802;
  assign n52088 = ~pi3068 & n52087;
  assign n52089 = ~n12415 & n51802;
  assign po3386 = n52088 | n52089;
  assign n52091 = ~pi3069 & ~n51153;
  assign n52092 = pi0858 & n51153;
  assign po3387 = n52091 | n52092;
  assign n52094 = ~pi3070 & ~n51446;
  assign n52095 = pi0855 & n51446;
  assign po3388 = n52094 | n52095;
  assign n52097 = ~pi3071 & ~n51217;
  assign n52098 = pi0856 & n51217;
  assign po3389 = n52097 | n52098;
  assign n52100 = ~pi3072 & ~n51534;
  assign n52101 = pi0938 & n51534;
  assign po3390 = n52100 | n52101;
  assign n52103 = ~pi3073 & ~n51534;
  assign n52104 = pi0860 & n51534;
  assign po3391 = n52103 | n52104;
  assign n52106 = ~n25699 & n51386;
  assign n52107 = pi3074 & ~n51386;
  assign po3392 = n52106 | n52107;
  assign n52109 = ~n24744 & n51386;
  assign n52110 = pi3075 & ~n51386;
  assign po3393 = n52109 | n52110;
  assign n52112 = pi3076 & ~n51730;
  assign n52113 = ~pi1827 & n51730;
  assign n52114 = ~n52112 & ~n52113;
  assign po3394 = po3627 & ~n52114;
  assign n52116 = ~pi3077 & ~n51321;
  assign n52117 = pi0857 & n51321;
  assign po3395 = n52116 | n52117;
  assign n52119 = ~pi3078 & ~n51446;
  assign n52120 = pi0857 & n51446;
  assign po3396 = n52119 | n52120;
  assign n52122 = ~n27570 & n51184;
  assign n52123 = pi3079 & ~n51184;
  assign po3397 = n52122 | n52123;
  assign n52125 = ~pi3080 & ~n51153;
  assign n52126 = pi0856 & n51153;
  assign po3398 = n52125 | n52126;
  assign n52128 = ~pi3081 & ~n51446;
  assign n52129 = pi0823 & n51446;
  assign po3399 = n52128 | n52129;
  assign n52131 = ~pi3082 & ~n51217;
  assign n52132 = pi0853 & n51217;
  assign po3400 = n52131 | n52132;
  assign n52134 = ~pi3083 & ~n51446;
  assign n52135 = pi0853 & n51446;
  assign po3401 = n52134 | n52135;
  assign n52137 = ~n30540 & n50627;
  assign n52138 = pi3084 & ~n50627;
  assign po3402 = n52137 | n52138;
  assign n52140 = ~pi3085 & ~n51321;
  assign n52141 = pi0858 & n51321;
  assign po3403 = n52140 | n52141;
  assign n52143 = n38779 & po3574;
  assign n52144 = pi0853 & n52143;
  assign po3404 = pi3086 & n52144;
  assign n52146 = ~pi3087 & ~n51446;
  assign n52147 = pi0859 & n51446;
  assign po3405 = n52146 | n52147;
  assign n52149 = ~pi3088 & ~n51213;
  assign n52150 = pi0857 & n51213;
  assign po3406 = n52149 | n52150;
  assign n52152 = ~pi3089 & ~n51217;
  assign n52153 = pi0785 & n51217;
  assign po3407 = n52152 | n52153;
  assign n52155 = ~pi3090 & ~n51446;
  assign n52156 = pi0730 & n51446;
  assign po3408 = n52155 | n52156;
  assign n52158 = ~n15426 & n50201;
  assign n52159 = pi3091 & ~n50201;
  assign po3409 = n52158 | n52159;
  assign n52161 = ~pi3092 & ~n51213;
  assign n52162 = pi0731 & n51213;
  assign po3410 = n52161 | n52162;
  assign n52164 = ~n38443 & n50298;
  assign n52165 = pi3093 & ~n50298;
  assign po3411 = n52164 | n52165;
  assign n52167 = ~pi3094 & ~n51321;
  assign n52168 = pi0856 & n51321;
  assign po3412 = n52167 | n52168;
  assign n52170 = ~pi3095 & ~n51196;
  assign n52171 = pi0859 & n51196;
  assign po3413 = n52170 | n52171;
  assign n52173 = ~n38428 & n50298;
  assign n52174 = pi3096 & ~n50298;
  assign po3414 = n52173 | n52174;
  assign n52176 = ~n17368 & n50201;
  assign n52177 = pi3097 & ~n50201;
  assign po3415 = n52176 | n52177;
  assign n52179 = pi0825 & n51452;
  assign n52180 = ~pi3098 & ~n51452;
  assign po3417 = n52179 | n52180;
  assign n52182 = ~n15115 & n50201;
  assign n52183 = pi3099 & ~n50201;
  assign po3418 = n52182 | n52183;
  assign n52185 = ~n14816 & n50201;
  assign n52186 = pi3100 & ~n50201;
  assign po3419 = n52185 | n52186;
  assign n52188 = ~n13701 & n50201;
  assign n52189 = pi3101 & ~n50201;
  assign po3420 = n52188 | n52189;
  assign n52191 = pi3102 & ~n39893;
  assign n52192 = pi3687 & n39893;
  assign po3421 = n52191 | n52192;
  assign n52194 = ~pi3103 & ~n51213;
  assign n52195 = pi0859 & n51213;
  assign po3422 = n52194 | n52195;
  assign n52197 = pi3104 & ~n39893;
  assign n52198 = pi3685 & n39893;
  assign po3423 = n52197 | n52198;
  assign n52200 = pi3105 & ~n39893;
  assign n52201 = pi3684 & n39893;
  assign po3424 = n52200 | n52201;
  assign n52203 = pi3106 & ~n39893;
  assign n52204 = pi3683 & n39893;
  assign po3425 = n52203 | n52204;
  assign n52206 = ~n12726 & n50201;
  assign n52207 = pi3107 & ~n50201;
  assign po3426 = n52206 | n52207;
  assign n52209 = ~pi3108 & ~n51196;
  assign n52210 = pi0938 & n51196;
  assign po3427 = n52209 | n52210;
  assign n52212 = pi3109 & ~n39893;
  assign n52213 = pi3688 & n39893;
  assign po3428 = n52212 | n52213;
  assign n52215 = ~pi3110 & ~n51153;
  assign n52216 = pi0938 & n51153;
  assign po3429 = n52215 | n52216;
  assign n52218 = pi3111 & ~n39893;
  assign n52219 = pi3689 & n39893;
  assign po3430 = n52218 | n52219;
  assign n52221 = pi3112 & ~n39893;
  assign n52222 = pi3690 & n39893;
  assign po3431 = n52221 | n52222;
  assign n52224 = ~n25999 & n51184;
  assign n52225 = pi3113 & ~n51184;
  assign po3432 = n52224 | n52225;
  assign n52227 = ~pi2029 & n50149;
  assign n52228 = ~pi2047 & ~n50149;
  assign n52229 = ~n52227 & ~n52228;
  assign n52230 = n51730 & ~n52229;
  assign n52231 = pi3114 & ~n51730;
  assign po3433 = n52230 | n52231;
  assign n52233 = pi3115 & ~n51730;
  assign n52234 = ~pi2045 & ~n50149;
  assign n52235 = n51730 & n52234;
  assign po3434 = n52233 | n52235;
  assign n52237 = pi3116 & ~n51730;
  assign n52238 = ~pi2065 & ~n50149;
  assign n52239 = n51730 & n52238;
  assign po3435 = n52237 | n52239;
  assign n52241 = pi3117 & ~n51730;
  assign n52242 = ~pi2037 & ~n50149;
  assign n52243 = n51730 & n52242;
  assign po3436 = n52241 | n52243;
  assign n52245 = ~pi2030 & n50149;
  assign n52246 = ~pi2046 & ~n50149;
  assign n52247 = ~n52245 & ~n52246;
  assign n52248 = n51730 & ~n52247;
  assign n52249 = pi3118 & ~n51730;
  assign po3437 = n52248 | n52249;
  assign n52251 = n24251 & n25554;
  assign n52252 = ~n30321 & n52251;
  assign n52253 = pi3119 & ~n52251;
  assign po3438 = n52252 | n52253;
  assign n52255 = pi3120 & n36128;
  assign n52256 = n36060 & n36091;
  assign po3439 = n52255 | n52256;
  assign n52258 = pi3121 & n8561;
  assign n52259 = ~n50151 & ~n52258;
  assign po3440 = po3627 & ~n52259;
  assign n52261 = ~n24289 & n52251;
  assign n52262 = pi3122 & ~n52251;
  assign po3441 = n52261 | n52262;
  assign n52264 = ~n24446 & n52251;
  assign n52265 = pi3123 & ~n52251;
  assign po3442 = n52264 | n52265;
  assign n52267 = pi3124 & ~n51730;
  assign n52268 = ~pi2062 & ~n50149;
  assign n52269 = n51730 & n52268;
  assign po3443 = n52267 | n52269;
  assign n52271 = ~n24744 & n52251;
  assign n52272 = pi3125 & ~n52251;
  assign po3444 = n52271 | n52272;
  assign n52274 = ~n30267 & n52251;
  assign n52275 = pi3126 & ~n52251;
  assign po3445 = n52274 | n52275;
  assign n52277 = n24251 & n25551;
  assign n52278 = ~n24488 & n52277;
  assign n52279 = pi3127 & ~n52277;
  assign po3446 = n52278 | n52279;
  assign n52281 = ~n24446 & n52277;
  assign n52282 = pi3128 & ~n52277;
  assign po3447 = n52281 | n52282;
  assign n52284 = ~pi3130 & n8561;
  assign n52285 = ~n8561 & n24826;
  assign po3449 = n52284 | n52285;
  assign n52287 = ~n24256 & n52277;
  assign n52288 = pi3131 & ~n52277;
  assign po3450 = n52287 | n52288;
  assign n52290 = ~n25718 & n52277;
  assign n52291 = pi3132 & ~n52277;
  assign po3451 = n52290 | n52291;
  assign n52293 = ~n24769 & n52277;
  assign n52294 = pi3133 & ~n52277;
  assign po3452 = n52293 | n52294;
  assign n52296 = ~n25699 & n52277;
  assign n52297 = pi3134 & ~n52277;
  assign po3453 = n52296 | n52297;
  assign n52299 = pi3135 & ~n51730;
  assign n52300 = ~pi2040 & ~n50149;
  assign n52301 = n51730 & n52300;
  assign po3454 = n52299 | n52301;
  assign n52303 = pi1755 & pi2107;
  assign n52304 = pi1760 & pi2110;
  assign n52305 = pi1752 & pi2104;
  assign n52306 = pi1751 & pi2103;
  assign n52307 = ~n52305 & ~n52306;
  assign n52308 = pi1754 & pi2106;
  assign n52309 = pi1753 & pi2105;
  assign n52310 = ~n52308 & ~n52309;
  assign n52311 = n52307 & n52310;
  assign n52312 = pi1759 & pi2123;
  assign n52313 = pi1758 & pi2109;
  assign n52314 = ~n52312 & ~n52313;
  assign n52315 = pi1750 & pi2102;
  assign n52316 = pi1749 & pi2101;
  assign n52317 = ~n52315 & ~n52316;
  assign n52318 = n52314 & n52317;
  assign n52319 = n52311 & n52318;
  assign n52320 = ~n52304 & n52319;
  assign n52321 = ~n52303 & n52320;
  assign n52322 = pi1757 & pi2108;
  assign n52323 = pi1756 & pi2141;
  assign n52324 = ~n52322 & ~n52323;
  assign po3456 = ~n52321 | ~n52324;
  assign n52326 = pi3138 & n9352;
  assign po3457 = n24340 | n52326;
  assign n52328 = pi3139 & ~n51730;
  assign n52329 = ~pi2041 & ~n50149;
  assign n52330 = n51730 & n52329;
  assign po3458 = n52328 | n52330;
  assign n52332 = ~n47724 & n50649;
  assign n52333 = pi3140 & ~n50649;
  assign po3459 = n52332 | n52333;
  assign n52335 = ~n30333 & n52251;
  assign n52336 = pi3143 & ~n52251;
  assign po3462 = n52335 | n52336;
  assign n52338 = pi2983 & n20522;
  assign n52339 = ~pi3145 & n9352;
  assign po3465 = n52338 | n52339;
  assign n52341 = ~pi3146 & n8561;
  assign po3466 = n51170 | n52341;
  assign n52343 = ~pi3147 & ~n39526;
  assign po3467 = n46822 | n52343;
  assign n52345 = ~pi3526 & ~po3831;
  assign n52346 = pi3148 & n52345;
  assign n52347 = ~po3948 & ~po3849;
  assign n52348 = n52346 & n52347;
  assign n52349 = ~pi3663 & ~n52345;
  assign po3468 = n52348 | n52349;
  assign n52351 = pi3692 & n51305;
  assign n52352 = pi3149 & ~n51305;
  assign po3469 = n52351 | n52352;
  assign n52354 = pi3691 & n51305;
  assign n52355 = pi3150 & ~n51305;
  assign po3470 = n52354 | n52355;
  assign n52357 = ~n47670 & n50608;
  assign n52358 = pi3151 & ~n50608;
  assign po3471 = n52357 | n52358;
  assign n52360 = ~n47679 & n50608;
  assign n52361 = pi3152 & ~n50608;
  assign po3472 = n52360 | n52361;
  assign n52363 = ~n47688 & n50608;
  assign n52364 = pi3153 & ~n50608;
  assign po3473 = n52363 | n52364;
  assign n52366 = ~n47697 & n50608;
  assign n52367 = pi3154 & ~n50608;
  assign po3474 = n52366 | n52367;
  assign n52369 = ~n47706 & n50608;
  assign n52370 = pi3155 & ~n50608;
  assign po3475 = n52369 | n52370;
  assign n52372 = ~n47715 & n50608;
  assign n52373 = pi3156 & ~n50608;
  assign po3476 = n52372 | n52373;
  assign n52375 = ~n46897 & n50608;
  assign n52376 = pi3157 & ~n50608;
  assign po3477 = n52375 | n52376;
  assign n52378 = ~n47724 & n50608;
  assign n52379 = pi3158 & ~n50608;
  assign po3478 = n52378 | n52379;
  assign n52381 = ~n30540 & n50608;
  assign n52382 = pi3159 & ~n50608;
  assign po3479 = n52381 | n52382;
  assign n52384 = ~n47670 & n50649;
  assign n52385 = pi3160 & ~n50649;
  assign po3480 = n52384 | n52385;
  assign n52387 = ~n47679 & n50649;
  assign n52388 = pi3161 & ~n50649;
  assign po3481 = n52387 | n52388;
  assign n52390 = ~n47688 & n50649;
  assign n52391 = pi3162 & ~n50649;
  assign po3482 = n52390 | n52391;
  assign n52393 = ~n47706 & n50649;
  assign n52394 = pi3163 & ~n50649;
  assign po3483 = n52393 | n52394;
  assign n52396 = ~n47715 & n50649;
  assign n52397 = pi3164 & ~n50649;
  assign po3484 = n52396 | n52397;
  assign n52399 = ~n46897 & n50649;
  assign n52400 = pi3165 & ~n50649;
  assign po3485 = n52399 | n52400;
  assign n52402 = ~n30540 & n50649;
  assign n52403 = pi3166 & ~n50649;
  assign po3486 = n52402 | n52403;
  assign n52405 = ~n30267 & n52277;
  assign n52406 = pi3167 & ~n52277;
  assign po3487 = n52405 | n52406;
  assign n52408 = ~n30288 & n52277;
  assign n52409 = pi3168 & ~n52277;
  assign po3488 = n52408 | n52409;
  assign n52411 = ~n24744 & n52277;
  assign n52412 = pi3169 & ~n52277;
  assign po3489 = n52411 | n52412;
  assign n52414 = ~n24289 & n52277;
  assign n52415 = pi3170 & ~n52277;
  assign po3490 = n52414 | n52415;
  assign n52417 = ~n24265 & n52277;
  assign n52418 = pi3171 & ~n52277;
  assign po3491 = n52417 | n52418;
  assign n52420 = ~n30309 & n52277;
  assign n52421 = pi3172 & ~n52277;
  assign po3492 = n52420 | n52421;
  assign n52423 = ~n30321 & n52277;
  assign n52424 = pi3173 & ~n52277;
  assign po3493 = n52423 | n52424;
  assign n52426 = ~n30333 & n52277;
  assign n52427 = pi3174 & ~n52277;
  assign po3494 = n52426 | n52427;
  assign n52429 = ~n27570 & n52277;
  assign n52430 = pi3175 & ~n52277;
  assign po3495 = n52429 | n52430;
  assign n52432 = ~n25999 & n52277;
  assign n52433 = pi3176 & ~n52277;
  assign po3496 = n52432 | n52433;
  assign n52435 = ~n30288 & n52251;
  assign n52436 = pi3177 & ~n52251;
  assign po3497 = n52435 | n52436;
  assign n52438 = ~n24769 & n52251;
  assign n52439 = pi3178 & ~n52251;
  assign po3498 = n52438 | n52439;
  assign n52441 = ~n25699 & n52251;
  assign n52442 = pi3179 & ~n52251;
  assign po3499 = n52441 | n52442;
  assign n52444 = ~n25718 & n52251;
  assign n52445 = pi3180 & ~n52251;
  assign po3500 = n52444 | n52445;
  assign n52447 = ~n24256 & n52251;
  assign n52448 = pi3181 & ~n52251;
  assign po3501 = n52447 | n52448;
  assign n52450 = ~n24265 & n52251;
  assign n52451 = pi3182 & ~n52251;
  assign po3502 = n52450 | n52451;
  assign n52453 = ~n30309 & n52251;
  assign n52454 = pi3183 & ~n52251;
  assign po3503 = n52453 | n52454;
  assign n52456 = ~n27570 & n52251;
  assign n52457 = pi3184 & ~n52251;
  assign po3504 = n52456 | n52457;
  assign n52459 = ~n25999 & n52251;
  assign n52460 = pi3185 & ~n52251;
  assign po3505 = n52459 | n52460;
  assign n52462 = pi3226 & ~n51802;
  assign n52463 = ~pi3186 & n52462;
  assign n52464 = ~n14403 & n51802;
  assign po3506 = n52463 | n52464;
  assign n52466 = pi3187 & ~n51730;
  assign n52467 = ~pi2064 & ~n50149;
  assign n52468 = n51730 & n52467;
  assign po3507 = n52466 | n52468;
  assign n52470 = pi0854 & pi3188;
  assign po3508 = n51452 & n52470;
  assign n52472 = pi3238 & ~n51802;
  assign n52473 = ~pi3189 & n52472;
  assign n52474 = ~n13701 & n51802;
  assign po3509 = n52473 | n52474;
  assign n52476 = ~pi0408 & po3627;
  assign n52477 = n9345 & n34040;
  assign n52478 = ~n8561 & n52477;
  assign n52479 = n52476 & n52478;
  assign n52480 = pi3190 & n36128;
  assign po3510 = n52479 | n52480;
  assign n52482 = n36060 & n36112;
  assign n52483 = ~pi3191 & n36128;
  assign po3511 = n52482 | n52483;
  assign n52485 = pi3192 & ~n51730;
  assign n52486 = ~pi2038 & ~n50149;
  assign n52487 = n51730 & n52486;
  assign po3512 = n52485 | n52487;
  assign n52489 = pi3193 & ~n51730;
  assign n52490 = ~pi2039 & ~n50149;
  assign n52491 = n51730 & n52490;
  assign po3513 = n52489 | n52491;
  assign n52493 = pi3194 & ~n51730;
  assign n52494 = ~pi2042 & ~n50149;
  assign n52495 = n51730 & n52494;
  assign po3514 = n52493 | n52495;
  assign n52497 = pi3195 & ~n51730;
  assign n52498 = ~pi2050 & ~n50149;
  assign n52499 = n51730 & n52498;
  assign po3515 = n52497 | n52499;
  assign n52501 = pi3196 & ~n51730;
  assign n52502 = ~pi2043 & ~n50149;
  assign n52503 = n51730 & n52502;
  assign po3516 = n52501 | n52503;
  assign n52505 = pi3197 & ~n51730;
  assign n52506 = ~pi2044 & ~n50149;
  assign n52507 = n51730 & n52506;
  assign po3517 = n52505 | n52507;
  assign n52509 = pi3198 & ~n51730;
  assign n52510 = ~pi2060 & ~n50149;
  assign n52511 = n51730 & n52510;
  assign po3518 = n52509 | n52511;
  assign n52513 = ~pi3199 & ~n48192;
  assign n52514 = ~pi3199 & ~n48194;
  assign n52515 = ~n48195 & ~n52514;
  assign n52516 = n48192 & ~n52515;
  assign n52517 = ~n52513 & ~n52516;
  assign po3519 = ~n36174 & n52517;
  assign n52519 = pi0856 & pi3200;
  assign po3520 = n51452 & n52519;
  assign n52521 = ~n47697 & n50649;
  assign n52522 = pi3201 & ~n50649;
  assign po3521 = n52521 | n52522;
  assign n52524 = ~n24488 & n52251;
  assign n52525 = pi3202 & ~n52251;
  assign po3522 = n52524 | n52525;
  assign n52527 = ~pi2487 & ~n9352;
  assign n52528 = pi3510 & n52527;
  assign n52529 = pi3511 & n52528;
  assign n52530 = ~pi3203 & ~n52528;
  assign po3523 = n52529 | n52530;
  assign n52532 = n34979 & n37340;
  assign n52533 = ~pi3204 & n52532;
  assign n52534 = pi0615 & n52533;
  assign po3524 = pi3204 | n52534;
  assign n52536 = pi0785 & pi3205;
  assign po3525 = n51452 & n52536;
  assign n52538 = pi3206 & ~n51730;
  assign n52539 = ~pi1954 & n50149;
  assign n52540 = ~pi2034 & ~n50149;
  assign n52541 = ~n52539 & ~n52540;
  assign n52542 = n51730 & ~n52541;
  assign po3526 = n52538 | n52542;
  assign n52544 = pi3207 & ~n51730;
  assign n52545 = ~pi2027 & n50149;
  assign n52546 = ~pi2066 & ~n50149;
  assign n52547 = ~n52545 & ~n52546;
  assign n52548 = n51730 & ~n52547;
  assign po3527 = n52544 | n52548;
  assign n52550 = pi3208 & ~n51730;
  assign n52551 = ~pi1970 & n50149;
  assign n52552 = ~pi2036 & ~n50149;
  assign n52553 = ~n52551 & ~n52552;
  assign n52554 = n51730 & ~n52553;
  assign po3528 = n52550 | n52554;
  assign n52556 = pi3209 & ~n51730;
  assign n52557 = ~pi2022 & n50149;
  assign n52558 = ~pi2031 & ~n50149;
  assign n52559 = ~n52557 & ~n52558;
  assign n52560 = n51730 & ~n52559;
  assign po3529 = n52556 | n52560;
  assign n52562 = pi0408 & po3627;
  assign n52563 = n50144 & n52562;
  assign n52564 = pi3210 & n36128;
  assign po3530 = n52563 | n52564;
  assign n52566 = ~pi3211 & n8561;
  assign n52567 = ~n50144 & ~n52566;
  assign po3531 = po3627 & ~n52567;
  assign n52569 = pi3212 & ~pi3534;
  assign n52570 = ~pi3488 & ~n52569;
  assign n52571 = ~pi3212 & pi3534;
  assign po3532 = n52570 | n52571;
  assign n52573 = pi3213 & ~pi3532;
  assign n52574 = ~pi3486 & ~n52573;
  assign n52575 = ~pi3213 & pi3532;
  assign po3533 = n52574 | n52575;
  assign n52577 = pi3214 & ~pi3531;
  assign n52578 = ~pi3485 & ~n52577;
  assign n52579 = ~pi3214 & pi3531;
  assign po3534 = n52578 | n52579;
  assign n52581 = ~n8621 & n8622;
  assign n52582 = n10740 & ~n10762;
  assign n52583 = ~n52581 & ~n52582;
  assign n52584 = n9345 & ~n52583;
  assign n52585 = ~pi3426 & n52584;
  assign n52586 = ~n8561 & n52585;
  assign n52587 = pi3215 & n8561;
  assign po3535 = n52586 | n52587;
  assign n52589 = ~n36433 & n49693;
  assign n52590 = pi3216 & n8561;
  assign po3536 = n52589 | n52590;
  assign n52592 = ~pi3217 & ~n51802;
  assign n52593 = pi3068 & n52592;
  assign n52594 = ~n13988 & n51802;
  assign po3537 = n52593 | n52594;
  assign n52596 = ~pi3218 & n41964;
  assign n52597 = pi3218 & ~pi3998;
  assign n52598 = ~pi3218 & pi3998;
  assign n52599 = pi3325 & ~n52598;
  assign n52600 = ~n52597 & ~n52599;
  assign n52601 = ~n41964 & n52600;
  assign po3538 = n52596 | n52601;
  assign n52603 = ~pi3219 & n41503;
  assign n52604 = pi3219 & ~pi4003;
  assign n52605 = ~pi3219 & pi4003;
  assign n52606 = pi3356 & ~n52605;
  assign n52607 = ~n52604 & ~n52606;
  assign n52608 = ~n41503 & n52607;
  assign po3539 = n52603 | n52608;
  assign n52610 = ~pi3220 & n41942;
  assign n52611 = ~pi3220 & pi4001;
  assign n52612 = pi3341 & ~n52611;
  assign n52613 = pi3220 & ~pi4001;
  assign n52614 = ~n52612 & ~n52613;
  assign n52615 = ~n41942 & n52614;
  assign po3540 = n52610 | n52615;
  assign n52617 = ~pi3221 & n41953;
  assign n52618 = ~pi3221 & pi3999;
  assign n52619 = pi3301 & ~n52618;
  assign n52620 = pi3221 & ~pi3999;
  assign n52621 = ~n52619 & ~n52620;
  assign n52622 = ~n41953 & n52621;
  assign po3541 = n52617 | n52622;
  assign n52624 = ~pi3222 & n41964;
  assign n52625 = ~pi3222 & pi3997;
  assign n52626 = pi3327 & ~n52625;
  assign n52627 = pi3222 & ~pi3997;
  assign n52628 = ~n52626 & ~n52627;
  assign n52629 = ~n41964 & n52628;
  assign po3542 = n52624 | n52629;
  assign n52631 = ~pi3223 & n41975;
  assign n52632 = pi3223 & ~pi3996;
  assign n52633 = ~pi3223 & pi3996;
  assign n52634 = pi3334 & ~n52633;
  assign n52635 = ~n52632 & ~n52634;
  assign n52636 = ~n41975 & n52635;
  assign po3543 = n52631 | n52636;
  assign n52638 = ~pi3224 & n41986;
  assign n52639 = pi3224 & ~pi4006;
  assign n52640 = ~pi3224 & pi4006;
  assign n52641 = pi3335 & ~n52640;
  assign n52642 = ~n52639 & ~n52641;
  assign n52643 = ~n41986 & n52642;
  assign po3544 = n52638 | n52643;
  assign n52645 = ~pi3225 & n41975;
  assign n52646 = ~pi3225 & pi3995;
  assign n52647 = pi3333 & ~n52646;
  assign n52648 = pi3225 & ~pi3995;
  assign n52649 = ~n52647 & ~n52648;
  assign n52650 = ~n41975 & n52649;
  assign po3545 = n52645 | n52650;
  assign n52652 = ~pi3226 & ~n51802;
  assign n52653 = pi3186 & n52652;
  assign n52654 = ~n15426 & n51802;
  assign po3546 = n52653 | n52654;
  assign n52656 = ~pi3227 & ~n51802;
  assign n52657 = pi2976 & n52656;
  assign n52658 = ~n12061 & n51802;
  assign po3547 = n52657 | n52658;
  assign n52660 = pi3228 & ~n51730;
  assign n52661 = ~pi2023 & n50149;
  assign n52662 = ~pi2032 & ~n50149;
  assign n52663 = ~n52661 & ~n52662;
  assign n52664 = n51730 & ~n52663;
  assign po3548 = n52660 | n52664;
  assign n52666 = pi3229 & ~n51730;
  assign n52667 = ~pi2024 & n50149;
  assign n52668 = ~pi1863 & ~n50149;
  assign n52669 = ~n52667 & ~n52668;
  assign n52670 = n51730 & ~n52669;
  assign po3549 = n52666 | n52670;
  assign n52672 = pi3230 & ~n51730;
  assign n52673 = ~pi2025 & n50149;
  assign n52674 = ~pi2033 & ~n50149;
  assign n52675 = ~n52673 & ~n52674;
  assign n52676 = n51730 & ~n52675;
  assign po3550 = n52672 | n52676;
  assign n52678 = pi3231 & ~n51730;
  assign n52679 = ~pi2026 & n50149;
  assign n52680 = ~pi1968 & ~n50149;
  assign n52681 = ~n52679 & ~n52680;
  assign n52682 = n51730 & ~n52681;
  assign po3551 = n52678 | n52682;
  assign n52684 = pi3232 & ~pi3533;
  assign n52685 = ~pi3487 & ~n52684;
  assign n52686 = ~pi3232 & pi3533;
  assign po3552 = n52685 | n52686;
  assign n52688 = pi3233 & n8561;
  assign n52689 = ~n8561 & ~n37737;
  assign po3553 = n52688 | n52689;
  assign n52691 = pi3234 & ~n51730;
  assign n52692 = ~pi1969 & n50149;
  assign n52693 = ~pi2035 & ~n50149;
  assign n52694 = ~n52692 & ~n52693;
  assign n52695 = n51730 & ~n52694;
  assign po3554 = n52691 | n52695;
  assign n52697 = pi3235 & ~n51730;
  assign n52698 = ~pi2028 & n50149;
  assign n52699 = ~pi2063 & ~n50149;
  assign n52700 = ~n52698 & ~n52699;
  assign n52701 = n51730 & ~n52700;
  assign po3555 = n52697 | n52701;
  assign n52703 = n9373 & n15588;
  assign n52704 = ~n8561 & n52703;
  assign n52705 = po3627 & n52704;
  assign n52706 = ~pi3641 & n52705;
  assign n52707 = pi3236 & n36128;
  assign po3556 = n52706 | n52707;
  assign n52709 = ~pi3237 & ~n51802;
  assign n52710 = pi2974 & n52709;
  assign n52711 = ~n13121 & n51802;
  assign po3557 = n52710 | n52711;
  assign n52713 = ~pi3238 & ~n51802;
  assign n52714 = pi3189 & n52713;
  assign n52715 = ~n12726 & n51802;
  assign po3558 = n52714 | n52715;
  assign n52717 = ~pi3239 & ~n51802;
  assign n52718 = pi2975 & n52717;
  assign n52719 = ~n14816 & n51802;
  assign po3559 = n52718 | n52719;
  assign n52721 = ~pi3240 & n41986;
  assign n52722 = ~pi3240 & pi4005;
  assign n52723 = pi3336 & ~n52722;
  assign n52724 = pi3240 & ~pi4005;
  assign n52725 = ~n52723 & ~n52724;
  assign n52726 = ~n41986 & n52725;
  assign po3560 = n52721 | n52726;
  assign n52728 = ~pi3241 & n41942;
  assign n52729 = pi3241 & ~pi4002;
  assign n52730 = ~pi3241 & pi4002;
  assign n52731 = pi3339 & ~n52730;
  assign n52732 = ~n52729 & ~n52731;
  assign n52733 = ~n41942 & n52732;
  assign po3561 = n52728 | n52733;
  assign n52735 = ~pi3242 & n41953;
  assign n52736 = pi3242 & ~pi4000;
  assign n52737 = ~pi3242 & pi4000;
  assign n52738 = pi3338 & ~n52737;
  assign n52739 = ~n52736 & ~n52738;
  assign n52740 = ~n41953 & n52739;
  assign po3562 = n52735 | n52740;
  assign n52742 = ~pi3243 & n41503;
  assign n52743 = pi3243 & ~pi4004;
  assign n52744 = ~pi3243 & pi4004;
  assign n52745 = pi3342 & ~n52744;
  assign n52746 = ~n52743 & ~n52745;
  assign n52747 = ~n41503 & n52746;
  assign po3563 = n52742 | n52747;
  assign n52749 = ~n8561 & ~n35466;
  assign n52750 = ~pi3244 & n8561;
  assign po3564 = n52749 | n52750;
  assign n52752 = pi3245 & n8561;
  assign n52753 = ~n35887 & ~n52752;
  assign po3565 = po3627 & ~n52753;
  assign n52755 = ~n38723 & ~n38742;
  assign n52756 = n38732 & n52755;
  assign n52757 = pi3266 & n52756;
  assign n52758 = pi3246 & ~n52756;
  assign po3566 = n52757 | n52758;
  assign n52760 = ~pi3247 & ~n42536;
  assign n52761 = ~pi3247 & pi3290;
  assign n52762 = pi3247 & ~pi3290;
  assign n52763 = ~n52761 & ~n52762;
  assign n52764 = n42536 & ~n52763;
  assign po3567 = n52760 | n52764;
  assign n52766 = pi3248 & n8561;
  assign n52767 = ~pi0427 & ~n8561;
  assign n52768 = ~n52766 & ~n52767;
  assign po3568 = ~po3897 & ~n52768;
  assign n52770 = pi3343 & pi3585;
  assign n52771 = pi3281 & n52770;
  assign n52772 = pi3099 & n52771;
  assign n52773 = ~pi3199 & n52772;
  assign n52774 = ~pi2049 & ~pi2759;
  assign po3572 = n52773 & n52774;
  assign n52776 = pi3682 & ~n8307;
  assign n52777 = n8211 & n52776;
  assign n52778 = ~pi3253 & ~n52777;
  assign n52779 = pi3994 & n52777;
  assign po3573 = n52778 | n52779;
  assign n52781 = pi3678 & n52756;
  assign n52782 = pi3255 & ~n52756;
  assign po3575 = n52781 | n52782;
  assign n52784 = ~n8621 & n49693;
  assign po3576 = n9349 | n52784;
  assign n52786 = ~n10762 & n49693;
  assign po3577 = n10766 | n52786;
  assign n52788 = ~pi3258 & ~n52777;
  assign n52789 = pi3692 & n52777;
  assign po3578 = n52788 | n52789;
  assign n52791 = ~pi3259 & ~n52777;
  assign n52792 = pi3691 & n52777;
  assign po3579 = n52791 | n52792;
  assign n52794 = ~pi3260 & ~n52777;
  assign n52795 = pi3686 & n52777;
  assign po3580 = n52794 | n52795;
  assign n52797 = ~pi3261 & ~n52777;
  assign n52798 = pi3992 & n52777;
  assign po3581 = n52797 | n52798;
  assign n52800 = ~pi3262 & ~n52777;
  assign n52801 = pi3684 & n52777;
  assign po3582 = n52800 | n52801;
  assign n52803 = ~pi3263 & ~n52777;
  assign n52804 = pi3989 & n52777;
  assign po3583 = n52803 | n52804;
  assign n52806 = ~pi3264 & ~n52777;
  assign n52807 = pi3987 & n52777;
  assign po3584 = n52806 | n52807;
  assign n52809 = ~pi3265 & ~n52777;
  assign n52810 = pi3693 & n52777;
  assign po3585 = n52809 | n52810;
  assign n52812 = pi3271 & n52756;
  assign n52813 = pi3266 & ~n52756;
  assign po3586 = n52812 | n52813;
  assign n52815 = pi3267 & n8561;
  assign n52816 = ~pi0407 & ~n8561;
  assign n52817 = ~n52815 & ~n52816;
  assign po3587 = ~po3897 & ~n52817;
  assign n52819 = ~pi2193 & ~n8561;
  assign n52820 = ~pi3268 & n8561;
  assign n52821 = ~n52819 & ~n52820;
  assign po3588 = po3627 & n52821;
  assign n52823 = n38253 & n38262;
  assign n52824 = pi3269 & ~n38262;
  assign po3589 = n52823 | n52824;
  assign po3590 = ~pi3424 & ~pi3639;
  assign n52827 = n42751 & ~n42778;
  assign n52828 = n42749 & n42772;
  assign n52829 = ~n42753 & ~n52828;
  assign po3896 = n52827 | ~n52829;
  assign n52831 = pi3647 & po3896;
  assign po3759 = ~pi3588 & n52831;
  assign n52833 = pi1735 & po3759;
  assign po3591 = ~pi3270 | n52833;
  assign n52835 = pi3255 & n52756;
  assign n52836 = pi3271 & ~n52756;
  assign po3592 = n52835 | n52836;
  assign n52838 = ~pi3272 & ~n52777;
  assign n52839 = pi3993 & n52777;
  assign po3593 = n52838 | n52839;
  assign n52841 = ~pi3273 & ~n52777;
  assign n52842 = pi3990 & n52777;
  assign po3594 = n52841 | n52842;
  assign n52844 = ~pi3274 & ~n52777;
  assign n52845 = pi3698 & n52777;
  assign po3595 = n52844 | n52845;
  assign n52847 = ~pi3275 & ~n52777;
  assign n52848 = pi3695 & n52777;
  assign po3596 = n52847 | n52848;
  assign n52850 = ~pi3276 & ~n52777;
  assign n52851 = pi3694 & n52777;
  assign po3597 = n52850 | n52851;
  assign n52853 = ~pi3277 & ~n52777;
  assign n52854 = pi3683 & n52777;
  assign po3598 = n52853 | n52854;
  assign po3599 = ~pi3427 & ~pi3638;
  assign n52857 = n44448 & ~n44475;
  assign n52858 = n44446 & n44469;
  assign n52859 = ~n44450 & ~n52858;
  assign po3879 = n52857 | ~n52859;
  assign n52861 = pi3635 & po3879;
  assign po3746 = ~pi3554 & n52861;
  assign n52863 = pi1444 & po3746;
  assign po3600 = ~pi3278 | n52863;
  assign n52865 = ~pi3279 & ~n52777;
  assign n52866 = pi3696 & n52777;
  assign po3601 = n52865 | n52866;
  assign n52868 = ~pi3280 & ~n52777;
  assign n52869 = pi3697 & n52777;
  assign po3602 = n52868 | n52869;
  assign n52871 = pi3281 & ~n48192;
  assign n52872 = ~pi3281 & pi3343;
  assign n52873 = pi3281 & ~pi3343;
  assign n52874 = ~n52872 & ~n52873;
  assign n52875 = n48192 & ~n52874;
  assign n52876 = ~n52871 & ~n52875;
  assign po3603 = ~n36174 & ~n52876;
  assign n52878 = ~pi3282 & ~n52777;
  assign n52879 = pi3988 & n52777;
  assign po3604 = n52878 | n52879;
  assign n52881 = ~pi3283 & ~n52777;
  assign n52882 = pi3991 & n52777;
  assign po3605 = n52881 | n52882;
  assign n52884 = ~pi3284 & ~n52777;
  assign n52885 = pi3685 & n52777;
  assign po3606 = n52884 | n52885;
  assign n52887 = n15594 & n46577;
  assign n52888 = ~pi1797 & n52887;
  assign n52889 = ~pi3285 & n52888;
  assign po3607 = pi3285 | n52889;
  assign n52891 = ~pi3286 & ~n52777;
  assign n52892 = pi3690 & n52777;
  assign po3608 = n52891 | n52892;
  assign n52894 = ~pi3287 & ~n52777;
  assign n52895 = pi3689 & n52777;
  assign po3609 = n52894 | n52895;
  assign n52897 = ~pi3288 & ~n52777;
  assign n52898 = pi3687 & n52777;
  assign po3610 = n52897 | n52898;
  assign n52900 = ~pi3289 & ~n52777;
  assign n52901 = pi3688 & n52777;
  assign po3611 = n52900 | n52901;
  assign n52903 = ~pi3290 & ~n42536;
  assign n52904 = pi3290 & n42536;
  assign po3612 = n52903 | n52904;
  assign n52906 = pi3291 & n15546;
  assign n52907 = po3831 & po3627;
  assign n52908 = ~pi1823 & n9345;
  assign n52909 = n52907 & n52908;
  assign po3613 = n52906 | n52909;
  assign n52911 = ~n8561 & ~n35482;
  assign n52912 = ~pi3292 & n8561;
  assign po3614 = n52911 | n52912;
  assign n52914 = ~pi0834 & ~n9352;
  assign n52915 = ~n12415 & n52914;
  assign n52916 = pi3293 & ~n52914;
  assign po3615 = n52915 | n52916;
  assign n52918 = po3841 & ~n9352;
  assign n52919 = pi3216 & ~n16904;
  assign n52920 = ~pi3216 & ~n15419;
  assign n52921 = ~n52919 & ~n52920;
  assign n52922 = n52918 & ~n52921;
  assign n52923 = pi3295 & ~n52918;
  assign po3617 = n52922 | n52923;
  assign n52925 = pi3216 & ~n16940;
  assign n52926 = ~pi3216 & ~n10601;
  assign n52927 = ~n52925 & ~n52926;
  assign n52928 = n52918 & ~n52927;
  assign n52929 = pi3296 & ~n52918;
  assign po3618 = n52928 | n52929;
  assign n52931 = pi3216 & ~n16581;
  assign n52932 = ~pi3216 & ~n15088;
  assign n52933 = ~n52931 & ~n52932;
  assign n52934 = n52918 & ~n52933;
  assign n52935 = pi3297 & ~n52918;
  assign po3619 = n52934 | n52935;
  assign n52937 = pi3216 & ~n16725;
  assign n52938 = ~pi3216 & ~n13371;
  assign n52939 = ~n52937 & ~n52938;
  assign n52940 = n52918 & ~n52939;
  assign n52941 = pi3298 & ~n52918;
  assign po3620 = n52940 | n52941;
  assign n52943 = pi3299 & n8561;
  assign n52944 = pi0415 & ~n8561;
  assign n52945 = ~n52943 & ~n52944;
  assign po3621 = ~po3897 & ~n52945;
  assign n52947 = ~pi3301 & n41953;
  assign n52948 = pi3999 & ~n41953;
  assign po3623 = n52947 | n52948;
  assign po3624 = pi3647 & n50482;
  assign n52951 = pi0890 & pi1931;
  assign n52952 = pi3569 & n52951;
  assign po3626 = ~pi3270 | n52952;
  assign n52954 = ~pi0418 & ~n8561;
  assign n52955 = n15550 & n52954;
  assign n52956 = pi3305 & n8561;
  assign po3628 = n52955 | n52956;
  assign n52958 = pi3216 & ~n16832;
  assign n52959 = ~pi3216 & ~n12700;
  assign n52960 = ~n52958 & ~n52959;
  assign n52961 = n52918 & ~n52960;
  assign n52962 = pi3306 & ~n52918;
  assign po3629 = n52961 | n52962;
  assign n52964 = pi3216 & ~n16796;
  assign n52965 = ~pi3216 & ~n13694;
  assign n52966 = ~n52964 & ~n52965;
  assign n52967 = n52918 & ~n52966;
  assign n52968 = pi3307 & ~n52918;
  assign po3630 = n52967 | n52968;
  assign n52970 = pi3216 & ~n16761;
  assign n52971 = ~pi3216 & ~n13114;
  assign n52972 = ~n52970 & ~n52971;
  assign n52973 = n52918 & ~n52972;
  assign n52974 = pi3308 & ~n52918;
  assign po3631 = n52973 | n52974;
  assign n52976 = pi3216 & ~n16689;
  assign n52977 = ~pi3216 & ~n13981;
  assign n52978 = ~n52976 & ~n52977;
  assign n52979 = n52918 & ~n52978;
  assign n52980 = pi3309 & ~n52918;
  assign po3632 = n52979 | n52980;
  assign n52982 = pi3216 & ~n16653;
  assign n52983 = ~pi3216 & ~n12408;
  assign n52984 = ~n52982 & ~n52983;
  assign n52985 = n52918 & ~n52984;
  assign n52986 = pi3310 & ~n52918;
  assign po3633 = n52985 | n52986;
  assign n52988 = pi3216 & ~n16617;
  assign n52989 = ~pi3216 & ~n14809;
  assign n52990 = ~n52988 & ~n52989;
  assign n52991 = n52918 & ~n52990;
  assign n52992 = pi3311 & ~n52918;
  assign po3634 = n52991 | n52992;
  assign n52994 = pi3216 & ~n16545;
  assign n52995 = ~pi3216 & ~n12034;
  assign n52996 = ~n52994 & ~n52995;
  assign n52997 = n52918 & ~n52996;
  assign n52998 = pi3312 & ~n52918;
  assign po3635 = n52997 | n52998;
  assign n53000 = pi3216 & ~n17374;
  assign n53001 = ~pi3216 & ~n17341;
  assign n53002 = ~n53000 & ~n53001;
  assign n53003 = n52918 & ~n53002;
  assign n53004 = pi3313 & ~n52918;
  assign po3636 = n53003 | n53004;
  assign n53006 = pi3216 & ~n17082;
  assign n53007 = ~pi3216 & ~n17172;
  assign n53008 = ~n53006 & ~n53007;
  assign n53009 = n52918 & ~n53008;
  assign n53010 = pi3314 & ~n52918;
  assign po3637 = n53009 | n53010;
  assign n53012 = pi3216 & ~n16868;
  assign n53013 = ~pi3216 & ~n14396;
  assign n53014 = ~n53012 & ~n53013;
  assign n53015 = n52918 & ~n53014;
  assign n53016 = pi3315 & ~n52918;
  assign po3638 = n53015 | n53016;
  assign n53018 = pi3216 & ~n16470;
  assign n53019 = ~pi3216 & ~n11174;
  assign n53020 = ~n53018 & ~n53019;
  assign n53021 = n52918 & ~n53020;
  assign n53022 = pi3316 & ~n52918;
  assign po3639 = n53021 | n53022;
  assign n53024 = ~pi3317 & n41503;
  assign po3640 = n41504 | n53024;
  assign n53026 = ~pi3318 & n41503;
  assign po3641 = n41933 | n53026;
  assign n53028 = ~pi3319 & n41964;
  assign n53029 = ~pi3222 & ~n41964;
  assign po3642 = n53028 | n53029;
  assign n53031 = ~pi3320 & n41975;
  assign po3643 = n41976 | n53031;
  assign n53033 = ~pi3321 & n41975;
  assign n53034 = ~pi3225 & ~n41975;
  assign po3644 = n53033 | n53034;
  assign n53036 = ~pi3325 & n41964;
  assign n53037 = pi3998 & ~n41964;
  assign po3648 = n53036 | n53037;
  assign n53039 = pi3326 & n8561;
  assign n53040 = pi0414 & ~n8561;
  assign n53041 = ~n53039 & ~n53040;
  assign po3649 = ~po3897 & ~n53041;
  assign n53043 = ~pi3327 & n41964;
  assign n53044 = pi3997 & ~n41964;
  assign po3650 = n53043 | n53044;
  assign n53046 = ~n15115 & n52914;
  assign n53047 = pi3328 & ~n52914;
  assign po3651 = n53046 | n53047;
  assign n53049 = ~n8561 & n36075;
  assign n53050 = pi3329 & n8561;
  assign po3652 = n53049 | n53050;
  assign n53052 = ~pi3330 & n8561;
  assign po3653 = n52816 | n53052;
  assign n53054 = pi1930 & ~n9352;
  assign n53055 = pi3402 & n53054;
  assign n53056 = pi3331 & ~n53054;
  assign po3654 = n53055 | n53056;
  assign n53058 = pi3400 & n53054;
  assign n53059 = pi3332 & ~n53054;
  assign po3655 = n53058 | n53059;
  assign n53061 = ~pi3333 & n41975;
  assign n53062 = pi3995 & ~n41975;
  assign po3656 = n53061 | n53062;
  assign n53064 = ~pi3334 & n41975;
  assign n53065 = pi3996 & ~n41975;
  assign po3657 = n53064 | n53065;
  assign n53067 = ~pi3335 & n41986;
  assign n53068 = pi4006 & ~n41986;
  assign po3658 = n53067 | n53068;
  assign n53070 = ~pi3336 & n41986;
  assign n53071 = pi4005 & ~n41986;
  assign po3659 = n53070 | n53071;
  assign n53073 = ~pi3337 & n50163;
  assign n53074 = ~pi3337 & pi3389;
  assign n53075 = pi3337 & ~pi3389;
  assign n53076 = ~n53074 & ~n53075;
  assign n53077 = ~n50163 & ~n53076;
  assign po3660 = n53073 | n53077;
  assign n53079 = ~pi3338 & n41953;
  assign n53080 = pi4000 & ~n41953;
  assign po3661 = n53079 | n53080;
  assign n53082 = ~pi3339 & n41942;
  assign n53083 = pi4002 & ~n41942;
  assign po3662 = n53082 | n53083;
  assign n53085 = ~pi3340 & n41986;
  assign n53086 = ~pi3240 & ~n41986;
  assign po3663 = n53085 | n53086;
  assign n53088 = ~pi3341 & n41942;
  assign n53089 = pi4001 & ~n41942;
  assign po3664 = n53088 | n53089;
  assign n53091 = ~pi3342 & n41503;
  assign n53092 = pi4004 & ~n41503;
  assign po3665 = n53091 | n53092;
  assign n53094 = ~pi3343 & ~n48192;
  assign n53095 = pi3343 & n48192;
  assign n53096 = ~n53094 & ~n53095;
  assign po3666 = ~n36174 & n53096;
  assign n53098 = pi3344 & n8561;
  assign n53099 = ~n36558 & ~n53098;
  assign po3667 = po3627 & ~n53099;
  assign n53101 = ~pi3345 & n41953;
  assign n53102 = ~pi3221 & ~n41953;
  assign po3668 = n53101 | n53102;
  assign n53104 = ~pi3346 & n41953;
  assign po3669 = n41954 | n53104;
  assign n53106 = pi3403 & n53054;
  assign n53107 = pi3347 & ~n53054;
  assign po3670 = n53106 | n53107;
  assign n53109 = ~pi3348 & n41964;
  assign po3671 = n41965 | n53109;
  assign n53111 = ~pi3349 & n41942;
  assign n53112 = ~pi3220 & ~n41942;
  assign po3672 = n53111 | n53112;
  assign n53114 = pi3682 & n8388;
  assign n53115 = pi3350 & ~n53114;
  assign po3934 = ~pi3682 | ~n48401;
  assign po3673 = n53115 | ~po3934;
  assign n53118 = ~pi3351 & n41942;
  assign po3674 = n41943 | n53118;
  assign n53120 = pi3404 & n53054;
  assign n53121 = pi3352 & ~n53054;
  assign po3675 = n53120 | n53121;
  assign n53123 = po0279 & n53054;
  assign n53124 = pi3353 & ~n53054;
  assign po3676 = n53123 | n53124;
  assign n53126 = pi3414 & n53054;
  assign n53127 = pi3354 & ~n53054;
  assign po3677 = n53126 | n53127;
  assign n53129 = po0278 & n53054;
  assign n53130 = pi3355 & ~n53054;
  assign po3678 = n53129 | n53130;
  assign n53132 = ~pi3356 & n41503;
  assign n53133 = pi4003 & ~n41503;
  assign po3679 = n53132 | n53133;
  assign n53135 = ~pi3357 & n41986;
  assign po3680 = n41987 | n53135;
  assign n53137 = pi3216 & ~n16976;
  assign n53138 = ~pi3216 & ~n9762;
  assign n53139 = ~n53137 & ~n53138;
  assign n53140 = n52918 & ~n53139;
  assign n53141 = pi3358 & ~n52918;
  assign po3681 = n53140 | n53141;
  assign n53143 = ~n8567 & ~n10777;
  assign n53144 = n10767 & ~n53143;
  assign po3682 = n15504 & ~n53144;
  assign n53146 = pi3360 & ~n52914;
  assign n53147 = ~n12061 & n52914;
  assign po3683 = n53146 | n53147;
  assign n53149 = pi3361 & ~n52914;
  assign n53150 = ~n11181 & n52914;
  assign po3684 = n53149 | n53150;
  assign po3686 = n15508 & ~n53144;
  assign po3687 = n15513 & ~n53144;
  assign po3688 = n15515 & ~n53144;
  assign n53155 = ~n8567 & ~n8595;
  assign n53156 = n9350 & ~n53155;
  assign po3689 = n10699 & ~n53156;
  assign n53158 = ~n8561 & n9381;
  assign n53159 = pi3367 & n8561;
  assign po3690 = n53158 | n53159;
  assign po3691 = n10709 & ~n53156;
  assign po3692 = n10704 & ~n53156;
  assign n53163 = pi3370 & ~pi3481;
  assign n53164 = n9352 & n53163;
  assign n53165 = pi3216 & ~n9352;
  assign po3693 = n53164 | n53165;
  assign n53167 = ~pi0540 & ~n9352;
  assign n53168 = ~pi3371 & n9352;
  assign n53169 = ~n53167 & ~n53168;
  assign po3694 = po3627 & n53169;
  assign po3695 = ~n17199 & n51802;
  assign po3696 = ~n9825 & n51802;
  assign po3697 = ~n10608 & n51802;
  assign po3698 = ~n17368 & n51802;
  assign n53175 = pi0796 & pi2111;
  assign n53176 = pi3570 & n53175;
  assign po3699 = ~pi3278 | n53176;
  assign n53178 = ~pi1771 & ~pi3377;
  assign n53179 = ~pi0491 & n53178;
  assign po3700 = n35295 | n53179;
  assign n53181 = pi3378 & ~pi3481;
  assign n53182 = n9352 & n53181;
  assign po3701 = n38276 | n53182;
  assign po3702 = n10717 & ~n53156;
  assign po3703 = n10715 & ~n53156;
  assign po3704 = n10713 & ~n53156;
  assign po3705 = po1234 & n50163;
  assign n53188 = pi3382 & ~pi3410;
  assign po3706 = pi3481 & ~n53188;
  assign po3707 = n10702 & ~n53156;
  assign po3708 = n10696 & ~n53156;
  assign po3709 = n15511 & ~n53144;
  assign po3710 = n15502 & ~n53144;
  assign po3711 = n15497 & ~n53144;
  assign po3712 = n15463 & ~n53144;
  assign n53196 = ~pi3389 & n50163;
  assign n53197 = pi3389 & ~n50163;
  assign po3713 = n53196 | n53197;
  assign n53199 = ~n8561 & n15550;
  assign n53200 = pi3390 & n8561;
  assign po3714 = n53199 | n53200;
  assign n53202 = ~n8561 & ~n9384;
  assign n53203 = pi3391 & n8561;
  assign po3715 = n53202 | n53203;
  assign n53205 = pi3392 & n8561;
  assign po3716 = n52944 | n53205;
  assign n53207 = pi3393 & n8561;
  assign n53208 = pi0419 & ~n8561;
  assign po3717 = n53207 | n53208;
  assign n53210 = ~pi3394 & n8561;
  assign po3718 = n52767 | n53210;
  assign n53212 = pi3395 & n8627;
  assign n53213 = ~n17561 & ~n53212;
  assign po3720 = ~pi3395 & ~n53213;
  assign n53215 = pi3396 & n8561;
  assign n53216 = pi0420 & ~n8561;
  assign po3721 = n53215 | n53216;
  assign n53218 = pi3397 & ~pi3583;
  assign n53219 = pi3481 & n53218;
  assign po3722 = n50167 | n53219;
  assign n53221 = pi3398 & n8561;
  assign po3723 = n53040 | n53221;
  assign po3724 = n15494 & ~n53144;
  assign n53224 = pi2516 & po3831;
  assign n53225 = pi3400 & ~po3831;
  assign po3725 = n53224 | n53225;
  assign n53227 = pi3401 & ~po3831;
  assign n53228 = pi2517 & po3831;
  assign po3726 = n53227 | n53228;
  assign n53230 = pi2482 & po3831;
  assign n53231 = pi3402 & ~po3831;
  assign po3727 = n53230 | n53231;
  assign n53233 = pi2483 & po3831;
  assign n53234 = pi3403 & ~po3831;
  assign po3728 = n53233 | n53234;
  assign n53236 = pi2481 & po3831;
  assign n53237 = pi3404 & ~po3831;
  assign po3729 = n53236 | n53237;
  assign n53239 = pi3405 & ~po3831;
  assign n53240 = pi2479 & po3831;
  assign po3730 = n53239 | n53240;
  assign n53242 = pi3406 & ~po3831;
  assign n53243 = pi2477 & po3831;
  assign po3731 = n53242 | n53243;
  assign po3732 = pi3407 & ~n52914;
  assign n53246 = ~n9342 & ~n9352;
  assign n53247 = pi3408 & n9352;
  assign po3733 = n53246 | n53247;
  assign n53249 = ~pi0783 & ~po3627;
  assign po3734 = ~po0493 | n53249;
  assign n53251 = pi3411 & ~po3831;
  assign n53252 = pi2476 & po3831;
  assign po3737 = n53251 | n53252;
  assign n53254 = ~n8623 & ~n10744;
  assign n53255 = ~n9352 & ~n53254;
  assign n53256 = pi3412 & n9352;
  assign po3738 = n53255 | n53256;
  assign n53258 = pi3413 & ~po3831;
  assign n53259 = pi2478 & po3831;
  assign po3739 = n53258 | n53259;
  assign n53261 = pi2480 & po3831;
  assign n53262 = pi3414 & ~po3831;
  assign po3740 = n53261 | n53262;
  assign n53264 = ~pi0936 & pi3415;
  assign n53265 = pi2492 & ~pi3415;
  assign po3742 = n53264 | n53265;
  assign n53267 = ~pi1046 & pi3481;
  assign n53268 = pi3416 & n53267;
  assign n53269 = ~pi3398 & ~pi3481;
  assign n53270 = po3850 & n53269;
  assign po3744 = n53268 | n53270;
  assign n53272 = n8577 & ~n8628;
  assign po3747 = ~pi3419 & n53272;
  assign n53274 = pi3420 & ~po3831;
  assign n53275 = pi2475 & po3831;
  assign po3748 = n53274 | n53275;
  assign n53277 = pi3421 & ~po3831;
  assign n53278 = pi2485 & po3831;
  assign po3749 = n53277 | n53278;
  assign n53280 = pi3422 & ~po3831;
  assign n53281 = pi2518 & po3831;
  assign po3750 = n53280 | n53281;
  assign n53283 = ~pi1930 & pi3423;
  assign n53284 = po0290 & po0307;
  assign n53285 = pi1930 & ~n53284;
  assign po3751 = n53283 | n53285;
  assign n53287 = ~pi3424 & n8627;
  assign n53288 = ~n8627 & ~n9420;
  assign n53289 = ~n53287 & ~n53288;
  assign po3752 = ~pi3424 & n53289;
  assign po3753 = po0767 & ~n38723;
  assign n53292 = pi3426 & n8561;
  assign n53293 = ~n8561 & ~n9345;
  assign po3754 = n53292 | n53293;
  assign n53295 = ~pi3427 & n8627;
  assign n53296 = ~n8568 & ~n8627;
  assign n53297 = ~n53295 & ~n53296;
  assign po3755 = ~pi3427 & n53297;
  assign n53299 = pi3428 & n8589;
  assign n53300 = pi3641 & n8628;
  assign po3756 = n53299 & ~n53300;
  assign n53302 = ~pi3429 & n8627;
  assign n53303 = ~n8627 & ~n9419;
  assign n53304 = ~n53302 & ~n53303;
  assign po3757 = ~pi3429 & n53304;
  assign n53306 = pi3430 & ~po3831;
  assign n53307 = pi2484 & po3831;
  assign po3758 = n53306 | n53307;
  assign n53309 = ~n15546 & ~n19018;
  assign n53310 = pi3432 & n15546;
  assign po3760 = n53309 | n53310;
  assign n53312 = ~n15546 & ~n18737;
  assign n53313 = pi3434 & n15546;
  assign po3762 = n53312 | n53313;
  assign n53315 = pi3435 & ~po3841;
  assign n53316 = po3841 & ~n9440;
  assign po3763 = n53315 | n53316;
  assign n53318 = pi3436 & ~po3841;
  assign n53319 = po3841 & ~n9433;
  assign po3764 = n53318 | n53319;
  assign n53321 = pi1908 & pi3415;
  assign po3769 = pi2492 & n53321;
  assign n53323 = ~pi3674 & pi3708;
  assign n53324 = ~pi3445 & pi3674;
  assign po3773 = n53323 | n53324;
  assign n53326 = ~pi3674 & pi3702;
  assign n53327 = ~pi3446 & pi3674;
  assign po3774 = n53326 | n53327;
  assign n53329 = ~pi3674 & pi3711;
  assign n53330 = ~pi3447 & pi3674;
  assign po3775 = n53329 | n53330;
  assign n53332 = ~pi3674 & pi3709;
  assign n53333 = ~pi3448 & pi3674;
  assign po3776 = n53332 | n53333;
  assign n53335 = pi3449 & po3934;
  assign n53336 = po0242 & ~po3934;
  assign po3777 = n53335 | n53336;
  assign n53338 = ~n15546 & ~n16110;
  assign n53339 = pi3450 & n15546;
  assign po3778 = n53338 | n53339;
  assign n53341 = po3841 & ~n9447;
  assign n53342 = pi3451 & ~po3841;
  assign po3779 = n53341 | n53342;
  assign n53344 = ~po3852 & ~po3849;
  assign po3780 = pi3148 & n53344;
  assign n53346 = ~n15546 & ~n18950;
  assign n53347 = pi3453 & n15546;
  assign po3781 = n53346 | n53347;
  assign n53349 = ~n15546 & ~n18882;
  assign n53350 = pi3454 & n15546;
  assign po3782 = n53349 | n53350;
  assign n53352 = ~n15546 & ~n18807;
  assign n53353 = pi3455 & n15546;
  assign po3783 = n53352 | n53353;
  assign n53355 = ~n15546 & ~n16025;
  assign n53356 = pi3458 & n15546;
  assign po3786 = n53355 | n53356;
  assign n53358 = ~n15546 & ~n19087;
  assign n53359 = pi3459 & n15546;
  assign po3787 = n53358 | n53359;
  assign n53361 = pi3473 & po3896;
  assign n53362 = pi2576 & ~po3896;
  assign po3789 = n53361 | n53362;
  assign n53364 = ~pi3674 & pi3701;
  assign n53365 = ~pi3462 & pi3674;
  assign po3790 = n53364 | n53365;
  assign n53367 = ~pi3674 & pi3710;
  assign n53368 = ~pi3463 & pi3674;
  assign po3791 = n53367 | n53368;
  assign n53370 = ~pi3674 & pi3699;
  assign n53371 = ~pi3464 & pi3674;
  assign po3792 = n53370 | n53371;
  assign n53373 = ~pi3674 & pi3713;
  assign n53374 = ~pi3465 & pi3674;
  assign po3793 = n53373 | n53374;
  assign n53376 = ~pi3674 & pi3712;
  assign n53377 = ~pi3466 & pi3674;
  assign po3794 = n53376 | n53377;
  assign n53379 = ~pi3674 & pi3714;
  assign n53380 = ~pi3467 & pi3674;
  assign po3795 = n53379 | n53380;
  assign n53382 = ~pi3674 & pi3700;
  assign n53383 = ~pi3468 & pi3674;
  assign po3796 = n53382 | n53383;
  assign n53385 = ~pi3674 & pi3703;
  assign n53386 = ~pi3470 & pi3674;
  assign po3798 = n53385 | n53386;
  assign n53388 = ~pi3597 & po3896;
  assign n53389 = pi2578 & ~po3896;
  assign po3799 = n53388 | n53389;
  assign n53391 = pi3471 & po3896;
  assign n53392 = pi2577 & ~po3896;
  assign po3801 = n53391 | n53392;
  assign n53394 = ~pi3674 & pi3707;
  assign n53395 = ~pi3474 & pi3674;
  assign po3802 = n53394 | n53395;
  assign n53397 = ~pi3674 & pi3704;
  assign n53398 = ~pi3475 & pi3674;
  assign po3803 = n53397 | n53398;
  assign n53400 = ~pi3674 & pi3705;
  assign n53401 = ~pi3476 & pi3674;
  assign po3804 = n53400 | n53401;
  assign n53403 = ~pi3674 & pi3706;
  assign n53404 = ~pi3477 & pi3674;
  assign po3805 = n53403 | n53404;
  assign n53406 = ~n15546 & ~n19160;
  assign n53407 = pi3478 & n15546;
  assign po3806 = n53406 | n53407;
  assign po3807 = ~po3627 | ~po0493;
  assign n53410 = ~pi3505 & ~pi3524;
  assign po3809 = pi3515 & ~n53410;
  assign n53412 = pi3489 & po3934;
  assign n53413 = po0236 & ~po3934;
  assign po3815 = n53412 | n53413;
  assign n53415 = pi3491 & po3934;
  assign n53416 = po0239 & ~po3934;
  assign po3817 = n53415 | n53416;
  assign n53418 = pi3492 & po3934;
  assign n53419 = po0237 & ~po3934;
  assign po3818 = n53418 | n53419;
  assign n53421 = pi3494 & po3934;
  assign n53422 = po0240 & ~po3934;
  assign po3820 = n53421 | n53422;
  assign n53424 = pi3495 & po3934;
  assign n53425 = po0232 & ~po3934;
  assign po3821 = n53424 | n53425;
  assign n53427 = pi3496 & po3934;
  assign n53428 = po0230 & ~po3934;
  assign po3822 = n53427 | n53428;
  assign n53430 = pi3497 & po3934;
  assign n53431 = po0231 & ~po3934;
  assign po3823 = n53430 | n53431;
  assign n53433 = pi3498 & po3934;
  assign n53434 = po0241 & ~po3934;
  assign po3824 = n53433 | n53434;
  assign n53436 = pi3499 & po3934;
  assign n53437 = po0234 & ~po3934;
  assign po3825 = n53436 | n53437;
  assign n53439 = pi3500 & po3934;
  assign n53440 = po0233 & ~po3934;
  assign po3826 = n53439 | n53440;
  assign n53442 = pi3501 & po3934;
  assign n53443 = po0238 & ~po3934;
  assign po3827 = n53442 | n53443;
  assign po3828 = po0767 & ~n38732;
  assign n53446 = pi3503 & po3934;
  assign n53447 = po0235 & ~po3934;
  assign po3829 = n53446 | n53447;
  assign po3832 = po0767 & ~n38742;
  assign po3833 = ~pi3673 & ~pi3674;
  assign n53451 = po3646 & ~po3616;
  assign n53452 = n48403 & n53451;
  assign n53453 = n8374 & n48400;
  assign n53454 = ~n53452 & ~n53453;
  assign n53455 = n48400 & n53451;
  assign po3894 = ~n53454 | n53455;
  assign n53457 = pi1897 & ~po3879;
  assign n53458 = ~pi3593 & po3879;
  assign po3900 = n53457 | n53458;
  assign n53460 = pi1866 & ~po3879;
  assign n53461 = pi3594 & po3879;
  assign po3901 = n53460 | n53461;
  assign n53463 = pi1743 & ~po3879;
  assign n53464 = pi3595 & po3879;
  assign po3902 = n53463 | n53464;
  assign n53466 = pi1744 & ~po3879;
  assign n53467 = pi3596 & po3879;
  assign po3903 = n53466 | n53467;
  assign n53469 = pi1714 & ~po3879;
  assign n53470 = pi3598 & po3879;
  assign po3904 = n53469 | n53470;
  assign n53472 = pi2579 & ~po3896;
  assign n53473 = pi3600 & po3896;
  assign po3905 = n53472 | n53473;
  assign n53475 = pi1745 & ~po3879;
  assign n53476 = pi3599 & po3879;
  assign po3906 = n53475 | n53476;
  assign n53478 = pi1742 & ~po3879;
  assign n53479 = pi3601 & po3879;
  assign po3907 = n53478 | n53479;
  assign n53481 = pi2580 & ~po3896;
  assign n53482 = pi3602 & po3896;
  assign po3908 = n53481 | n53482;
  assign n53484 = pi1741 & ~po3879;
  assign n53485 = pi3603 & po3879;
  assign po3909 = n53484 | n53485;
  assign n53487 = pi2581 & ~po3896;
  assign n53488 = pi3604 & po3896;
  assign po3910 = n53487 | n53488;
  assign n53490 = pi1867 & ~po3879;
  assign n53491 = pi3605 & po3879;
  assign po3911 = n53490 | n53491;
  assign n53493 = pi2768 & ~po3896;
  assign n53494 = pi3606 & po3896;
  assign po3912 = n53493 | n53494;
  assign n53496 = pi0368 & ~po3879;
  assign n53497 = pi3607 & po3879;
  assign po3913 = n53496 | n53497;
  assign n53499 = pi2568 & ~po3896;
  assign n53500 = pi3608 & po3896;
  assign po3914 = n53499 | n53500;
  assign n53502 = pi0314 & ~po3879;
  assign n53503 = pi3609 & po3879;
  assign po3915 = n53502 | n53503;
  assign n53505 = pi2569 & ~po3896;
  assign n53506 = pi3610 & po3896;
  assign po3916 = n53505 | n53506;
  assign n53508 = pi0330 & ~po3879;
  assign n53509 = pi3611 & po3879;
  assign po3917 = n53508 | n53509;
  assign n53511 = pi2570 & ~po3896;
  assign n53512 = pi3612 & po3896;
  assign po3918 = n53511 | n53512;
  assign n53514 = pi0072 & ~po3879;
  assign n53515 = pi3613 & po3879;
  assign po3919 = n53514 | n53515;
  assign n53517 = pi2571 & ~po3896;
  assign n53518 = pi3614 & po3896;
  assign po3920 = n53517 | n53518;
  assign n53520 = pi0127 & ~po3879;
  assign n53521 = pi3615 & po3879;
  assign po3921 = n53520 | n53521;
  assign n53523 = pi2572 & ~po3896;
  assign n53524 = pi3616 & po3896;
  assign po3922 = n53523 | n53524;
  assign n53526 = pi0073 & ~po3879;
  assign n53527 = pi3618 & po3879;
  assign po3923 = n53526 | n53527;
  assign n53529 = pi2573 & ~po3896;
  assign n53530 = pi3617 & po3896;
  assign po3924 = n53529 | n53530;
  assign n53532 = pi2574 & ~po3896;
  assign n53533 = pi3619 & po3896;
  assign po3925 = n53532 | n53533;
  assign po3926 = pi0128 & ~po3879;
  assign n53536 = pi2575 & ~po3896;
  assign n53537 = pi3623 & po3896;
  assign po3927 = n53536 | n53537;
  assign n53539 = n8390 & n48404;
  assign n53540 = pi2795 & n8375;
  assign n53541 = pi2789 & n8375;
  assign n53542 = ~pi2789 & ~pi2795;
  assign n53543 = n8196 & ~n53542;
  assign n53544 = ~n53541 & ~n53543;
  assign po3933 = n53540 | ~n53544;
  assign n53546 = n8211 & n8390;
  assign n53547 = ~po3933 & ~n53546;
  assign n53548 = pi3216 & n8232;
  assign n53549 = pi3216 & n8381;
  assign po3932 = n53548 | n53549;
  assign n53551 = n53547 & ~po3932;
  assign po3928 = n53539 | ~n53551;
  assign n53553 = ~n8390 & n48404;
  assign n53554 = pi2779 & n8375;
  assign n53555 = ~n53553 & ~n53554;
  assign n53556 = pi3257 & n8375;
  assign n53557 = pi3256 & n8381;
  assign n53558 = ~n53556 & ~n53557;
  assign n53559 = n53555 & n53558;
  assign n53560 = ~n53455 & n53559;
  assign n53561 = pi3099 & n53455;
  assign po3929 = n53560 | n53561;
  assign n53563 = ~n53540 & ~n53541;
  assign n53564 = ~n53549 & n53563;
  assign po3930 = ~n53539 & n53564;
  assign po3931 = pi2582 & ~po3896;
  assign n53567 = pi0565 & pi3362;
  assign n53568 = ~pi2813 & pi3528;
  assign po3947 = n53567 | n53568;
  assign n53570 = ~po3878 & ~po3947;
  assign n53571 = pi3641 & ~n53570;
  assign n53572 = ~n44985 & ~n53571;
  assign n53573 = ~n44984 & n53572;
  assign po3938 = n36128 & ~n53573;
  assign po3939 = n38798 | n38800;
  assign po3940 = pi2143 | po3897;
  assign n53577 = ~pi0044 & ~pi0048;
  assign n53578 = ~pi0057 & n53577;
  assign n53579 = ~pi0043 & n53578;
  assign n53580 = ~pi0061 & n53579;
  assign n53581 = ~pi0083 & n53580;
  assign n53582 = ~pi0082 & n53581;
  assign n53583 = ~pi0084 & n53582;
  assign n53584 = ~pi0060 & n53583;
  assign n53585 = pi0044 & pi0057;
  assign n53586 = pi0048 & n53585;
  assign n53587 = pi0043 & pi0084;
  assign n53588 = pi0060 & n53587;
  assign n53589 = n53586 & n53588;
  assign n53590 = pi0083 & n53589;
  assign n53591 = pi0061 & n53590;
  assign n53592 = pi0082 & n53591;
  assign n53593 = ~n53584 & ~n53592;
  assign n53594 = pi3138 & n53593;
  assign n53595 = ~pi1025 & ~n53594;
  assign po3941 = ~po3897 & ~n53595;
  assign po3949 = ~pi3672 & ~pi3674;
  assign po0053 = 1'b1;
  assign po0054 = 1'b1;
  assign po0055 = 1'b1;
  assign po0056 = 1'b1;
  assign po0057 = 1'b1;
  assign po0058 = 1'b1;
  assign po0059 = 1'b1;
  assign po0060 = 1'b1;
  assign po0071 = 1'b1;
  assign po0072 = 1'b1;
  assign po0073 = 1'b1;
  assign po0074 = 1'b1;
  assign po0075 = 1'b1;
  assign po0076 = 1'b1;
  assign po0077 = 1'b1;
  assign po0078 = 1'b1;
  assign po0079 = 1'b1;
  assign po0090 = 1'b1;
  assign po0091 = 1'b1;
  assign po0092 = 1'b1;
  assign po0093 = 1'b1;
  assign po0094 = 1'b1;
  assign po0095 = 1'b1;
  assign po0096 = 1'b1;
  assign po0097 = 1'b1;
  assign po0098 = 1'b1;
  assign po0292 = 1'b1;
  assign po0000 = ~po3853;
  assign po0012 = ~pi3452;
  assign po0024 = ~pi3350;
  assign po0757 = ~pi3589;
  assign po0770 = ~po0739;
  assign po0779 = ~po0896;
  assign po0886 = ~pi3639;
  assign po0888 = ~pi3638;
  assign po1115 = ~pi3556;
  assign po1123 = ~pi3587;
  assign po3460 = ~pi3300;
  assign po3463 = ~pi3303;
  assign po3736 = ~pi3382;
  assign po3766 = ~pi3472;
  assign po3767 = ~pi3469;
  assign po3770 = ~pi3537;
  assign po3771 = ~pi3536;
  assign po3797 = ~pi1882;
  assign po3800 = ~pi2099;
  assign po3810 = ~pi3571;
  assign po3851 = ~po0767;
  assign po3856 = ~pi0582;
  assign po3857 = ~pi3660;
  assign po3858 = ~pi3657;
  assign po3859 = ~pi3658;
  assign po3860 = ~pi3659;
  assign po3861 = ~pi0581;
  assign po3862 = ~pi3661;
  assign po3863 = ~pi3656;
  assign po3864 = ~pi3214;
  assign po3865 = ~pi1596;
  assign po3866 = ~pi3200;
  assign po3867 = ~pi3213;
  assign po3868 = ~pi3232;
  assign po3869 = ~pi3212;
  assign po3870 = ~pi3662;
  assign po3875 = ~pi2399;
  assign po3876 = ~pi2387;
  assign po3877 = ~pi3098;
  assign po3880 = ~po0493;
  assign po3951 = ~pi3676;
  assign po0001 = po0000;
  assign po0002 = po0000;
  assign po0003 = po0000;
  assign po0004 = po0000;
  assign po0005 = po0000;
  assign po0006 = po0000;
  assign po0007 = po0000;
  assign po0008 = po0000;
  assign po0010 = pi3397;
  assign po0016 = pi3626;
  assign po0019 = pi3621;
  assign po0025 = pi3627;
  assign po0029 = pi0959;
  assign po0031 = pi0887;
  assign po0033 = pi0941;
  assign po0035 = pi0792;
  assign po0037 = pi0790;
  assign po0039 = pi0738;
  assign po0040 = pi1771;
  assign po0042 = pi3648;
  assign po0178 = pi1769;
  assign po0179 = pi1767;
  assign po0180 = pi1766;
  assign po0181 = pi1858;
  assign po0182 = pi1765;
  assign po0183 = pi1764;
  assign po0184 = pi1763;
  assign po0185 = pi1857;
  assign po0186 = pi1762;
  assign po0187 = pi1761;
  assign po0188 = pi1854;
  assign po0189 = pi1768;
  assign po0190 = pi1103;
  assign po0191 = pi1023;
  assign po0192 = pi1101;
  assign po0193 = pi1022;
  assign po0194 = pi1100;
  assign po0195 = pi1021;
  assign po0196 = pi1099;
  assign po0197 = pi1020;
  assign po0198 = pi1019;
  assign po0199 = pi0974;
  assign po0200 = pi1102;
  assign po0201 = pi1024;
  assign po0273 = pi3400;
  assign po0274 = pi3403;
  assign po0275 = pi3402;
  assign po0276 = pi3404;
  assign po0277 = pi3414;
  assign po0676 = pi3561;
  assign po0769 = pi3647;
  assign po0778 = pi3635;
  assign po0786 = pi3584;
  assign po0793 = pi3558;
  assign po0806 = pi3483;
  assign po0867 = pi0635;
  assign po0868 = pi0633;
  assign po0898 = pi3479;
  assign po0974 = pi3482;
  assign po0978 = pi3525;
  assign po0980 = pi3562;
  assign po1023 = pi3676;
  assign po1280 = pi0979;
  assign po1402 = pi1641;
  assign po1770 = pi3409;
  assign po1950 = pi1875;
  assign po2080 = pi3557;
  assign po2879 = pi3137;
  assign po2882 = pi3142;
  assign po2915 = pi3129;
  assign po3416 = pi3527;
  assign po3461 = pi3254;
  assign po3464 = pi3205;
  assign po3622 = pi3418;
  assign po3625 = pi3431;
  assign po3719 = pi3555;
  assign po3735 = pi1609;
  assign po3761 = po0270;
  assign po3765 = po0269;
  assign po3768 = pi3507;
  assign po3772 = pi0827;
  assign po3784 = po0272;
  assign po3785 = po0271;
  assign po3788 = po0268;
  assign po3808 = pi3549;
  assign po3811 = pi3531;
  assign po3812 = pi3532;
  assign po3813 = pi3533;
  assign po3814 = pi3534;
  assign po3816 = pi3544;
  assign po3819 = pi3550;
  assign po3854 = pi3551;
  assign po3881 = pi2385;
  assign po3883 = pi1931;
  assign po3884 = pi2111;
  assign po3885 = pi0939;
  assign po3886 = pi3645;
  assign po3887 = pi3679;
  assign po3888 = pi3674;
  assign po3889 = pi3675;
  assign po3890 = pi3673;
  assign po3891 = pi3672;
  assign po3892 = pi0565;
  assign po3895 = pi3591;
  assign po3898 = pi3585;
  assign po3899 = pi0936;
  assign po3935 = pi3629;
  assign po3936 = pi3630;
  assign po3942 = pi3637;
  assign po3944 = pi3640;
  assign po3952 = pi0853;
endmodule


