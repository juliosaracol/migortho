module pci_spoci_ctrl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21, pi22, pi23,
    pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47,
    pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81, pi82, pi83,
    pi84,
    po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10, po11,
    po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22, po23,
    po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46, po47,
    po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19, pi20, pi21,
    pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33,
    pi34, pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44, pi45,
    pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57,
    pi58, pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80, pi81,
    pi82, pi83, pi84;
  output po00, po01, po02, po03, po04, po05, po06, po07, po08, po09, po10,
    po11, po12, po13, po14, po15, po16, po17, po18, po19, po20, po21, po22,
    po23, po24, po25, po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43, po44, po45, po46,
    po47, po48, po49, po50, po51, po52, po53, po54, po55, po56, po57, po58,
    po59, po60, po61, po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75;
  wire n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
    n331, n332, n333, n335, n336, n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411, n412, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n485, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522, n524, n525, n526, n527, n528,
    n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559, n560, n561, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
    n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
    n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n631, n632, n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n729, n730, n731, n732, n733, n734, n735, n736, n737,
    n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n810, n811,
    n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
    n848, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n950, n951, n952, n953, n954, n955, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002, n1004, n1005, n1006, n1007,
    n1008, n1010, n1011, n1012, n1013, n1014, n1015, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1036, n1037, n1038, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
    n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
    n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
    n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
    n1304, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1440, n1441, n1442,
    n1443, n1444, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
    n1454, n1455, n1456, n1457, n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1467, n1468, n1469, n1470, n1471, n1472, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1487,
    n1488, n1489, n1490, n1492, n1493, n1494, n1495, n1496, n1498, n1499,
    n1500, n1501, n1502, n1504, n1505, n1506, n1507, n1508, n1510, n1511,
    n1512, n1513, n1514, n1516, n1517, n1518, n1519, n1520, n1522, n1523,
    n1524, n1525, n1526, n1528, n1529, n1530, n1531, n1532, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1542, n1543, n1544, n1545, n1546,
    n1547;
  assign n163 = ~pi13 & ~pi14;
  assign n164 = ~pi11 & n163;
  assign n165 = pi19 & n164;
  assign n166 = ~pi26 & n165;
  assign n167 = ~pi19 & pi26;
  assign n168 = n164 & n167;
  assign n169 = ~pi19 & ~pi26;
  assign n170 = ~pi11 & n169;
  assign n171 = ~pi13 & n170;
  assign n172 = pi14 & n171;
  assign n173 = pi11 & n169;
  assign n174 = n163 & n173;
  assign n175 = ~n172 & ~n174;
  assign n176 = ~n168 & n175;
  assign n177 = ~n166 & n176;
  assign n178 = pi00 & n177;
  assign n179 = pi00 & pi12;
  assign n180 = pi00 & ~pi28;
  assign n181 = ~pi17 & pi21;
  assign n182 = ~pi18 & pi22;
  assign n183 = pi16 & ~pi24;
  assign n184 = n182 & n183;
  assign n185 = pi20 & ~pi23;
  assign n186 = n184 & n185;
  assign n187 = n181 & n186;
  assign n188 = pi25 & n187;
  assign n189 = pi32 & ~pi38;
  assign n190 = ~pi35 & ~pi42;
  assign n191 = ~pi30 & n190;
  assign n192 = ~pi36 & n191;
  assign n193 = ~pi15 & ~pi44;
  assign n194 = ~pi37 & n193;
  assign n195 = n192 & n194;
  assign n196 = n189 & n195;
  assign n197 = n188 & n196;
  assign n198 = ~pi27 & ~n197;
  assign n199 = n180 & n198;
  assign n200 = ~pi32 & ~pi38;
  assign n201 = ~pi58 & n200;
  assign n202 = ~pi24 & ~pi25;
  assign n203 = ~pi20 & pi21;
  assign n204 = pi16 & pi23;
  assign n205 = n203 & n204;
  assign n206 = pi18 & pi22;
  assign n207 = pi17 & n206;
  assign n208 = n205 & n207;
  assign n209 = n202 & n208;
  assign n210 = ~pi15 & pi44;
  assign n211 = ~pi37 & n210;
  assign n212 = n192 & n211;
  assign n213 = n209 & n212;
  assign n214 = n201 & n213;
  assign n215 = pi00 & pi27;
  assign n216 = ~pi28 & n215;
  assign n217 = n214 & n216;
  assign n218 = ~n199 & ~n217;
  assign n219 = pi00 & pi28;
  assign n220 = pi27 & ~pi28;
  assign n221 = ~pi58 & n202;
  assign n222 = n200 & n221;
  assign n223 = n208 & n222;
  assign n224 = n212 & n223;
  assign n225 = pi00 & ~n224;
  assign n226 = n192 & n200;
  assign n227 = n211 & n226;
  assign n228 = n209 & n227;
  assign n229 = pi58 & n228;
  assign n230 = ~n214 & n229;
  assign n231 = ~n225 & ~n230;
  assign n232 = n220 & ~n231;
  assign n233 = ~n219 & ~n232;
  assign n234 = n218 & n233;
  assign n235 = ~pi12 & ~n234;
  assign n236 = ~n179 & ~n235;
  assign n237 = n174 & ~n236;
  assign n238 = ~n178 & ~n237;
  assign n239 = pi00 & pi10;
  assign n240 = ~pi46 & ~pi49;
  assign n241 = ~n197 & n240;
  assign n242 = pi00 & n241;
  assign n243 = ~pi46 & pi49;
  assign n244 = pi00 & n243;
  assign n245 = ~n242 & ~n244;
  assign n246 = ~pi10 & ~n245;
  assign n247 = ~pi23 & ~pi25;
  assign n248 = pi17 & ~pi20;
  assign n249 = pi21 & pi24;
  assign n250 = ~pi16 & n249;
  assign n251 = n248 & n250;
  assign n252 = n182 & n251;
  assign n253 = n247 & n252;
  assign n254 = ~pi32 & pi38;
  assign n255 = n194 & n254;
  assign n256 = n192 & n255;
  assign n257 = n253 & n256;
  assign n258 = ~pi00 & ~n257;
  assign n259 = ~pi10 & pi46;
  assign n260 = ~n258 & n259;
  assign n261 = ~n246 & ~n260;
  assign n262 = ~n239 & n261;
  assign n263 = n166 & ~n262;
  assign n264 = ~n199 & ~n219;
  assign n265 = pi27 & n224;
  assign n266 = pi27 & n229;
  assign n267 = ~n215 & ~n266;
  assign n268 = ~n265 & n267;
  assign n269 = ~pi28 & ~n268;
  assign n270 = n264 & ~n269;
  assign n271 = n172 & ~n270;
  assign n272 = n218 & ~n232;
  assign n273 = ~n219 & n272;
  assign n274 = n168 & ~n273;
  assign n275 = ~n271 & ~n274;
  assign n276 = ~n263 & n275;
  assign po16 = ~n238 | ~n276;
  assign n278 = pi13 & ~pi14;
  assign n279 = n170 & n278;
  assign n280 = n176 & ~n279;
  assign n281 = pi01 & n280;
  assign n282 = pi75 & n279;
  assign n283 = ~pi27 & ~pi28;
  assign n284 = pi01 & n283;
  assign n285 = ~pi37 & ~pi44;
  assign n286 = ~pi35 & n200;
  assign n287 = ~pi30 & n286;
  assign n288 = n285 & n287;
  assign n289 = ~pi15 & n288;
  assign n290 = pi42 & n289;
  assign n291 = ~pi36 & n290;
  assign n292 = n253 & n291;
  assign n293 = ~pi05 & n292;
  assign n294 = ~pi01 & ~n292;
  assign n295 = pi28 & ~n294;
  assign n296 = ~n293 & n295;
  assign n297 = ~n284 & ~n296;
  assign n298 = pi01 & ~n214;
  assign n299 = pi50 & n224;
  assign n300 = pi79 & n299;
  assign n301 = ~pi45 & ~pi47;
  assign n302 = ~pi50 & n224;
  assign n303 = pi01 & n302;
  assign n304 = n301 & n303;
  assign n305 = ~n300 & ~n304;
  assign n306 = ~n298 & n305;
  assign n307 = ~pi28 & ~n306;
  assign n308 = pi27 & n307;
  assign n309 = n297 & ~n308;
  assign n310 = n168 & ~n309;
  assign n311 = ~n282 & ~n310;
  assign n312 = pi01 & ~pi28;
  assign n313 = ~n296 & ~n312;
  assign n314 = n172 & ~n313;
  assign n315 = n311 & ~n314;
  assign n316 = ~n281 & n315;
  assign n317 = ~pi12 & n296;
  assign n318 = pi31 & ~pi50;
  assign n319 = n224 & ~n318;
  assign n320 = pi68 & n319;
  assign n321 = n214 & n318;
  assign n322 = pi01 & n321;
  assign n323 = ~n320 & ~n322;
  assign n324 = ~n298 & n323;
  assign n325 = pi27 & n324;
  assign n326 = ~pi01 & ~pi27;
  assign n327 = ~pi12 & ~pi28;
  assign n328 = ~n326 & n327;
  assign n329 = ~n325 & n328;
  assign n330 = ~n317 & ~n329;
  assign n331 = pi01 & pi12;
  assign n332 = n330 & ~n331;
  assign n333 = n174 & ~n332;
  assign po17 = ~n316 | n333;
  assign n335 = pi02 & ~pi27;
  assign n336 = n327 & n335;
  assign n337 = pi02 & ~n224;
  assign n338 = pi02 & n321;
  assign n339 = ~n337 & ~n338;
  assign n340 = pi70 & ~n318;
  assign n341 = n224 & n340;
  assign n342 = n339 & ~n341;
  assign n343 = pi27 & n327;
  assign n344 = ~n342 & n343;
  assign n345 = ~n336 & ~n344;
  assign n346 = pi02 & pi12;
  assign n347 = ~pi06 & n292;
  assign n348 = ~pi02 & ~n292;
  assign n349 = ~n347 & ~n348;
  assign n350 = pi28 & n349;
  assign n351 = ~pi12 & n350;
  assign n352 = ~n346 & ~n351;
  assign n353 = n345 & n352;
  assign n354 = n174 & ~n353;
  assign n355 = pi02 & n280;
  assign n356 = pi02 & n302;
  assign n357 = n301 & n356;
  assign n358 = pi81 & n214;
  assign n359 = pi50 & n358;
  assign n360 = ~n337 & ~n359;
  assign n361 = ~n357 & n360;
  assign n362 = ~pi28 & ~n361;
  assign n363 = pi27 & n362;
  assign n364 = ~pi28 & n335;
  assign n365 = ~n350 & ~n364;
  assign n366 = ~n363 & n365;
  assign n367 = n168 & ~n366;
  assign n368 = ~n355 & ~n367;
  assign n369 = ~n354 & n368;
  assign n370 = pi02 & ~pi28;
  assign n371 = ~n350 & ~n370;
  assign n372 = n172 & ~n371;
  assign po18 = ~n369 | n372;
  assign n374 = pi12 & n174;
  assign n375 = pi03 & n374;
  assign n376 = pi03 & n280;
  assign n377 = ~n375 & ~n376;
  assign n378 = ~pi03 & ~n292;
  assign n379 = ~pi08 & n292;
  assign n380 = ~n378 & ~n379;
  assign n381 = pi28 & n380;
  assign n382 = pi03 & ~pi28;
  assign n383 = ~n381 & ~n382;
  assign n384 = n172 & ~n383;
  assign n385 = n168 & n381;
  assign n386 = pi03 & n283;
  assign n387 = pi83 & n214;
  assign n388 = pi50 & n387;
  assign n389 = pi03 & ~n224;
  assign n390 = ~pi50 & n301;
  assign n391 = pi03 & n224;
  assign n392 = n390 & n391;
  assign n393 = ~n389 & ~n392;
  assign n394 = ~n388 & n393;
  assign n395 = ~pi28 & ~n394;
  assign n396 = pi27 & n395;
  assign n397 = ~n386 & ~n396;
  assign n398 = n168 & ~n397;
  assign n399 = ~n385 & ~n398;
  assign n400 = ~pi27 & n327;
  assign n401 = pi03 & n400;
  assign n402 = ~pi12 & n381;
  assign n403 = n318 & n391;
  assign n404 = ~n389 & ~n403;
  assign n405 = pi72 & n319;
  assign n406 = n404 & ~n405;
  assign n407 = n343 & ~n406;
  assign n408 = ~n402 & ~n407;
  assign n409 = ~n401 & n408;
  assign n410 = n174 & ~n409;
  assign n411 = n399 & ~n410;
  assign n412 = ~n384 & n411;
  assign po19 = ~n377 | ~n412;
  assign n414 = pi04 & ~n220;
  assign n415 = pi04 & n321;
  assign n416 = pi66 & n319;
  assign n417 = ~n415 & ~n416;
  assign n418 = pi04 & ~n224;
  assign n419 = n417 & ~n418;
  assign n420 = ~pi28 & ~n419;
  assign n421 = pi27 & n420;
  assign n422 = ~n414 & ~n421;
  assign n423 = ~pi12 & ~n422;
  assign n424 = pi04 & pi12;
  assign n425 = ~n423 & ~n424;
  assign n426 = n174 & ~n425;
  assign n427 = ~n172 & ~n280;
  assign n428 = pi04 & ~n427;
  assign n429 = ~n426 & ~n428;
  assign n430 = ~pi50 & ~n301;
  assign n431 = pi04 & ~pi50;
  assign n432 = ~n430 & ~n431;
  assign n433 = n214 & ~n432;
  assign n434 = pi77 & n299;
  assign n435 = ~n433 & ~n434;
  assign n436 = ~n418 & n435;
  assign n437 = pi27 & ~n436;
  assign n438 = ~pi28 & n437;
  assign n439 = pi04 & n283;
  assign n440 = ~n438 & ~n439;
  assign n441 = pi04 & pi28;
  assign n442 = n440 & ~n441;
  assign n443 = n168 & ~n442;
  assign po20 = ~n429 | n443;
  assign n445 = n224 & n390;
  assign n446 = pi05 & n445;
  assign n447 = pi78 & n299;
  assign n448 = ~n446 & ~n447;
  assign n449 = pi27 & ~n448;
  assign n450 = pi05 & ~n214;
  assign n451 = pi27 & n450;
  assign n452 = ~n449 & ~n451;
  assign n453 = ~pi28 & ~n452;
  assign n454 = ~pi04 & n292;
  assign n455 = ~pi05 & ~n292;
  assign n456 = pi28 & ~n455;
  assign n457 = ~n454 & n456;
  assign n458 = pi05 & n283;
  assign n459 = ~n457 & ~n458;
  assign n460 = ~n453 & n459;
  assign n461 = n168 & ~n460;
  assign n462 = pi74 & n279;
  assign n463 = pi05 & n280;
  assign n464 = ~n462 & ~n463;
  assign n465 = pi05 & ~pi28;
  assign n466 = ~n457 & ~n465;
  assign n467 = n172 & ~n466;
  assign n468 = n464 & ~n467;
  assign n469 = ~n461 & n468;
  assign n470 = ~pi05 & ~pi27;
  assign n471 = ~pi28 & ~n470;
  assign n472 = pi67 & n319;
  assign n473 = pi27 & ~n450;
  assign n474 = pi05 & n321;
  assign n475 = n473 & ~n474;
  assign n476 = ~n472 & n475;
  assign n477 = ~pi12 & ~n476;
  assign n478 = n471 & n477;
  assign n479 = ~pi12 & n457;
  assign n480 = ~n478 & ~n479;
  assign n481 = pi05 & pi12;
  assign n482 = n480 & ~n481;
  assign n483 = n174 & ~n482;
  assign po21 = ~n469 | n483;
  assign n485 = pi76 & n279;
  assign n486 = pi06 & n280;
  assign n487 = ~n485 & ~n486;
  assign n488 = pi06 & n301;
  assign n489 = n302 & n488;
  assign n490 = pi80 & n299;
  assign n491 = ~n489 & ~n490;
  assign n492 = pi27 & ~n491;
  assign n493 = pi06 & ~n214;
  assign n494 = pi27 & n493;
  assign n495 = ~n492 & ~n494;
  assign n496 = ~pi28 & ~n495;
  assign n497 = ~pi01 & n292;
  assign n498 = ~pi06 & ~n292;
  assign n499 = pi28 & ~n498;
  assign n500 = ~n497 & n499;
  assign n501 = pi06 & n283;
  assign n502 = ~n500 & ~n501;
  assign n503 = ~n496 & n502;
  assign n504 = n168 & ~n503;
  assign n505 = pi06 & ~pi28;
  assign n506 = ~n500 & ~n505;
  assign n507 = n172 & ~n506;
  assign n508 = ~n504 & ~n507;
  assign n509 = n487 & n508;
  assign n510 = ~pi12 & n500;
  assign n511 = pi06 & ~pi27;
  assign n512 = pi06 & n321;
  assign n513 = pi69 & n319;
  assign n514 = ~n493 & ~n513;
  assign n515 = ~n512 & n514;
  assign n516 = pi27 & ~n515;
  assign n517 = ~n511 & ~n516;
  assign n518 = n327 & ~n517;
  assign n519 = ~n510 & ~n518;
  assign n520 = pi06 & pi12;
  assign n521 = n519 & ~n520;
  assign n522 = n174 & ~n521;
  assign po22 = ~n509 | n522;
  assign n524 = pi07 & n280;
  assign n525 = ~n279 & ~n524;
  assign n526 = ~pi03 & n292;
  assign n527 = ~pi07 & ~n292;
  assign n528 = pi28 & ~n527;
  assign n529 = ~n526 & n528;
  assign n530 = pi07 & ~pi28;
  assign n531 = ~n529 & ~n530;
  assign n532 = n172 & ~n531;
  assign n533 = n525 & ~n532;
  assign n534 = pi07 & ~pi50;
  assign n535 = ~n430 & ~n534;
  assign n536 = n214 & ~n535;
  assign n537 = pi84 & n299;
  assign n538 = ~n536 & ~n537;
  assign n539 = pi27 & ~n538;
  assign n540 = pi07 & ~n224;
  assign n541 = pi27 & n540;
  assign n542 = ~n539 & ~n541;
  assign n543 = ~pi28 & ~n542;
  assign n544 = pi07 & n283;
  assign n545 = ~n529 & ~n544;
  assign n546 = ~n543 & n545;
  assign n547 = n168 & ~n546;
  assign n548 = n533 & ~n547;
  assign n549 = ~pi07 & ~pi27;
  assign n550 = pi07 & n321;
  assign n551 = pi73 & n319;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n540 & n552;
  assign n554 = pi27 & n553;
  assign n555 = ~n549 & ~n554;
  assign n556 = n327 & n555;
  assign n557 = ~pi12 & n529;
  assign n558 = ~n556 & ~n557;
  assign n559 = pi07 & pi12;
  assign n560 = n558 & ~n559;
  assign n561 = n174 & ~n560;
  assign po23 = ~n548 | n561;
  assign n563 = pi08 & ~pi27;
  assign n564 = pi08 & ~n214;
  assign n565 = pi71 & ~n318;
  assign n566 = n224 & n565;
  assign n567 = ~n564 & ~n566;
  assign n568 = pi08 & n321;
  assign n569 = n567 & ~n568;
  assign n570 = pi27 & ~n569;
  assign n571 = ~n563 & ~n570;
  assign n572 = n327 & ~n571;
  assign n573 = ~pi02 & n292;
  assign n574 = ~pi08 & ~n292;
  assign n575 = ~n573 & ~n574;
  assign n576 = pi28 & n575;
  assign n577 = ~pi12 & n576;
  assign n578 = ~n279 & ~n577;
  assign n579 = ~n572 & n578;
  assign n580 = ~n174 & ~n279;
  assign n581 = ~n579 & ~n580;
  assign n582 = pi08 & pi12;
  assign n583 = n174 & n582;
  assign n584 = pi08 & ~pi28;
  assign n585 = ~n576 & ~n584;
  assign n586 = n172 & ~n585;
  assign n587 = pi08 & n283;
  assign n588 = ~n576 & ~n587;
  assign n589 = pi27 & n564;
  assign n590 = pi08 & ~pi50;
  assign n591 = ~n430 & ~n590;
  assign n592 = n214 & ~n591;
  assign n593 = pi82 & n299;
  assign n594 = ~n592 & ~n593;
  assign n595 = pi27 & ~n594;
  assign n596 = ~n589 & ~n595;
  assign n597 = ~pi28 & ~n596;
  assign n598 = n588 & ~n597;
  assign n599 = n168 & ~n598;
  assign n600 = pi08 & n280;
  assign n601 = ~n599 & ~n600;
  assign n602 = ~n586 & n601;
  assign n603 = ~n583 & n602;
  assign po24 = n581 | ~n603;
  assign n605 = pi09 & pi12;
  assign n606 = pi09 & pi28;
  assign n607 = pi09 & ~n224;
  assign n608 = ~n230 & ~n607;
  assign n609 = pi27 & ~n608;
  assign n610 = ~pi00 & ~pi27;
  assign n611 = pi09 & n610;
  assign n612 = pi09 & pi27;
  assign n613 = n224 & n612;
  assign n614 = ~n611 & ~n613;
  assign n615 = ~n609 & n614;
  assign n616 = ~pi28 & ~n615;
  assign n617 = ~n606 & ~n616;
  assign n618 = ~pi12 & ~n617;
  assign n619 = ~n605 & ~n618;
  assign n620 = n174 & ~n619;
  assign n621 = n168 & ~n617;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~n611 & ~n612;
  assign n624 = ~n266 & n623;
  assign n625 = ~pi28 & ~n624;
  assign n626 = ~n606 & ~n625;
  assign n627 = n172 & ~n626;
  assign n628 = pi09 & n176;
  assign n629 = ~n627 & ~n628;
  assign po25 = ~n622 | ~n629;
  assign n631 = ~pi12 & pi28;
  assign n632 = pi10 & n631;
  assign n633 = pi10 & n283;
  assign n634 = pi10 & n214;
  assign n635 = ~n321 & ~n634;
  assign n636 = pi27 & ~n635;
  assign n637 = pi27 & ~n224;
  assign n638 = pi10 & n637;
  assign n639 = ~n636 & ~n638;
  assign n640 = ~pi28 & ~n639;
  assign n641 = ~n633 & ~n640;
  assign n642 = ~pi12 & ~n641;
  assign n643 = pi10 & pi12;
  assign n644 = ~n642 & ~n643;
  assign n645 = ~n632 & n644;
  assign n646 = n174 & ~n645;
  assign n647 = ~n166 & ~n174;
  assign n648 = pi10 & n647;
  assign n649 = n192 & n193;
  assign n650 = pi37 & n200;
  assign n651 = n649 & n650;
  assign n652 = n253 & n651;
  assign n653 = ~pi10 & ~n652;
  assign n654 = pi49 & ~n653;
  assign n655 = pi63 & n654;
  assign n656 = pi10 & pi49;
  assign n657 = ~pi63 & n656;
  assign n658 = ~pi10 & ~n657;
  assign n659 = ~n655 & n658;
  assign n660 = ~pi33 & ~pi34;
  assign n661 = ~pi39 & n660;
  assign n662 = pi40 & n661;
  assign n663 = pi10 & n662;
  assign n664 = ~n259 & ~n663;
  assign n665 = ~n659 & n664;
  assign n666 = n166 & n665;
  assign n667 = ~n648 & ~n666;
  assign po26 = n646 | ~n667;
  assign n669 = pi15 & ~pi30;
  assign n670 = n200 & n285;
  assign n671 = n190 & n670;
  assign n672 = ~pi36 & ~pi47;
  assign n673 = ~pi50 & n672;
  assign n674 = ~pi45 & n673;
  assign n675 = n671 & n674;
  assign n676 = n669 & n675;
  assign n677 = ~pi62 & ~pi64;
  assign n678 = ~pi63 & n677;
  assign n679 = n676 & ~n678;
  assign n680 = pi11 & n676;
  assign n681 = ~n679 & ~n680;
  assign n682 = pi11 & ~n676;
  assign n683 = n681 & ~n682;
  assign n684 = n279 & ~n683;
  assign n685 = pi00 & n197;
  assign n686 = pi11 & n283;
  assign n687 = ~n685 & n686;
  assign n688 = pi11 & pi28;
  assign n689 = ~n687 & ~n688;
  assign n690 = ~pi11 & n301;
  assign n691 = ~pi50 & ~n690;
  assign n692 = n265 & n691;
  assign n693 = pi11 & n637;
  assign n694 = ~n692 & ~n693;
  assign n695 = ~pi28 & ~n694;
  assign n696 = n689 & ~n695;
  assign n697 = n168 & ~n696;
  assign n698 = ~n684 & ~n697;
  assign n699 = ~pi10 & ~pi46;
  assign n700 = pi11 & ~n699;
  assign n701 = pi11 & ~n685;
  assign n702 = ~pi49 & n701;
  assign n703 = pi11 & pi49;
  assign n704 = ~n702 & ~n703;
  assign n705 = n699 & ~n704;
  assign n706 = ~n700 & ~n705;
  assign n707 = n166 & ~n706;
  assign n708 = n698 & ~n707;
  assign n709 = pi11 & n220;
  assign n710 = ~n687 & ~n709;
  assign n711 = ~n688 & n710;
  assign n712 = n172 & ~n711;
  assign n713 = pi11 & pi12;
  assign n714 = n174 & n713;
  assign n715 = ~pi12 & n174;
  assign n716 = ~pi27 & n701;
  assign n717 = ~n693 & ~n716;
  assign n718 = ~pi28 & ~n717;
  assign n719 = ~n688 & ~n718;
  assign n720 = n715 & ~n719;
  assign n721 = ~n714 & ~n720;
  assign n722 = ~n168 & ~n279;
  assign n723 = ~n166 & n722;
  assign n724 = n175 & n723;
  assign n725 = pi11 & n724;
  assign n726 = n721 & ~n725;
  assign n727 = ~n712 & n726;
  assign po27 = ~n708 | ~n727;
  assign n729 = ~pi16 & ~pi17;
  assign n730 = pi23 & ~pi25;
  assign n731 = ~pi22 & n730;
  assign n732 = pi20 & n249;
  assign n733 = n731 & n732;
  assign n734 = pi18 & n733;
  assign n735 = n729 & n734;
  assign n736 = ~pi15 & ~pi42;
  assign n737 = ~pi36 & n736;
  assign n738 = n670 & n737;
  assign n739 = pi30 & n738;
  assign n740 = ~pi35 & n739;
  assign n741 = n735 & n740;
  assign n742 = n374 & ~n741;
  assign n743 = pi12 & ~n174;
  assign n744 = ~n168 & n743;
  assign n745 = ~n279 & n744;
  assign n746 = ~n742 & ~n745;
  assign n747 = pi12 & ~n676;
  assign n748 = pi12 & n676;
  assign n749 = ~n679 & ~n748;
  assign n750 = ~n747 & n749;
  assign n751 = n279 & ~n750;
  assign n752 = n746 & ~n751;
  assign n753 = pi12 & pi50;
  assign n754 = pi12 & ~pi50;
  assign n755 = ~n430 & ~n754;
  assign n756 = ~n753 & n755;
  assign n757 = n214 & ~n756;
  assign n758 = pi27 & n757;
  assign n759 = pi12 & n637;
  assign n760 = ~n758 & ~n759;
  assign n761 = ~pi28 & ~n760;
  assign n762 = pi12 & n283;
  assign n763 = ~n761 & ~n762;
  assign n764 = pi12 & pi28;
  assign n765 = n763 & ~n764;
  assign n766 = n168 & ~n765;
  assign po28 = ~n752 | n766;
  assign n768 = ~pi13 & ~n685;
  assign n769 = n283 & ~n768;
  assign n770 = pi13 & pi28;
  assign n771 = pi13 & n220;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n769 & n772;
  assign n774 = n172 & ~n773;
  assign n775 = pi13 & pi27;
  assign n776 = ~n224 & n775;
  assign n777 = ~pi27 & ~n768;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~pi28 & ~n778;
  assign n780 = ~n770 & ~n779;
  assign n781 = n715 & ~n780;
  assign n782 = ~n774 & ~n781;
  assign n783 = n214 & n775;
  assign n784 = n390 & n783;
  assign n785 = ~n776 & ~n784;
  assign n786 = ~pi28 & ~n785;
  assign n787 = ~n769 & ~n786;
  assign n788 = ~n770 & n787;
  assign n789 = n168 & ~n788;
  assign n790 = n782 & ~n789;
  assign n791 = n279 & n676;
  assign n792 = n678 & n791;
  assign n793 = n279 & ~n676;
  assign n794 = ~n792 & ~n793;
  assign n795 = pi13 & ~n794;
  assign n796 = pi13 & n724;
  assign n797 = pi12 & pi13;
  assign n798 = n174 & n797;
  assign n799 = ~n796 & ~n798;
  assign n800 = ~n795 & n799;
  assign n801 = pi13 & ~n699;
  assign n802 = ~pi49 & ~n768;
  assign n803 = pi13 & pi49;
  assign n804 = ~n802 & ~n803;
  assign n805 = n699 & ~n804;
  assign n806 = ~n801 & ~n805;
  assign n807 = n166 & ~n806;
  assign n808 = n800 & ~n807;
  assign po29 = ~n790 | ~n808;
  assign n810 = pi14 & n724;
  assign n811 = pi14 & pi28;
  assign n812 = pi14 & n220;
  assign n813 = pi14 & n283;
  assign n814 = ~n685 & n813;
  assign n815 = ~n812 & ~n814;
  assign n816 = ~n811 & n815;
  assign n817 = n172 & ~n816;
  assign n818 = pi14 & ~n699;
  assign n819 = pi14 & ~n685;
  assign n820 = ~pi49 & n819;
  assign n821 = pi14 & pi49;
  assign n822 = ~n820 & ~n821;
  assign n823 = n699 & ~n822;
  assign n824 = ~n818 & ~n823;
  assign n825 = n166 & ~n824;
  assign n826 = pi12 & pi14;
  assign n827 = n174 & n826;
  assign n828 = pi14 & n637;
  assign n829 = ~pi27 & n819;
  assign n830 = ~n828 & ~n829;
  assign n831 = ~pi28 & ~n830;
  assign n832 = ~n811 & ~n831;
  assign n833 = n715 & ~n832;
  assign n834 = ~n827 & ~n833;
  assign n835 = ~n825 & n834;
  assign n836 = ~n817 & n835;
  assign n837 = ~n810 & n836;
  assign n838 = pi14 & ~n794;
  assign n839 = ~n811 & ~n814;
  assign n840 = pi14 & n301;
  assign n841 = n214 & n840;
  assign n842 = ~n299 & ~n841;
  assign n843 = pi27 & ~n842;
  assign n844 = ~n828 & ~n843;
  assign n845 = ~pi28 & ~n844;
  assign n846 = n839 & ~n845;
  assign n847 = n168 & ~n846;
  assign n848 = ~n838 & ~n847;
  assign po30 = ~n837 | ~n848;
  assign n850 = ~pi30 & pi35;
  assign n851 = n738 & n850;
  assign n852 = ~n651 & ~n851;
  assign n853 = n192 & n670;
  assign n854 = pi15 & n853;
  assign n855 = ~n740 & ~n854;
  assign n856 = ~n291 & n855;
  assign n857 = n288 & n736;
  assign n858 = pi36 & n857;
  assign n859 = ~n196 & ~n858;
  assign n860 = ~n227 & ~n256;
  assign n861 = n859 & n860;
  assign n862 = n856 & n861;
  assign n863 = n852 & n862;
  assign n864 = ~pi12 & n854;
  assign n865 = ~n863 & ~n864;
  assign n866 = pi15 & ~n865;
  assign n867 = pi15 & ~n188;
  assign n868 = n740 & n867;
  assign n869 = ~pi10 & n240;
  assign n870 = pi10 & pi15;
  assign n871 = ~n869 & ~n870;
  assign n872 = n188 & n851;
  assign n873 = ~n871 & n872;
  assign n874 = n188 & n740;
  assign n875 = ~pi28 & n874;
  assign n876 = ~n873 & ~n875;
  assign n877 = ~n868 & n876;
  assign n878 = ~pi00 & n188;
  assign n879 = ~n867 & ~n878;
  assign n880 = n256 & ~n879;
  assign n881 = pi15 & n196;
  assign n882 = ~n197 & ~n881;
  assign n883 = n851 & n867;
  assign n884 = n882 & ~n883;
  assign n885 = ~n880 & n884;
  assign n886 = ~pi00 & ~pi28;
  assign n887 = ~pi12 & n886;
  assign n888 = ~pi10 & n188;
  assign n889 = n227 & n888;
  assign n890 = n887 & n889;
  assign n891 = n227 & n867;
  assign n892 = ~n890 & ~n891;
  assign n893 = pi15 & pi28;
  assign n894 = ~n283 & ~n893;
  assign n895 = n188 & n291;
  assign n896 = ~n894 & n895;
  assign n897 = n291 & n867;
  assign n898 = ~n896 & ~n897;
  assign n899 = n892 & n898;
  assign n900 = n885 & n899;
  assign n901 = n877 & n900;
  assign n902 = ~pi12 & n735;
  assign n903 = pi15 & ~n735;
  assign n904 = ~n902 & ~n903;
  assign n905 = n858 & ~n904;
  assign n906 = ~n867 & ~n888;
  assign n907 = n651 & ~n906;
  assign n908 = ~n905 & ~n907;
  assign n909 = n901 & n908;
  assign po31 = n866 | ~n909;
  assign n911 = pi36 & n671;
  assign n912 = pi37 & ~pi44;
  assign n913 = n200 & n912;
  assign n914 = ~pi44 & ~n189;
  assign n915 = ~n254 & n914;
  assign n916 = pi44 & ~n200;
  assign n917 = ~n915 & ~n916;
  assign n918 = ~pi37 & n917;
  assign n919 = ~n913 & ~n918;
  assign n920 = n190 & ~n919;
  assign n921 = ~pi35 & pi42;
  assign n922 = n670 & n921;
  assign n923 = pi35 & n285;
  assign n924 = n200 & n923;
  assign n925 = ~pi42 & n924;
  assign n926 = ~n922 & ~n925;
  assign n927 = ~n920 & n926;
  assign n928 = ~pi36 & ~n927;
  assign n929 = ~n911 & ~n928;
  assign n930 = ~pi30 & ~n929;
  assign n931 = pi30 & ~pi36;
  assign n932 = n671 & n931;
  assign n933 = ~n930 & ~n932;
  assign n934 = ~pi15 & ~n933;
  assign n935 = pi16 & n732;
  assign n936 = ~pi16 & ~n732;
  assign n937 = ~n935 & ~n936;
  assign n938 = n934 & n937;
  assign n939 = pi16 & ~n934;
  assign n940 = ~n938 & ~n939;
  assign n941 = pi12 & n854;
  assign n942 = ~n895 & ~n941;
  assign n943 = n735 & n858;
  assign n944 = n852 & n860;
  assign n945 = n188 & ~n944;
  assign n946 = ~n943 & ~n945;
  assign n947 = ~n874 & n946;
  assign n948 = n942 & n947;
  assign po32 = ~n940 & n948;
  assign n950 = pi17 & n935;
  assign n951 = ~pi17 & ~n935;
  assign n952 = ~n950 & ~n951;
  assign n953 = n934 & n952;
  assign n954 = pi17 & ~n934;
  assign n955 = ~n953 & ~n954;
  assign po33 = n948 & ~n955;
  assign n957 = pi16 & pi17;
  assign n958 = pi20 & pi21;
  assign n959 = n957 & n958;
  assign n960 = pi24 & n959;
  assign n961 = ~pi18 & n960;
  assign n962 = pi18 & ~n960;
  assign n963 = ~n961 & ~n962;
  assign n964 = n934 & ~n963;
  assign n965 = pi18 & ~n934;
  assign n966 = ~n964 & ~n965;
  assign po34 = n948 & ~n966;
  assign n968 = pi19 & pi28;
  assign n969 = pi19 & ~n685;
  assign n970 = n283 & n969;
  assign n971 = pi19 & ~pi28;
  assign n972 = pi27 & n971;
  assign n973 = ~n970 & ~n972;
  assign n974 = ~n968 & n973;
  assign n975 = n172 & ~n974;
  assign n976 = pi19 & n724;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n968 & ~n970;
  assign n979 = pi19 & ~n214;
  assign n980 = ~n321 & ~n979;
  assign n981 = n220 & ~n980;
  assign n982 = n978 & ~n981;
  assign n983 = n715 & ~n982;
  assign n984 = pi12 & pi19;
  assign n985 = n174 & n984;
  assign n986 = ~n983 & ~n985;
  assign n987 = n214 & ~n390;
  assign n988 = pi27 & ~n987;
  assign n989 = n971 & n988;
  assign n990 = n978 & ~n989;
  assign n991 = n168 & ~n990;
  assign n992 = pi19 & ~n794;
  assign n993 = ~n991 & ~n992;
  assign n994 = pi19 & ~n699;
  assign n995 = ~pi49 & n969;
  assign n996 = pi19 & pi49;
  assign n997 = ~n995 & ~n996;
  assign n998 = n699 & ~n997;
  assign n999 = ~n994 & ~n998;
  assign n1000 = n166 & ~n999;
  assign n1001 = n993 & ~n1000;
  assign n1002 = n986 & n1001;
  assign po35 = ~n977 | ~n1002;
  assign n1004 = ~pi20 & ~n249;
  assign n1005 = ~n732 & ~n1004;
  assign n1006 = n934 & n1005;
  assign n1007 = pi20 & ~n934;
  assign n1008 = ~n1006 & ~n1007;
  assign po36 = n948 & ~n1008;
  assign n1010 = pi21 & ~pi24;
  assign n1011 = ~pi21 & pi24;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = n934 & ~n1012;
  assign n1014 = pi21 & ~n934;
  assign n1015 = ~n1013 & ~n1014;
  assign po37 = n948 & ~n1015;
  assign n1017 = n249 & n957;
  assign n1018 = pi20 & n1017;
  assign n1019 = pi18 & n1018;
  assign n1020 = ~pi22 & n1019;
  assign n1021 = pi22 & ~n1019;
  assign n1022 = ~n1020 & ~n1021;
  assign n1023 = n934 & ~n1022;
  assign n1024 = pi22 & ~n934;
  assign n1025 = ~n1023 & ~n1024;
  assign po38 = n948 & ~n1025;
  assign n1027 = n206 & n957;
  assign n1028 = n732 & n1027;
  assign n1029 = pi23 & n1028;
  assign n1030 = ~pi23 & ~n1028;
  assign n1031 = ~n1029 & ~n1030;
  assign n1032 = n934 & n1031;
  assign n1033 = pi23 & ~n934;
  assign n1034 = ~n1032 & ~n1033;
  assign po39 = n948 & ~n1034;
  assign n1036 = pi24 & n934;
  assign n1037 = ~pi24 & ~n934;
  assign n1038 = ~n1036 & ~n1037;
  assign po40 = n948 & n1038;
  assign n1040 = pi17 & pi23;
  assign n1041 = pi18 & n935;
  assign n1042 = pi22 & n1041;
  assign n1043 = n1040 & n1042;
  assign n1044 = pi25 & n1043;
  assign n1045 = ~pi25 & ~n1043;
  assign n1046 = ~n1044 & ~n1045;
  assign n1047 = n934 & n1046;
  assign n1048 = pi25 & ~n934;
  assign n1049 = ~n1047 & ~n1048;
  assign po41 = n948 & ~n1049;
  assign n1051 = pi26 & pi28;
  assign n1052 = pi26 & ~n685;
  assign n1053 = n283 & n1052;
  assign n1054 = pi26 & ~pi28;
  assign n1055 = pi27 & n1054;
  assign n1056 = ~n1053 & ~n1055;
  assign n1057 = ~n1051 & n1056;
  assign n1058 = n172 & ~n1057;
  assign n1059 = pi26 & n724;
  assign n1060 = ~n1058 & ~n1059;
  assign n1061 = ~n1051 & ~n1053;
  assign n1062 = pi26 & ~n214;
  assign n1063 = ~n319 & ~n1062;
  assign n1064 = n220 & ~n1063;
  assign n1065 = n1061 & ~n1064;
  assign n1066 = n715 & ~n1065;
  assign n1067 = pi12 & pi26;
  assign n1068 = n174 & n1067;
  assign n1069 = ~n1066 & ~n1068;
  assign n1070 = n988 & n1054;
  assign n1071 = n1061 & ~n1070;
  assign n1072 = n168 & ~n1071;
  assign n1073 = pi26 & ~n794;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = pi26 & ~n699;
  assign n1076 = ~pi49 & n1052;
  assign n1077 = pi26 & pi49;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = n699 & ~n1078;
  assign n1080 = ~n1075 & ~n1079;
  assign n1081 = n166 & ~n1080;
  assign n1082 = n1074 & ~n1081;
  assign n1083 = n1069 & n1082;
  assign po42 = ~n1060 | ~n1083;
  assign n1085 = n220 & ~n229;
  assign n1086 = ~n214 & n1085;
  assign n1087 = ~pi27 & ~n662;
  assign n1088 = pi28 & ~n1087;
  assign n1089 = ~n1086 & ~n1088;
  assign n1090 = n172 & ~n1089;
  assign n1091 = n168 & ~n1089;
  assign n1092 = pi27 & n176;
  assign n1093 = ~n1091 & ~n1092;
  assign n1094 = pi12 & pi27;
  assign n1095 = ~pi12 & ~n1089;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = n174 & ~n1096;
  assign n1098 = n1093 & ~n1097;
  assign po43 = n1090 | ~n1098;
  assign n1100 = ~pi28 & ~n741;
  assign n1101 = n374 & ~n1100;
  assign n1102 = pi28 & n176;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = pi28 & ~n662;
  assign n1105 = ~pi27 & pi28;
  assign n1106 = ~pi28 & ~n319;
  assign n1107 = pi27 & ~n1106;
  assign n1108 = ~n1105 & ~n1107;
  assign n1109 = ~pi28 & ~n1108;
  assign n1110 = ~n1104 & ~n1109;
  assign n1111 = n715 & ~n1110;
  assign n1112 = ~pi28 & ~n299;
  assign n1113 = pi27 & ~n1112;
  assign n1114 = ~n1105 & ~n1113;
  assign n1115 = ~pi28 & ~n1114;
  assign n1116 = ~n1104 & ~n1115;
  assign n1117 = n168 & ~n1116;
  assign n1118 = n172 & n1104;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1111 & n1119;
  assign po44 = ~n1103 | ~n1120;
  assign n1122 = ~pi28 & n188;
  assign n1123 = n740 & ~n1122;
  assign n1124 = ~pi07 & n253;
  assign n1125 = n291 & n1124;
  assign n1126 = ~pi28 & ~n220;
  assign n1127 = n188 & ~n1126;
  assign n1128 = n1125 & n1127;
  assign n1129 = ~n188 & n1125;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n188 & n253;
  assign n1132 = pi28 & n188;
  assign n1133 = n253 & n1132;
  assign n1134 = ~pi28 & n253;
  assign n1135 = ~n283 & ~n1134;
  assign n1136 = n188 & ~n1135;
  assign n1137 = ~n1133 & ~n1136;
  assign n1138 = ~n1131 & n1137;
  assign n1139 = n291 & ~n1138;
  assign n1140 = pi28 & ~n735;
  assign n1141 = n874 & ~n1140;
  assign n1142 = ~n188 & n741;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = ~n851 & ~n858;
  assign n1145 = n253 & ~n1144;
  assign n1146 = ~n197 & ~n1145;
  assign n1147 = ~n196 & n860;
  assign n1148 = n253 & ~n1147;
  assign n1149 = n1146 & ~n1148;
  assign n1150 = pi10 & ~n253;
  assign n1151 = n188 & ~n1150;
  assign n1152 = ~n1131 & ~n1151;
  assign n1153 = n651 & ~n1152;
  assign n1154 = n1149 & ~n1153;
  assign n1155 = n1143 & n1154;
  assign n1156 = ~n1139 & n1155;
  assign n1157 = pi10 & n188;
  assign n1158 = n253 & n1157;
  assign n1159 = ~n1131 & ~n1158;
  assign n1160 = n651 & ~n1159;
  assign n1161 = n196 & n1131;
  assign n1162 = ~n1160 & ~n1161;
  assign n1163 = ~n1156 & n1162;
  assign n1164 = n1130 & n1163;
  assign n1165 = ~n1123 & n1164;
  assign n1166 = pi29 & n1156;
  assign po45 = n1165 | n1166;
  assign n1168 = pi30 & ~n188;
  assign n1169 = pi30 & n1157;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = n851 & ~n1170;
  assign n1172 = ~n854 & ~n863;
  assign n1173 = pi30 & ~n1172;
  assign n1174 = ~n941 & ~n1173;
  assign n1175 = n740 & n1168;
  assign n1176 = ~n860 & n1168;
  assign n1177 = pi28 & pi30;
  assign n1178 = n188 & n1177;
  assign n1179 = ~n1168 & ~n1178;
  assign n1180 = n291 & ~n1179;
  assign n1181 = ~n1176 & ~n1180;
  assign n1182 = ~n1175 & n1181;
  assign n1183 = n1174 & n1182;
  assign n1184 = ~n1171 & n1183;
  assign n1185 = ~pi30 & ~n735;
  assign n1186 = ~n902 & ~n1185;
  assign n1187 = n858 & n1186;
  assign n1188 = n651 & n1168;
  assign n1189 = ~n1187 & ~n1188;
  assign po46 = ~n1184 | ~n1189;
  assign n1191 = pi31 & n722;
  assign n1192 = pi27 & pi31;
  assign n1193 = ~n265 & ~n1192;
  assign n1194 = ~pi28 & ~n1193;
  assign n1195 = pi31 & n283;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = pi28 & pi31;
  assign n1198 = n1196 & ~n1197;
  assign n1199 = n168 & ~n1198;
  assign po47 = n1191 | n1199;
  assign n1201 = pi32 & ~n188;
  assign n1202 = pi00 & n188;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = n256 & ~n1203;
  assign n1205 = pi32 & n863;
  assign n1206 = ~n1204 & ~n1205;
  assign n1207 = n188 & n227;
  assign n1208 = ~pi10 & n1207;
  assign n1209 = n180 & n1208;
  assign n1210 = pi32 & n1157;
  assign n1211 = ~n1201 & ~n1210;
  assign n1212 = n851 & ~n1211;
  assign n1213 = pi28 & pi32;
  assign n1214 = n188 & n1213;
  assign n1215 = ~n1201 & ~n1214;
  assign n1216 = n291 & ~n1215;
  assign n1217 = ~n1212 & ~n1216;
  assign n1218 = ~n196 & ~n651;
  assign n1219 = n1201 & ~n1218;
  assign n1220 = n1217 & ~n1219;
  assign n1221 = ~n1209 & n1220;
  assign po48 = ~n1206 | ~n1221;
  assign n1223 = pi33 & ~n292;
  assign n1224 = ~pi33 & n292;
  assign n1225 = ~n1223 & ~n1224;
  assign n1226 = pi28 & ~n1225;
  assign n1227 = pi33 & n283;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n172 & ~n715;
  assign n1230 = ~n168 & n1229;
  assign n1231 = ~n1228 & ~n1230;
  assign n1232 = pi33 & n177;
  assign n1233 = n209 & n851;
  assign n1234 = pi33 & ~n1233;
  assign n1235 = ~pi33 & n1233;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = pi10 & ~n1236;
  assign n1238 = pi33 & n869;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = n166 & ~n1239;
  assign n1241 = ~n1232 & ~n1240;
  assign po49 = n1231 | ~n1241;
  assign n1243 = pi34 & ~n292;
  assign n1244 = pi33 & pi39;
  assign n1245 = ~pi34 & n1244;
  assign n1246 = pi34 & ~n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = n292 & ~n1247;
  assign n1249 = ~n1243 & ~n1248;
  assign n1250 = pi28 & ~n1249;
  assign n1251 = pi34 & n283;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1230 & ~n1252;
  assign n1254 = pi34 & n177;
  assign n1255 = pi34 & ~n1233;
  assign n1256 = n1233 & ~n1247;
  assign n1257 = ~n1255 & ~n1256;
  assign n1258 = pi10 & ~n1257;
  assign n1259 = pi34 & n869;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = n166 & ~n1260;
  assign n1262 = ~n1254 & ~n1261;
  assign po50 = n1253 | ~n1262;
  assign n1264 = pi35 & ~n188;
  assign n1265 = pi35 & n1157;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = n851 & ~n1266;
  assign n1268 = pi10 & ~pi28;
  assign n1269 = n188 & n1268;
  assign n1270 = ~n1264 & ~n1269;
  assign n1271 = n227 & ~n1270;
  assign n1272 = ~n1267 & ~n1271;
  assign n1273 = pi35 & n863;
  assign n1274 = pi28 & pi35;
  assign n1275 = n188 & n1274;
  assign n1276 = ~n1264 & ~n1275;
  assign n1277 = n291 & ~n1276;
  assign n1278 = ~n1273 & ~n1277;
  assign n1279 = ~n1157 & ~n1264;
  assign n1280 = n651 & ~n1279;
  assign n1281 = n740 & n1264;
  assign n1282 = ~n1280 & ~n1281;
  assign n1283 = n1278 & n1282;
  assign po51 = ~n1272 | ~n1283;
  assign n1285 = pi12 & n886;
  assign n1286 = n889 & n1285;
  assign n1287 = pi36 & ~n188;
  assign n1288 = n227 & n1287;
  assign n1289 = ~n1286 & ~n1288;
  assign n1290 = pi36 & n1157;
  assign n1291 = ~n1287 & ~n1290;
  assign n1292 = n851 & ~n1291;
  assign n1293 = pi36 & n863;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~n735 & n858;
  assign n1296 = pi36 & n1295;
  assign n1297 = pi28 & pi36;
  assign n1298 = n188 & n1297;
  assign n1299 = ~n1287 & ~n1298;
  assign n1300 = n291 & ~n1299;
  assign n1301 = n651 & n1287;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~n1296 & n1302;
  assign n1304 = n1294 & n1303;
  assign po52 = ~n1289 | ~n1304;
  assign n1306 = pi37 & ~n188;
  assign n1307 = n851 & n1306;
  assign n1308 = ~pi10 & pi49;
  assign n1309 = pi10 & pi37;
  assign n1310 = ~n1308 & ~n1309;
  assign n1311 = n872 & ~n1310;
  assign n1312 = ~n1307 & ~n1311;
  assign n1313 = ~n1147 & n1306;
  assign n1314 = n1312 & ~n1313;
  assign n1315 = pi37 & n863;
  assign n1316 = pi28 & pi37;
  assign n1317 = n188 & n1316;
  assign n1318 = ~n1306 & ~n1317;
  assign n1319 = n291 & ~n1318;
  assign n1320 = ~n1315 & ~n1319;
  assign n1321 = n1314 & n1320;
  assign n1322 = n651 & n1306;
  assign po53 = ~n1321 | n1322;
  assign n1324 = pi38 & ~n188;
  assign n1325 = pi10 & pi38;
  assign n1326 = n188 & n1325;
  assign n1327 = pi46 & n188;
  assign n1328 = ~pi10 & ~pi49;
  assign n1329 = n1327 & n1328;
  assign n1330 = ~n1326 & ~n1329;
  assign n1331 = ~n1324 & n1330;
  assign n1332 = n851 & ~n1331;
  assign n1333 = pi38 & n863;
  assign n1334 = ~n1332 & ~n1333;
  assign n1335 = ~n860 & n1324;
  assign n1336 = pi28 & pi38;
  assign n1337 = n188 & n1336;
  assign n1338 = ~n1324 & ~n1337;
  assign n1339 = n291 & ~n1338;
  assign n1340 = ~n1335 & ~n1339;
  assign n1341 = n651 & n1324;
  assign n1342 = n1340 & ~n1341;
  assign po54 = ~n1334 | ~n1342;
  assign n1344 = pi39 & ~n292;
  assign n1345 = ~pi33 & pi39;
  assign n1346 = pi33 & ~pi39;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = n292 & ~n1347;
  assign n1349 = ~n1344 & ~n1348;
  assign n1350 = pi28 & ~n1349;
  assign n1351 = pi39 & n283;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = ~n1230 & ~n1352;
  assign n1354 = pi39 & n177;
  assign n1355 = pi39 & ~n1233;
  assign n1356 = n1233 & ~n1347;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = pi10 & ~n1357;
  assign n1359 = pi39 & n869;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = n166 & ~n1360;
  assign n1362 = ~n1354 & ~n1361;
  assign po55 = n1353 | ~n1362;
  assign n1364 = pi40 & ~n292;
  assign n1365 = pi34 & n1244;
  assign n1366 = pi40 & ~n1365;
  assign n1367 = ~pi40 & n1365;
  assign n1368 = ~n1366 & ~n1367;
  assign n1369 = n292 & ~n1368;
  assign n1370 = ~n1364 & ~n1369;
  assign n1371 = pi28 & ~n1370;
  assign n1372 = pi40 & n283;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = ~n1230 & ~n1373;
  assign n1375 = pi40 & n177;
  assign n1376 = pi40 & ~n1233;
  assign n1377 = n1233 & ~n1368;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = pi10 & ~n1378;
  assign n1380 = pi40 & n869;
  assign n1381 = ~n1379 & ~n1380;
  assign n1382 = n166 & ~n1381;
  assign n1383 = ~n1375 & ~n1382;
  assign po56 = n1374 | ~n1383;
  assign n1385 = ~n291 & n852;
  assign n1386 = n861 & n1385;
  assign n1387 = ~pi18 & ~pi22;
  assign n1388 = n729 & n1387;
  assign n1389 = n247 & n1388;
  assign n1390 = ~pi24 & n1389;
  assign n1391 = ~pi20 & ~pi21;
  assign n1392 = n1390 & n1391;
  assign n1393 = ~n735 & ~n1392;
  assign n1394 = ~n1386 & ~n1393;
  assign n1395 = pi41 & ~n1394;
  assign n1396 = ~n1386 & n1392;
  assign n1397 = ~n735 & n1396;
  assign n1398 = n1394 & ~n1397;
  assign po57 = n1395 | n1398;
  assign n1400 = pi42 & ~n188;
  assign n1401 = pi42 & n1157;
  assign n1402 = ~n1400 & ~n1401;
  assign n1403 = n851 & ~n1402;
  assign n1404 = pi28 & pi42;
  assign n1405 = n188 & n1404;
  assign n1406 = ~n1400 & ~n1405;
  assign n1407 = n291 & ~n1406;
  assign n1408 = ~n1403 & ~n1407;
  assign n1409 = ~n1132 & ~n1400;
  assign n1410 = n740 & ~n1409;
  assign n1411 = n651 & n1400;
  assign n1412 = ~n1410 & ~n1411;
  assign n1413 = pi42 & n863;
  assign n1414 = n227 & ~n1409;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = n1412 & n1415;
  assign po58 = ~n1408 | ~n1416;
  assign n1418 = ~pi28 & n172;
  assign n1419 = pi43 & ~n1418;
  assign n1420 = pi00 & ~pi27;
  assign n1421 = pi43 & ~n1420;
  assign n1422 = ~n265 & ~n1421;
  assign n1423 = n172 & ~n1422;
  assign n1424 = ~pi28 & n1423;
  assign po59 = n1419 | n1424;
  assign n1426 = pi28 & pi44;
  assign n1427 = ~n220 & ~n1426;
  assign n1428 = n895 & ~n1427;
  assign n1429 = pi44 & ~n188;
  assign n1430 = n651 & n1429;
  assign n1431 = pi44 & n863;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = pi44 & n1157;
  assign n1434 = ~n1429 & ~n1433;
  assign n1435 = n851 & ~n1434;
  assign n1436 = ~n860 & n1429;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = n1432 & n1437;
  assign po60 = n1428 | ~n1438;
  assign n1440 = pi45 & ~n279;
  assign n1441 = ~pi45 & ~pi62;
  assign n1442 = ~pi64 & n279;
  assign n1443 = n676 & n1442;
  assign n1444 = ~n1441 & n1443;
  assign po61 = n1440 | n1444;
  assign n1446 = pi46 & ~n166;
  assign n1447 = ~pi45 & ~pi46;
  assign n1448 = n663 & ~n1447;
  assign n1449 = pi46 & ~n662;
  assign n1450 = pi10 & n1449;
  assign n1451 = ~n257 & n259;
  assign n1452 = ~pi46 & n1308;
  assign n1453 = ~pi63 & n1452;
  assign n1454 = ~n1451 & ~n1453;
  assign n1455 = ~n1450 & n1454;
  assign n1456 = ~n1448 & n1455;
  assign n1457 = n166 & ~n1456;
  assign po62 = n1446 | n1457;
  assign n1459 = ~pi47 & ~pi63;
  assign n1460 = n677 & ~n1459;
  assign n1461 = pi47 & pi62;
  assign n1462 = ~pi64 & n1461;
  assign n1463 = ~n1460 & ~n1462;
  assign n1464 = n791 & ~n1463;
  assign n1465 = pi47 & ~n279;
  assign po63 = n1464 | n1465;
  assign n1467 = pi10 & n166;
  assign n1468 = pi48 & ~n1467;
  assign n1469 = pi48 & ~n1233;
  assign n1470 = pi53 & n1233;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = n1467 & ~n1471;
  assign po64 = n1468 | n1472;
  assign n1474 = pi45 & ~pi49;
  assign n1475 = n663 & ~n1474;
  assign n1476 = n656 & ~n662;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = n166 & ~n1477;
  assign n1479 = pi49 & ~n166;
  assign n1480 = ~n1478 & ~n1479;
  assign n1481 = pi63 & ~n652;
  assign n1482 = n1452 & n1481;
  assign n1483 = pi46 & n1308;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = n166 & ~n1484;
  assign po65 = ~n1480 | n1485;
  assign n1487 = pi50 & ~n279;
  assign n1488 = pi64 & n279;
  assign n1489 = ~pi50 & ~n1488;
  assign n1490 = n676 & ~n1489;
  assign po66 = n1487 | n1490;
  assign n1492 = pi51 & ~n1467;
  assign n1493 = pi51 & ~n1233;
  assign n1494 = pi57 & n1233;
  assign n1495 = ~n1493 & ~n1494;
  assign n1496 = n1467 & ~n1495;
  assign po67 = n1492 | n1496;
  assign n1498 = pi52 & ~n1467;
  assign n1499 = pi52 & ~n1233;
  assign n1500 = pi51 & n1233;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = n1467 & ~n1501;
  assign po68 = n1498 | n1502;
  assign n1504 = pi53 & ~n1467;
  assign n1505 = pi53 & ~n1233;
  assign n1506 = pi52 & n1233;
  assign n1507 = ~n1505 & ~n1506;
  assign n1508 = n1467 & ~n1507;
  assign po69 = n1504 | n1508;
  assign n1510 = pi54 & ~n1467;
  assign n1511 = pi54 & ~n1233;
  assign n1512 = pi48 & n1233;
  assign n1513 = ~n1511 & ~n1512;
  assign n1514 = n1467 & ~n1513;
  assign po70 = n1510 | n1514;
  assign n1516 = pi55 & ~n1467;
  assign n1517 = pi55 & ~n1233;
  assign n1518 = pi54 & n1233;
  assign n1519 = ~n1517 & ~n1518;
  assign n1520 = n1467 & ~n1519;
  assign po71 = n1516 | n1520;
  assign n1522 = pi56 & ~n1467;
  assign n1523 = pi56 & ~n1233;
  assign n1524 = pi55 & n1233;
  assign n1525 = ~n1523 & ~n1524;
  assign n1526 = n1467 & ~n1525;
  assign po72 = n1522 | n1526;
  assign n1528 = pi57 & ~n1467;
  assign n1529 = pi57 & ~n1233;
  assign n1530 = pi58 & n1233;
  assign n1531 = ~n1529 & ~n1530;
  assign n1532 = n1467 & ~n1531;
  assign po73 = n1528 | n1532;
  assign n1534 = pi44 & n286;
  assign n1535 = ~pi37 & n1534;
  assign n1536 = ~n924 & ~n1535;
  assign n1537 = n737 & ~n1536;
  assign n1538 = ~pi30 & n1537;
  assign n1539 = pi58 & ~n1538;
  assign n1540 = pi65 & n1538;
  assign po74 = n1539 | n1540;
  assign n1542 = pi59 & n240;
  assign n1543 = ~pi10 & ~n1542;
  assign n1544 = ~pi59 & ~n662;
  assign n1545 = ~n1543 & ~n1544;
  assign n1546 = n166 & n1545;
  assign n1547 = pi59 & ~n166;
  assign po75 = n1546 | n1547;
  assign po14 = 1'b1;
  assign po13 = ~pi60;
  assign po00 = pi43;
  assign po01 = pi59;
  assign po02 = pi09;
  assign po03 = pi29;
  assign po04 = pi41;
  assign po05 = pi57;
  assign po06 = pi51;
  assign po07 = pi52;
  assign po08 = pi53;
  assign po09 = pi48;
  assign po10 = pi54;
  assign po11 = pi55;
  assign po12 = pi56;
  assign po15 = pi61;
endmodule


