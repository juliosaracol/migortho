module top (
            pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, 
            po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129);
input pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511;
output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009, po010, po011, po012, po013, po014, po015, po016, po017, po018, po019, po020, po021, po022, po023, po024, po025, po026, po027, po028, po029, po030, po031, po032, po033, po034, po035, po036, po037, po038, po039, po040, po041, po042, po043, po044, po045, po046, po047, po048, po049, po050, po051, po052, po053, po054, po055, po056, po057, po058, po059, po060, po061, po062, po063, po064, po065, po066, po067, po068, po069, po070, po071, po072, po073, po074, po075, po076, po077, po078, po079, po080, po081, po082, po083, po084, po085, po086, po087, po088, po089, po090, po091, po092, po093, po094, po095, po096, po097, po098, po099, po100, po101, po102, po103, po104, po105, po106, po107, po108, po109, po110, po111, po112, po113, po114, po115, po116, po117, po118, po119, po120, po121, po122, po123, po124, po125, po126, po127, po128, po129;
wire w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209;
assign w0 = pi024 & ~pi152;
assign w1 = pi016 & ~pi144;
assign w2 = pi006 & ~pi134;
assign w3 = ~pi005 & pi133;
assign w4 = pi001 & ~pi129;
assign w5 = pi000 & ~pi128;
assign w6 = ~w4 & ~w5;
assign w7 = ~pi001 & pi129;
assign w8 = ~pi002 & pi130;
assign w9 = ~w7 & ~w8;
assign w10 = ~w6 & w9;
assign w11 = pi003 & ~pi131;
assign w12 = pi002 & ~pi130;
assign w13 = ~w11 & ~w12;
assign w14 = ~pi004 & pi132;
assign w15 = ~pi003 & pi131;
assign w16 = ~w14 & ~w15;
assign w17 = (w16 & w10) | (w16 & w2743) | (w10 & w2743);
assign w18 = pi004 & ~pi132;
assign w19 = pi005 & ~pi133;
assign w20 = ~w18 & ~w19;
assign w21 = ~pi006 & pi134;
assign w22 = ~pi007 & pi135;
assign w23 = ~w21 & ~w22;
assign w24 = (w17 & w3647) | (w17 & w3648) | (w3647 & w3648);
assign w25 = pi008 & ~pi136;
assign w26 = pi007 & ~pi135;
assign w27 = ~w25 & ~w26;
assign w28 = ~pi008 & pi136;
assign w29 = ~pi010 & pi138;
assign w30 = ~pi009 & pi137;
assign w31 = ~w28 & ~w29;
assign w32 = ~w30 & w31;
assign w33 = pi011 & ~pi139;
assign w34 = pi010 & ~pi138;
assign w35 = pi009 & ~pi137;
assign w36 = ~w29 & w35;
assign w37 = ~w33 & ~w34;
assign w38 = ~w36 & w37;
assign w39 = (~w24 & w3932) | (~w24 & w3933) | (w3932 & w3933);
assign w40 = ~pi012 & pi140;
assign w41 = ~pi014 & pi142;
assign w42 = ~pi013 & pi141;
assign w43 = ~w41 & ~w42;
assign w44 = ~pi011 & pi139;
assign w45 = ~w40 & ~w44;
assign w46 = w43 & w45;
assign w47 = pi014 & ~pi142;
assign w48 = pi013 & ~pi141;
assign w49 = pi012 & ~pi140;
assign w50 = ~w48 & ~w49;
assign w51 = w43 & ~w50;
assign w52 = pi015 & ~pi143;
assign w53 = ~w47 & ~w52;
assign w54 = ~w51 & w53;
assign w55 = ~pi015 & pi143;
assign w56 = ~pi016 & pi144;
assign w57 = ~w55 & ~w56;
assign w58 = ~pi018 & pi146;
assign w59 = ~pi017 & pi145;
assign w60 = ~w58 & ~w59;
assign w61 = pi019 & ~pi147;
assign w62 = pi018 & ~pi146;
assign w63 = pi017 & ~pi145;
assign w64 = ~w58 & w63;
assign w65 = ~w61 & ~w62;
assign w66 = ~w64 & w65;
assign w67 = (w39 & w3990) | (w39 & w3991) | (w3990 & w3991);
assign w68 = ~pi019 & pi147;
assign w69 = ~pi022 & pi150;
assign w70 = ~pi021 & pi149;
assign w71 = ~pi020 & pi148;
assign w72 = ~w68 & ~w69;
assign w73 = ~w70 & ~w71;
assign w74 = w72 & w73;
assign w75 = pi022 & ~pi150;
assign w76 = pi023 & ~pi151;
assign w77 = pi021 & ~pi149;
assign w78 = pi020 & ~pi148;
assign w79 = ~w70 & w78;
assign w80 = (~w69 & w79) | (~w69 & w4056) | (w79 & w4056);
assign w81 = ~w75 & ~w76;
assign w82 = ~pi023 & pi151;
assign w83 = ~pi024 & pi152;
assign w84 = ~w82 & ~w83;
assign w85 = ~pi026 & pi154;
assign w86 = ~pi025 & pi153;
assign w87 = ~w85 & ~w86;
assign w88 = pi027 & ~pi155;
assign w89 = pi026 & ~pi154;
assign w90 = pi025 & ~pi153;
assign w91 = ~w85 & w90;
assign w92 = ~w88 & ~w89;
assign w93 = ~w91 & w92;
assign w94 = ~pi029 & pi157;
assign w95 = ~pi028 & pi156;
assign w96 = ~pi027 & pi155;
assign w97 = ~w94 & ~w95;
assign w98 = ~w96 & w97;
assign w99 = pi030 & ~pi158;
assign w100 = pi029 & ~pi157;
assign w101 = pi028 & ~pi156;
assign w102 = ~w94 & w101;
assign w103 = ~w99 & ~w100;
assign w104 = ~w102 & w103;
assign w105 = (w67 & w4040) | (w67 & w4041) | (w4040 & w4041);
assign w106 = ~pi036 & pi164;
assign w107 = ~pi039 & pi167;
assign w108 = ~pi038 & pi166;
assign w109 = ~pi037 & pi165;
assign w110 = ~w107 & ~w108;
assign w111 = ~w109 & w110;
assign w112 = ~pi033 & pi161;
assign w113 = ~pi160 & ~w112;
assign w114 = pi032 & ~w112;
assign w115 = ~w113 & ~w114;
assign w116 = ~pi035 & pi163;
assign w117 = ~pi034 & pi162;
assign w118 = ~w116 & ~w117;
assign w119 = ~pi030 & pi158;
assign w120 = ~pi031 & pi159;
assign w121 = ~w106 & ~w119;
assign w122 = ~w120 & w121;
assign w123 = w118 & w122;
assign w124 = w111 & ~w115;
assign w125 = w123 & w124;
assign w126 = ~w105 & w125;
assign w127 = pi038 & ~pi166;
assign w128 = ~w107 & w127;
assign w129 = ~pi047 & pi175;
assign w130 = pi046 & ~pi174;
assign w131 = ~w129 & w130;
assign w132 = pi047 & ~pi175;
assign w133 = ~pi046 & pi174;
assign w134 = ~pi045 & pi173;
assign w135 = ~w129 & ~w133;
assign w136 = ~w134 & w135;
assign w137 = pi044 & ~pi172;
assign w138 = pi045 & ~pi173;
assign w139 = ~pi044 & pi172;
assign w140 = pi043 & ~pi171;
assign w141 = ~pi043 & pi171;
assign w142 = ~pi042 & pi170;
assign w143 = ~w141 & ~w142;
assign w144 = pi042 & ~pi170;
assign w145 = pi041 & ~pi169;
assign w146 = ~pi041 & pi169;
assign w147 = pi040 & ~pi168;
assign w148 = ~w146 & w147;
assign w149 = ~w144 & ~w145;
assign w150 = ~w148 & w149;
assign w151 = (~w140 & w150) | (~w140 & w4024) | (w150 & w4024);
assign w152 = ~w137 & ~w138;
assign w153 = (w152 & w151) | (w152 & w4042) | (w151 & w4042);
assign w154 = w136 & ~w153;
assign w155 = ~w131 & ~w132;
assign w156 = ~w154 & w155;
assign w157 = pi039 & ~pi167;
assign w158 = pi036 & ~pi164;
assign w159 = pi037 & ~pi165;
assign w160 = pi035 & ~pi163;
assign w161 = pi034 & ~pi162;
assign w162 = pi033 & ~pi161;
assign w163 = ~w112 & w4025;
assign w164 = pi031 & ~pi159;
assign w165 = ~w115 & w164;
assign w166 = ~w161 & ~w162;
assign w167 = ~w163 & w166;
assign w168 = (w118 & w165) | (w118 & w4026) | (w165 & w4026);
assign w169 = ~w158 & ~w159;
assign w170 = w169 & w4202;
assign w171 = w111 & ~w170;
assign w172 = ~w128 & ~w157;
assign w173 = ~w154 & w4044;
assign w174 = ~w171 & w173;
assign w175 = ~w126 & w174;
assign w176 = ~pi040 & pi168;
assign w177 = ~w139 & ~w146;
assign w178 = ~w176 & w177;
assign w179 = w143 & w178;
assign w180 = w136 & w179;
assign w181 = w156 & ~w180;
assign w182 = ~pi059 & pi187;
assign w183 = ~pi058 & pi186;
assign w184 = ~w182 & ~w183;
assign w185 = ~pi057 & pi185;
assign w186 = ~pi056 & pi184;
assign w187 = ~w185 & ~w186;
assign w188 = w184 & w187;
assign w189 = ~pi051 & pi179;
assign w190 = ~pi050 & pi178;
assign w191 = ~w189 & ~w190;
assign w192 = ~pi054 & pi182;
assign w193 = ~pi055 & pi183;
assign w194 = ~w192 & ~w193;
assign w195 = ~pi053 & pi181;
assign w196 = ~pi052 & pi180;
assign w197 = ~w195 & ~w196;
assign w198 = ~pi049 & pi177;
assign w199 = ~pi060 & pi188;
assign w200 = ~pi063 & pi191;
assign w201 = ~pi062 & pi190;
assign w202 = ~pi061 & pi189;
assign w203 = ~w200 & ~w201;
assign w204 = ~w202 & w203;
assign w205 = ~w199 & w204;
assign w206 = ~pi048 & pi176;
assign w207 = ~w198 & ~w206;
assign w208 = w191 & w207;
assign w209 = w194 & w197;
assign w210 = w208 & w209;
assign w211 = w188 & w210;
assign w212 = w205 & w211;
assign w213 = ~w181 & w212;
assign w214 = ~w175 & w213;
assign w215 = pi063 & ~pi191;
assign w216 = pi057 & ~pi185;
assign w217 = pi058 & ~pi186;
assign w218 = pi056 & ~pi184;
assign w219 = ~w185 & w218;
assign w220 = ~w216 & ~w217;
assign w221 = ~w219 & w220;
assign w222 = w184 & ~w221;
assign w223 = pi059 & ~pi187;
assign w224 = pi055 & ~pi183;
assign w225 = pi054 & ~pi182;
assign w226 = pi053 & ~pi181;
assign w227 = pi051 & ~pi179;
assign w228 = pi052 & ~pi180;
assign w229 = pi050 & ~pi178;
assign w230 = pi049 & ~pi177;
assign w231 = pi048 & ~pi176;
assign w232 = ~w198 & w231;
assign w233 = ~w229 & ~w230;
assign w234 = ~w232 & w233;
assign w235 = ~w227 & ~w228;
assign w236 = (w235 & w234) | (w235 & w4027) | (w234 & w4027);
assign w237 = ~w225 & ~w226;
assign w238 = w194 & w4203;
assign w239 = (w188 & w238) | (w188 & w4065) | (w238 & w4065);
assign w240 = ~w222 & ~w223;
assign w241 = (w205 & w239) | (w205 & w4076) | (w239 & w4076);
assign w242 = pi067 & ~pi195;
assign w243 = ~pi067 & pi195;
assign w244 = ~pi066 & pi194;
assign w245 = ~w243 & ~w244;
assign w246 = pi065 & ~pi193;
assign w247 = pi066 & ~pi194;
assign w248 = ~pi065 & pi193;
assign w249 = pi064 & ~pi192;
assign w250 = ~w248 & w249;
assign w251 = ~w246 & ~w247;
assign w252 = ~w250 & w251;
assign w253 = (~w242 & w252) | (~w242 & w4066) | (w252 & w4066);
assign w254 = pi061 & ~pi189;
assign w255 = pi060 & ~pi188;
assign w256 = ~w254 & ~w255;
assign w257 = w204 & ~w256;
assign w258 = pi062 & ~pi190;
assign w259 = ~w200 & w258;
assign w260 = ~w215 & ~w259;
assign w261 = ~w257 & w260;
assign w262 = w253 & w261;
assign w263 = ~pi075 & pi203;
assign w264 = ~pi074 & pi202;
assign w265 = ~w263 & ~w264;
assign w266 = ~pi064 & pi192;
assign w267 = ~w248 & ~w266;
assign w268 = w245 & w267;
assign w269 = w253 & ~w268;
assign w270 = ~pi070 & pi198;
assign w271 = ~pi069 & pi197;
assign w272 = ~w270 & ~w271;
assign w273 = ~pi068 & pi196;
assign w274 = ~pi071 & pi199;
assign w275 = ~pi073 & pi201;
assign w276 = ~pi072 & pi200;
assign w277 = ~w274 & ~w275;
assign w278 = ~w276 & w277;
assign w279 = w265 & ~w273;
assign w280 = w272 & w279;
assign w281 = w278 & w280;
assign w282 = ~w269 & w281;
assign w283 = pi075 & ~pi203;
assign w284 = pi070 & ~pi198;
assign w285 = pi071 & ~pi199;
assign w286 = pi069 & ~pi197;
assign w287 = pi068 & ~pi196;
assign w288 = ~w286 & ~w287;
assign w289 = w272 & ~w288;
assign w290 = ~w284 & ~w285;
assign w291 = ~w289 & w290;
assign w292 = pi074 & ~pi202;
assign w293 = pi073 & ~pi201;
assign w294 = pi072 & ~pi200;
assign w295 = ~w275 & w294;
assign w296 = ~w292 & ~w293;
assign w297 = ~w295 & w296;
assign w298 = (w297 & w291) | (w297 & w4067) | (w291 & w4067);
assign w299 = w265 & ~w298;
assign w300 = pi079 & ~pi207;
assign w301 = pi077 & ~pi205;
assign w302 = pi076 & ~pi204;
assign w303 = ~w301 & ~w302;
assign w304 = ~pi079 & pi207;
assign w305 = ~pi078 & pi206;
assign w306 = ~pi077 & pi205;
assign w307 = ~w304 & ~w305;
assign w308 = ~w306 & w307;
assign w309 = ~w303 & w308;
assign w310 = pi078 & ~pi206;
assign w311 = ~w304 & w310;
assign w312 = ~w300 & ~w311;
assign w313 = ~w309 & w312;
assign w314 = ~w309 & w4077;
assign w315 = ~w299 & w314;
assign w316 = ~pi080 & pi208;
assign w317 = ~pi076 & pi204;
assign w318 = w308 & ~w317;
assign w319 = w313 & ~w318;
assign w320 = ~pi081 & pi209;
assign w321 = ~pi082 & pi210;
assign w322 = ~pi084 & pi212;
assign w323 = ~pi086 & pi214;
assign w324 = ~pi087 & pi215;
assign w325 = ~pi085 & pi213;
assign w326 = ~w323 & ~w324;
assign w327 = ~w325 & w326;
assign w328 = ~w322 & w327;
assign w329 = ~pi083 & pi211;
assign w330 = ~w321 & ~w329;
assign w331 = w328 & w330;
assign w332 = ~w316 & ~w320;
assign w333 = w331 & w332;
assign w334 = ~w319 & w333;
assign w335 = pi087 & ~pi215;
assign w336 = pi082 & ~pi210;
assign w337 = pi081 & ~pi209;
assign w338 = pi080 & ~pi208;
assign w339 = ~w320 & w338;
assign w340 = ~w336 & ~w337;
assign w341 = ~w339 & w340;
assign w342 = w331 & ~w341;
assign w343 = pi083 & ~pi211;
assign w344 = w328 & w343;
assign w345 = pi091 & ~pi219;
assign w346 = ~pi091 & pi219;
assign w347 = ~pi090 & pi218;
assign w348 = ~w346 & ~w347;
assign w349 = pi089 & ~pi217;
assign w350 = pi090 & ~pi218;
assign w351 = ~pi089 & pi217;
assign w352 = pi088 & ~pi216;
assign w353 = ~w351 & w352;
assign w354 = ~w349 & ~w350;
assign w355 = ~w353 & w354;
assign w356 = w348 & ~w355;
assign w357 = ~w345 & ~w356;
assign w358 = pi085 & ~pi213;
assign w359 = pi084 & ~pi212;
assign w360 = ~w358 & ~w359;
assign w361 = w327 & ~w360;
assign w362 = pi086 & ~pi214;
assign w363 = ~w324 & w362;
assign w364 = ~w335 & ~w363;
assign w365 = ~w361 & w364;
assign w366 = ~w344 & w365;
assign w367 = w357 & w366;
assign w368 = ~w342 & w367;
assign w369 = ~pi099 & pi227;
assign w370 = ~pi098 & pi226;
assign w371 = ~w369 & ~w370;
assign w372 = ~pi088 & pi216;
assign w373 = ~w351 & ~w372;
assign w374 = w348 & w373;
assign w375 = w357 & ~w374;
assign w376 = ~pi094 & pi222;
assign w377 = ~pi093 & pi221;
assign w378 = ~w376 & ~w377;
assign w379 = ~pi092 & pi220;
assign w380 = ~pi095 & pi223;
assign w381 = ~pi097 & pi225;
assign w382 = ~pi096 & pi224;
assign w383 = ~w380 & ~w381;
assign w384 = ~w382 & w383;
assign w385 = w371 & ~w379;
assign w386 = w378 & w385;
assign w387 = w384 & w386;
assign w388 = ~w375 & w387;
assign w389 = (w214 & w4068) | (w214 & w4069) | (w4068 & w4069);
assign w390 = pi099 & ~pi227;
assign w391 = pi094 & ~pi222;
assign w392 = pi095 & ~pi223;
assign w393 = pi093 & ~pi221;
assign w394 = pi092 & ~pi220;
assign w395 = ~w393 & ~w394;
assign w396 = w378 & ~w395;
assign w397 = ~w391 & ~w392;
assign w398 = ~w396 & w397;
assign w399 = w384 & ~w398;
assign w400 = pi098 & ~pi226;
assign w401 = pi097 & ~pi225;
assign w402 = pi096 & ~pi224;
assign w403 = ~w381 & w402;
assign w404 = ~w400 & ~w401;
assign w405 = ~w403 & w404;
assign w406 = ~w399 & w405;
assign w407 = w371 & ~w406;
assign w408 = pi103 & ~pi231;
assign w409 = pi101 & ~pi229;
assign w410 = pi100 & ~pi228;
assign w411 = ~w409 & ~w410;
assign w412 = ~pi103 & pi231;
assign w413 = ~pi102 & pi230;
assign w414 = ~pi101 & pi229;
assign w415 = ~w412 & ~w413;
assign w416 = ~w414 & w415;
assign w417 = ~w411 & w416;
assign w418 = pi102 & ~pi230;
assign w419 = ~w412 & w418;
assign w420 = ~w408 & ~w419;
assign w421 = ~w417 & w420;
assign w422 = ~w390 & w421;
assign w423 = ~w407 & w422;
assign w424 = ~pi104 & pi232;
assign w425 = ~pi100 & pi228;
assign w426 = w416 & ~w425;
assign w427 = w421 & ~w426;
assign w428 = ~pi105 & pi233;
assign w429 = ~pi106 & pi234;
assign w430 = ~pi108 & pi236;
assign w431 = ~pi110 & pi238;
assign w432 = ~pi111 & pi239;
assign w433 = ~pi109 & pi237;
assign w434 = ~w431 & ~w432;
assign w435 = ~w433 & w434;
assign w436 = ~w430 & w435;
assign w437 = ~pi107 & pi235;
assign w438 = ~w429 & ~w437;
assign w439 = w436 & w438;
assign w440 = ~w424 & ~w428;
assign w441 = w439 & w440;
assign w442 = ~w427 & w441;
assign w443 = pi111 & ~pi239;
assign w444 = pi106 & ~pi234;
assign w445 = pi105 & ~pi233;
assign w446 = pi104 & ~pi232;
assign w447 = ~w428 & w446;
assign w448 = ~w444 & ~w445;
assign w449 = ~w447 & w448;
assign w450 = w439 & ~w449;
assign w451 = pi107 & ~pi235;
assign w452 = w436 & w451;
assign w453 = pi115 & ~pi243;
assign w454 = ~pi115 & pi243;
assign w455 = ~pi114 & pi242;
assign w456 = ~w454 & ~w455;
assign w457 = pi113 & ~pi241;
assign w458 = pi114 & ~pi242;
assign w459 = ~pi113 & pi241;
assign w460 = pi112 & ~pi240;
assign w461 = ~w459 & w460;
assign w462 = ~w457 & ~w458;
assign w463 = ~w461 & w462;
assign w464 = w456 & ~w463;
assign w465 = ~w453 & ~w464;
assign w466 = pi109 & ~pi237;
assign w467 = pi108 & ~pi236;
assign w468 = ~w466 & ~w467;
assign w469 = w435 & ~w468;
assign w470 = pi110 & ~pi238;
assign w471 = ~w432 & w470;
assign w472 = ~w443 & ~w471;
assign w473 = ~w469 & w472;
assign w474 = ~w452 & w473;
assign w475 = w465 & w474;
assign w476 = ~w450 & w475;
assign w477 = ~pi112 & pi240;
assign w478 = ~w459 & ~w477;
assign w479 = w456 & w478;
assign w480 = w465 & ~w479;
assign w481 = ~pi119 & pi247;
assign w482 = ~pi120 & pi248;
assign w483 = ~w481 & ~w482;
assign w484 = ~pi116 & pi244;
assign w485 = ~pi118 & pi246;
assign w486 = ~pi117 & pi245;
assign w487 = ~w485 & ~w486;
assign w488 = ~pi123 & pi251;
assign w489 = ~pi122 & pi250;
assign w490 = ~pi121 & pi249;
assign w491 = ~w489 & ~w490;
assign w492 = ~w484 & ~w488;
assign w493 = w483 & w492;
assign w494 = w487 & w491;
assign w495 = w493 & w494;
assign w496 = ~w480 & w495;
assign w497 = pi123 & ~pi251;
assign w498 = pi121 & ~pi249;
assign w499 = pi119 & ~pi247;
assign w500 = pi117 & ~pi245;
assign w501 = pi116 & ~pi244;
assign w502 = ~w500 & ~w501;
assign w503 = w487 & ~w502;
assign w504 = pi118 & ~pi246;
assign w505 = ~w499 & ~w504;
assign w506 = ~w503 & w505;
assign w507 = w483 & ~w506;
assign w508 = pi120 & ~pi248;
assign w509 = ~w498 & ~w508;
assign w510 = ~w507 & w509;
assign w511 = w491 & ~w510;
assign w512 = pi122 & ~pi250;
assign w513 = ~w511 & ~w512;
assign w514 = ~w488 & ~w513;
assign w515 = ~w497 & ~w514;
assign w516 = (~w389 & w4088) | (~w389 & w4089) | (w4088 & w4089);
assign w517 = ~pi124 & pi252;
assign w518 = pi127 & ~pi255;
assign w519 = ~pi126 & pi254;
assign w520 = ~pi125 & pi253;
assign w521 = ~w518 & ~w519;
assign w522 = ~w520 & w521;
assign w523 = ~w517 & w522;
assign w524 = (w389 & w4198) | (w389 & w4199) | (w4198 & w4199);
assign w525 = pi125 & ~pi253;
assign w526 = pi124 & ~pi252;
assign w527 = ~w525 & ~w526;
assign w528 = w522 & ~w527;
assign w529 = pi126 & ~pi254;
assign w530 = ~w518 & w529;
assign w531 = ~w528 & ~w530;
assign w532 = (w531 & w4090) | (w531 & w516) | (w4090 & w516);
assign w533 = ~pi127 & pi255;
assign w534 = w532 & ~w533;
assign w535 = (pi000 & ~w532) | (pi000 & w4200) | (~w532 & w4200);
assign w536 = w532 & w4201;
assign w537 = ~w535 & ~w536;
assign w538 = pi280 & ~pi408;
assign w539 = pi272 & ~pi400;
assign w540 = pi262 & ~pi390;
assign w541 = ~pi261 & pi389;
assign w542 = pi257 & ~pi385;
assign w543 = pi256 & ~pi384;
assign w544 = ~w542 & ~w543;
assign w545 = ~pi257 & pi385;
assign w546 = ~pi258 & pi386;
assign w547 = ~w545 & ~w546;
assign w548 = ~w544 & w547;
assign w549 = pi259 & ~pi387;
assign w550 = pi258 & ~pi386;
assign w551 = ~w549 & ~w550;
assign w552 = ~pi260 & pi388;
assign w553 = ~pi259 & pi387;
assign w554 = ~w552 & ~w553;
assign w555 = (w554 & w548) | (w554 & w2744) | (w548 & w2744);
assign w556 = pi260 & ~pi388;
assign w557 = pi261 & ~pi389;
assign w558 = ~w556 & ~w557;
assign w559 = ~pi262 & pi390;
assign w560 = ~pi263 & pi391;
assign w561 = ~w559 & ~w560;
assign w562 = pi264 & ~pi392;
assign w563 = pi263 & ~pi391;
assign w564 = ~w562 & ~w563;
assign w565 = (~w555 & w3649) | (~w555 & w3650) | (w3649 & w3650);
assign w566 = ~pi264 & pi392;
assign w567 = ~pi266 & pi394;
assign w568 = ~pi265 & pi393;
assign w569 = ~w566 & ~w567;
assign w570 = ~w568 & w569;
assign w571 = pi267 & ~pi395;
assign w572 = pi266 & ~pi394;
assign w573 = pi265 & ~pi393;
assign w574 = ~w567 & w573;
assign w575 = ~w571 & ~w572;
assign w576 = ~w574 & w575;
assign w577 = ~pi267 & pi395;
assign w578 = ~pi270 & pi398;
assign w579 = ~pi269 & pi397;
assign w580 = ~w578 & ~w579;
assign w581 = ~pi268 & pi396;
assign w582 = ~w577 & ~w581;
assign w583 = w580 & w582;
assign w584 = (~w565 & w3782) | (~w565 & w3783) | (w3782 & w3783);
assign w585 = pi270 & ~pi398;
assign w586 = pi269 & ~pi397;
assign w587 = pi268 & ~pi396;
assign w588 = ~w586 & ~w587;
assign w589 = w580 & ~w588;
assign w590 = pi271 & ~pi399;
assign w591 = ~w585 & ~w590;
assign w592 = ~w589 & w591;
assign w593 = ~pi271 & pi399;
assign w594 = ~pi272 & pi400;
assign w595 = ~w593 & ~w594;
assign w596 = (~w584 & w3934) | (~w584 & w3935) | (w3934 & w3935);
assign w597 = ~pi274 & pi402;
assign w598 = ~pi273 & pi401;
assign w599 = ~w597 & ~w598;
assign w600 = pi275 & ~pi403;
assign w601 = pi274 & ~pi402;
assign w602 = pi273 & ~pi401;
assign w603 = ~w597 & w602;
assign w604 = ~w600 & ~w601;
assign w605 = ~w603 & w604;
assign w606 = ~pi275 & pi403;
assign w607 = ~pi278 & pi406;
assign w608 = ~pi277 & pi405;
assign w609 = ~pi276 & pi404;
assign w610 = ~w606 & ~w607;
assign w611 = ~w608 & ~w609;
assign w612 = w610 & w611;
assign w613 = pi278 & ~pi406;
assign w614 = pi279 & ~pi407;
assign w615 = pi277 & ~pi405;
assign w616 = pi276 & ~pi404;
assign w617 = ~w608 & w616;
assign w618 = (~w607 & w617) | (~w607 & w3993) | (w617 & w3993);
assign w619 = ~w613 & ~w614;
assign w620 = ~w618 & w619;
assign w621 = ~pi279 & pi407;
assign w622 = ~pi280 & pi408;
assign w623 = ~w621 & ~w622;
assign w624 = (~w596 & w3986) | (~w596 & w3987) | (w3986 & w3987);
assign w625 = ~pi282 & pi410;
assign w626 = ~pi281 & pi409;
assign w627 = ~w625 & ~w626;
assign w628 = pi283 & ~pi411;
assign w629 = pi282 & ~pi410;
assign w630 = pi281 & ~pi409;
assign w631 = ~w625 & w630;
assign w632 = ~w628 & ~w629;
assign w633 = ~w631 & w632;
assign w634 = ~pi285 & pi413;
assign w635 = ~pi284 & pi412;
assign w636 = ~pi283 & pi411;
assign w637 = ~w634 & ~w635;
assign w638 = ~w636 & w637;
assign w639 = pi286 & ~pi414;
assign w640 = pi285 & ~pi413;
assign w641 = pi284 & ~pi412;
assign w642 = ~w634 & w641;
assign w643 = ~w639 & ~w640;
assign w644 = ~w642 & w643;
assign w645 = ~pi292 & pi420;
assign w646 = ~pi295 & pi423;
assign w647 = ~pi294 & pi422;
assign w648 = ~pi293 & pi421;
assign w649 = ~w646 & ~w647;
assign w650 = ~w648 & w649;
assign w651 = ~pi289 & pi417;
assign w652 = ~pi416 & ~w651;
assign w653 = pi288 & ~w651;
assign w654 = ~w652 & ~w653;
assign w655 = ~pi291 & pi419;
assign w656 = ~pi290 & pi418;
assign w657 = ~w655 & ~w656;
assign w658 = ~pi286 & pi414;
assign w659 = ~pi287 & pi415;
assign w660 = ~w645 & ~w658;
assign w661 = ~w659 & w660;
assign w662 = w657 & w661;
assign w663 = w650 & ~w654;
assign w664 = w662 & w663;
assign w665 = (w624 & w4011) | (w624 & w4012) | (w4011 & w4012);
assign w666 = pi294 & ~pi422;
assign w667 = ~w646 & w666;
assign w668 = ~pi303 & pi431;
assign w669 = pi302 & ~pi430;
assign w670 = ~w668 & w669;
assign w671 = pi303 & ~pi431;
assign w672 = ~pi302 & pi430;
assign w673 = ~pi301 & pi429;
assign w674 = ~w668 & ~w672;
assign w675 = ~w673 & w674;
assign w676 = pi300 & ~pi428;
assign w677 = pi301 & ~pi429;
assign w678 = ~pi300 & pi428;
assign w679 = pi299 & ~pi427;
assign w680 = ~pi299 & pi427;
assign w681 = ~pi298 & pi426;
assign w682 = ~w680 & ~w681;
assign w683 = pi298 & ~pi426;
assign w684 = pi297 & ~pi425;
assign w685 = ~pi297 & pi425;
assign w686 = pi296 & ~pi424;
assign w687 = ~w685 & w686;
assign w688 = ~w683 & ~w684;
assign w689 = ~w687 & w688;
assign w690 = (~w679 & w689) | (~w679 & w4002) | (w689 & w4002);
assign w691 = ~w676 & ~w677;
assign w692 = (~w690 & w4029) | (~w690 & w4030) | (w4029 & w4030);
assign w693 = ~w670 & ~w671;
assign w694 = ~w692 & w693;
assign w695 = pi295 & ~pi423;
assign w696 = pi292 & ~pi420;
assign w697 = pi293 & ~pi421;
assign w698 = pi291 & ~pi419;
assign w699 = pi290 & ~pi418;
assign w700 = pi289 & ~pi417;
assign w701 = ~w651 & w4003;
assign w702 = pi287 & ~pi415;
assign w703 = ~w654 & w702;
assign w704 = ~w699 & ~w700;
assign w705 = ~w701 & w704;
assign w706 = (w657 & w703) | (w657 & w4004) | (w703 & w4004);
assign w707 = ~w696 & ~w697;
assign w708 = (w706 & w4047) | (w706 & w4048) | (w4047 & w4048);
assign w709 = ~w667 & ~w695;
assign w710 = ~w692 & w4049;
assign w711 = ~w708 & w710;
assign w712 = ~pi296 & pi424;
assign w713 = ~w678 & ~w685;
assign w714 = ~w712 & w713;
assign w715 = w682 & w714;
assign w716 = w675 & w715;
assign w717 = w694 & ~w716;
assign w718 = ~pi315 & pi443;
assign w719 = ~pi314 & pi442;
assign w720 = ~w718 & ~w719;
assign w721 = ~pi313 & pi441;
assign w722 = ~pi312 & pi440;
assign w723 = ~w721 & ~w722;
assign w724 = w720 & w723;
assign w725 = ~pi307 & pi435;
assign w726 = ~pi306 & pi434;
assign w727 = ~w725 & ~w726;
assign w728 = ~pi310 & pi438;
assign w729 = ~pi311 & pi439;
assign w730 = ~w728 & ~w729;
assign w731 = ~pi309 & pi437;
assign w732 = ~pi308 & pi436;
assign w733 = ~w731 & ~w732;
assign w734 = ~pi305 & pi433;
assign w735 = ~pi316 & pi444;
assign w736 = ~pi319 & pi447;
assign w737 = ~pi318 & pi446;
assign w738 = ~pi317 & pi445;
assign w739 = ~w736 & ~w737;
assign w740 = ~w738 & w739;
assign w741 = ~w735 & w740;
assign w742 = ~pi304 & pi432;
assign w743 = ~w734 & ~w742;
assign w744 = w727 & w743;
assign w745 = w730 & w733;
assign w746 = w744 & w745;
assign w747 = w724 & w746;
assign w748 = w741 & w747;
assign w749 = ~w717 & w748;
assign w750 = (w749 & w665) | (w749 & w4033) | (w665 & w4033);
assign w751 = pi319 & ~pi447;
assign w752 = pi313 & ~pi441;
assign w753 = pi314 & ~pi442;
assign w754 = pi312 & ~pi440;
assign w755 = ~w721 & w754;
assign w756 = ~w752 & ~w753;
assign w757 = ~w755 & w756;
assign w758 = pi315 & ~pi443;
assign w759 = pi311 & ~pi439;
assign w760 = pi310 & ~pi438;
assign w761 = pi309 & ~pi437;
assign w762 = pi307 & ~pi435;
assign w763 = pi308 & ~pi436;
assign w764 = pi306 & ~pi434;
assign w765 = pi305 & ~pi433;
assign w766 = pi304 & ~pi432;
assign w767 = ~w734 & w766;
assign w768 = ~w764 & ~w765;
assign w769 = ~w767 & w768;
assign w770 = ~w762 & ~w763;
assign w771 = (w770 & w769) | (w770 & w4005) | (w769 & w4005);
assign w772 = ~w760 & ~w761;
assign w773 = (~w771 & w4015) | (~w771 & w4016) | (w4015 & w4016);
assign w774 = (w724 & w773) | (w724 & w4017) | (w773 & w4017);
assign w775 = (~w758 & w757) | (~w758 & w4050) | (w757 & w4050);
assign w776 = (w741 & w774) | (w741 & w4034) | (w774 & w4034);
assign w777 = pi323 & ~pi451;
assign w778 = ~pi323 & pi451;
assign w779 = ~pi322 & pi450;
assign w780 = ~w778 & ~w779;
assign w781 = pi321 & ~pi449;
assign w782 = pi322 & ~pi450;
assign w783 = ~pi321 & pi449;
assign w784 = pi320 & ~pi448;
assign w785 = ~w783 & w784;
assign w786 = ~w781 & ~w782;
assign w787 = ~w785 & w786;
assign w788 = w780 & ~w787;
assign w789 = ~w777 & ~w788;
assign w790 = pi317 & ~pi445;
assign w791 = pi316 & ~pi444;
assign w792 = ~w790 & ~w791;
assign w793 = w740 & ~w792;
assign w794 = pi318 & ~pi446;
assign w795 = ~w736 & w794;
assign w796 = ~w751 & ~w795;
assign w797 = ~w793 & w796;
assign w798 = w789 & w797;
assign w799 = ~w776 & w798;
assign w800 = ~pi331 & pi459;
assign w801 = ~pi330 & pi458;
assign w802 = ~w800 & ~w801;
assign w803 = ~pi320 & pi448;
assign w804 = ~w783 & ~w803;
assign w805 = w780 & w804;
assign w806 = w789 & ~w805;
assign w807 = ~pi326 & pi454;
assign w808 = ~pi325 & pi453;
assign w809 = ~w807 & ~w808;
assign w810 = ~pi324 & pi452;
assign w811 = ~pi327 & pi455;
assign w812 = ~pi329 & pi457;
assign w813 = ~pi328 & pi456;
assign w814 = ~w811 & ~w812;
assign w815 = ~w813 & w814;
assign w816 = w802 & ~w810;
assign w817 = w809 & w816;
assign w818 = w815 & w817;
assign w819 = ~w806 & w818;
assign w820 = pi331 & ~pi459;
assign w821 = pi326 & ~pi454;
assign w822 = pi327 & ~pi455;
assign w823 = pi325 & ~pi453;
assign w824 = pi324 & ~pi452;
assign w825 = ~w823 & ~w824;
assign w826 = w809 & ~w825;
assign w827 = ~w821 & ~w822;
assign w828 = ~w826 & w827;
assign w829 = w815 & ~w828;
assign w830 = pi330 & ~pi458;
assign w831 = pi329 & ~pi457;
assign w832 = pi328 & ~pi456;
assign w833 = ~w812 & w832;
assign w834 = ~w830 & ~w831;
assign w835 = ~w833 & w834;
assign w836 = ~w829 & w835;
assign w837 = w802 & ~w836;
assign w838 = pi335 & ~pi463;
assign w839 = pi333 & ~pi461;
assign w840 = pi332 & ~pi460;
assign w841 = ~w839 & ~w840;
assign w842 = ~pi335 & pi463;
assign w843 = ~pi334 & pi462;
assign w844 = ~pi333 & pi461;
assign w845 = ~w842 & ~w843;
assign w846 = ~w844 & w845;
assign w847 = ~w841 & w846;
assign w848 = pi334 & ~pi462;
assign w849 = ~w842 & w848;
assign w850 = ~w838 & ~w849;
assign w851 = ~w847 & w850;
assign w852 = ~w820 & w851;
assign w853 = ~w837 & w852;
assign w854 = (~w750 & w4018) | (~w750 & w4019) | (w4018 & w4019);
assign w855 = ~pi336 & pi464;
assign w856 = ~pi332 & pi460;
assign w857 = w846 & ~w856;
assign w858 = w851 & ~w857;
assign w859 = ~pi337 & pi465;
assign w860 = ~pi338 & pi466;
assign w861 = ~pi340 & pi468;
assign w862 = ~pi342 & pi470;
assign w863 = ~pi343 & pi471;
assign w864 = ~pi341 & pi469;
assign w865 = ~w862 & ~w863;
assign w866 = ~w864 & w865;
assign w867 = w865 & w4060;
assign w868 = ~pi339 & pi467;
assign w869 = ~w860 & ~w868;
assign w870 = w867 & w869;
assign w871 = ~w855 & ~w859;
assign w872 = w870 & w871;
assign w873 = ~w858 & w872;
assign w874 = pi343 & ~pi471;
assign w875 = pi338 & ~pi466;
assign w876 = pi337 & ~pi465;
assign w877 = pi336 & ~pi464;
assign w878 = ~w859 & w877;
assign w879 = ~w875 & ~w876;
assign w880 = ~w878 & w879;
assign w881 = w870 & ~w880;
assign w882 = pi339 & ~pi467;
assign w883 = w867 & w882;
assign w884 = pi347 & ~pi475;
assign w885 = ~pi347 & pi475;
assign w886 = ~pi346 & pi474;
assign w887 = ~w885 & ~w886;
assign w888 = pi345 & ~pi473;
assign w889 = pi346 & ~pi474;
assign w890 = ~pi345 & pi473;
assign w891 = pi344 & ~pi472;
assign w892 = ~w890 & w891;
assign w893 = ~w888 & ~w889;
assign w894 = ~w892 & w893;
assign w895 = (~w884 & w894) | (~w884 & w4071) | (w894 & w4071);
assign w896 = pi341 & ~pi469;
assign w897 = pi340 & ~pi468;
assign w898 = ~w896 & ~w897;
assign w899 = w866 & ~w898;
assign w900 = pi342 & ~pi470;
assign w901 = ~w863 & w900;
assign w902 = ~w874 & ~w901;
assign w903 = ~w899 & w902;
assign w904 = ~w883 & w903;
assign w905 = w904 & w4061;
assign w906 = ~pi355 & pi483;
assign w907 = ~pi354 & pi482;
assign w908 = ~w906 & ~w907;
assign w909 = ~pi344 & pi472;
assign w910 = ~w890 & ~w909;
assign w911 = w887 & w910;
assign w912 = w895 & ~w911;
assign w913 = ~pi350 & pi478;
assign w914 = ~pi349 & pi477;
assign w915 = ~w913 & ~w914;
assign w916 = ~pi348 & pi476;
assign w917 = ~pi351 & pi479;
assign w918 = ~pi353 & pi481;
assign w919 = ~pi352 & pi480;
assign w920 = ~w917 & ~w918;
assign w921 = ~w919 & w920;
assign w922 = w908 & ~w916;
assign w923 = w915 & w922;
assign w924 = w921 & w923;
assign w925 = ~w912 & w924;
assign w926 = pi355 & ~pi483;
assign w927 = pi350 & ~pi478;
assign w928 = pi351 & ~pi479;
assign w929 = pi349 & ~pi477;
assign w930 = pi348 & ~pi476;
assign w931 = ~w929 & ~w930;
assign w932 = w915 & ~w931;
assign w933 = ~w927 & ~w928;
assign w934 = ~w932 & w933;
assign w935 = w921 & ~w934;
assign w936 = pi353 & ~pi481;
assign w937 = pi354 & ~pi482;
assign w938 = pi352 & ~pi480;
assign w939 = ~w918 & w938;
assign w940 = ~w936 & ~w937;
assign w941 = ~w939 & w940;
assign w942 = ~w935 & w941;
assign w943 = w908 & ~w942;
assign w944 = pi359 & ~pi487;
assign w945 = pi357 & ~pi485;
assign w946 = pi356 & ~pi484;
assign w947 = ~w945 & ~w946;
assign w948 = ~pi359 & pi487;
assign w949 = ~pi358 & pi486;
assign w950 = ~pi357 & pi485;
assign w951 = ~w948 & ~w949;
assign w952 = ~w950 & w951;
assign w953 = ~w947 & w952;
assign w954 = pi358 & ~pi486;
assign w955 = ~w948 & w954;
assign w956 = ~w944 & ~w955;
assign w957 = ~w953 & w956;
assign w958 = ~w926 & w957;
assign w959 = ~w943 & w958;
assign w960 = ~pi360 & pi488;
assign w961 = ~pi356 & pi484;
assign w962 = w952 & ~w961;
assign w963 = w957 & ~w962;
assign w964 = ~pi361 & pi489;
assign w965 = ~pi362 & pi490;
assign w966 = ~pi364 & pi492;
assign w967 = ~pi366 & pi494;
assign w968 = ~pi367 & pi495;
assign w969 = ~pi365 & pi493;
assign w970 = ~w967 & ~w968;
assign w971 = ~w969 & w970;
assign w972 = w970 & w4091;
assign w973 = ~pi363 & pi491;
assign w974 = ~w965 & ~w973;
assign w975 = w972 & w974;
assign w976 = ~w960 & ~w964;
assign w977 = w975 & w976;
assign w978 = ~w963 & w977;
assign w979 = (~w854 & w4062) | (~w854 & w4063) | (w4062 & w4063);
assign w980 = pi367 & ~pi495;
assign w981 = pi362 & ~pi490;
assign w982 = pi361 & ~pi489;
assign w983 = pi360 & ~pi488;
assign w984 = ~w964 & w983;
assign w985 = ~w981 & ~w982;
assign w986 = ~w984 & w985;
assign w987 = w975 & ~w986;
assign w988 = pi363 & ~pi491;
assign w989 = w972 & w988;
assign w990 = pi371 & ~pi499;
assign w991 = ~pi371 & pi499;
assign w992 = ~pi370 & pi498;
assign w993 = ~w991 & ~w992;
assign w994 = pi369 & ~pi497;
assign w995 = pi370 & ~pi498;
assign w996 = ~pi369 & pi497;
assign w997 = pi368 & ~pi496;
assign w998 = ~w996 & w997;
assign w999 = ~w994 & ~w995;
assign w1000 = ~w998 & w999;
assign w1001 = w993 & ~w1000;
assign w1002 = ~w990 & ~w1001;
assign w1003 = pi365 & ~pi493;
assign w1004 = pi364 & ~pi492;
assign w1005 = ~w1003 & ~w1004;
assign w1006 = w971 & ~w1005;
assign w1007 = pi366 & ~pi494;
assign w1008 = ~w968 & w1007;
assign w1009 = ~w980 & ~w1008;
assign w1010 = ~w1006 & w1009;
assign w1011 = ~w989 & w1010;
assign w1012 = w1011 & w4092;
assign w1013 = ~pi368 & pi496;
assign w1014 = ~w996 & ~w1013;
assign w1015 = w993 & w1014;
assign w1016 = w1002 & ~w1015;
assign w1017 = ~pi375 & pi503;
assign w1018 = ~pi376 & pi504;
assign w1019 = ~w1017 & ~w1018;
assign w1020 = ~pi372 & pi500;
assign w1021 = ~pi374 & pi502;
assign w1022 = ~pi373 & pi501;
assign w1023 = ~w1021 & ~w1022;
assign w1024 = ~pi379 & pi507;
assign w1025 = ~pi378 & pi506;
assign w1026 = ~pi377 & pi505;
assign w1027 = ~w1025 & ~w1026;
assign w1028 = ~w1020 & ~w1024;
assign w1029 = w1019 & w1028;
assign w1030 = w1023 & w1027;
assign w1031 = w1029 & w1030;
assign w1032 = ~w1016 & w1031;
assign w1033 = pi379 & ~pi507;
assign w1034 = pi377 & ~pi505;
assign w1035 = pi375 & ~pi503;
assign w1036 = pi373 & ~pi501;
assign w1037 = pi372 & ~pi500;
assign w1038 = ~w1036 & ~w1037;
assign w1039 = w1023 & ~w1038;
assign w1040 = pi374 & ~pi502;
assign w1041 = ~w1035 & ~w1040;
assign w1042 = (w1019 & w1039) | (w1019 & w4081) | (w1039 & w4081);
assign w1043 = pi376 & ~pi504;
assign w1044 = ~w1034 & ~w1043;
assign w1045 = (w1027 & w1042) | (w1027 & w4093) | (w1042 & w4093);
assign w1046 = pi378 & ~pi506;
assign w1047 = ~w1045 & ~w1046;
assign w1048 = ~w1024 & ~w1047;
assign w1049 = ~w1033 & ~w1048;
assign w1050 = ~pi380 & pi508;
assign w1051 = pi383 & ~pi511;
assign w1052 = ~pi382 & pi510;
assign w1053 = ~pi381 & pi509;
assign w1054 = ~w1051 & ~w1052;
assign w1055 = ~w1053 & w1054;
assign w1056 = ~w1050 & w1055;
assign w1057 = pi381 & ~pi509;
assign w1058 = pi380 & ~pi508;
assign w1059 = ~w1057 & ~w1058;
assign w1060 = w1055 & ~w1059;
assign w1061 = pi382 & ~pi510;
assign w1062 = ~w1051 & w1061;
assign w1063 = ~w1060 & ~w1062;
assign w1064 = w1063 & w4204;
assign w1065 = ~pi511 & w1064;
assign w1066 = pi383 & ~w1065;
assign w1067 = ~pi255 & w532;
assign w1068 = pi127 & ~w1067;
assign w1069 = ~w1066 & w1068;
assign w1070 = (pi010 & ~w532) | (pi010 & w3058) | (~w532 & w3058);
assign w1071 = w532 & w3059;
assign w1072 = ~w1070 & ~w1071;
assign w1073 = ~pi383 & pi511;
assign w1074 = (~w979 & w4094) | (~w979 & w4095) | (w4094 & w4095);
assign w1075 = pi266 & ~w1074;
assign w1076 = pi394 & w1074;
assign w1077 = ~w1075 & ~w1076;
assign w1078 = w1072 & ~w1077;
assign w1079 = pi009 & ~w534;
assign w1080 = pi137 & w534;
assign w1081 = ~w1079 & ~w1080;
assign w1082 = pi265 & ~w1074;
assign w1083 = pi393 & w1074;
assign w1084 = ~w1082 & ~w1083;
assign w1085 = ~w1081 & w1084;
assign w1086 = pi007 & ~w534;
assign w1087 = pi135 & w534;
assign w1088 = ~w1086 & ~w1087;
assign w1089 = pi263 & ~w1074;
assign w1090 = pi391 & w1074;
assign w1091 = ~w1089 & ~w1090;
assign w1092 = w1088 & ~w1091;
assign w1093 = pi006 & ~w534;
assign w1094 = pi134 & w534;
assign w1095 = ~w1093 & ~w1094;
assign w1096 = pi262 & ~w1074;
assign w1097 = pi390 & w1074;
assign w1098 = ~w1096 & ~w1097;
assign w1099 = ~w1095 & w1098;
assign w1100 = (pi001 & ~w532) | (pi001 & w2745) | (~w532 & w2745);
assign w1101 = w532 & w2746;
assign w1102 = ~w1100 & ~w1101;
assign w1103 = pi257 & ~w1074;
assign w1104 = pi385 & w1074;
assign w1105 = ~w1103 & ~w1104;
assign w1106 = ~w1102 & w1105;
assign w1107 = pi256 & ~w1074;
assign w1108 = pi384 & w1074;
assign w1109 = ~w1107 & ~w1108;
assign w1110 = ~w537 & w1109;
assign w1111 = ~w1106 & ~w1110;
assign w1112 = w1102 & ~w1105;
assign w1113 = (pi002 & ~w532) | (pi002 & w2747) | (~w532 & w2747);
assign w1114 = w532 & w2748;
assign w1115 = ~w1113 & ~w1114;
assign w1116 = pi258 & ~w1074;
assign w1117 = pi386 & w1074;
assign w1118 = ~w1116 & ~w1117;
assign w1119 = w1115 & ~w1118;
assign w1120 = ~w1112 & ~w1119;
assign w1121 = ~w1111 & w1120;
assign w1122 = (pi003 & ~w532) | (pi003 & w3060) | (~w532 & w3060);
assign w1123 = w532 & w3061;
assign w1124 = ~w1122 & ~w1123;
assign w1125 = pi259 & ~w1074;
assign w1126 = pi387 & w1074;
assign w1127 = ~w1125 & ~w1126;
assign w1128 = ~w1124 & w1127;
assign w1129 = ~w1115 & w1118;
assign w1130 = ~w1128 & ~w1129;
assign w1131 = (pi004 & ~w532) | (pi004 & w3062) | (~w532 & w3062);
assign w1132 = w532 & w3063;
assign w1133 = ~w1131 & ~w1132;
assign w1134 = pi260 & ~w1074;
assign w1135 = pi388 & w1074;
assign w1136 = ~w1134 & ~w1135;
assign w1137 = w1133 & ~w1136;
assign w1138 = w1124 & ~w1127;
assign w1139 = ~w1137 & ~w1138;
assign w1140 = (w1139 & w1121) | (w1139 & w2749) | (w1121 & w2749);
assign w1141 = ~w1133 & w1136;
assign w1142 = pi005 & ~w534;
assign w1143 = pi133 & w534;
assign w1144 = ~w1142 & ~w1143;
assign w1145 = pi261 & ~w1074;
assign w1146 = pi389 & w1074;
assign w1147 = ~w1145 & ~w1146;
assign w1148 = ~w1144 & w1147;
assign w1149 = ~w1141 & ~w1148;
assign w1150 = w1095 & ~w1098;
assign w1151 = w1144 & ~w1147;
assign w1152 = ~w1150 & ~w1151;
assign w1153 = (w1152 & w1140) | (w1152 & w2750) | (w1140 & w2750);
assign w1154 = pi264 & ~w1074;
assign w1155 = pi392 & w1074;
assign w1156 = ~w1154 & ~w1155;
assign w1157 = pi008 & ~w534;
assign w1158 = pi136 & w534;
assign w1159 = ~w1157 & ~w1158;
assign w1160 = w1156 & ~w1159;
assign w1161 = ~w1088 & w1091;
assign w1162 = ~w1160 & ~w1161;
assign w1163 = ~w1156 & w1159;
assign w1164 = w1081 & ~w1084;
assign w1165 = ~w1163 & ~w1164;
assign w1166 = (w1153 & w2754) | (w1153 & w2755) | (w2754 & w2755);
assign w1167 = (pi011 & ~w532) | (pi011 & w3064) | (~w532 & w3064);
assign w1168 = w532 & w3065;
assign w1169 = ~w1167 & ~w1168;
assign w1170 = pi267 & ~w1074;
assign w1171 = pi395 & w1074;
assign w1172 = ~w1170 & ~w1171;
assign w1173 = ~w1169 & w1172;
assign w1174 = ~w1072 & w1077;
assign w1175 = ~w1173 & ~w1174;
assign w1176 = (pi013 & ~w532) | (pi013 & w3066) | (~w532 & w3066);
assign w1177 = w532 & w3067;
assign w1178 = ~w1176 & ~w1177;
assign w1179 = pi269 & ~w1074;
assign w1180 = pi397 & w1074;
assign w1181 = ~w1179 & ~w1180;
assign w1182 = w1178 & ~w1181;
assign w1183 = pi268 & ~w1074;
assign w1184 = pi396 & w1074;
assign w1185 = ~w1183 & ~w1184;
assign w1186 = (pi012 & ~w532) | (pi012 & w3068) | (~w532 & w3068);
assign w1187 = w532 & w3069;
assign w1188 = ~w1186 & ~w1187;
assign w1189 = ~w1185 & w1188;
assign w1190 = w1169 & ~w1172;
assign w1191 = ~w1182 & ~w1189;
assign w1192 = ~w1190 & w1191;
assign w1193 = ~w1178 & w1181;
assign w1194 = pi014 & ~w534;
assign w1195 = pi142 & w534;
assign w1196 = ~w1194 & ~w1195;
assign w1197 = pi270 & ~w1074;
assign w1198 = pi398 & w1074;
assign w1199 = ~w1197 & ~w1198;
assign w1200 = ~w1196 & w1199;
assign w1201 = w1185 & ~w1188;
assign w1202 = ~w1182 & w1201;
assign w1203 = ~w1193 & ~w1200;
assign w1204 = ~w1202 & w1203;
assign w1205 = (pi015 & ~w532) | (pi015 & w3785) | (~w532 & w3785);
assign w1206 = w532 & w3786;
assign w1207 = ~w1205 & ~w1206;
assign w1208 = pi271 & ~w1074;
assign w1209 = pi399 & w1074;
assign w1210 = ~w1208 & ~w1209;
assign w1211 = w1207 & ~w1210;
assign w1212 = w1196 & ~w1199;
assign w1213 = ~w1211 & ~w1212;
assign w1214 = (w1166 & w2762) | (w1166 & w2763) | (w2762 & w2763);
assign w1215 = ~w1207 & w1210;
assign w1216 = (w524 & w3787) | (w524 & w3788) | (w3787 & w3788);
assign w1217 = ~w524 & w3789;
assign w1218 = ~w1216 & ~w1217;
assign w1219 = pi272 & ~w1074;
assign w1220 = pi400 & w1074;
assign w1221 = ~w1219 & ~w1220;
assign w1222 = ~w1218 & w1221;
assign w1223 = ~w1215 & ~w1222;
assign w1224 = w1218 & ~w1221;
assign w1225 = (w524 & w3790) | (w524 & w3791) | (w3790 & w3791);
assign w1226 = ~w524 & w3792;
assign w1227 = ~w1225 & ~w1226;
assign w1228 = pi274 & ~w1074;
assign w1229 = pi402 & w1074;
assign w1230 = ~w1228 & ~w1229;
assign w1231 = w1227 & ~w1230;
assign w1232 = (w524 & w3793) | (w524 & w3794) | (w3793 & w3794);
assign w1233 = ~w524 & w3795;
assign w1234 = ~w1232 & ~w1233;
assign w1235 = pi273 & ~w1074;
assign w1236 = pi401 & w1074;
assign w1237 = ~w1235 & ~w1236;
assign w1238 = w1234 & ~w1237;
assign w1239 = ~w1224 & ~w1231;
assign w1240 = ~w1238 & w1239;
assign w1241 = (w524 & w3796) | (w524 & w3797) | (w3796 & w3797);
assign w1242 = ~w524 & w3798;
assign w1243 = ~w1241 & ~w1242;
assign w1244 = pi275 & ~w1074;
assign w1245 = pi403 & w1074;
assign w1246 = ~w1244 & ~w1245;
assign w1247 = ~w1243 & w1246;
assign w1248 = ~w1227 & w1230;
assign w1249 = ~w1234 & w1237;
assign w1250 = ~w1231 & w1249;
assign w1251 = ~w1247 & ~w1248;
assign w1252 = ~w1250 & w1251;
assign w1253 = w1243 & ~w1246;
assign w1254 = (w524 & w3799) | (w524 & w3800) | (w3799 & w3800);
assign w1255 = ~w524 & w3801;
assign w1256 = ~w1254 & ~w1255;
assign w1257 = pi277 & ~w1074;
assign w1258 = pi405 & w1074;
assign w1259 = ~w1257 & ~w1258;
assign w1260 = w1256 & ~w1259;
assign w1261 = (pi020 & ~w532) | (pi020 & w3802) | (~w532 & w3802);
assign w1262 = w532 & w3803;
assign w1263 = ~w1261 & ~w1262;
assign w1264 = pi276 & ~w1074;
assign w1265 = pi404 & w1074;
assign w1266 = ~w1264 & ~w1265;
assign w1267 = w1263 & ~w1266;
assign w1268 = ~w1253 & ~w1260;
assign w1269 = ~w1267 & w1268;
assign w1270 = (w524 & w3804) | (w524 & w3805) | (w3804 & w3805);
assign w1271 = ~w524 & w3806;
assign w1272 = ~w1270 & ~w1271;
assign w1273 = pi278 & ~w1074;
assign w1274 = pi406 & w1074;
assign w1275 = ~w1273 & ~w1274;
assign w1276 = ~w1272 & w1275;
assign w1277 = ~w1256 & w1259;
assign w1278 = ~w1263 & w1266;
assign w1279 = ~w1260 & w1278;
assign w1280 = ~w1276 & ~w1277;
assign w1281 = ~w1279 & w1280;
assign w1282 = (w524 & w3807) | (w524 & w3808) | (w3807 & w3808);
assign w1283 = ~w524 & w3809;
assign w1284 = ~w1282 & ~w1283;
assign w1285 = pi279 & ~w1074;
assign w1286 = pi407 & w1074;
assign w1287 = ~w1285 & ~w1286;
assign w1288 = w1284 & ~w1287;
assign w1289 = w1272 & ~w1275;
assign w1290 = ~w1288 & ~w1289;
assign w1291 = (w524 & w3810) | (w524 & w3811) | (w3810 & w3811);
assign w1292 = ~w524 & w3812;
assign w1293 = ~w1291 & ~w1292;
assign w1294 = pi280 & ~w1074;
assign w1295 = pi408 & w1074;
assign w1296 = ~w1294 & ~w1295;
assign w1297 = ~w1293 & w1296;
assign w1298 = ~w1284 & w1287;
assign w1299 = ~w1297 & ~w1298;
assign w1300 = (w524 & w3813) | (w524 & w3814) | (w3813 & w3814);
assign w1301 = ~w524 & w3815;
assign w1302 = ~w1300 & ~w1301;
assign w1303 = pi282 & ~w1074;
assign w1304 = pi410 & w1074;
assign w1305 = ~w1303 & ~w1304;
assign w1306 = w1302 & ~w1305;
assign w1307 = (w524 & w3816) | (w524 & w3817) | (w3816 & w3817);
assign w1308 = ~w524 & w3818;
assign w1309 = ~w1307 & ~w1308;
assign w1310 = pi281 & ~w1074;
assign w1311 = pi409 & w1074;
assign w1312 = ~w1310 & ~w1311;
assign w1313 = w1309 & ~w1312;
assign w1314 = w1293 & ~w1296;
assign w1315 = ~w1306 & ~w1313;
assign w1316 = ~w1314 & w1315;
assign w1317 = (pi027 & ~w532) | (pi027 & w3819) | (~w532 & w3819);
assign w1318 = w532 & w3820;
assign w1319 = ~w1317 & ~w1318;
assign w1320 = pi283 & ~w1074;
assign w1321 = pi411 & w1074;
assign w1322 = ~w1320 & ~w1321;
assign w1323 = ~w1319 & w1322;
assign w1324 = ~w1302 & w1305;
assign w1325 = ~w1309 & w1312;
assign w1326 = ~w1306 & w1325;
assign w1327 = ~w1323 & ~w1324;
assign w1328 = ~w1326 & w1327;
assign w1329 = w1319 & ~w1322;
assign w1330 = (pi029 & ~w532) | (pi029 & w3821) | (~w532 & w3821);
assign w1331 = w532 & w3822;
assign w1332 = ~w1330 & ~w1331;
assign w1333 = pi285 & ~w1074;
assign w1334 = pi413 & w1074;
assign w1335 = ~w1333 & ~w1334;
assign w1336 = w1332 & ~w1335;
assign w1337 = pi028 & ~w534;
assign w1338 = pi156 & w534;
assign w1339 = ~w1337 & ~w1338;
assign w1340 = pi284 & ~w1074;
assign w1341 = pi412 & w1074;
assign w1342 = ~w1340 & ~w1341;
assign w1343 = w1339 & ~w1342;
assign w1344 = ~w1329 & ~w1336;
assign w1345 = ~w1343 & w1344;
assign w1346 = pi030 & ~w534;
assign w1347 = pi158 & w534;
assign w1348 = ~w1346 & ~w1347;
assign w1349 = pi286 & ~w1074;
assign w1350 = pi414 & w1074;
assign w1351 = ~w1349 & ~w1350;
assign w1352 = ~w1348 & w1351;
assign w1353 = ~w1332 & w1335;
assign w1354 = ~w1339 & w1342;
assign w1355 = ~w1336 & w1354;
assign w1356 = ~w1352 & ~w1353;
assign w1357 = ~w1355 & w1356;
assign w1358 = (w389 & w4096) | (w389 & w4097) | (w4096 & w4097);
assign w1359 = (~w389 & w4098) | (~w389 & w4099) | (w4098 & w4099);
assign w1360 = ~w1358 & ~w1359;
assign w1361 = (w979 & w4100) | (w979 & w4101) | (w4100 & w4101);
assign w1362 = (~w979 & w4102) | (~w979 & w4103) | (w4102 & w4103);
assign w1363 = ~w1361 & ~w1362;
assign w1364 = w1360 & ~w1363;
assign w1365 = pi290 & ~w1074;
assign w1366 = pi418 & w1074;
assign w1367 = ~w1365 & ~w1366;
assign w1368 = (~w516 & w3941) | (~w516 & w3942) | (w3941 & w3942);
assign w1369 = (w3826 & w516) | (w3826 & w3943) | (w516 & w3943);
assign w1370 = ~w1368 & ~w1369;
assign w1371 = ~w1367 & w1370;
assign w1372 = ~w1364 & ~w1371;
assign w1373 = pi294 & ~w1074;
assign w1374 = pi422 & w1074;
assign w1375 = ~w1373 & ~w1374;
assign w1376 = pi038 & ~w534;
assign w1377 = pi166 & w534;
assign w1378 = ~w1376 & ~w1377;
assign w1379 = ~w1375 & w1378;
assign w1380 = (pi037 & ~w532) | (pi037 & w3944) | (~w532 & w3944);
assign w1381 = w532 & w3945;
assign w1382 = ~w1380 & ~w1381;
assign w1383 = pi293 & ~w1074;
assign w1384 = pi421 & w1074;
assign w1385 = ~w1383 & ~w1384;
assign w1386 = w1382 & ~w1385;
assign w1387 = ~w1379 & ~w1386;
assign w1388 = (~w516 & w3946) | (~w516 & w3947) | (w3946 & w3947);
assign w1389 = (w3827 & w516) | (w3827 & w3948) | (w516 & w3948);
assign w1390 = ~w1388 & ~w1389;
assign w1391 = pi292 & ~w1074;
assign w1392 = pi420 & w1074;
assign w1393 = ~w1391 & ~w1392;
assign w1394 = w1390 & ~w1393;
assign w1395 = (~w516 & w3949) | (~w516 & w3950) | (w3949 & w3950);
assign w1396 = (w3828 & w516) | (w3828 & w3951) | (w516 & w3951);
assign w1397 = ~w1395 & ~w1396;
assign w1398 = pi291 & ~w1074;
assign w1399 = pi419 & w1074;
assign w1400 = ~w1398 & ~w1399;
assign w1401 = w1397 & ~w1400;
assign w1402 = ~w1394 & ~w1401;
assign w1403 = w1348 & ~w1351;
assign w1404 = pi039 & ~w534;
assign w1405 = pi167 & w534;
assign w1406 = ~w1404 & ~w1405;
assign w1407 = pi295 & ~w1074;
assign w1408 = pi423 & w1074;
assign w1409 = ~w1407 & ~w1408;
assign w1410 = w1406 & ~w1409;
assign w1411 = (w979 & w4104) | (w979 & w4105) | (w4104 & w4105);
assign w1412 = (~w979 & w4106) | (~w979 & w4107) | (w4106 & w4107);
assign w1413 = ~w1411 & ~w1412;
assign w1414 = (w389 & w4108) | (w389 & w4109) | (w4108 & w4109);
assign w1415 = (~w389 & w4110) | (~w389 & w4111) | (w4110 & w4111);
assign w1416 = ~w1414 & ~w1415;
assign w1417 = ~w1413 & w1416;
assign w1418 = (w389 & w4112) | (w389 & w4113) | (w4112 & w4113);
assign w1419 = (~w389 & w4114) | (~w389 & w4115) | (w4114 & w4115);
assign w1420 = ~w1418 & ~w1419;
assign w1421 = (w979 & w4116) | (w979 & w4117) | (w4116 & w4117);
assign w1422 = (~w979 & w4118) | (~w979 & w4119) | (w4118 & w4119);
assign w1423 = ~w1421 & ~w1422;
assign w1424 = w1420 & ~w1423;
assign w1425 = ~w1403 & ~w1410;
assign w1426 = ~w1417 & ~w1424;
assign w1427 = w1425 & w1426;
assign w1428 = w1372 & w1387;
assign w1429 = w1402 & w1428;
assign w1430 = w1427 & w1429;
assign w1431 = (w1214 & w3681) | (w1214 & w3682) | (w3681 & w3682);
assign w1432 = ~w1406 & w1409;
assign w1433 = ~w1382 & w1385;
assign w1434 = ~w1390 & w1393;
assign w1435 = w1367 & ~w1370;
assign w1436 = ~w1397 & w1400;
assign w1437 = ~w1360 & w1363;
assign w1438 = w1413 & ~w1416;
assign w1439 = ~w1420 & w1423;
assign w1440 = ~w1417 & w1439;
assign w1441 = ~w1437 & ~w1438;
assign w1442 = ~w1440 & w1441;
assign w1443 = w1372 & ~w1442;
assign w1444 = ~w1435 & ~w1436;
assign w1445 = (w1402 & w1443) | (w1402 & w3081) | (w1443 & w3081);
assign w1446 = ~w1433 & ~w1434;
assign w1447 = ~w1445 & w1446;
assign w1448 = w1375 & ~w1378;
assign w1449 = (~w1448 & w1447) | (~w1448 & w4120) | (w1447 & w4120);
assign w1450 = ~w1410 & ~w1449;
assign w1451 = pi302 & ~w1074;
assign w1452 = pi430 & w1074;
assign w1453 = ~w1451 & ~w1452;
assign w1454 = (pi047 & ~w532) | (pi047 & w3960) | (~w532 & w3960);
assign w1455 = w532 & w3961;
assign w1456 = ~w1454 & ~w1455;
assign w1457 = pi303 & ~w1074;
assign w1458 = pi431 & w1074;
assign w1459 = ~w1457 & ~w1458;
assign w1460 = w1456 & ~w1459;
assign w1461 = (pi046 & ~w532) | (pi046 & w3962) | (~w532 & w3962);
assign w1462 = w532 & w3963;
assign w1463 = ~w1461 & ~w1462;
assign w1464 = w1453 & ~w1463;
assign w1465 = ~w1460 & w1464;
assign w1466 = ~w1456 & w1459;
assign w1467 = (pi045 & ~w532) | (pi045 & w3964) | (~w532 & w3964);
assign w1468 = w532 & w3965;
assign w1469 = ~w1467 & ~w1468;
assign w1470 = pi301 & ~w1074;
assign w1471 = pi429 & w1074;
assign w1472 = ~w1470 & ~w1471;
assign w1473 = w1469 & ~w1472;
assign w1474 = ~w1453 & w1463;
assign w1475 = ~w1460 & ~w1473;
assign w1476 = ~w1474 & w1475;
assign w1477 = (~w516 & w4121) | (~w516 & w4122) | (w4121 & w4122);
assign w1478 = (w3966 & w516) | (w3966 & w4123) | (w516 & w4123);
assign w1479 = ~w1477 & ~w1478;
assign w1480 = pi300 & ~w1074;
assign w1481 = pi428 & w1074;
assign w1482 = ~w1480 & ~w1481;
assign w1483 = ~w1479 & w1482;
assign w1484 = ~w1469 & w1472;
assign w1485 = w1479 & ~w1482;
assign w1486 = (~w516 & w4124) | (~w516 & w4125) | (w4124 & w4125);
assign w1487 = (w3967 & w516) | (w3967 & w4126) | (w516 & w4126);
assign w1488 = ~w1486 & ~w1487;
assign w1489 = pi299 & ~w1074;
assign w1490 = pi427 & w1074;
assign w1491 = ~w1489 & ~w1490;
assign w1492 = w1488 & ~w1491;
assign w1493 = (~w516 & w4127) | (~w516 & w4128) | (w4127 & w4128);
assign w1494 = (w3968 & w516) | (w3968 & w4129) | (w516 & w4129);
assign w1495 = ~w1493 & ~w1494;
assign w1496 = pi298 & ~w1074;
assign w1497 = pi426 & w1074;
assign w1498 = ~w1496 & ~w1497;
assign w1499 = w1495 & ~w1498;
assign w1500 = ~w1485 & ~w1492;
assign w1501 = ~w1499 & w1500;
assign w1502 = (~w516 & w4130) | (~w516 & w4131) | (w4130 & w4131);
assign w1503 = (w3969 & w516) | (w3969 & w4132) | (w516 & w4132);
assign w1504 = ~w1502 & ~w1503;
assign w1505 = pi297 & ~w1074;
assign w1506 = pi425 & w1074;
assign w1507 = ~w1505 & ~w1506;
assign w1508 = w1504 & ~w1507;
assign w1509 = pi296 & ~w1074;
assign w1510 = pi424 & w1074;
assign w1511 = ~w1509 & ~w1510;
assign w1512 = (~w516 & w4133) | (~w516 & w4134) | (w4133 & w4134);
assign w1513 = (w3970 & w516) | (w3970 & w4135) | (w516 & w4135);
assign w1514 = ~w1512 & ~w1513;
assign w1515 = w1511 & ~w1514;
assign w1516 = ~w1508 & w1515;
assign w1517 = ~w1495 & w1498;
assign w1518 = ~w1504 & w1507;
assign w1519 = ~w1517 & ~w1518;
assign w1520 = ~w1516 & w1519;
assign w1521 = w1501 & ~w1520;
assign w1522 = ~w1488 & w1491;
assign w1523 = ~w1485 & w1522;
assign w1524 = ~w1483 & ~w1484;
assign w1525 = ~w1523 & w1524;
assign w1526 = ~w1521 & w1525;
assign w1527 = ~w1465 & ~w1466;
assign w1528 = (w1527 & w1526) | (w1527 & w3693) | (w1526 & w3693);
assign w1529 = ~w1432 & w1528;
assign w1530 = ~w1450 & w1529;
assign w1531 = ~w1511 & w1514;
assign w1532 = ~w1508 & ~w1531;
assign w1533 = w1476 & w1532;
assign w1534 = w1501 & w1533;
assign w1535 = w1528 & ~w1534;
assign w1536 = (pi057 & ~w532) | (pi057 & w3971) | (~w532 & w3971);
assign w1537 = w532 & w3972;
assign w1538 = ~w1536 & ~w1537;
assign w1539 = pi313 & ~w1074;
assign w1540 = pi441 & w1074;
assign w1541 = ~w1539 & ~w1540;
assign w1542 = w1538 & ~w1541;
assign w1543 = pi056 & ~w534;
assign w1544 = pi184 & w534;
assign w1545 = ~w1543 & ~w1544;
assign w1546 = ~w1542 & ~w1545;
assign w1547 = pi312 & ~w1074;
assign w1548 = pi440 & w1074;
assign w1549 = ~w1547 & ~w1548;
assign w1550 = ~w1542 & w1549;
assign w1551 = ~w1546 & ~w1550;
assign w1552 = (~w516 & w3694) | (~w516 & w3695) | (w3694 & w3695);
assign w1553 = (w3082 & w516) | (w3082 & w3696) | (w516 & w3696);
assign w1554 = ~w1552 & ~w1553;
assign w1555 = (w979 & w4136) | (w979 & w4137) | (w4136 & w4137);
assign w1556 = w3084 & w4205;
assign w1557 = ~w1555 & ~w1556;
assign w1558 = w1554 & ~w1557;
assign w1559 = (w979 & w4138) | (w979 & w4139) | (w4138 & w4139);
assign w1560 = w3086 & w4205;
assign w1561 = ~w1559 & ~w1560;
assign w1562 = (~w516 & w3697) | (~w516 & w3698) | (w3697 & w3698);
assign w1563 = (w3087 & w516) | (w3087 & w3699) | (w516 & w3699);
assign w1564 = ~w1562 & ~w1563;
assign w1565 = ~w1561 & w1564;
assign w1566 = ~w1558 & ~w1565;
assign w1567 = (pi059 & ~w532) | (pi059 & w3973) | (~w532 & w3973);
assign w1568 = w532 & w3974;
assign w1569 = ~w1567 & ~w1568;
assign w1570 = pi315 & ~w1074;
assign w1571 = pi443 & w1074;
assign w1572 = ~w1570 & ~w1571;
assign w1573 = w1569 & ~w1572;
assign w1574 = (pi058 & ~w532) | (pi058 & w3975) | (~w532 & w3975);
assign w1575 = w532 & w3976;
assign w1576 = ~w1574 & ~w1575;
assign w1577 = pi314 & ~w1074;
assign w1578 = pi442 & w1074;
assign w1579 = ~w1577 & ~w1578;
assign w1580 = w1576 & ~w1579;
assign w1581 = ~w1573 & ~w1580;
assign w1582 = (~w516 & w4140) | (~w516 & w4141) | (w4140 & w4141);
assign w1583 = (w3700 & w516) | (w3700 & w4142) | (w516 & w4142);
assign w1584 = ~w1582 & ~w1583;
assign w1585 = pi309 & ~w1074;
assign w1586 = pi437 & w1074;
assign w1587 = ~w1585 & ~w1586;
assign w1588 = w1584 & ~w1587;
assign w1589 = pi308 & ~w1074;
assign w1590 = pi436 & w1074;
assign w1591 = ~w1589 & ~w1590;
assign w1592 = (~w516 & w4143) | (~w516 & w4144) | (w4143 & w4144);
assign w1593 = (w3701 & w516) | (w3701 & w4145) | (w516 & w4145);
assign w1594 = ~w1592 & ~w1593;
assign w1595 = ~w1591 & w1594;
assign w1596 = (w3702 & w3703) | (w3702 & w4206) | (w3703 & w4206);
assign w1597 = (w3704 & w516) | (w3704 & w4146) | (w516 & w4146);
assign w1598 = ~w1596 & ~w1597;
assign w1599 = pi307 & ~w1074;
assign w1600 = pi435 & w1074;
assign w1601 = ~w1599 & ~w1600;
assign w1602 = w1598 & ~w1601;
assign w1603 = ~w1588 & ~w1595;
assign w1604 = ~w1602 & w1603;
assign w1605 = pi060 & ~w534;
assign w1606 = pi188 & w534;
assign w1607 = ~w1605 & ~w1606;
assign w1608 = pi316 & ~w1074;
assign w1609 = pi444 & w1074;
assign w1610 = ~w1608 & ~w1609;
assign w1611 = w1607 & ~w1610;
assign w1612 = pi063 & ~w534;
assign w1613 = pi191 & w534;
assign w1614 = ~w1612 & ~w1613;
assign w1615 = pi319 & ~w1074;
assign w1616 = pi447 & w1074;
assign w1617 = ~w1615 & ~w1616;
assign w1618 = w1614 & ~w1617;
assign w1619 = pi318 & ~w1074;
assign w1620 = pi446 & w1074;
assign w1621 = ~w1619 & ~w1620;
assign w1622 = pi062 & ~w534;
assign w1623 = pi190 & w534;
assign w1624 = ~w1622 & ~w1623;
assign w1625 = ~w1621 & w1624;
assign w1626 = pi061 & ~w534;
assign w1627 = pi189 & w534;
assign w1628 = ~w1626 & ~w1627;
assign w1629 = pi317 & ~w1074;
assign w1630 = pi445 & w1074;
assign w1631 = ~w1629 & ~w1630;
assign w1632 = w1628 & ~w1631;
assign w1633 = ~w1618 & ~w1625;
assign w1634 = ~w1632 & w1633;
assign w1635 = ~w1611 & w1634;
assign w1636 = pi310 & ~w1074;
assign w1637 = pi438 & w1074;
assign w1638 = ~w1636 & ~w1637;
assign w1639 = (~w516 & w4147) | (~w516 & w4148) | (w4147 & w4148);
assign w1640 = (w3705 & w516) | (w3705 & w4149) | (w516 & w4149);
assign w1641 = ~w1639 & ~w1640;
assign w1642 = ~w1638 & w1641;
assign w1643 = pi311 & ~w1074;
assign w1644 = pi439 & w1074;
assign w1645 = ~w1643 & ~w1644;
assign w1646 = (pi055 & ~w532) | (pi055 & w3706) | (~w532 & w3706);
assign w1647 = w532 & w3707;
assign w1648 = ~w1646 & ~w1647;
assign w1649 = ~w1645 & w1648;
assign w1650 = ~w1642 & ~w1649;
assign w1651 = (w979 & w4150) | (w979 & w4151) | (w4150 & w4151);
assign w1652 = w3097 & w4205;
assign w1653 = ~w1651 & ~w1652;
assign w1654 = (~w516 & w3708) | (~w516 & w3709) | (w3708 & w3709);
assign w1655 = (w3098 & w516) | (w3098 & w3710) | (w516 & w3710);
assign w1656 = ~w1654 & ~w1655;
assign w1657 = ~w1653 & w1656;
assign w1658 = w1566 & ~w1657;
assign w1659 = w1581 & w1650;
assign w1660 = w1658 & w1659;
assign w1661 = ~w1551 & w1604;
assign w1662 = w1660 & w1661;
assign w1663 = w1635 & w1662;
assign w1664 = ~w1535 & w1663;
assign w1665 = (w1664 & w1431) | (w1664 & w3835) | (w1431 & w3835);
assign w1666 = ~w1614 & w1617;
assign w1667 = ~w1569 & w1572;
assign w1668 = w1546 & w1549;
assign w1669 = ~w1576 & w1579;
assign w1670 = ~w1538 & w1541;
assign w1671 = w1645 & ~w1648;
assign w1672 = ~w1584 & w1587;
assign w1673 = w1638 & ~w1641;
assign w1674 = ~w1598 & w1601;
assign w1675 = ~w1554 & w1557;
assign w1676 = w1653 & ~w1656;
assign w1677 = ~w1675 & ~w1676;
assign w1678 = w1566 & ~w1677;
assign w1679 = w1561 & ~w1564;
assign w1680 = ~w1674 & ~w1679;
assign w1681 = ~w1678 & w1680;
assign w1682 = w1604 & ~w1681;
assign w1683 = w1591 & ~w1594;
assign w1684 = ~w1588 & w1683;
assign w1685 = ~w1672 & ~w1673;
assign w1686 = ~w1684 & w1685;
assign w1687 = (~w1682 & w4152) | (~w1682 & w4153) | (w4152 & w4153);
assign w1688 = ~w1551 & ~w1687;
assign w1689 = ~w1669 & ~w1670;
assign w1690 = ~w1668 & w1689;
assign w1691 = (w1581 & w1688) | (w1581 & w3836) | (w1688 & w3836);
assign w1692 = ~w1667 & ~w1691;
assign w1693 = (pi067 & ~w532) | (pi067 & w3837) | (~w532 & w3837);
assign w1694 = w532 & w3838;
assign w1695 = ~w1693 & ~w1694;
assign w1696 = pi323 & ~w1074;
assign w1697 = pi451 & w1074;
assign w1698 = ~w1696 & ~w1697;
assign w1699 = ~w1695 & w1698;
assign w1700 = w1695 & ~w1698;
assign w1701 = pi322 & ~w1074;
assign w1702 = pi450 & w1074;
assign w1703 = ~w1701 & ~w1702;
assign w1704 = (~w516 & w4154) | (~w516 & w4155) | (w4154 & w4155);
assign w1705 = (w3839 & w516) | (w3839 & w4156) | (w516 & w4156);
assign w1706 = ~w1704 & ~w1705;
assign w1707 = ~w1703 & w1706;
assign w1708 = ~w1700 & ~w1707;
assign w1709 = (~w516 & w4157) | (~w516 & w4158) | (w4157 & w4158);
assign w1710 = (w3840 & w516) | (w3840 & w4159) | (w516 & w4159);
assign w1711 = ~w1709 & ~w1710;
assign w1712 = pi321 & ~w1074;
assign w1713 = pi449 & w1074;
assign w1714 = ~w1712 & ~w1713;
assign w1715 = ~w1711 & w1714;
assign w1716 = w1703 & ~w1706;
assign w1717 = pi320 & ~w1074;
assign w1718 = pi448 & w1074;
assign w1719 = ~w1717 & ~w1718;
assign w1720 = w1711 & ~w1714;
assign w1721 = (~w516 & w4160) | (~w516 & w4161) | (w4160 & w4161);
assign w1722 = (w3841 & w516) | (w3841 & w4162) | (w516 & w4162);
assign w1723 = ~w1721 & ~w1722;
assign w1724 = w1719 & ~w1723;
assign w1725 = ~w1720 & w1724;
assign w1726 = ~w1715 & ~w1716;
assign w1727 = ~w1725 & w1726;
assign w1728 = w1708 & ~w1727;
assign w1729 = ~w1699 & ~w1728;
assign w1730 = ~w1628 & w1631;
assign w1731 = ~w1607 & w1610;
assign w1732 = ~w1730 & ~w1731;
assign w1733 = w1634 & ~w1732;
assign w1734 = w1621 & ~w1624;
assign w1735 = ~w1618 & w1734;
assign w1736 = ~w1666 & ~w1735;
assign w1737 = ~w1733 & w3842;
assign w1738 = pi075 & ~w534;
assign w1739 = w532 & w3843;
assign w1740 = ~w1738 & ~w1739;
assign w1741 = pi331 & ~w1074;
assign w1742 = pi459 & w1074;
assign w1743 = ~w1741 & ~w1742;
assign w1744 = ~w1738 & w3844;
assign w1745 = pi330 & ~w1074;
assign w1746 = pi458 & w1074;
assign w1747 = ~w1745 & ~w1746;
assign w1748 = (pi074 & ~w532) | (pi074 & w3845) | (~w532 & w3845);
assign w1749 = w532 & w3846;
assign w1750 = ~w1748 & ~w1749;
assign w1751 = ~w1747 & w1750;
assign w1752 = ~w1744 & ~w1751;
assign w1753 = ~w1719 & w1723;
assign w1754 = ~w1720 & ~w1753;
assign w1755 = w1708 & w1754;
assign w1756 = w1729 & ~w1755;
assign w1757 = pi326 & ~w1074;
assign w1758 = pi454 & w1074;
assign w1759 = ~w1757 & ~w1758;
assign w1760 = (~w516 & w3847) | (~w516 & w3848) | (w3847 & w3848);
assign w1761 = (w3717 & w516) | (w3717 & w3849) | (w516 & w3849);
assign w1762 = ~w1760 & ~w1761;
assign w1763 = ~w1759 & w1762;
assign w1764 = (~w516 & w3850) | (~w516 & w3851) | (w3850 & w3851);
assign w1765 = (w3718 & w516) | (w3718 & w3852) | (w516 & w3852);
assign w1766 = ~w1764 & ~w1765;
assign w1767 = pi325 & ~w1074;
assign w1768 = pi453 & w1074;
assign w1769 = ~w1767 & ~w1768;
assign w1770 = w1766 & ~w1769;
assign w1771 = ~w1763 & ~w1770;
assign w1772 = (~w516 & w3853) | (~w516 & w3854) | (w3853 & w3854);
assign w1773 = (w3719 & w516) | (w3719 & w3855) | (w516 & w3855);
assign w1774 = ~w1772 & ~w1773;
assign w1775 = pi324 & ~w1074;
assign w1776 = pi452 & w1074;
assign w1777 = ~w1775 & ~w1776;
assign w1778 = w1774 & ~w1777;
assign w1779 = (w3856 & w3857) | (w3856 & w4206) | (w3857 & w4206);
assign w1780 = (w3858 & w516) | (w3858 & w4163) | (w516 & w4163);
assign w1781 = ~w1779 & ~w1780;
assign w1782 = pi329 & ~w1074;
assign w1783 = pi457 & w1074;
assign w1784 = ~w1782 & ~w1783;
assign w1785 = w1781 & ~w1784;
assign w1786 = pi328 & ~w1074;
assign w1787 = pi456 & w1074;
assign w1788 = ~w1786 & ~w1787;
assign w1789 = (w3859 & w3860) | (w3859 & w4206) | (w3860 & w4206);
assign w1790 = (w3861 & w516) | (w3861 & w4164) | (w516 & w4164);
assign w1791 = ~w1789 & ~w1790;
assign w1792 = ~w1788 & w1791;
assign w1793 = (w3862 & w3863) | (w3862 & w4206) | (w3863 & w4206);
assign w1794 = (w3864 & w516) | (w3864 & w4165) | (w516 & w4165);
assign w1795 = ~w1793 & ~w1794;
assign w1796 = pi327 & ~w1074;
assign w1797 = pi455 & w1074;
assign w1798 = ~w1796 & ~w1797;
assign w1799 = w1795 & ~w1798;
assign w1800 = ~w1785 & ~w1792;
assign w1801 = ~w1799 & w1800;
assign w1802 = w1752 & ~w1778;
assign w1803 = w1771 & w1802;
assign w1804 = w1801 & w1803;
assign w1805 = ~w1756 & w1804;
assign w1806 = (w1805 & w1665) | (w1805 & w2781) | (w1665 & w2781);
assign w1807 = ~w1740 & w1743;
assign w1808 = w1759 & ~w1762;
assign w1809 = ~w1795 & w1798;
assign w1810 = ~w1766 & w1769;
assign w1811 = ~w1774 & w1777;
assign w1812 = ~w1810 & ~w1811;
assign w1813 = w1771 & ~w1812;
assign w1814 = ~w1808 & ~w1809;
assign w1815 = ~w1813 & w1814;
assign w1816 = w1801 & ~w1815;
assign w1817 = w1747 & ~w1750;
assign w1818 = ~w1781 & w1784;
assign w1819 = w1788 & ~w1791;
assign w1820 = ~w1785 & w1819;
assign w1821 = ~w1817 & ~w1818;
assign w1822 = ~w1820 & w1821;
assign w1823 = (w1752 & w1816) | (w1752 & w4166) | (w1816 & w4166);
assign w1824 = (~w516 & w3865) | (~w516 & w3866) | (w3865 & w3866);
assign w1825 = (w3726 & w516) | (w3726 & w3867) | (w516 & w3867);
assign w1826 = ~w1824 & ~w1825;
assign w1827 = pi335 & ~w1074;
assign w1828 = pi463 & w1074;
assign w1829 = ~w1827 & ~w1828;
assign w1830 = ~w1826 & w1829;
assign w1831 = (w3868 & w3869) | (w3868 & w4206) | (w3869 & w4206);
assign w1832 = (w3870 & w516) | (w3870 & w4167) | (w516 & w4167);
assign w1833 = ~w1831 & ~w1832;
assign w1834 = pi333 & ~w1074;
assign w1835 = pi461 & w1074;
assign w1836 = ~w1834 & ~w1835;
assign w1837 = ~w1833 & w1836;
assign w1838 = pi332 & ~w1074;
assign w1839 = pi460 & w1074;
assign w1840 = ~w1838 & ~w1839;
assign w1841 = (w3871 & w3872) | (w3871 & w4206) | (w3872 & w4206);
assign w1842 = (w3873 & w516) | (w3873 & w4168) | (w516 & w4168);
assign w1843 = ~w1841 & ~w1842;
assign w1844 = w1840 & ~w1843;
assign w1845 = ~w1837 & ~w1844;
assign w1846 = w1826 & ~w1829;
assign w1847 = (~w516 & w3874) | (~w516 & w3875) | (w3874 & w3875);
assign w1848 = (w3731 & w516) | (w3731 & w3876) | (w516 & w3876);
assign w1849 = ~w1847 & ~w1848;
assign w1850 = pi334 & ~w1074;
assign w1851 = pi462 & w1074;
assign w1852 = ~w1850 & ~w1851;
assign w1853 = w1849 & ~w1852;
assign w1854 = w1833 & ~w1836;
assign w1855 = ~w1846 & ~w1853;
assign w1856 = ~w1854 & w1855;
assign w1857 = ~w1845 & w1856;
assign w1858 = ~w1849 & w1852;
assign w1859 = ~w1846 & w1858;
assign w1860 = ~w1830 & ~w1859;
assign w1861 = ~w1857 & w1860;
assign w1862 = ~w1807 & w1861;
assign w1863 = ~w1823 & w1862;
assign w1864 = pi336 & ~w1074;
assign w1865 = pi464 & w1074;
assign w1866 = ~w1864 & ~w1865;
assign w1867 = (w3732 & w3733) | (w3732 & w4206) | (w3733 & w4206);
assign w1868 = (w3734 & w516) | (w3734 & w3877) | (w516 & w3877);
assign w1869 = ~w1867 & ~w1868;
assign w1870 = ~w1866 & w1869;
assign w1871 = ~w1840 & w1843;
assign w1872 = w1856 & ~w1871;
assign w1873 = w1861 & ~w1872;
assign w1874 = (w3878 & w3879) | (w3878 & w4206) | (w3879 & w4206);
assign w1875 = (w3880 & w516) | (w3880 & w4169) | (w516 & w4169);
assign w1876 = ~w1874 & ~w1875;
assign w1877 = pi341 & ~w1074;
assign w1878 = pi469 & w1074;
assign w1879 = ~w1877 & ~w1878;
assign w1880 = w1876 & ~w1879;
assign w1881 = (w3881 & w3882) | (w3881 & w4206) | (w3882 & w4206);
assign w1882 = (w3883 & w516) | (w3883 & w4170) | (w516 & w4170);
assign w1883 = ~w1881 & ~w1882;
assign w1884 = pi343 & ~w1074;
assign w1885 = pi471 & w1074;
assign w1886 = ~w1884 & ~w1885;
assign w1887 = w1883 & ~w1886;
assign w1888 = pi342 & ~w1074;
assign w1889 = pi470 & w1074;
assign w1890 = ~w1888 & ~w1889;
assign w1891 = (pi086 & ~w532) | (pi086 & w3884) | (~w532 & w3884);
assign w1892 = w532 & w3885;
assign w1893 = ~w1891 & ~w1892;
assign w1894 = ~w1890 & w1893;
assign w1895 = ~w1880 & ~w1887;
assign w1896 = ~w1894 & w1895;
assign w1897 = pi338 & ~w1074;
assign w1898 = pi466 & w1074;
assign w1899 = ~w1897 & ~w1898;
assign w1900 = (w3739 & w3740) | (w3739 & w4206) | (w3740 & w4206);
assign w1901 = (w3741 & w516) | (w3741 & w3886) | (w516 & w3886);
assign w1902 = ~w1900 & ~w1901;
assign w1903 = ~w1899 & w1902;
assign w1904 = (w3742 & w3743) | (w3742 & w4206) | (w3743 & w4206);
assign w1905 = (w3744 & w516) | (w3744 & w3887) | (w516 & w3887);
assign w1906 = ~w1904 & ~w1905;
assign w1907 = pi340 & ~w1074;
assign w1908 = pi468 & w1074;
assign w1909 = ~w1907 & ~w1908;
assign w1910 = w1906 & ~w1909;
assign w1911 = (w3888 & w3889) | (w3888 & w4206) | (w3889 & w4206);
assign w1912 = (w3890 & w516) | (w3890 & w4171) | (w516 & w4171);
assign w1913 = ~w1911 & ~w1912;
assign w1914 = pi339 & ~w1074;
assign w1915 = pi467 & w1074;
assign w1916 = ~w1914 & ~w1915;
assign w1917 = w1913 & ~w1916;
assign w1918 = ~w1903 & ~w1910;
assign w1919 = ~w1917 & w1918;
assign w1920 = (w3747 & w3748) | (w3747 & w4206) | (w3748 & w4206);
assign w1921 = (w3749 & w516) | (w3749 & w3891) | (w516 & w3891);
assign w1922 = ~w1920 & ~w1921;
assign w1923 = pi337 & ~w1074;
assign w1924 = pi465 & w1074;
assign w1925 = ~w1923 & ~w1924;
assign w1926 = w1922 & ~w1925;
assign w1927 = ~w1870 & ~w1926;
assign w1928 = w1896 & w1927;
assign w1929 = w1919 & w1928;
assign w1930 = ~w1873 & w1929;
assign w1931 = w1890 & ~w1893;
assign w1932 = ~w1887 & w1931;
assign w1933 = (w3892 & w3893) | (w3892 & w4206) | (w3893 & w4206);
assign w1934 = (w3894 & w516) | (w3894 & w4172) | (w516 & w4172);
assign w1935 = ~w1933 & ~w1934;
assign w1936 = pi347 & ~w1074;
assign w1937 = pi475 & w1074;
assign w1938 = ~w1936 & ~w1937;
assign w1939 = ~w1935 & w1938;
assign w1940 = w1935 & ~w1938;
assign w1941 = pi346 & ~w1074;
assign w1942 = pi474 & w1074;
assign w1943 = ~w1941 & ~w1942;
assign w1944 = (w3752 & w3753) | (w3752 & w4206) | (w3753 & w4206);
assign w1945 = (w3754 & w516) | (w3754 & w3895) | (w516 & w3895);
assign w1946 = ~w1944 & ~w1945;
assign w1947 = ~w1943 & w1946;
assign w1948 = ~w1940 & ~w1947;
assign w1949 = (w3755 & w3756) | (w3755 & w4206) | (w3756 & w4206);
assign w1950 = (w3757 & w516) | (w3757 & w3896) | (w516 & w3896);
assign w1951 = ~w1949 & ~w1950;
assign w1952 = pi345 & ~w1074;
assign w1953 = pi473 & w1074;
assign w1954 = ~w1952 & ~w1953;
assign w1955 = ~w1951 & w1954;
assign w1956 = w1943 & ~w1946;
assign w1957 = pi344 & ~w1074;
assign w1958 = pi472 & w1074;
assign w1959 = ~w1957 & ~w1958;
assign w1960 = w1951 & ~w1954;
assign w1961 = (w3758 & w3759) | (w3758 & w4206) | (w3759 & w4206);
assign w1962 = (w3760 & w516) | (w3760 & w3897) | (w516 & w3897);
assign w1963 = ~w1961 & ~w1962;
assign w1964 = w1959 & ~w1963;
assign w1965 = ~w1960 & w1964;
assign w1966 = ~w1955 & ~w1956;
assign w1967 = ~w1965 & w1966;
assign w1968 = (~w1939 & w1967) | (~w1939 & w4173) | (w1967 & w4173);
assign w1969 = ~w1883 & w1886;
assign w1970 = ~w1906 & w1909;
assign w1971 = ~w1876 & w1879;
assign w1972 = ~w1922 & w1925;
assign w1973 = w1899 & ~w1902;
assign w1974 = w1866 & ~w1869;
assign w1975 = ~w1926 & w1974;
assign w1976 = ~w1972 & ~w1973;
assign w1977 = ~w1975 & w1976;
assign w1978 = w1919 & ~w1977;
assign w1979 = ~w1913 & w1916;
assign w1980 = ~w1910 & w1979;
assign w1981 = ~w1970 & ~w1971;
assign w1982 = ~w1980 & w1981;
assign w1983 = (w1896 & w1978) | (w1896 & w4174) | (w1978 & w4174);
assign w1984 = ~w1932 & ~w1969;
assign w1985 = w1968 & w1984;
assign w1986 = ~w1983 & w1985;
assign w1987 = (pi099 & ~w532) | (pi099 & w3898) | (~w532 & w3898);
assign w1988 = w532 & w3899;
assign w1989 = ~w1987 & ~w1988;
assign w1990 = pi355 & ~w1074;
assign w1991 = pi483 & w1074;
assign w1992 = ~w1990 & ~w1991;
assign w1993 = w1989 & ~w1992;
assign w1994 = pi354 & ~w1074;
assign w1995 = pi482 & w1074;
assign w1996 = ~w1994 & ~w1995;
assign w1997 = (pi098 & ~w532) | (pi098 & w3900) | (~w532 & w3900);
assign w1998 = w532 & w3901;
assign w1999 = ~w1997 & ~w1998;
assign w2000 = ~w1996 & w1999;
assign w2001 = ~w1993 & ~w2000;
assign w2002 = ~w1959 & w1963;
assign w2003 = ~w1960 & ~w2002;
assign w2004 = w1948 & w2003;
assign w2005 = w1968 & ~w2004;
assign w2006 = (~w516 & w4175) | (~w516 & w4176) | (w4175 & w4176);
assign w2007 = (w3902 & w516) | (w3902 & w4177) | (w516 & w4177);
assign w2008 = ~w2006 & ~w2007;
assign w2009 = pi349 & ~w1074;
assign w2010 = pi477 & w1074;
assign w2011 = ~w2009 & ~w2010;
assign w2012 = w2008 & ~w2011;
assign w2013 = pi350 & ~w1074;
assign w2014 = pi478 & w1074;
assign w2015 = ~w2013 & ~w2014;
assign w2016 = (~w516 & w4178) | (~w516 & w4179) | (w4178 & w4179);
assign w2017 = (w3903 & w516) | (w3903 & w4180) | (w516 & w4180);
assign w2018 = ~w2016 & ~w2017;
assign w2019 = ~w2015 & w2018;
assign w2020 = ~w2012 & ~w2019;
assign w2021 = (~w516 & w4181) | (~w516 & w4182) | (w4181 & w4182);
assign w2022 = (w3904 & w516) | (w3904 & w4183) | (w516 & w4183);
assign w2023 = ~w2021 & ~w2022;
assign w2024 = pi348 & ~w1074;
assign w2025 = pi476 & w1074;
assign w2026 = ~w2024 & ~w2025;
assign w2027 = w2023 & ~w2026;
assign w2028 = (pi095 & ~w532) | (pi095 & w3905) | (~w532 & w3905);
assign w2029 = w532 & w3906;
assign w2030 = ~w2028 & ~w2029;
assign w2031 = pi351 & ~w1074;
assign w2032 = pi479 & w1074;
assign w2033 = ~w2031 & ~w2032;
assign w2034 = w2030 & ~w2033;
assign w2035 = (pi097 & ~w532) | (pi097 & w3907) | (~w532 & w3907);
assign w2036 = w532 & w3908;
assign w2037 = ~w2035 & ~w2036;
assign w2038 = pi353 & ~w1074;
assign w2039 = pi481 & w1074;
assign w2040 = ~w2038 & ~w2039;
assign w2041 = w2037 & ~w2040;
assign w2042 = pi352 & ~w1074;
assign w2043 = pi480 & w1074;
assign w2044 = ~w2042 & ~w2043;
assign w2045 = pi096 & ~w534;
assign w2046 = pi224 & w534;
assign w2047 = ~w2045 & ~w2046;
assign w2048 = ~w2044 & w2047;
assign w2049 = ~w2034 & ~w2041;
assign w2050 = ~w2048 & w2049;
assign w2051 = w2001 & ~w2027;
assign w2052 = w2020 & w2051;
assign w2053 = w2050 & w2052;
assign w2054 = ~w2005 & w2053;
assign w2055 = ~w1989 & w1992;
assign w2056 = w2015 & ~w2018;
assign w2057 = ~w2030 & w2033;
assign w2058 = ~w2008 & w2011;
assign w2059 = ~w2023 & w2026;
assign w2060 = ~w2058 & ~w2059;
assign w2061 = w2020 & ~w2060;
assign w2062 = ~w2056 & ~w2057;
assign w2063 = ~w2061 & w2062;
assign w2064 = w2050 & ~w2063;
assign w2065 = w1996 & ~w1999;
assign w2066 = ~w2037 & w2040;
assign w2067 = w2044 & ~w2047;
assign w2068 = ~w2041 & w2067;
assign w2069 = ~w2065 & ~w2066;
assign w2070 = ~w2068 & w2069;
assign w2071 = ~w2064 & w2070;
assign w2072 = w2001 & ~w2071;
assign w2073 = (pi103 & ~w532) | (pi103 & w3909) | (~w532 & w3909);
assign w2074 = w532 & w3910;
assign w2075 = ~w2073 & ~w2074;
assign w2076 = pi359 & ~w1074;
assign w2077 = pi487 & w1074;
assign w2078 = ~w2076 & ~w2077;
assign w2079 = ~w2075 & w2078;
assign w2080 = pi101 & ~w534;
assign w2081 = pi229 & w534;
assign w2082 = ~w2080 & ~w2081;
assign w2083 = pi357 & ~w1074;
assign w2084 = pi485 & w1074;
assign w2085 = ~w2083 & ~w2084;
assign w2086 = ~w2082 & w2085;
assign w2087 = pi356 & ~w1074;
assign w2088 = pi484 & w1074;
assign w2089 = ~w2087 & ~w2088;
assign w2090 = pi100 & ~w534;
assign w2091 = pi228 & w534;
assign w2092 = ~w2090 & ~w2091;
assign w2093 = w2089 & ~w2092;
assign w2094 = ~w2086 & ~w2093;
assign w2095 = w2075 & ~w2078;
assign w2096 = (pi102 & ~w532) | (pi102 & w3911) | (~w532 & w3911);
assign w2097 = w532 & w3912;
assign w2098 = ~w2096 & ~w2097;
assign w2099 = pi358 & ~w1074;
assign w2100 = pi486 & w1074;
assign w2101 = ~w2099 & ~w2100;
assign w2102 = w2098 & ~w2101;
assign w2103 = w2082 & ~w2085;
assign w2104 = ~w2095 & ~w2102;
assign w2105 = ~w2103 & w2104;
assign w2106 = ~w2094 & w2105;
assign w2107 = ~w2098 & w2101;
assign w2108 = ~w2095 & w2107;
assign w2109 = ~w2079 & ~w2108;
assign w2110 = ~w2106 & w2109;
assign w2111 = ~w2055 & w2110;
assign w2112 = ~w2072 & w2111;
assign w2113 = pi360 & ~w1074;
assign w2114 = pi488 & w1074;
assign w2115 = ~w2113 & ~w2114;
assign w2116 = pi104 & ~w534;
assign w2117 = pi232 & w534;
assign w2118 = ~w2116 & ~w2117;
assign w2119 = ~w2115 & w2118;
assign w2120 = ~w2089 & w2092;
assign w2121 = w2105 & ~w2120;
assign w2122 = w2110 & ~w2121;
assign w2123 = pi109 & ~w534;
assign w2124 = pi237 & w534;
assign w2125 = ~w2123 & ~w2124;
assign w2126 = pi365 & ~w1074;
assign w2127 = pi493 & w1074;
assign w2128 = ~w2126 & ~w2127;
assign w2129 = w2125 & ~w2128;
assign w2130 = pi111 & ~w534;
assign w2131 = pi239 & w534;
assign w2132 = ~w2130 & ~w2131;
assign w2133 = pi367 & ~w1074;
assign w2134 = pi495 & w1074;
assign w2135 = ~w2133 & ~w2134;
assign w2136 = w2132 & ~w2135;
assign w2137 = pi366 & ~w1074;
assign w2138 = pi494 & w1074;
assign w2139 = ~w2137 & ~w2138;
assign w2140 = pi110 & ~w534;
assign w2141 = pi238 & w534;
assign w2142 = ~w2140 & ~w2141;
assign w2143 = ~w2139 & w2142;
assign w2144 = ~w2129 & ~w2136;
assign w2145 = ~w2143 & w2144;
assign w2146 = pi362 & ~w1074;
assign w2147 = pi490 & w1074;
assign w2148 = ~w2146 & ~w2147;
assign w2149 = pi106 & ~w534;
assign w2150 = pi234 & w534;
assign w2151 = ~w2149 & ~w2150;
assign w2152 = ~w2148 & w2151;
assign w2153 = pi108 & ~w534;
assign w2154 = pi236 & w534;
assign w2155 = ~w2153 & ~w2154;
assign w2156 = pi364 & ~w1074;
assign w2157 = pi492 & w1074;
assign w2158 = ~w2156 & ~w2157;
assign w2159 = w2155 & ~w2158;
assign w2160 = pi107 & ~w534;
assign w2161 = pi235 & w534;
assign w2162 = ~w2160 & ~w2161;
assign w2163 = pi363 & ~w1074;
assign w2164 = pi491 & w1074;
assign w2165 = ~w2163 & ~w2164;
assign w2166 = w2162 & ~w2165;
assign w2167 = ~w2152 & ~w2159;
assign w2168 = ~w2166 & w2167;
assign w2169 = pi105 & ~w534;
assign w2170 = pi233 & w534;
assign w2171 = ~w2169 & ~w2170;
assign w2172 = pi361 & ~w1074;
assign w2173 = pi489 & w1074;
assign w2174 = ~w2172 & ~w2173;
assign w2175 = w2171 & ~w2174;
assign w2176 = ~w2119 & ~w2175;
assign w2177 = w2145 & w2176;
assign w2178 = w2168 & w2177;
assign w2179 = ~w2122 & w2178;
assign w2180 = w2139 & ~w2142;
assign w2181 = ~w2136 & w2180;
assign w2182 = (pi115 & ~w532) | (pi115 & w3913) | (~w532 & w3913);
assign w2183 = w532 & w3914;
assign w2184 = ~w2182 & ~w2183;
assign w2185 = pi371 & ~w1074;
assign w2186 = pi499 & w1074;
assign w2187 = ~w2185 & ~w2186;
assign w2188 = ~w2184 & w2187;
assign w2189 = w2184 & ~w2187;
assign w2190 = pi370 & ~w1074;
assign w2191 = pi498 & w1074;
assign w2192 = ~w2190 & ~w2191;
assign w2193 = (~w516 & w4184) | (~w516 & w4185) | (w4184 & w4185);
assign w2194 = (w3915 & w516) | (w3915 & w4186) | (w516 & w4186);
assign w2195 = ~w2193 & ~w2194;
assign w2196 = ~w2192 & w2195;
assign w2197 = ~w2189 & ~w2196;
assign w2198 = (~w516 & w4187) | (~w516 & w4188) | (w4187 & w4188);
assign w2199 = (w3916 & w516) | (w3916 & w4189) | (w516 & w4189);
assign w2200 = ~w2198 & ~w2199;
assign w2201 = pi369 & ~w1074;
assign w2202 = pi497 & w1074;
assign w2203 = ~w2201 & ~w2202;
assign w2204 = ~w2200 & w2203;
assign w2205 = w2192 & ~w2195;
assign w2206 = pi368 & ~w1074;
assign w2207 = pi496 & w1074;
assign w2208 = ~w2206 & ~w2207;
assign w2209 = w2200 & ~w2203;
assign w2210 = (~w516 & w4190) | (~w516 & w4191) | (w4190 & w4191);
assign w2211 = (w3917 & w516) | (w3917 & w4192) | (w516 & w4192);
assign w2212 = ~w2210 & ~w2211;
assign w2213 = w2208 & ~w2212;
assign w2214 = ~w2209 & w2213;
assign w2215 = ~w2204 & ~w2205;
assign w2216 = ~w2214 & w2215;
assign w2217 = w2197 & ~w2216;
assign w2218 = ~w2188 & ~w2217;
assign w2219 = ~w2132 & w2135;
assign w2220 = ~w2155 & w2158;
assign w2221 = ~w2125 & w2128;
assign w2222 = ~w2171 & w2174;
assign w2223 = w2148 & ~w2151;
assign w2224 = w2115 & ~w2118;
assign w2225 = ~w2175 & w2224;
assign w2226 = ~w2222 & ~w2223;
assign w2227 = ~w2225 & w2226;
assign w2228 = w2168 & ~w2227;
assign w2229 = ~w2162 & w2165;
assign w2230 = ~w2159 & w2229;
assign w2231 = ~w2220 & ~w2221;
assign w2232 = ~w2230 & w2231;
assign w2233 = ~w2228 & w2232;
assign w2234 = w2145 & ~w2233;
assign w2235 = ~w2181 & ~w2219;
assign w2236 = w2218 & w2235;
assign w2237 = ~w2234 & w2236;
assign w2238 = (~w1806 & w2787) | (~w1806 & w2788) | (w2787 & w2788);
assign w2239 = pi123 & ~w534;
assign w2240 = pi251 & w534;
assign w2241 = ~w2239 & ~w2240;
assign w2242 = pi379 & ~w1074;
assign w2243 = pi507 & w1074;
assign w2244 = ~w2242 & ~w2243;
assign w2245 = w2241 & ~w2244;
assign w2246 = pi378 & ~w1074;
assign w2247 = pi506 & w1074;
assign w2248 = ~w2246 & ~w2247;
assign w2249 = pi122 & ~w534;
assign w2250 = pi250 & w534;
assign w2251 = ~w2249 & ~w2250;
assign w2252 = ~w2248 & w2251;
assign w2253 = ~w2245 & ~w2252;
assign w2254 = ~w2208 & w2212;
assign w2255 = ~w2209 & ~w2254;
assign w2256 = w2197 & w2255;
assign w2257 = w2218 & ~w2256;
assign w2258 = pi121 & ~w534;
assign w2259 = pi249 & w534;
assign w2260 = ~w2258 & ~w2259;
assign w2261 = pi377 & ~w1074;
assign w2262 = pi505 & w1074;
assign w2263 = ~w2261 & ~w2262;
assign w2264 = w2260 & ~w2263;
assign w2265 = pi372 & ~w1074;
assign w2266 = pi500 & w1074;
assign w2267 = ~w2265 & ~w2266;
assign w2268 = (~w516 & w3918) | (~w516 & w3919) | (w3918 & w3919);
assign w2269 = (w3773 & w516) | (w3773 & w3920) | (w516 & w3920);
assign w2270 = ~w2268 & ~w2269;
assign w2271 = ~w2267 & w2270;
assign w2272 = (w3921 & w3922) | (w3921 & w4206) | (w3922 & w4206);
assign w2273 = (w3923 & w516) | (w3923 & w4193) | (w516 & w4193);
assign w2274 = ~w2272 & ~w2273;
assign w2275 = pi375 & ~w1074;
assign w2276 = pi503 & w1074;
assign w2277 = ~w2275 & ~w2276;
assign w2278 = w2274 & ~w2277;
assign w2279 = pi376 & ~w1074;
assign w2280 = pi504 & w1074;
assign w2281 = ~w2279 & ~w2280;
assign w2282 = (pi120 & ~w532) | (pi120 & w3924) | (~w532 & w3924);
assign w2283 = w532 & w3925;
assign w2284 = ~w2282 & ~w2283;
assign w2285 = ~w2281 & w2284;
assign w2286 = ~w2278 & ~w2285;
assign w2287 = pi374 & ~w1074;
assign w2288 = pi502 & w1074;
assign w2289 = ~w2287 & ~w2288;
assign w2290 = (~w516 & w3926) | (~w516 & w3927) | (w3926 & w3927);
assign w2291 = (w3776 & w516) | (w3776 & w3928) | (w516 & w3928);
assign w2292 = ~w2290 & ~w2291;
assign w2293 = ~w2289 & w2292;
assign w2294 = (~w516 & w3929) | (~w516 & w3930) | (w3929 & w3930);
assign w2295 = (w3777 & w516) | (w3777 & w3931) | (w516 & w3931);
assign w2296 = ~w2294 & ~w2295;
assign w2297 = pi373 & ~w1074;
assign w2298 = pi501 & w1074;
assign w2299 = ~w2297 & ~w2298;
assign w2300 = w2296 & ~w2299;
assign w2301 = ~w2293 & ~w2300;
assign w2302 = ~w2264 & ~w2271;
assign w2303 = w2253 & w2302;
assign w2304 = w2286 & w2301;
assign w2305 = w2303 & w2304;
assign w2306 = ~w2257 & w2305;
assign w2307 = ~w2241 & w2244;
assign w2308 = ~w2260 & w2263;
assign w2309 = w2248 & ~w2251;
assign w2310 = w2281 & ~w2284;
assign w2311 = ~w2274 & w2277;
assign w2312 = w2289 & ~w2292;
assign w2313 = ~w2296 & w2299;
assign w2314 = w2267 & ~w2270;
assign w2315 = ~w2313 & ~w2314;
assign w2316 = w2301 & ~w2315;
assign w2317 = ~w2311 & ~w2312;
assign w2318 = ~w2316 & w2317;
assign w2319 = (~w2310 & w2318) | (~w2310 & w4194) | (w2318 & w4194);
assign w2320 = ~w2264 & ~w2319;
assign w2321 = ~w2308 & ~w2309;
assign w2322 = ~w2320 & w2321;
assign w2323 = w2253 & ~w2322;
assign w2324 = ~w2307 & ~w2323;
assign w2325 = pi126 & ~w534;
assign w2326 = pi254 & w534;
assign w2327 = ~w2325 & ~w2326;
assign w2328 = pi382 & ~w1074;
assign w2329 = pi510 & w1074;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = w2327 & ~w2330;
assign w2332 = pi125 & ~w534;
assign w2333 = pi253 & w534;
assign w2334 = ~w2332 & ~w2333;
assign w2335 = pi381 & ~w1074;
assign w2336 = pi509 & w1074;
assign w2337 = ~w2335 & ~w2336;
assign w2338 = w2334 & ~w2337;
assign w2339 = ~w2331 & ~w2338;
assign w2340 = pi124 & ~w534;
assign w2341 = pi252 & w534;
assign w2342 = ~w2340 & ~w2341;
assign w2343 = pi380 & ~w1074;
assign w2344 = pi508 & w1074;
assign w2345 = ~w2343 & ~w2344;
assign w2346 = w2342 & ~w2345;
assign w2347 = w2339 & ~w2346;
assign w2348 = ~w2327 & w2330;
assign w2349 = ~w2334 & w2337;
assign w2350 = ~w2342 & w2345;
assign w2351 = ~w2349 & ~w2350;
assign w2352 = w2339 & ~w2351;
assign w2353 = w1066 & ~w1068;
assign w2354 = ~w2348 & ~w2353;
assign w2355 = ~w2352 & w2354;
assign w2356 = (~w1806 & w3778) | (~w1806 & w3779) | (w3778 & w3779);
assign w2357 = ~w1069 & ~w2356;
assign w2358 = (~w2238 & w3129) | (~w2238 & w3130) | (w3129 & w3130);
assign w2359 = (w2238 & w3131) | (w2238 & w3132) | (w3131 & w3132);
assign w2360 = ~w2358 & ~w2359;
assign w2361 = (w2238 & w3133) | (w2238 & w3134) | (w3133 & w3134);
assign w2362 = (~w2238 & w3135) | (~w2238 & w3136) | (w3135 & w3136);
assign w2363 = ~w2361 & ~w2362;
assign w2364 = (w2238 & w3137) | (w2238 & w3138) | (w3137 & w3138);
assign w2365 = (~w2238 & w3139) | (~w2238 & w3140) | (w3139 & w3140);
assign w2366 = ~w2364 & ~w2365;
assign w2367 = (w2238 & w3141) | (w2238 & w3142) | (w3141 & w3142);
assign w2368 = (~w2238 & w3143) | (~w2238 & w3144) | (w3143 & w3144);
assign w2369 = ~w2367 & ~w2368;
assign w2370 = (w2238 & w3145) | (w2238 & w3146) | (w3145 & w3146);
assign w2371 = (~w2238 & w3147) | (~w2238 & w3148) | (w3147 & w3148);
assign w2372 = ~w2370 & ~w2371;
assign w2373 = (w2238 & w3149) | (w2238 & w3150) | (w3149 & w3150);
assign w2374 = (~w2238 & w3151) | (~w2238 & w3152) | (w3151 & w3152);
assign w2375 = ~w2373 & ~w2374;
assign w2376 = (w2238 & w3153) | (w2238 & w3154) | (w3153 & w3154);
assign w2377 = (~w2238 & w3155) | (~w2238 & w3156) | (w3155 & w3156);
assign w2378 = ~w2376 & ~w2377;
assign w2379 = (w2238 & w3157) | (w2238 & w3158) | (w3157 & w3158);
assign w2380 = (~w2238 & w3159) | (~w2238 & w3160) | (w3159 & w3160);
assign w2381 = ~w2379 & ~w2380;
assign w2382 = (w2238 & w3161) | (w2238 & w3162) | (w3161 & w3162);
assign w2383 = (~w2238 & w3163) | (~w2238 & w3164) | (w3163 & w3164);
assign w2384 = ~w2382 & ~w2383;
assign w2385 = (w2238 & w3165) | (w2238 & w3166) | (w3165 & w3166);
assign w2386 = (~w2238 & w3167) | (~w2238 & w3168) | (w3167 & w3168);
assign w2387 = ~w2385 & ~w2386;
assign w2388 = (w2238 & w3169) | (w2238 & w3170) | (w3169 & w3170);
assign w2389 = (~w2238 & w3171) | (~w2238 & w3172) | (w3171 & w3172);
assign w2390 = ~w2388 & ~w2389;
assign w2391 = (w2238 & w3173) | (w2238 & w3174) | (w3173 & w3174);
assign w2392 = (~w2238 & w3175) | (~w2238 & w3176) | (w3175 & w3176);
assign w2393 = ~w2391 & ~w2392;
assign w2394 = (w2238 & w3177) | (w2238 & w3178) | (w3177 & w3178);
assign w2395 = (~w2238 & w3179) | (~w2238 & w3180) | (w3179 & w3180);
assign w2396 = ~w2394 & ~w2395;
assign w2397 = (w2238 & w3181) | (w2238 & w3182) | (w3181 & w3182);
assign w2398 = (~w2238 & w3183) | (~w2238 & w3184) | (w3183 & w3184);
assign w2399 = ~w2397 & ~w2398;
assign w2400 = (w2238 & w3185) | (w2238 & w3186) | (w3185 & w3186);
assign w2401 = (~w2238 & w3187) | (~w2238 & w3188) | (w3187 & w3188);
assign w2402 = ~w2400 & ~w2401;
assign w2403 = (w2238 & w3189) | (w2238 & w3190) | (w3189 & w3190);
assign w2404 = (~w2238 & w3191) | (~w2238 & w3192) | (w3191 & w3192);
assign w2405 = ~w2403 & ~w2404;
assign w2406 = (w2238 & w3193) | (w2238 & w3194) | (w3193 & w3194);
assign w2407 = (~w2238 & w3195) | (~w2238 & w3196) | (w3195 & w3196);
assign w2408 = ~w2406 & ~w2407;
assign w2409 = (w2238 & w3197) | (w2238 & w3198) | (w3197 & w3198);
assign w2410 = (~w2238 & w3199) | (~w2238 & w3200) | (w3199 & w3200);
assign w2411 = ~w2409 & ~w2410;
assign w2412 = (w2238 & w3201) | (w2238 & w3202) | (w3201 & w3202);
assign w2413 = (~w2238 & w3203) | (~w2238 & w3204) | (w3203 & w3204);
assign w2414 = ~w2412 & ~w2413;
assign w2415 = (w2238 & w3205) | (w2238 & w3206) | (w3205 & w3206);
assign w2416 = (~w2238 & w3207) | (~w2238 & w3208) | (w3207 & w3208);
assign w2417 = ~w2415 & ~w2416;
assign w2418 = (w2238 & w3209) | (w2238 & w3210) | (w3209 & w3210);
assign w2419 = (~w2238 & w3211) | (~w2238 & w3212) | (w3211 & w3212);
assign w2420 = ~w2418 & ~w2419;
assign w2421 = (w2238 & w3213) | (w2238 & w3214) | (w3213 & w3214);
assign w2422 = (~w2238 & w3215) | (~w2238 & w3216) | (w3215 & w3216);
assign w2423 = ~w2421 & ~w2422;
assign w2424 = (w2238 & w3217) | (w2238 & w3218) | (w3217 & w3218);
assign w2425 = (~w2238 & w3219) | (~w2238 & w3220) | (w3219 & w3220);
assign w2426 = ~w2424 & ~w2425;
assign w2427 = (w2238 & w3221) | (w2238 & w3222) | (w3221 & w3222);
assign w2428 = (~w2238 & w3223) | (~w2238 & w3224) | (w3223 & w3224);
assign w2429 = ~w2427 & ~w2428;
assign w2430 = (w2238 & w3225) | (w2238 & w3226) | (w3225 & w3226);
assign w2431 = (~w2238 & w3227) | (~w2238 & w3228) | (w3227 & w3228);
assign w2432 = ~w2430 & ~w2431;
assign w2433 = (w2238 & w3229) | (w2238 & w3230) | (w3229 & w3230);
assign w2434 = (~w2238 & w3231) | (~w2238 & w3232) | (w3231 & w3232);
assign w2435 = ~w2433 & ~w2434;
assign w2436 = (w2238 & w3233) | (w2238 & w3234) | (w3233 & w3234);
assign w2437 = (~w2238 & w3235) | (~w2238 & w3236) | (w3235 & w3236);
assign w2438 = ~w2436 & ~w2437;
assign w2439 = (w2238 & w3237) | (w2238 & w3238) | (w3237 & w3238);
assign w2440 = (~w2238 & w3239) | (~w2238 & w3240) | (w3239 & w3240);
assign w2441 = ~w2439 & ~w2440;
assign w2442 = (w2238 & w3241) | (w2238 & w3242) | (w3241 & w3242);
assign w2443 = (~w2238 & w3243) | (~w2238 & w3244) | (w3243 & w3244);
assign w2444 = ~w2442 & ~w2443;
assign w2445 = (w2238 & w3245) | (w2238 & w3246) | (w3245 & w3246);
assign w2446 = (~w2238 & w3247) | (~w2238 & w3248) | (w3247 & w3248);
assign w2447 = ~w2445 & ~w2446;
assign w2448 = (w2238 & w3249) | (w2238 & w3250) | (w3249 & w3250);
assign w2449 = (~w2238 & w3251) | (~w2238 & w3252) | (w3251 & w3252);
assign w2450 = ~w2448 & ~w2449;
assign w2451 = (w2238 & w3253) | (w2238 & w3254) | (w3253 & w3254);
assign w2452 = (~w2238 & w3255) | (~w2238 & w3256) | (w3255 & w3256);
assign w2453 = ~w2451 & ~w2452;
assign w2454 = (w2238 & w3257) | (w2238 & w3258) | (w3257 & w3258);
assign w2455 = (~w2238 & w3259) | (~w2238 & w3260) | (w3259 & w3260);
assign w2456 = ~w2454 & ~w2455;
assign w2457 = (w2238 & w3261) | (w2238 & w3262) | (w3261 & w3262);
assign w2458 = (~w2238 & w3263) | (~w2238 & w3264) | (w3263 & w3264);
assign w2459 = ~w2457 & ~w2458;
assign w2460 = (w2238 & w3265) | (w2238 & w3266) | (w3265 & w3266);
assign w2461 = (~w2238 & w3267) | (~w2238 & w3268) | (w3267 & w3268);
assign w2462 = ~w2460 & ~w2461;
assign w2463 = (w2238 & w3269) | (w2238 & w3270) | (w3269 & w3270);
assign w2464 = (~w2238 & w3271) | (~w2238 & w3272) | (w3271 & w3272);
assign w2465 = ~w2463 & ~w2464;
assign w2466 = (w2238 & w3273) | (w2238 & w3274) | (w3273 & w3274);
assign w2467 = (~w2238 & w3275) | (~w2238 & w3276) | (w3275 & w3276);
assign w2468 = ~w2466 & ~w2467;
assign w2469 = (w2238 & w3277) | (w2238 & w3278) | (w3277 & w3278);
assign w2470 = (~w2238 & w3279) | (~w2238 & w3280) | (w3279 & w3280);
assign w2471 = ~w2469 & ~w2470;
assign w2472 = (w2238 & w3281) | (w2238 & w3282) | (w3281 & w3282);
assign w2473 = (~w2238 & w3283) | (~w2238 & w3284) | (w3283 & w3284);
assign w2474 = ~w2472 & ~w2473;
assign w2475 = (w2238 & w3285) | (w2238 & w3286) | (w3285 & w3286);
assign w2476 = (~w2238 & w3287) | (~w2238 & w3288) | (w3287 & w3288);
assign w2477 = ~w2475 & ~w2476;
assign w2478 = (w2238 & w3289) | (w2238 & w3290) | (w3289 & w3290);
assign w2479 = (~w2238 & w3291) | (~w2238 & w3292) | (w3291 & w3292);
assign w2480 = ~w2478 & ~w2479;
assign w2481 = (w2238 & w3293) | (w2238 & w3294) | (w3293 & w3294);
assign w2482 = (~w2238 & w3295) | (~w2238 & w3296) | (w3295 & w3296);
assign w2483 = ~w2481 & ~w2482;
assign w2484 = (w2238 & w3297) | (w2238 & w3298) | (w3297 & w3298);
assign w2485 = (~w2238 & w3299) | (~w2238 & w3300) | (w3299 & w3300);
assign w2486 = ~w2484 & ~w2485;
assign w2487 = (w2238 & w3301) | (w2238 & w3302) | (w3301 & w3302);
assign w2488 = (~w2238 & w3303) | (~w2238 & w3304) | (w3303 & w3304);
assign w2489 = ~w2487 & ~w2488;
assign w2490 = (w2238 & w3305) | (w2238 & w3306) | (w3305 & w3306);
assign w2491 = (~w2238 & w3307) | (~w2238 & w3308) | (w3307 & w3308);
assign w2492 = ~w2490 & ~w2491;
assign w2493 = (w2238 & w3309) | (w2238 & w3310) | (w3309 & w3310);
assign w2494 = (~w2238 & w3311) | (~w2238 & w3312) | (w3311 & w3312);
assign w2495 = ~w2493 & ~w2494;
assign w2496 = (w2238 & w3313) | (w2238 & w3314) | (w3313 & w3314);
assign w2497 = (~w2238 & w3315) | (~w2238 & w3316) | (w3315 & w3316);
assign w2498 = ~w2496 & ~w2497;
assign w2499 = (w2238 & w3317) | (w2238 & w3318) | (w3317 & w3318);
assign w2500 = (~w2238 & w3319) | (~w2238 & w3320) | (w3319 & w3320);
assign w2501 = ~w2499 & ~w2500;
assign w2502 = (w2238 & w3321) | (w2238 & w3322) | (w3321 & w3322);
assign w2503 = (~w2238 & w3323) | (~w2238 & w3324) | (w3323 & w3324);
assign w2504 = ~w2502 & ~w2503;
assign w2505 = (w2238 & w3325) | (w2238 & w3326) | (w3325 & w3326);
assign w2506 = (~w2238 & w3327) | (~w2238 & w3328) | (w3327 & w3328);
assign w2507 = ~w2505 & ~w2506;
assign w2508 = (w2238 & w3329) | (w2238 & w3330) | (w3329 & w3330);
assign w2509 = (~w2238 & w3331) | (~w2238 & w3332) | (w3331 & w3332);
assign w2510 = ~w2508 & ~w2509;
assign w2511 = (w2238 & w3333) | (w2238 & w3334) | (w3333 & w3334);
assign w2512 = (~w2238 & w3335) | (~w2238 & w3336) | (w3335 & w3336);
assign w2513 = ~w2511 & ~w2512;
assign w2514 = (w2238 & w3337) | (w2238 & w3338) | (w3337 & w3338);
assign w2515 = (~w2238 & w3339) | (~w2238 & w3340) | (w3339 & w3340);
assign w2516 = ~w2514 & ~w2515;
assign w2517 = (w2238 & w3341) | (w2238 & w3342) | (w3341 & w3342);
assign w2518 = (~w2238 & w3343) | (~w2238 & w3344) | (w3343 & w3344);
assign w2519 = ~w2517 & ~w2518;
assign w2520 = (w2238 & w3345) | (w2238 & w3346) | (w3345 & w3346);
assign w2521 = (~w2238 & w3347) | (~w2238 & w3348) | (w3347 & w3348);
assign w2522 = ~w2520 & ~w2521;
assign w2523 = (w2238 & w3349) | (w2238 & w3350) | (w3349 & w3350);
assign w2524 = (~w2238 & w3351) | (~w2238 & w3352) | (w3351 & w3352);
assign w2525 = ~w2523 & ~w2524;
assign w2526 = (w2238 & w3353) | (w2238 & w3354) | (w3353 & w3354);
assign w2527 = (~w2238 & w3355) | (~w2238 & w3356) | (w3355 & w3356);
assign w2528 = ~w2526 & ~w2527;
assign w2529 = (w2238 & w3357) | (w2238 & w3358) | (w3357 & w3358);
assign w2530 = (~w2238 & w3359) | (~w2238 & w3360) | (w3359 & w3360);
assign w2531 = ~w2529 & ~w2530;
assign w2532 = (w2238 & w3361) | (w2238 & w3362) | (w3361 & w3362);
assign w2533 = (~w2238 & w3363) | (~w2238 & w3364) | (w3363 & w3364);
assign w2534 = ~w2532 & ~w2533;
assign w2535 = (w2238 & w3365) | (w2238 & w3366) | (w3365 & w3366);
assign w2536 = (~w2238 & w3367) | (~w2238 & w3368) | (w3367 & w3368);
assign w2537 = ~w2535 & ~w2536;
assign w2538 = (w2238 & w3369) | (w2238 & w3370) | (w3369 & w3370);
assign w2539 = (~w2238 & w3371) | (~w2238 & w3372) | (w3371 & w3372);
assign w2540 = ~w2538 & ~w2539;
assign w2541 = (w2238 & w3373) | (w2238 & w3374) | (w3373 & w3374);
assign w2542 = (~w2238 & w3375) | (~w2238 & w3376) | (w3375 & w3376);
assign w2543 = ~w2541 & ~w2542;
assign w2544 = (w2238 & w3377) | (w2238 & w3378) | (w3377 & w3378);
assign w2545 = (~w2238 & w3379) | (~w2238 & w3380) | (w3379 & w3380);
assign w2546 = ~w2544 & ~w2545;
assign w2547 = (w2238 & w3381) | (w2238 & w3382) | (w3381 & w3382);
assign w2548 = (~w2238 & w3383) | (~w2238 & w3384) | (w3383 & w3384);
assign w2549 = ~w2547 & ~w2548;
assign w2550 = (w2238 & w3385) | (w2238 & w3386) | (w3385 & w3386);
assign w2551 = (~w2238 & w3387) | (~w2238 & w3388) | (w3387 & w3388);
assign w2552 = ~w2550 & ~w2551;
assign w2553 = (w2238 & w3389) | (w2238 & w3390) | (w3389 & w3390);
assign w2554 = (~w2238 & w3391) | (~w2238 & w3392) | (w3391 & w3392);
assign w2555 = ~w2553 & ~w2554;
assign w2556 = (w2238 & w3393) | (w2238 & w3394) | (w3393 & w3394);
assign w2557 = (~w2238 & w3395) | (~w2238 & w3396) | (w3395 & w3396);
assign w2558 = ~w2556 & ~w2557;
assign w2559 = (w2238 & w3397) | (w2238 & w3398) | (w3397 & w3398);
assign w2560 = (~w2238 & w3399) | (~w2238 & w3400) | (w3399 & w3400);
assign w2561 = ~w2559 & ~w2560;
assign w2562 = (w2238 & w3401) | (w2238 & w3402) | (w3401 & w3402);
assign w2563 = (~w2238 & w3403) | (~w2238 & w3404) | (w3403 & w3404);
assign w2564 = ~w2562 & ~w2563;
assign w2565 = (w2238 & w3405) | (w2238 & w3406) | (w3405 & w3406);
assign w2566 = (~w2238 & w3407) | (~w2238 & w3408) | (w3407 & w3408);
assign w2567 = ~w2565 & ~w2566;
assign w2568 = (w2238 & w3409) | (w2238 & w3410) | (w3409 & w3410);
assign w2569 = (~w2238 & w3411) | (~w2238 & w3412) | (w3411 & w3412);
assign w2570 = ~w2568 & ~w2569;
assign w2571 = (w2238 & w3413) | (w2238 & w3414) | (w3413 & w3414);
assign w2572 = (~w2238 & w3415) | (~w2238 & w3416) | (w3415 & w3416);
assign w2573 = ~w2571 & ~w2572;
assign w2574 = (w2238 & w3417) | (w2238 & w3418) | (w3417 & w3418);
assign w2575 = (~w2238 & w3419) | (~w2238 & w3420) | (w3419 & w3420);
assign w2576 = ~w2574 & ~w2575;
assign w2577 = (w2238 & w3421) | (w2238 & w3422) | (w3421 & w3422);
assign w2578 = (~w2238 & w3423) | (~w2238 & w3424) | (w3423 & w3424);
assign w2579 = ~w2577 & ~w2578;
assign w2580 = (w2238 & w3425) | (w2238 & w3426) | (w3425 & w3426);
assign w2581 = (~w2238 & w3427) | (~w2238 & w3428) | (w3427 & w3428);
assign w2582 = ~w2580 & ~w2581;
assign w2583 = (w2238 & w3429) | (w2238 & w3430) | (w3429 & w3430);
assign w2584 = (~w2238 & w3431) | (~w2238 & w3432) | (w3431 & w3432);
assign w2585 = ~w2583 & ~w2584;
assign w2586 = (w2238 & w3433) | (w2238 & w3434) | (w3433 & w3434);
assign w2587 = (~w2238 & w3435) | (~w2238 & w3436) | (w3435 & w3436);
assign w2588 = ~w2586 & ~w2587;
assign w2589 = (w2238 & w3437) | (w2238 & w3438) | (w3437 & w3438);
assign w2590 = (~w2238 & w3439) | (~w2238 & w3440) | (w3439 & w3440);
assign w2591 = ~w2589 & ~w2590;
assign w2592 = (w2238 & w3441) | (w2238 & w3442) | (w3441 & w3442);
assign w2593 = (~w2238 & w3443) | (~w2238 & w3444) | (w3443 & w3444);
assign w2594 = ~w2592 & ~w2593;
assign w2595 = (w2238 & w3445) | (w2238 & w3446) | (w3445 & w3446);
assign w2596 = (~w2238 & w3447) | (~w2238 & w3448) | (w3447 & w3448);
assign w2597 = ~w2595 & ~w2596;
assign w2598 = (w2238 & w3449) | (w2238 & w3450) | (w3449 & w3450);
assign w2599 = (~w2238 & w3451) | (~w2238 & w3452) | (w3451 & w3452);
assign w2600 = ~w2598 & ~w2599;
assign w2601 = (w2238 & w3453) | (w2238 & w3454) | (w3453 & w3454);
assign w2602 = (~w2238 & w3455) | (~w2238 & w3456) | (w3455 & w3456);
assign w2603 = ~w2601 & ~w2602;
assign w2604 = (w2238 & w3457) | (w2238 & w3458) | (w3457 & w3458);
assign w2605 = (~w2238 & w3459) | (~w2238 & w3460) | (w3459 & w3460);
assign w2606 = ~w2604 & ~w2605;
assign w2607 = (w2238 & w3461) | (w2238 & w3462) | (w3461 & w3462);
assign w2608 = (~w2238 & w3463) | (~w2238 & w3464) | (w3463 & w3464);
assign w2609 = ~w2607 & ~w2608;
assign w2610 = (w2238 & w3465) | (w2238 & w3466) | (w3465 & w3466);
assign w2611 = (~w2238 & w3467) | (~w2238 & w3468) | (w3467 & w3468);
assign w2612 = ~w2610 & ~w2611;
assign w2613 = (w2238 & w3469) | (w2238 & w3470) | (w3469 & w3470);
assign w2614 = (~w2238 & w3471) | (~w2238 & w3472) | (w3471 & w3472);
assign w2615 = ~w2613 & ~w2614;
assign w2616 = (w2238 & w3473) | (w2238 & w3474) | (w3473 & w3474);
assign w2617 = (~w2238 & w3475) | (~w2238 & w3476) | (w3475 & w3476);
assign w2618 = ~w2616 & ~w2617;
assign w2619 = (w2238 & w3477) | (w2238 & w3478) | (w3477 & w3478);
assign w2620 = (~w2238 & w3479) | (~w2238 & w3480) | (w3479 & w3480);
assign w2621 = ~w2619 & ~w2620;
assign w2622 = (w2238 & w3481) | (w2238 & w3482) | (w3481 & w3482);
assign w2623 = (~w2238 & w3483) | (~w2238 & w3484) | (w3483 & w3484);
assign w2624 = ~w2622 & ~w2623;
assign w2625 = (w2238 & w3485) | (w2238 & w3486) | (w3485 & w3486);
assign w2626 = (~w2238 & w3487) | (~w2238 & w3488) | (w3487 & w3488);
assign w2627 = ~w2625 & ~w2626;
assign w2628 = (w2238 & w3489) | (w2238 & w3490) | (w3489 & w3490);
assign w2629 = (~w2238 & w3491) | (~w2238 & w3492) | (w3491 & w3492);
assign w2630 = ~w2628 & ~w2629;
assign w2631 = (w2238 & w3493) | (w2238 & w3494) | (w3493 & w3494);
assign w2632 = (~w2238 & w3495) | (~w2238 & w3496) | (w3495 & w3496);
assign w2633 = ~w2631 & ~w2632;
assign w2634 = (w2238 & w3497) | (w2238 & w3498) | (w3497 & w3498);
assign w2635 = (~w2238 & w3499) | (~w2238 & w3500) | (w3499 & w3500);
assign w2636 = ~w2634 & ~w2635;
assign w2637 = (w2238 & w3501) | (w2238 & w3502) | (w3501 & w3502);
assign w2638 = (~w2238 & w3503) | (~w2238 & w3504) | (w3503 & w3504);
assign w2639 = ~w2637 & ~w2638;
assign w2640 = (w2238 & w3505) | (w2238 & w3506) | (w3505 & w3506);
assign w2641 = (~w2238 & w3507) | (~w2238 & w3508) | (w3507 & w3508);
assign w2642 = ~w2640 & ~w2641;
assign w2643 = (w2238 & w3509) | (w2238 & w3510) | (w3509 & w3510);
assign w2644 = (~w2238 & w3511) | (~w2238 & w3512) | (w3511 & w3512);
assign w2645 = ~w2643 & ~w2644;
assign w2646 = (w2238 & w3513) | (w2238 & w3514) | (w3513 & w3514);
assign w2647 = (~w2238 & w3515) | (~w2238 & w3516) | (w3515 & w3516);
assign w2648 = ~w2646 & ~w2647;
assign w2649 = (w2238 & w3517) | (w2238 & w3518) | (w3517 & w3518);
assign w2650 = (~w2238 & w3519) | (~w2238 & w3520) | (w3519 & w3520);
assign w2651 = ~w2649 & ~w2650;
assign w2652 = (w2238 & w3521) | (w2238 & w3522) | (w3521 & w3522);
assign w2653 = (~w2238 & w3523) | (~w2238 & w3524) | (w3523 & w3524);
assign w2654 = ~w2652 & ~w2653;
assign w2655 = (w2238 & w3525) | (w2238 & w3526) | (w3525 & w3526);
assign w2656 = (~w2238 & w3527) | (~w2238 & w3528) | (w3527 & w3528);
assign w2657 = ~w2655 & ~w2656;
assign w2658 = (w2238 & w3529) | (w2238 & w3530) | (w3529 & w3530);
assign w2659 = (~w2238 & w3531) | (~w2238 & w3532) | (w3531 & w3532);
assign w2660 = ~w2658 & ~w2659;
assign w2661 = (w2238 & w3533) | (w2238 & w3534) | (w3533 & w3534);
assign w2662 = (~w2238 & w3535) | (~w2238 & w3536) | (w3535 & w3536);
assign w2663 = ~w2661 & ~w2662;
assign w2664 = (w2238 & w3537) | (w2238 & w3538) | (w3537 & w3538);
assign w2665 = (~w2238 & w3539) | (~w2238 & w3540) | (w3539 & w3540);
assign w2666 = ~w2664 & ~w2665;
assign w2667 = (w2238 & w3541) | (w2238 & w3542) | (w3541 & w3542);
assign w2668 = (~w2238 & w3543) | (~w2238 & w3544) | (w3543 & w3544);
assign w2669 = ~w2667 & ~w2668;
assign w2670 = (w2238 & w3545) | (w2238 & w3546) | (w3545 & w3546);
assign w2671 = (~w2238 & w3547) | (~w2238 & w3548) | (w3547 & w3548);
assign w2672 = ~w2670 & ~w2671;
assign w2673 = (w2238 & w3549) | (w2238 & w3550) | (w3549 & w3550);
assign w2674 = (~w2238 & w3551) | (~w2238 & w3552) | (w3551 & w3552);
assign w2675 = ~w2673 & ~w2674;
assign w2676 = (w2238 & w3553) | (w2238 & w3554) | (w3553 & w3554);
assign w2677 = (~w2238 & w3555) | (~w2238 & w3556) | (w3555 & w3556);
assign w2678 = ~w2676 & ~w2677;
assign w2679 = (w2238 & w3557) | (w2238 & w3558) | (w3557 & w3558);
assign w2680 = (~w2238 & w3559) | (~w2238 & w3560) | (w3559 & w3560);
assign w2681 = ~w2679 & ~w2680;
assign w2682 = (w2238 & w3561) | (w2238 & w3562) | (w3561 & w3562);
assign w2683 = (~w2238 & w3563) | (~w2238 & w3564) | (w3563 & w3564);
assign w2684 = ~w2682 & ~w2683;
assign w2685 = (w2238 & w3565) | (w2238 & w3566) | (w3565 & w3566);
assign w2686 = (~w2238 & w3567) | (~w2238 & w3568) | (w3567 & w3568);
assign w2687 = ~w2685 & ~w2686;
assign w2688 = (w2238 & w3569) | (w2238 & w3570) | (w3569 & w3570);
assign w2689 = (~w2238 & w3571) | (~w2238 & w3572) | (w3571 & w3572);
assign w2690 = ~w2688 & ~w2689;
assign w2691 = (w2238 & w3573) | (w2238 & w3574) | (w3573 & w3574);
assign w2692 = (~w2238 & w3575) | (~w2238 & w3576) | (w3575 & w3576);
assign w2693 = ~w2691 & ~w2692;
assign w2694 = (w2238 & w3577) | (w2238 & w3578) | (w3577 & w3578);
assign w2695 = (~w2238 & w3579) | (~w2238 & w3580) | (w3579 & w3580);
assign w2696 = ~w2694 & ~w2695;
assign w2697 = (w2238 & w3581) | (w2238 & w3582) | (w3581 & w3582);
assign w2698 = (~w2238 & w3583) | (~w2238 & w3584) | (w3583 & w3584);
assign w2699 = ~w2697 & ~w2698;
assign w2700 = (w2238 & w3585) | (w2238 & w3586) | (w3585 & w3586);
assign w2701 = (~w2238 & w3587) | (~w2238 & w3588) | (w3587 & w3588);
assign w2702 = ~w2700 & ~w2701;
assign w2703 = (w2238 & w3589) | (w2238 & w3590) | (w3589 & w3590);
assign w2704 = (~w2238 & w3591) | (~w2238 & w3592) | (w3591 & w3592);
assign w2705 = ~w2703 & ~w2704;
assign w2706 = (w2238 & w3593) | (w2238 & w3594) | (w3593 & w3594);
assign w2707 = (~w2238 & w3595) | (~w2238 & w3596) | (w3595 & w3596);
assign w2708 = ~w2706 & ~w2707;
assign w2709 = (w2238 & w3597) | (w2238 & w3598) | (w3597 & w3598);
assign w2710 = (~w2238 & w3599) | (~w2238 & w3600) | (w3599 & w3600);
assign w2711 = ~w2709 & ~w2710;
assign w2712 = (w2238 & w3601) | (w2238 & w3602) | (w3601 & w3602);
assign w2713 = (~w2238 & w3603) | (~w2238 & w3604) | (w3603 & w3604);
assign w2714 = ~w2712 & ~w2713;
assign w2715 = (w2238 & w3605) | (w2238 & w3606) | (w3605 & w3606);
assign w2716 = (~w2238 & w3607) | (~w2238 & w3608) | (w3607 & w3608);
assign w2717 = ~w2715 & ~w2716;
assign w2718 = (w2238 & w3609) | (w2238 & w3610) | (w3609 & w3610);
assign w2719 = (~w2238 & w3611) | (~w2238 & w3612) | (w3611 & w3612);
assign w2720 = ~w2718 & ~w2719;
assign w2721 = (w2238 & w3613) | (w2238 & w3614) | (w3613 & w3614);
assign w2722 = (~w2238 & w3615) | (~w2238 & w3616) | (w3615 & w3616);
assign w2723 = ~w2721 & ~w2722;
assign w2724 = (w2238 & w3617) | (w2238 & w3618) | (w3617 & w3618);
assign w2725 = (~w2238 & w3619) | (~w2238 & w3620) | (w3619 & w3620);
assign w2726 = ~w2724 & ~w2725;
assign w2727 = (w2238 & w3621) | (w2238 & w3622) | (w3621 & w3622);
assign w2728 = (~w2238 & w3623) | (~w2238 & w3624) | (w3623 & w3624);
assign w2729 = ~w2727 & ~w2728;
assign w2730 = (w2238 & w3625) | (w2238 & w3626) | (w3625 & w3626);
assign w2731 = (~w2238 & w3627) | (~w2238 & w3628) | (w3627 & w3628);
assign w2732 = ~w2730 & ~w2731;
assign w2733 = (w2238 & w3629) | (w2238 & w3630) | (w3629 & w3630);
assign w2734 = (~w2238 & w3631) | (~w2238 & w3632) | (w3631 & w3632);
assign w2735 = ~w2733 & ~w2734;
assign w2736 = (w2238 & w3633) | (w2238 & w3634) | (w3633 & w3634);
assign w2737 = (~w2238 & w3635) | (~w2238 & w3636) | (w3635 & w3636);
assign w2738 = ~w2736 & ~w2737;
assign w2739 = w1066 & w1068;
assign w2740 = (w2238 & w3637) | (w2238 & w3638) | (w3637 & w3638);
assign w2741 = (~w2238 & w3639) | (~w2238 & w3640) | (w3639 & w3640);
assign w2742 = ~w2740 & ~w2741;
assign w2743 = ~w13 & w16;
assign w2744 = ~w551 & w554;
assign w2745 = w533 & pi001;
assign w2746 = ~w533 & pi129;
assign w2747 = w533 & pi002;
assign w2748 = ~w533 & pi130;
assign w2749 = ~w1130 & w1139;
assign w2750 = ~w1149 & w1152;
assign w2751 = w1099 & ~w1092;
assign w2752 = w1162 & w1092;
assign w2753 = w1162 & ~w2751;
assign w2754 = w1165 & ~w2753;
assign w2755 = w1165 & ~w2752;
assign w2756 = w1085 & ~w1078;
assign w2757 = w1175 & w1078;
assign w2758 = w1175 & ~w2756;
assign w2759 = w1192 & ~w2758;
assign w2760 = w1192 & ~w2757;
assign w2761 = w1204 & ~w2760;
assign w2762 = (w1213 & w2759) | (w1213 & w3050) | (w2759 & w3050);
assign w2763 = w1213 & ~w2761;
assign w2764 = ~w1223 & w1240;
assign w2765 = w1252 & ~w1240;
assign w2766 = (w1269 & w2764) | (w1269 & w3051) | (w2764 & w3051);
assign w2767 = (w1281 & w2765) | (w1281 & w3641) | (w2765 & w3641);
assign w2768 = w1281 & ~w2766;
assign w2769 = ~w1290 & w1299;
assign w2770 = w1316 & ~w1299;
assign w2771 = w1316 & ~w2769;
assign w2772 = (w1345 & w2770) | (w1345 & w3642) | (w2770 & w3642);
assign w2773 = (w1345 & w2771) | (w1345 & w3642) | (w2771 & w3642);
assign w2774 = w533 & pi049;
assign w2775 = ~w533 & pi177;
assign w2776 = w533 & pi050;
assign w2777 = ~w533 & pi178;
assign w2778 = w533 & pi048;
assign w2779 = ~w533 & pi176;
assign w2780 = ~w1686 & w1650;
assign w2781 = (~w1692 & w3643) | (~w1692 & w3644) | (w3643 & w3644);
assign w2782 = w1986 & ~w1930;
assign w2783 = w2054 & ~w2782;
assign w2784 = (~w2782 & w4195) | (~w2782 & w4196) | (w4195 & w4196);
assign w2785 = (w2179 & w2783) | (w2179 & w3645) | (w2783 & w3645);
assign w2786 = (w2179 & w2784) | (w2179 & w3645) | (w2784 & w3645);
assign w2787 = w2237 & ~w2785;
assign w2788 = w2237 & ~w2786;
assign w2789 = ~w2323 & w3646;
assign w2790 = w2347 & ~w2324;
assign w2791 = w2347 & ~w2789;
assign w2792 = w2355 & ~w2790;
assign w2793 = w2355 & ~w2791;
assign w2794 = ~w1069 & ~w537;
assign w2795 = w1069 & ~w1109;
assign w2796 = w1069 & ~w1105;
assign w2797 = ~w1069 & ~w1102;
assign w2798 = w1069 & ~w1118;
assign w2799 = ~w1069 & ~w1115;
assign w2800 = w1069 & ~w1127;
assign w2801 = ~w1069 & ~w1124;
assign w2802 = w1069 & ~w1136;
assign w2803 = ~w1069 & ~w1133;
assign w2804 = w1069 & ~w1147;
assign w2805 = ~w1069 & ~w1144;
assign w2806 = w1069 & ~w1098;
assign w2807 = ~w1069 & ~w1095;
assign w2808 = w1069 & ~w1091;
assign w2809 = ~w1069 & ~w1088;
assign w2810 = w1069 & w1156;
assign w2811 = ~w1069 & w1159;
assign w2812 = w1069 & ~w1084;
assign w2813 = ~w1069 & ~w1081;
assign w2814 = w1069 & ~w1077;
assign w2815 = ~w1069 & ~w1072;
assign w2816 = w1069 & ~w1172;
assign w2817 = ~w1069 & ~w1169;
assign w2818 = w1069 & w1185;
assign w2819 = ~w1069 & w1188;
assign w2820 = w1069 & ~w1181;
assign w2821 = ~w1069 & ~w1178;
assign w2822 = w1069 & ~w1199;
assign w2823 = ~w1069 & ~w1196;
assign w2824 = w1069 & ~w1210;
assign w2825 = ~w1069 & ~w1207;
assign w2826 = w1069 & ~w1221;
assign w2827 = ~w1069 & ~w1218;
assign w2828 = w1069 & ~w1237;
assign w2829 = ~w1069 & ~w1234;
assign w2830 = w1069 & ~w1230;
assign w2831 = ~w1069 & ~w1227;
assign w2832 = w1069 & ~w1246;
assign w2833 = ~w1069 & ~w1243;
assign w2834 = w1069 & ~w1266;
assign w2835 = ~w1069 & ~w1263;
assign w2836 = w1069 & ~w1259;
assign w2837 = ~w1069 & ~w1256;
assign w2838 = w1069 & ~w1275;
assign w2839 = ~w1069 & ~w1272;
assign w2840 = w1069 & ~w1287;
assign w2841 = ~w1069 & ~w1284;
assign w2842 = w1069 & ~w1296;
assign w2843 = ~w1069 & ~w1293;
assign w2844 = w1069 & ~w1312;
assign w2845 = ~w1069 & ~w1309;
assign w2846 = w1069 & ~w1305;
assign w2847 = ~w1069 & ~w1302;
assign w2848 = w1069 & ~w1322;
assign w2849 = ~w1069 & ~w1319;
assign w2850 = w1069 & ~w1342;
assign w2851 = ~w1069 & ~w1339;
assign w2852 = w1069 & ~w1335;
assign w2853 = ~w1069 & ~w1332;
assign w2854 = w1069 & ~w1351;
assign w2855 = ~w1069 & ~w1348;
assign w2856 = w1069 & ~w1423;
assign w2857 = ~w1069 & ~w1420;
assign w2858 = w1069 & w1413;
assign w2859 = ~w1069 & w1416;
assign w2860 = w1069 & ~w1363;
assign w2861 = ~w1069 & ~w1360;
assign w2862 = w1069 & w1367;
assign w2863 = ~w1069 & w1370;
assign w2864 = w1069 & ~w1400;
assign w2865 = ~w1069 & ~w1397;
assign w2866 = w1069 & ~w1393;
assign w2867 = ~w1069 & ~w1390;
assign w2868 = w1069 & ~w1385;
assign w2869 = ~w1069 & ~w1382;
assign w2870 = w1069 & w1375;
assign w2871 = ~w1069 & w1378;
assign w2872 = w1069 & ~w1409;
assign w2873 = ~w1069 & ~w1406;
assign w2874 = w1069 & w1511;
assign w2875 = ~w1069 & w1514;
assign w2876 = w1069 & ~w1507;
assign w2877 = ~w1069 & ~w1504;
assign w2878 = w1069 & ~w1498;
assign w2879 = ~w1069 & ~w1495;
assign w2880 = w1069 & ~w1491;
assign w2881 = ~w1069 & ~w1488;
assign w2882 = w1069 & ~w1482;
assign w2883 = ~w1069 & ~w1479;
assign w2884 = w1069 & ~w1472;
assign w2885 = ~w1069 & ~w1469;
assign w2886 = w1069 & ~w1453;
assign w2887 = ~w1069 & ~w1463;
assign w2888 = w1069 & ~w1459;
assign w2889 = ~w1069 & ~w1456;
assign w2890 = w1069 & w1653;
assign w2891 = ~w1069 & w1656;
assign w2892 = w1069 & ~w1557;
assign w2893 = ~w1069 & ~w1554;
assign w2894 = w1069 & w1561;
assign w2895 = ~w1069 & w1564;
assign w2896 = w1069 & ~w1601;
assign w2897 = ~w1069 & ~w1598;
assign w2898 = w1069 & w1591;
assign w2899 = ~w1069 & w1594;
assign w2900 = w1069 & ~w1587;
assign w2901 = ~w1069 & ~w1584;
assign w2902 = w1069 & w1638;
assign w2903 = ~w1069 & w1641;
assign w2904 = w1069 & w1645;
assign w2905 = ~w1069 & w1648;
assign w2906 = w1069 & w1549;
assign w2907 = ~w1069 & w1545;
assign w2908 = w1069 & ~w1541;
assign w2909 = ~w1069 & ~w1538;
assign w2910 = w1069 & ~w1579;
assign w2911 = ~w1069 & ~w1576;
assign w2912 = w1069 & ~w1572;
assign w2913 = ~w1069 & ~w1569;
assign w2914 = w1069 & ~w1610;
assign w2915 = ~w1069 & ~w1607;
assign w2916 = w1069 & ~w1631;
assign w2917 = ~w1069 & ~w1628;
assign w2918 = w1069 & w1621;
assign w2919 = ~w1069 & w1624;
assign w2920 = w1069 & ~w1617;
assign w2921 = ~w1069 & ~w1614;
assign w2922 = w1069 & w1719;
assign w2923 = ~w1069 & w1723;
assign w2924 = w1069 & ~w1714;
assign w2925 = ~w1069 & ~w1711;
assign w2926 = w1069 & w1703;
assign w2927 = ~w1069 & w1706;
assign w2928 = w1069 & ~w1698;
assign w2929 = ~w1069 & ~w1695;
assign w2930 = w1069 & ~w1777;
assign w2931 = ~w1069 & ~w1774;
assign w2932 = w1069 & ~w1769;
assign w2933 = ~w1069 & ~w1766;
assign w2934 = w1069 & w1759;
assign w2935 = ~w1069 & w1762;
assign w2936 = w1069 & ~w1798;
assign w2937 = ~w1069 & ~w1795;
assign w2938 = w1069 & w1788;
assign w2939 = ~w1069 & w1791;
assign w2940 = w1069 & ~w1784;
assign w2941 = ~w1069 & ~w1781;
assign w2942 = w1069 & w1747;
assign w2943 = ~w1069 & w1750;
assign w2944 = w1069 & ~w1743;
assign w2945 = ~w1069 & ~w1740;
assign w2946 = w1069 & w1840;
assign w2947 = ~w1069 & w1843;
assign w2948 = w1069 & ~w1836;
assign w2949 = ~w1069 & ~w1833;
assign w2950 = w1069 & ~w1852;
assign w2951 = ~w1069 & ~w1849;
assign w2952 = w1069 & ~w1829;
assign w2953 = ~w1069 & ~w1826;
assign w2954 = w1069 & w1866;
assign w2955 = ~w1069 & w1869;
assign w2956 = w1069 & ~w1925;
assign w2957 = ~w1069 & ~w1922;
assign w2958 = w1069 & w1899;
assign w2959 = ~w1069 & w1902;
assign w2960 = w1069 & ~w1916;
assign w2961 = ~w1069 & ~w1913;
assign w2962 = w1069 & ~w1909;
assign w2963 = ~w1069 & ~w1906;
assign w2964 = w1069 & ~w1879;
assign w2965 = ~w1069 & ~w1876;
assign w2966 = w1069 & w1890;
assign w2967 = ~w1069 & w1893;
assign w2968 = w1069 & ~w1886;
assign w2969 = ~w1069 & ~w1883;
assign w2970 = w1069 & w1959;
assign w2971 = ~w1069 & w1963;
assign w2972 = w1069 & ~w1954;
assign w2973 = ~w1069 & ~w1951;
assign w2974 = w1069 & w1943;
assign w2975 = ~w1069 & w1946;
assign w2976 = w1069 & ~w1938;
assign w2977 = ~w1069 & ~w1935;
assign w2978 = w1069 & ~w2026;
assign w2979 = ~w1069 & ~w2023;
assign w2980 = w1069 & ~w2011;
assign w2981 = ~w1069 & ~w2008;
assign w2982 = w1069 & w2015;
assign w2983 = ~w1069 & w2018;
assign w2984 = w1069 & ~w2033;
assign w2985 = ~w1069 & ~w2030;
assign w2986 = w1069 & w2044;
assign w2987 = ~w1069 & w2047;
assign w2988 = w1069 & ~w2040;
assign w2989 = ~w1069 & ~w2037;
assign w2990 = w1069 & w1996;
assign w2991 = ~w1069 & w1999;
assign w2992 = w1069 & ~w1992;
assign w2993 = ~w1069 & ~w1989;
assign w2994 = w1069 & w2089;
assign w2995 = ~w1069 & w2092;
assign w2996 = w1069 & ~w2085;
assign w2997 = ~w1069 & ~w2082;
assign w2998 = w1069 & ~w2101;
assign w2999 = ~w1069 & ~w2098;
assign w3000 = w1069 & ~w2078;
assign w3001 = ~w1069 & ~w2075;
assign w3002 = w1069 & w2115;
assign w3003 = ~w1069 & w2118;
assign w3004 = w1069 & ~w2174;
assign w3005 = ~w1069 & ~w2171;
assign w3006 = w1069 & w2148;
assign w3007 = ~w1069 & w2151;
assign w3008 = w1069 & ~w2165;
assign w3009 = ~w1069 & ~w2162;
assign w3010 = w1069 & ~w2158;
assign w3011 = ~w1069 & ~w2155;
assign w3012 = w1069 & ~w2128;
assign w3013 = ~w1069 & ~w2125;
assign w3014 = w1069 & w2139;
assign w3015 = ~w1069 & w2142;
assign w3016 = w1069 & ~w2135;
assign w3017 = ~w1069 & ~w2132;
assign w3018 = w1069 & w2208;
assign w3019 = ~w1069 & w2212;
assign w3020 = w1069 & ~w2203;
assign w3021 = ~w1069 & ~w2200;
assign w3022 = w1069 & w2192;
assign w3023 = ~w1069 & w2195;
assign w3024 = w1069 & ~w2187;
assign w3025 = ~w1069 & ~w2184;
assign w3026 = w1069 & w2267;
assign w3027 = ~w1069 & w2270;
assign w3028 = w1069 & ~w2299;
assign w3029 = ~w1069 & ~w2296;
assign w3030 = w1069 & w2289;
assign w3031 = ~w1069 & w2292;
assign w3032 = w1069 & ~w2277;
assign w3033 = ~w1069 & ~w2274;
assign w3034 = w1069 & w2281;
assign w3035 = ~w1069 & w2284;
assign w3036 = w1069 & ~w2263;
assign w3037 = ~w1069 & ~w2260;
assign w3038 = w1069 & w2248;
assign w3039 = ~w1069 & w2251;
assign w3040 = w1069 & ~w2244;
assign w3041 = ~w1069 & ~w2241;
assign w3042 = w1069 & ~w2345;
assign w3043 = ~w1069 & ~w2342;
assign w3044 = w1069 & ~w2337;
assign w3045 = ~w1069 & ~w2334;
assign w3046 = w1069 & ~w2330;
assign w3047 = ~w1069 & ~w2327;
assign w3048 = w1069 & w1074;
assign w3049 = ~w1069 & w534;
assign w3050 = ~w1204 & w1213;
assign w3051 = ~w1252 & w1269;
assign w3052 = ~w1737 & w1805;
assign w3053 = ~w20 & ~w3;
assign w3054 = w2 & w23;
assign w3055 = ~w540 & w541;
assign w3056 = (~w540 & w558) | (~w540 & w3055) | (w558 & w3055);
assign w3057 = ~w561 & w564;
assign w3058 = w533 & pi010;
assign w3059 = ~w533 & pi138;
assign w3060 = w533 & pi003;
assign w3061 = ~w533 & pi131;
assign w3062 = w533 & pi004;
assign w3063 = ~w533 & pi132;
assign w3064 = w533 & pi011;
assign w3065 = ~w533 & pi139;
assign w3066 = w533 & pi013;
assign w3067 = ~w533 & pi141;
assign w3068 = w533 & pi012;
assign w3069 = ~w533 & pi140;
assign w3070 = (w2773 & w2772) | (w2773 & ~w2768) | (w2772 & ~w2768);
assign w3071 = (w2773 & w2772) | (w2773 & ~w2767) | (w2772 & ~w2767);
assign w3072 = w533 & pi033;
assign w3073 = ~w533 & pi161;
assign w3074 = w533 & pi032;
assign w3075 = ~w533 & pi160;
assign w3076 = w533 & pi031;
assign w3077 = ~w533 & pi159;
assign w3078 = w1073 & pi287;
assign w3079 = ~w1073 & pi415;
assign w3080 = w1429 & w3780;
assign w3081 = ~w1444 & w1402;
assign w3082 = w531 & w2775;
assign w3083 = w1073 & pi305;
assign w3084 = ~w1073 & pi433;
assign w3085 = w1073 & pi306;
assign w3086 = ~w1073 & pi434;
assign w3087 = w531 & w2777;
assign w3088 = w533 & pi053;
assign w3089 = ~w533 & pi181;
assign w3090 = w533 & pi052;
assign w3091 = ~w533 & pi180;
assign w3092 = w533 & pi051;
assign w3093 = ~w533 & pi179;
assign w3094 = w533 & pi054;
assign w3095 = ~w533 & pi182;
assign w3096 = w1073 & pi304;
assign w3097 = ~w1073 & pi432;
assign w3098 = w531 & w2779;
assign w3099 = w533 & pi070;
assign w3100 = ~w533 & pi198;
assign w3101 = w533 & pi069;
assign w3102 = ~w533 & pi197;
assign w3103 = w533 & pi068;
assign w3104 = ~w533 & pi196;
assign w3105 = w533 & pi079;
assign w3106 = ~w533 & pi207;
assign w3107 = w533 & pi078;
assign w3108 = ~w533 & pi206;
assign w3109 = w533 & pi080;
assign w3110 = ~w533 & pi208;
assign w3111 = w533 & pi082;
assign w3112 = ~w533 & pi210;
assign w3113 = w533 & pi084;
assign w3114 = ~w533 & pi212;
assign w3115 = w533 & pi081;
assign w3116 = ~w533 & pi209;
assign w3117 = w533 & pi090;
assign w3118 = ~w533 & pi218;
assign w3119 = w533 & pi089;
assign w3120 = ~w533 & pi217;
assign w3121 = w533 & pi088;
assign w3122 = ~w533 & pi216;
assign w3123 = w533 & pi116;
assign w3124 = ~w533 & pi244;
assign w3125 = w533 & pi118;
assign w3126 = ~w533 & pi246;
assign w3127 = w533 & pi117;
assign w3128 = ~w533 & pi245;
assign w3129 = w2794 & ~w2792;
assign w3130 = w2794 & ~w2793;
assign w3131 = (~w1109 & w2795) | (~w1109 & w2792) | (w2795 & w2792);
assign w3132 = (~w1109 & w2795) | (~w1109 & w2793) | (w2795 & w2793);
assign w3133 = (~w1105 & w2796) | (~w1105 & w2792) | (w2796 & w2792);
assign w3134 = (~w1105 & w2796) | (~w1105 & w2793) | (w2796 & w2793);
assign w3135 = w2797 & ~w2792;
assign w3136 = w2797 & ~w2793;
assign w3137 = (~w1118 & w2798) | (~w1118 & w2792) | (w2798 & w2792);
assign w3138 = (~w1118 & w2798) | (~w1118 & w2793) | (w2798 & w2793);
assign w3139 = w2799 & ~w2792;
assign w3140 = w2799 & ~w2793;
assign w3141 = (~w1127 & w2800) | (~w1127 & w2792) | (w2800 & w2792);
assign w3142 = (~w1127 & w2800) | (~w1127 & w2793) | (w2800 & w2793);
assign w3143 = w2801 & ~w2792;
assign w3144 = w2801 & ~w2793;
assign w3145 = (~w1136 & w2802) | (~w1136 & w2792) | (w2802 & w2792);
assign w3146 = (~w1136 & w2802) | (~w1136 & w2793) | (w2802 & w2793);
assign w3147 = w2803 & ~w2792;
assign w3148 = w2803 & ~w2793;
assign w3149 = (~w1147 & w2804) | (~w1147 & w2792) | (w2804 & w2792);
assign w3150 = (~w1147 & w2804) | (~w1147 & w2793) | (w2804 & w2793);
assign w3151 = w2805 & ~w2792;
assign w3152 = w2805 & ~w2793;
assign w3153 = (~w1098 & w2806) | (~w1098 & w2792) | (w2806 & w2792);
assign w3154 = (~w1098 & w2806) | (~w1098 & w2793) | (w2806 & w2793);
assign w3155 = w2807 & ~w2792;
assign w3156 = w2807 & ~w2793;
assign w3157 = (~w1091 & w2808) | (~w1091 & w2792) | (w2808 & w2792);
assign w3158 = (~w1091 & w2808) | (~w1091 & w2793) | (w2808 & w2793);
assign w3159 = w2809 & ~w2792;
assign w3160 = w2809 & ~w2793;
assign w3161 = (w1156 & w2810) | (w1156 & w2792) | (w2810 & w2792);
assign w3162 = (w1156 & w2810) | (w1156 & w2793) | (w2810 & w2793);
assign w3163 = w2811 & ~w2792;
assign w3164 = w2811 & ~w2793;
assign w3165 = (~w1084 & w2812) | (~w1084 & w2792) | (w2812 & w2792);
assign w3166 = (~w1084 & w2812) | (~w1084 & w2793) | (w2812 & w2793);
assign w3167 = w2813 & ~w2792;
assign w3168 = w2813 & ~w2793;
assign w3169 = (~w1077 & w2814) | (~w1077 & w2792) | (w2814 & w2792);
assign w3170 = (~w1077 & w2814) | (~w1077 & w2793) | (w2814 & w2793);
assign w3171 = w2815 & ~w2792;
assign w3172 = w2815 & ~w2793;
assign w3173 = (~w1172 & w2816) | (~w1172 & w2792) | (w2816 & w2792);
assign w3174 = (~w1172 & w2816) | (~w1172 & w2793) | (w2816 & w2793);
assign w3175 = w2817 & ~w2792;
assign w3176 = w2817 & ~w2793;
assign w3177 = (w1185 & w2818) | (w1185 & w2792) | (w2818 & w2792);
assign w3178 = (w1185 & w2818) | (w1185 & w2793) | (w2818 & w2793);
assign w3179 = w2819 & ~w2792;
assign w3180 = w2819 & ~w2793;
assign w3181 = (~w1181 & w2820) | (~w1181 & w2792) | (w2820 & w2792);
assign w3182 = (~w1181 & w2820) | (~w1181 & w2793) | (w2820 & w2793);
assign w3183 = w2821 & ~w2792;
assign w3184 = w2821 & ~w2793;
assign w3185 = (~w1199 & w2822) | (~w1199 & w2792) | (w2822 & w2792);
assign w3186 = (~w1199 & w2822) | (~w1199 & w2793) | (w2822 & w2793);
assign w3187 = w2823 & ~w2792;
assign w3188 = w2823 & ~w2793;
assign w3189 = (~w1210 & w2824) | (~w1210 & w2792) | (w2824 & w2792);
assign w3190 = (~w1210 & w2824) | (~w1210 & w2793) | (w2824 & w2793);
assign w3191 = w2825 & ~w2792;
assign w3192 = w2825 & ~w2793;
assign w3193 = (~w1221 & w2826) | (~w1221 & w2792) | (w2826 & w2792);
assign w3194 = (~w1221 & w2826) | (~w1221 & w2793) | (w2826 & w2793);
assign w3195 = w2827 & ~w2792;
assign w3196 = w2827 & ~w2793;
assign w3197 = (~w1237 & w2828) | (~w1237 & w2792) | (w2828 & w2792);
assign w3198 = (~w1237 & w2828) | (~w1237 & w2793) | (w2828 & w2793);
assign w3199 = w2829 & ~w2792;
assign w3200 = w2829 & ~w2793;
assign w3201 = (~w1230 & w2830) | (~w1230 & w2792) | (w2830 & w2792);
assign w3202 = (~w1230 & w2830) | (~w1230 & w2793) | (w2830 & w2793);
assign w3203 = w2831 & ~w2792;
assign w3204 = w2831 & ~w2793;
assign w3205 = (~w1246 & w2832) | (~w1246 & w2792) | (w2832 & w2792);
assign w3206 = (~w1246 & w2832) | (~w1246 & w2793) | (w2832 & w2793);
assign w3207 = w2833 & ~w2792;
assign w3208 = w2833 & ~w2793;
assign w3209 = (~w1266 & w2834) | (~w1266 & w2792) | (w2834 & w2792);
assign w3210 = (~w1266 & w2834) | (~w1266 & w2793) | (w2834 & w2793);
assign w3211 = w2835 & ~w2792;
assign w3212 = w2835 & ~w2793;
assign w3213 = (~w1259 & w2836) | (~w1259 & w2792) | (w2836 & w2792);
assign w3214 = (~w1259 & w2836) | (~w1259 & w2793) | (w2836 & w2793);
assign w3215 = w2837 & ~w2792;
assign w3216 = w2837 & ~w2793;
assign w3217 = (~w1275 & w2838) | (~w1275 & w2792) | (w2838 & w2792);
assign w3218 = (~w1275 & w2838) | (~w1275 & w2793) | (w2838 & w2793);
assign w3219 = w2839 & ~w2792;
assign w3220 = w2839 & ~w2793;
assign w3221 = (~w1287 & w2840) | (~w1287 & w2792) | (w2840 & w2792);
assign w3222 = (~w1287 & w2840) | (~w1287 & w2793) | (w2840 & w2793);
assign w3223 = w2841 & ~w2792;
assign w3224 = w2841 & ~w2793;
assign w3225 = (~w1296 & w2842) | (~w1296 & w2792) | (w2842 & w2792);
assign w3226 = (~w1296 & w2842) | (~w1296 & w2793) | (w2842 & w2793);
assign w3227 = w2843 & ~w2792;
assign w3228 = w2843 & ~w2793;
assign w3229 = (~w1312 & w2844) | (~w1312 & w2792) | (w2844 & w2792);
assign w3230 = (~w1312 & w2844) | (~w1312 & w2793) | (w2844 & w2793);
assign w3231 = w2845 & ~w2792;
assign w3232 = w2845 & ~w2793;
assign w3233 = (~w1305 & w2846) | (~w1305 & w2792) | (w2846 & w2792);
assign w3234 = (~w1305 & w2846) | (~w1305 & w2793) | (w2846 & w2793);
assign w3235 = w2847 & ~w2792;
assign w3236 = w2847 & ~w2793;
assign w3237 = (~w1322 & w2848) | (~w1322 & w2792) | (w2848 & w2792);
assign w3238 = (~w1322 & w2848) | (~w1322 & w2793) | (w2848 & w2793);
assign w3239 = w2849 & ~w2792;
assign w3240 = w2849 & ~w2793;
assign w3241 = (~w1342 & w2850) | (~w1342 & w2792) | (w2850 & w2792);
assign w3242 = (~w1342 & w2850) | (~w1342 & w2793) | (w2850 & w2793);
assign w3243 = w2851 & ~w2792;
assign w3244 = w2851 & ~w2793;
assign w3245 = (~w1335 & w2852) | (~w1335 & w2792) | (w2852 & w2792);
assign w3246 = (~w1335 & w2852) | (~w1335 & w2793) | (w2852 & w2793);
assign w3247 = w2853 & ~w2792;
assign w3248 = w2853 & ~w2793;
assign w3249 = (~w1351 & w2854) | (~w1351 & w2792) | (w2854 & w2792);
assign w3250 = (~w1351 & w2854) | (~w1351 & w2793) | (w2854 & w2793);
assign w3251 = w2855 & ~w2792;
assign w3252 = w2855 & ~w2793;
assign w3253 = (~w1423 & w2856) | (~w1423 & w2792) | (w2856 & w2792);
assign w3254 = (~w1423 & w2856) | (~w1423 & w2793) | (w2856 & w2793);
assign w3255 = w2857 & ~w2792;
assign w3256 = w2857 & ~w2793;
assign w3257 = (w1413 & w2858) | (w1413 & w2792) | (w2858 & w2792);
assign w3258 = (w1413 & w2858) | (w1413 & w2793) | (w2858 & w2793);
assign w3259 = w2859 & ~w2792;
assign w3260 = w2859 & ~w2793;
assign w3261 = (~w1363 & w2860) | (~w1363 & w2792) | (w2860 & w2792);
assign w3262 = (~w1363 & w2860) | (~w1363 & w2793) | (w2860 & w2793);
assign w3263 = w2861 & ~w2792;
assign w3264 = w2861 & ~w2793;
assign w3265 = (w1367 & w2862) | (w1367 & w2792) | (w2862 & w2792);
assign w3266 = (w1367 & w2862) | (w1367 & w2793) | (w2862 & w2793);
assign w3267 = w2863 & ~w2792;
assign w3268 = w2863 & ~w2793;
assign w3269 = (~w1400 & w2864) | (~w1400 & w2792) | (w2864 & w2792);
assign w3270 = (~w1400 & w2864) | (~w1400 & w2793) | (w2864 & w2793);
assign w3271 = w2865 & ~w2792;
assign w3272 = w2865 & ~w2793;
assign w3273 = (~w1393 & w2866) | (~w1393 & w2792) | (w2866 & w2792);
assign w3274 = (~w1393 & w2866) | (~w1393 & w2793) | (w2866 & w2793);
assign w3275 = w2867 & ~w2792;
assign w3276 = w2867 & ~w2793;
assign w3277 = (~w1385 & w2868) | (~w1385 & w2792) | (w2868 & w2792);
assign w3278 = (~w1385 & w2868) | (~w1385 & w2793) | (w2868 & w2793);
assign w3279 = w2869 & ~w2792;
assign w3280 = w2869 & ~w2793;
assign w3281 = (w1375 & w2870) | (w1375 & w2792) | (w2870 & w2792);
assign w3282 = (w1375 & w2870) | (w1375 & w2793) | (w2870 & w2793);
assign w3283 = w2871 & ~w2792;
assign w3284 = w2871 & ~w2793;
assign w3285 = (~w1409 & w2872) | (~w1409 & w2792) | (w2872 & w2792);
assign w3286 = (~w1409 & w2872) | (~w1409 & w2793) | (w2872 & w2793);
assign w3287 = w2873 & ~w2792;
assign w3288 = w2873 & ~w2793;
assign w3289 = (w1511 & w2874) | (w1511 & w2792) | (w2874 & w2792);
assign w3290 = (w1511 & w2874) | (w1511 & w2793) | (w2874 & w2793);
assign w3291 = w2875 & ~w2792;
assign w3292 = w2875 & ~w2793;
assign w3293 = (~w1507 & w2876) | (~w1507 & w2792) | (w2876 & w2792);
assign w3294 = (~w1507 & w2876) | (~w1507 & w2793) | (w2876 & w2793);
assign w3295 = w2877 & ~w2792;
assign w3296 = w2877 & ~w2793;
assign w3297 = (~w1498 & w2878) | (~w1498 & w2792) | (w2878 & w2792);
assign w3298 = (~w1498 & w2878) | (~w1498 & w2793) | (w2878 & w2793);
assign w3299 = w2879 & ~w2792;
assign w3300 = w2879 & ~w2793;
assign w3301 = (~w1491 & w2880) | (~w1491 & w2792) | (w2880 & w2792);
assign w3302 = (~w1491 & w2880) | (~w1491 & w2793) | (w2880 & w2793);
assign w3303 = w2881 & ~w2792;
assign w3304 = w2881 & ~w2793;
assign w3305 = (~w1482 & w2882) | (~w1482 & w2792) | (w2882 & w2792);
assign w3306 = (~w1482 & w2882) | (~w1482 & w2793) | (w2882 & w2793);
assign w3307 = w2883 & ~w2792;
assign w3308 = w2883 & ~w2793;
assign w3309 = (~w1472 & w2884) | (~w1472 & w2792) | (w2884 & w2792);
assign w3310 = (~w1472 & w2884) | (~w1472 & w2793) | (w2884 & w2793);
assign w3311 = w2885 & ~w2792;
assign w3312 = w2885 & ~w2793;
assign w3313 = (~w1453 & w2886) | (~w1453 & w2792) | (w2886 & w2792);
assign w3314 = (~w1453 & w2886) | (~w1453 & w2793) | (w2886 & w2793);
assign w3315 = w2887 & ~w2792;
assign w3316 = w2887 & ~w2793;
assign w3317 = (~w1459 & w2888) | (~w1459 & w2792) | (w2888 & w2792);
assign w3318 = (~w1459 & w2888) | (~w1459 & w2793) | (w2888 & w2793);
assign w3319 = w2889 & ~w2792;
assign w3320 = w2889 & ~w2793;
assign w3321 = (w1653 & w2890) | (w1653 & w2792) | (w2890 & w2792);
assign w3322 = (w1653 & w2890) | (w1653 & w2793) | (w2890 & w2793);
assign w3323 = w2891 & ~w2792;
assign w3324 = w2891 & ~w2793;
assign w3325 = (~w1557 & w2892) | (~w1557 & w2792) | (w2892 & w2792);
assign w3326 = (~w1557 & w2892) | (~w1557 & w2793) | (w2892 & w2793);
assign w3327 = w2893 & ~w2792;
assign w3328 = w2893 & ~w2793;
assign w3329 = (w1561 & w2894) | (w1561 & w2792) | (w2894 & w2792);
assign w3330 = (w1561 & w2894) | (w1561 & w2793) | (w2894 & w2793);
assign w3331 = w2895 & ~w2792;
assign w3332 = w2895 & ~w2793;
assign w3333 = (~w1601 & w2896) | (~w1601 & w2792) | (w2896 & w2792);
assign w3334 = (~w1601 & w2896) | (~w1601 & w2793) | (w2896 & w2793);
assign w3335 = w2897 & ~w2792;
assign w3336 = w2897 & ~w2793;
assign w3337 = (w1591 & w2898) | (w1591 & w2792) | (w2898 & w2792);
assign w3338 = (w1591 & w2898) | (w1591 & w2793) | (w2898 & w2793);
assign w3339 = w2899 & ~w2792;
assign w3340 = w2899 & ~w2793;
assign w3341 = (~w1587 & w2900) | (~w1587 & w2792) | (w2900 & w2792);
assign w3342 = (~w1587 & w2900) | (~w1587 & w2793) | (w2900 & w2793);
assign w3343 = w2901 & ~w2792;
assign w3344 = w2901 & ~w2793;
assign w3345 = (w1638 & w2902) | (w1638 & w2792) | (w2902 & w2792);
assign w3346 = (w1638 & w2902) | (w1638 & w2793) | (w2902 & w2793);
assign w3347 = w2903 & ~w2792;
assign w3348 = w2903 & ~w2793;
assign w3349 = (w1645 & w2904) | (w1645 & w2792) | (w2904 & w2792);
assign w3350 = (w1645 & w2904) | (w1645 & w2793) | (w2904 & w2793);
assign w3351 = w2905 & ~w2792;
assign w3352 = w2905 & ~w2793;
assign w3353 = (w1549 & w2906) | (w1549 & w2792) | (w2906 & w2792);
assign w3354 = (w1549 & w2906) | (w1549 & w2793) | (w2906 & w2793);
assign w3355 = w2907 & ~w2792;
assign w3356 = w2907 & ~w2793;
assign w3357 = (~w1541 & w2908) | (~w1541 & w2792) | (w2908 & w2792);
assign w3358 = (~w1541 & w2908) | (~w1541 & w2793) | (w2908 & w2793);
assign w3359 = w2909 & ~w2792;
assign w3360 = w2909 & ~w2793;
assign w3361 = (~w1579 & w2910) | (~w1579 & w2792) | (w2910 & w2792);
assign w3362 = (~w1579 & w2910) | (~w1579 & w2793) | (w2910 & w2793);
assign w3363 = w2911 & ~w2792;
assign w3364 = w2911 & ~w2793;
assign w3365 = (~w1572 & w2912) | (~w1572 & w2792) | (w2912 & w2792);
assign w3366 = (~w1572 & w2912) | (~w1572 & w2793) | (w2912 & w2793);
assign w3367 = w2913 & ~w2792;
assign w3368 = w2913 & ~w2793;
assign w3369 = (~w1610 & w2914) | (~w1610 & w2792) | (w2914 & w2792);
assign w3370 = (~w1610 & w2914) | (~w1610 & w2793) | (w2914 & w2793);
assign w3371 = w2915 & ~w2792;
assign w3372 = w2915 & ~w2793;
assign w3373 = (~w1631 & w2916) | (~w1631 & w2792) | (w2916 & w2792);
assign w3374 = (~w1631 & w2916) | (~w1631 & w2793) | (w2916 & w2793);
assign w3375 = w2917 & ~w2792;
assign w3376 = w2917 & ~w2793;
assign w3377 = (w1621 & w2918) | (w1621 & w2792) | (w2918 & w2792);
assign w3378 = (w1621 & w2918) | (w1621 & w2793) | (w2918 & w2793);
assign w3379 = w2919 & ~w2792;
assign w3380 = w2919 & ~w2793;
assign w3381 = (~w1617 & w2920) | (~w1617 & w2792) | (w2920 & w2792);
assign w3382 = (~w1617 & w2920) | (~w1617 & w2793) | (w2920 & w2793);
assign w3383 = w2921 & ~w2792;
assign w3384 = w2921 & ~w2793;
assign w3385 = (w1719 & w2922) | (w1719 & w2792) | (w2922 & w2792);
assign w3386 = (w1719 & w2922) | (w1719 & w2793) | (w2922 & w2793);
assign w3387 = w2923 & ~w2792;
assign w3388 = w2923 & ~w2793;
assign w3389 = (~w1714 & w2924) | (~w1714 & w2792) | (w2924 & w2792);
assign w3390 = (~w1714 & w2924) | (~w1714 & w2793) | (w2924 & w2793);
assign w3391 = w2925 & ~w2792;
assign w3392 = w2925 & ~w2793;
assign w3393 = (w1703 & w2926) | (w1703 & w2792) | (w2926 & w2792);
assign w3394 = (w1703 & w2926) | (w1703 & w2793) | (w2926 & w2793);
assign w3395 = w2927 & ~w2792;
assign w3396 = w2927 & ~w2793;
assign w3397 = (~w1698 & w2928) | (~w1698 & w2792) | (w2928 & w2792);
assign w3398 = (~w1698 & w2928) | (~w1698 & w2793) | (w2928 & w2793);
assign w3399 = w2929 & ~w2792;
assign w3400 = w2929 & ~w2793;
assign w3401 = (~w1777 & w2930) | (~w1777 & w2792) | (w2930 & w2792);
assign w3402 = (~w1777 & w2930) | (~w1777 & w2793) | (w2930 & w2793);
assign w3403 = w2931 & ~w2792;
assign w3404 = w2931 & ~w2793;
assign w3405 = (~w1769 & w2932) | (~w1769 & w2792) | (w2932 & w2792);
assign w3406 = (~w1769 & w2932) | (~w1769 & w2793) | (w2932 & w2793);
assign w3407 = w2933 & ~w2792;
assign w3408 = w2933 & ~w2793;
assign w3409 = (w1759 & w2934) | (w1759 & w2792) | (w2934 & w2792);
assign w3410 = (w1759 & w2934) | (w1759 & w2793) | (w2934 & w2793);
assign w3411 = w2935 & ~w2792;
assign w3412 = w2935 & ~w2793;
assign w3413 = (~w1798 & w2936) | (~w1798 & w2792) | (w2936 & w2792);
assign w3414 = (~w1798 & w2936) | (~w1798 & w2793) | (w2936 & w2793);
assign w3415 = w2937 & ~w2792;
assign w3416 = w2937 & ~w2793;
assign w3417 = (w1788 & w2938) | (w1788 & w2792) | (w2938 & w2792);
assign w3418 = (w1788 & w2938) | (w1788 & w2793) | (w2938 & w2793);
assign w3419 = w2939 & ~w2792;
assign w3420 = w2939 & ~w2793;
assign w3421 = (~w1784 & w2940) | (~w1784 & w2792) | (w2940 & w2792);
assign w3422 = (~w1784 & w2940) | (~w1784 & w2793) | (w2940 & w2793);
assign w3423 = w2941 & ~w2792;
assign w3424 = w2941 & ~w2793;
assign w3425 = (w1747 & w2942) | (w1747 & w2792) | (w2942 & w2792);
assign w3426 = (w1747 & w2942) | (w1747 & w2793) | (w2942 & w2793);
assign w3427 = w2943 & ~w2792;
assign w3428 = w2943 & ~w2793;
assign w3429 = (~w1743 & w2944) | (~w1743 & w2792) | (w2944 & w2792);
assign w3430 = (~w1743 & w2944) | (~w1743 & w2793) | (w2944 & w2793);
assign w3431 = w2945 & ~w2792;
assign w3432 = w2945 & ~w2793;
assign w3433 = (w1840 & w2946) | (w1840 & w2792) | (w2946 & w2792);
assign w3434 = (w1840 & w2946) | (w1840 & w2793) | (w2946 & w2793);
assign w3435 = w2947 & ~w2792;
assign w3436 = w2947 & ~w2793;
assign w3437 = (~w1836 & w2948) | (~w1836 & w2792) | (w2948 & w2792);
assign w3438 = (~w1836 & w2948) | (~w1836 & w2793) | (w2948 & w2793);
assign w3439 = w2949 & ~w2792;
assign w3440 = w2949 & ~w2793;
assign w3441 = (~w1852 & w2950) | (~w1852 & w2792) | (w2950 & w2792);
assign w3442 = (~w1852 & w2950) | (~w1852 & w2793) | (w2950 & w2793);
assign w3443 = w2951 & ~w2792;
assign w3444 = w2951 & ~w2793;
assign w3445 = (~w1829 & w2952) | (~w1829 & w2792) | (w2952 & w2792);
assign w3446 = (~w1829 & w2952) | (~w1829 & w2793) | (w2952 & w2793);
assign w3447 = w2953 & ~w2792;
assign w3448 = w2953 & ~w2793;
assign w3449 = (w1866 & w2954) | (w1866 & w2792) | (w2954 & w2792);
assign w3450 = (w1866 & w2954) | (w1866 & w2793) | (w2954 & w2793);
assign w3451 = w2955 & ~w2792;
assign w3452 = w2955 & ~w2793;
assign w3453 = (~w1925 & w2956) | (~w1925 & w2792) | (w2956 & w2792);
assign w3454 = (~w1925 & w2956) | (~w1925 & w2793) | (w2956 & w2793);
assign w3455 = w2957 & ~w2792;
assign w3456 = w2957 & ~w2793;
assign w3457 = (w1899 & w2958) | (w1899 & w2792) | (w2958 & w2792);
assign w3458 = (w1899 & w2958) | (w1899 & w2793) | (w2958 & w2793);
assign w3459 = w2959 & ~w2792;
assign w3460 = w2959 & ~w2793;
assign w3461 = (~w1916 & w2960) | (~w1916 & w2792) | (w2960 & w2792);
assign w3462 = (~w1916 & w2960) | (~w1916 & w2793) | (w2960 & w2793);
assign w3463 = w2961 & ~w2792;
assign w3464 = w2961 & ~w2793;
assign w3465 = (~w1909 & w2962) | (~w1909 & w2792) | (w2962 & w2792);
assign w3466 = (~w1909 & w2962) | (~w1909 & w2793) | (w2962 & w2793);
assign w3467 = w2963 & ~w2792;
assign w3468 = w2963 & ~w2793;
assign w3469 = (~w1879 & w2964) | (~w1879 & w2792) | (w2964 & w2792);
assign w3470 = (~w1879 & w2964) | (~w1879 & w2793) | (w2964 & w2793);
assign w3471 = w2965 & ~w2792;
assign w3472 = w2965 & ~w2793;
assign w3473 = (w1890 & w2966) | (w1890 & w2792) | (w2966 & w2792);
assign w3474 = (w1890 & w2966) | (w1890 & w2793) | (w2966 & w2793);
assign w3475 = w2967 & ~w2792;
assign w3476 = w2967 & ~w2793;
assign w3477 = (~w1886 & w2968) | (~w1886 & w2792) | (w2968 & w2792);
assign w3478 = (~w1886 & w2968) | (~w1886 & w2793) | (w2968 & w2793);
assign w3479 = w2969 & ~w2792;
assign w3480 = w2969 & ~w2793;
assign w3481 = (w1959 & w2970) | (w1959 & w2792) | (w2970 & w2792);
assign w3482 = (w1959 & w2970) | (w1959 & w2793) | (w2970 & w2793);
assign w3483 = w2971 & ~w2792;
assign w3484 = w2971 & ~w2793;
assign w3485 = (~w1954 & w2972) | (~w1954 & w2792) | (w2972 & w2792);
assign w3486 = (~w1954 & w2972) | (~w1954 & w2793) | (w2972 & w2793);
assign w3487 = w2973 & ~w2792;
assign w3488 = w2973 & ~w2793;
assign w3489 = (w1943 & w2974) | (w1943 & w2792) | (w2974 & w2792);
assign w3490 = (w1943 & w2974) | (w1943 & w2793) | (w2974 & w2793);
assign w3491 = w2975 & ~w2792;
assign w3492 = w2975 & ~w2793;
assign w3493 = (~w1938 & w2976) | (~w1938 & w2792) | (w2976 & w2792);
assign w3494 = (~w1938 & w2976) | (~w1938 & w2793) | (w2976 & w2793);
assign w3495 = w2977 & ~w2792;
assign w3496 = w2977 & ~w2793;
assign w3497 = (~w2026 & w2978) | (~w2026 & w2792) | (w2978 & w2792);
assign w3498 = (~w2026 & w2978) | (~w2026 & w2793) | (w2978 & w2793);
assign w3499 = w2979 & ~w2792;
assign w3500 = w2979 & ~w2793;
assign w3501 = (~w2011 & w2980) | (~w2011 & w2792) | (w2980 & w2792);
assign w3502 = (~w2011 & w2980) | (~w2011 & w2793) | (w2980 & w2793);
assign w3503 = w2981 & ~w2792;
assign w3504 = w2981 & ~w2793;
assign w3505 = (w2015 & w2982) | (w2015 & w2792) | (w2982 & w2792);
assign w3506 = (w2015 & w2982) | (w2015 & w2793) | (w2982 & w2793);
assign w3507 = w2983 & ~w2792;
assign w3508 = w2983 & ~w2793;
assign w3509 = (~w2033 & w2984) | (~w2033 & w2792) | (w2984 & w2792);
assign w3510 = (~w2033 & w2984) | (~w2033 & w2793) | (w2984 & w2793);
assign w3511 = w2985 & ~w2792;
assign w3512 = w2985 & ~w2793;
assign w3513 = (w2044 & w2986) | (w2044 & w2792) | (w2986 & w2792);
assign w3514 = (w2044 & w2986) | (w2044 & w2793) | (w2986 & w2793);
assign w3515 = w2987 & ~w2792;
assign w3516 = w2987 & ~w2793;
assign w3517 = (~w2040 & w2988) | (~w2040 & w2792) | (w2988 & w2792);
assign w3518 = (~w2040 & w2988) | (~w2040 & w2793) | (w2988 & w2793);
assign w3519 = w2989 & ~w2792;
assign w3520 = w2989 & ~w2793;
assign w3521 = (w1996 & w2990) | (w1996 & w2792) | (w2990 & w2792);
assign w3522 = (w1996 & w2990) | (w1996 & w2793) | (w2990 & w2793);
assign w3523 = w2991 & ~w2792;
assign w3524 = w2991 & ~w2793;
assign w3525 = (~w1992 & w2992) | (~w1992 & w2792) | (w2992 & w2792);
assign w3526 = (~w1992 & w2992) | (~w1992 & w2793) | (w2992 & w2793);
assign w3527 = w2993 & ~w2792;
assign w3528 = w2993 & ~w2793;
assign w3529 = (w2089 & w2994) | (w2089 & w2792) | (w2994 & w2792);
assign w3530 = (w2089 & w2994) | (w2089 & w2793) | (w2994 & w2793);
assign w3531 = w2995 & ~w2792;
assign w3532 = w2995 & ~w2793;
assign w3533 = (~w2085 & w2996) | (~w2085 & w2792) | (w2996 & w2792);
assign w3534 = (~w2085 & w2996) | (~w2085 & w2793) | (w2996 & w2793);
assign w3535 = w2997 & ~w2792;
assign w3536 = w2997 & ~w2793;
assign w3537 = (~w2101 & w2998) | (~w2101 & w2792) | (w2998 & w2792);
assign w3538 = (~w2101 & w2998) | (~w2101 & w2793) | (w2998 & w2793);
assign w3539 = w2999 & ~w2792;
assign w3540 = w2999 & ~w2793;
assign w3541 = (~w2078 & w3000) | (~w2078 & w2792) | (w3000 & w2792);
assign w3542 = (~w2078 & w3000) | (~w2078 & w2793) | (w3000 & w2793);
assign w3543 = w3001 & ~w2792;
assign w3544 = w3001 & ~w2793;
assign w3545 = (w2115 & w3002) | (w2115 & w2792) | (w3002 & w2792);
assign w3546 = (w2115 & w3002) | (w2115 & w2793) | (w3002 & w2793);
assign w3547 = w3003 & ~w2792;
assign w3548 = w3003 & ~w2793;
assign w3549 = (~w2174 & w3004) | (~w2174 & w2792) | (w3004 & w2792);
assign w3550 = (~w2174 & w3004) | (~w2174 & w2793) | (w3004 & w2793);
assign w3551 = w3005 & ~w2792;
assign w3552 = w3005 & ~w2793;
assign w3553 = (w2148 & w3006) | (w2148 & w2792) | (w3006 & w2792);
assign w3554 = (w2148 & w3006) | (w2148 & w2793) | (w3006 & w2793);
assign w3555 = w3007 & ~w2792;
assign w3556 = w3007 & ~w2793;
assign w3557 = (~w2165 & w3008) | (~w2165 & w2792) | (w3008 & w2792);
assign w3558 = (~w2165 & w3008) | (~w2165 & w2793) | (w3008 & w2793);
assign w3559 = w3009 & ~w2792;
assign w3560 = w3009 & ~w2793;
assign w3561 = (~w2158 & w3010) | (~w2158 & w2792) | (w3010 & w2792);
assign w3562 = (~w2158 & w3010) | (~w2158 & w2793) | (w3010 & w2793);
assign w3563 = w3011 & ~w2792;
assign w3564 = w3011 & ~w2793;
assign w3565 = (~w2128 & w3012) | (~w2128 & w2792) | (w3012 & w2792);
assign w3566 = (~w2128 & w3012) | (~w2128 & w2793) | (w3012 & w2793);
assign w3567 = w3013 & ~w2792;
assign w3568 = w3013 & ~w2793;
assign w3569 = (w2139 & w3014) | (w2139 & w2792) | (w3014 & w2792);
assign w3570 = (w2139 & w3014) | (w2139 & w2793) | (w3014 & w2793);
assign w3571 = w3015 & ~w2792;
assign w3572 = w3015 & ~w2793;
assign w3573 = (~w2135 & w3016) | (~w2135 & w2792) | (w3016 & w2792);
assign w3574 = (~w2135 & w3016) | (~w2135 & w2793) | (w3016 & w2793);
assign w3575 = w3017 & ~w2792;
assign w3576 = w3017 & ~w2793;
assign w3577 = (w2208 & w3018) | (w2208 & w2792) | (w3018 & w2792);
assign w3578 = (w2208 & w3018) | (w2208 & w2793) | (w3018 & w2793);
assign w3579 = w3019 & ~w2792;
assign w3580 = w3019 & ~w2793;
assign w3581 = (~w2203 & w3020) | (~w2203 & w2792) | (w3020 & w2792);
assign w3582 = (~w2203 & w3020) | (~w2203 & w2793) | (w3020 & w2793);
assign w3583 = w3021 & ~w2792;
assign w3584 = w3021 & ~w2793;
assign w3585 = (w2192 & w3022) | (w2192 & w2792) | (w3022 & w2792);
assign w3586 = (w2192 & w3022) | (w2192 & w2793) | (w3022 & w2793);
assign w3587 = w3023 & ~w2792;
assign w3588 = w3023 & ~w2793;
assign w3589 = (~w2187 & w3024) | (~w2187 & w2792) | (w3024 & w2792);
assign w3590 = (~w2187 & w3024) | (~w2187 & w2793) | (w3024 & w2793);
assign w3591 = w3025 & ~w2792;
assign w3592 = w3025 & ~w2793;
assign w3593 = (w2267 & w3026) | (w2267 & w2792) | (w3026 & w2792);
assign w3594 = (w2267 & w3026) | (w2267 & w2793) | (w3026 & w2793);
assign w3595 = w3027 & ~w2792;
assign w3596 = w3027 & ~w2793;
assign w3597 = (~w2299 & w3028) | (~w2299 & w2792) | (w3028 & w2792);
assign w3598 = (~w2299 & w3028) | (~w2299 & w2793) | (w3028 & w2793);
assign w3599 = w3029 & ~w2792;
assign w3600 = w3029 & ~w2793;
assign w3601 = (w2289 & w3030) | (w2289 & w2792) | (w3030 & w2792);
assign w3602 = (w2289 & w3030) | (w2289 & w2793) | (w3030 & w2793);
assign w3603 = w3031 & ~w2792;
assign w3604 = w3031 & ~w2793;
assign w3605 = (~w2277 & w3032) | (~w2277 & w2792) | (w3032 & w2792);
assign w3606 = (~w2277 & w3032) | (~w2277 & w2793) | (w3032 & w2793);
assign w3607 = w3033 & ~w2792;
assign w3608 = w3033 & ~w2793;
assign w3609 = (w2281 & w3034) | (w2281 & w2792) | (w3034 & w2792);
assign w3610 = (w2281 & w3034) | (w2281 & w2793) | (w3034 & w2793);
assign w3611 = w3035 & ~w2792;
assign w3612 = w3035 & ~w2793;
assign w3613 = (~w2263 & w3036) | (~w2263 & w2792) | (w3036 & w2792);
assign w3614 = (~w2263 & w3036) | (~w2263 & w2793) | (w3036 & w2793);
assign w3615 = w3037 & ~w2792;
assign w3616 = w3037 & ~w2793;
assign w3617 = (w2248 & w3038) | (w2248 & w2792) | (w3038 & w2792);
assign w3618 = (w2248 & w3038) | (w2248 & w2793) | (w3038 & w2793);
assign w3619 = w3039 & ~w2792;
assign w3620 = w3039 & ~w2793;
assign w3621 = (~w2244 & w3040) | (~w2244 & w2792) | (w3040 & w2792);
assign w3622 = (~w2244 & w3040) | (~w2244 & w2793) | (w3040 & w2793);
assign w3623 = w3041 & ~w2792;
assign w3624 = w3041 & ~w2793;
assign w3625 = (~w2345 & w3042) | (~w2345 & w2792) | (w3042 & w2792);
assign w3626 = (~w2345 & w3042) | (~w2345 & w2793) | (w3042 & w2793);
assign w3627 = w3043 & ~w2792;
assign w3628 = w3043 & ~w2793;
assign w3629 = (~w2337 & w3044) | (~w2337 & w2792) | (w3044 & w2792);
assign w3630 = (~w2337 & w3044) | (~w2337 & w2793) | (w3044 & w2793);
assign w3631 = w3045 & ~w2792;
assign w3632 = w3045 & ~w2793;
assign w3633 = (~w2330 & w3046) | (~w2330 & w2792) | (w3046 & w2792);
assign w3634 = (~w2330 & w3046) | (~w2330 & w2793) | (w3046 & w2793);
assign w3635 = w3047 & ~w2792;
assign w3636 = w3047 & ~w2793;
assign w3637 = (w1074 & w3048) | (w1074 & w2792) | (w3048 & w2792);
assign w3638 = (w1074 & w3048) | (w1074 & w2793) | (w3048 & w2793);
assign w3639 = w3049 & ~w2792;
assign w3640 = w3049 & ~w2793;
assign w3641 = ~w1269 & w1281;
assign w3642 = ~w1328 & w1345;
assign w3643 = w3052 & w1805;
assign w3644 = (w1805 & w3052) | (w1805 & w1635) | (w3052 & w1635);
assign w3645 = ~w2112 & w2179;
assign w3646 = ~w2307 & ~w2306;
assign w3647 = (w23 & w3054) | (w23 & ~w3) | (w3054 & ~w3);
assign w3648 = (w23 & w3054) | (w23 & w3053) | (w3054 & w3053);
assign w3649 = (w564 & w3057) | (w564 & w3055) | (w3057 & w3055);
assign w3650 = (w564 & w3057) | (w564 & w3056) | (w3057 & w3056);
assign w3651 = ~w570 & w576;
assign w3652 = w533 & pi016;
assign w3653 = ~w533 & pi144;
assign w3654 = w533 & pi018;
assign w3655 = ~w533 & pi146;
assign w3656 = w533 & pi017;
assign w3657 = ~w533 & pi145;
assign w3658 = w533 & pi019;
assign w3659 = ~w533 & pi147;
assign w3660 = w533 & pi021;
assign w3661 = ~w533 & pi149;
assign w3662 = w533 & pi022;
assign w3663 = ~w533 & pi150;
assign w3664 = w533 & pi023;
assign w3665 = ~w533 & pi151;
assign w3666 = w533 & pi024;
assign w3667 = ~w533 & pi152;
assign w3668 = w533 & pi026;
assign w3669 = ~w533 & pi154;
assign w3670 = w533 & pi025;
assign w3671 = ~w533 & pi153;
assign w3672 = w531 & w3073;
assign w3673 = w533 & pi034;
assign w3674 = ~w533 & pi162;
assign w3675 = w533 & pi036;
assign w3676 = ~w533 & pi164;
assign w3677 = w533 & pi035;
assign w3678 = ~w533 & pi163;
assign w3679 = w531 & w3075;
assign w3680 = w531 & w3077;
assign w3681 = (w1430 & w3080) | (w1430 & w3071) | (w3080 & w3071);
assign w3682 = (w1430 & w3080) | (w1430 & w3070) | (w3080 & w3070);
assign w3683 = w533 & pi044;
assign w3684 = ~w533 & pi172;
assign w3685 = w533 & pi043;
assign w3686 = ~w533 & pi171;
assign w3687 = w533 & pi042;
assign w3688 = ~w533 & pi170;
assign w3689 = w533 & pi041;
assign w3690 = ~w533 & pi169;
assign w3691 = w533 & pi040;
assign w3692 = ~w533 & pi168;
assign w3693 = ~w1476 & w1527;
assign w3694 = (pi049 & w2774) | (pi049 & ~w531) | (w2774 & ~w531);
assign w3695 = (pi049 & w2774) | (pi049 & ~w4090) | (w2774 & ~w4090);
assign w3696 = ~w523 & w3082;
assign w3697 = (pi050 & w2776) | (pi050 & ~w531) | (w2776 & ~w531);
assign w3698 = (pi050 & w2776) | (pi050 & ~w4090) | (w2776 & ~w4090);
assign w3699 = ~w523 & w3087;
assign w3700 = w531 & w3089;
assign w3701 = w531 & w3091;
assign w3702 = w3092 | pi051;
assign w3703 = (pi051 & w3092) | (pi051 & ~w531) | (w3092 & ~w531);
assign w3704 = w531 & w3093;
assign w3705 = w531 & w3095;
assign w3706 = w533 & pi055;
assign w3707 = ~w533 & pi183;
assign w3708 = (pi048 & w2778) | (pi048 & ~w531) | (w2778 & ~w531);
assign w3709 = (pi048 & w2778) | (pi048 & ~w4090) | (w2778 & ~w4090);
assign w3710 = ~w523 & w3098;
assign w3711 = w533 & pi066;
assign w3712 = ~w533 & pi194;
assign w3713 = w533 & pi065;
assign w3714 = ~w533 & pi193;
assign w3715 = w533 & pi064;
assign w3716 = ~w533 & pi192;
assign w3717 = w531 & w3100;
assign w3718 = w531 & w3102;
assign w3719 = w531 & w3104;
assign w3720 = w533 & pi073;
assign w3721 = ~w533 & pi201;
assign w3722 = w533 & pi072;
assign w3723 = ~w533 & pi200;
assign w3724 = w533 & pi071;
assign w3725 = ~w533 & pi199;
assign w3726 = w531 & w3106;
assign w3727 = w533 & pi077;
assign w3728 = ~w533 & pi205;
assign w3729 = w533 & pi076;
assign w3730 = ~w533 & pi204;
assign w3731 = w531 & w3108;
assign w3732 = w3109 | pi080;
assign w3733 = (pi080 & w3109) | (pi080 & ~w531) | (w3109 & ~w531);
assign w3734 = w531 & w3110;
assign w3735 = w533 & pi085;
assign w3736 = ~w533 & pi213;
assign w3737 = w533 & pi087;
assign w3738 = ~w533 & pi215;
assign w3739 = w3111 | pi082;
assign w3740 = (pi082 & w3111) | (pi082 & ~w531) | (w3111 & ~w531);
assign w3741 = w531 & w3112;
assign w3742 = w3113 | pi084;
assign w3743 = (pi084 & w3113) | (pi084 & ~w531) | (w3113 & ~w531);
assign w3744 = w531 & w3114;
assign w3745 = w533 & pi083;
assign w3746 = ~w533 & pi211;
assign w3747 = w3115 | pi081;
assign w3748 = (pi081 & w3115) | (pi081 & ~w531) | (w3115 & ~w531);
assign w3749 = w531 & w3116;
assign w3750 = w533 & pi091;
assign w3751 = ~w533 & pi219;
assign w3752 = w3117 | pi090;
assign w3753 = (pi090 & w3117) | (pi090 & ~w531) | (w3117 & ~w531);
assign w3754 = w531 & w3118;
assign w3755 = w3119 | pi089;
assign w3756 = (pi089 & w3119) | (pi089 & ~w531) | (w3119 & ~w531);
assign w3757 = w531 & w3120;
assign w3758 = w3121 | pi088;
assign w3759 = (pi088 & w3121) | (pi088 & ~w531) | (w3121 & ~w531);
assign w3760 = w531 & w3122;
assign w3761 = w533 & pi093;
assign w3762 = ~w533 & pi221;
assign w3763 = w533 & pi094;
assign w3764 = ~w533 & pi222;
assign w3765 = w533 & pi092;
assign w3766 = ~w533 & pi220;
assign w3767 = w533 & pi114;
assign w3768 = ~w533 & pi242;
assign w3769 = w533 & pi113;
assign w3770 = ~w533 & pi241;
assign w3771 = w533 & pi112;
assign w3772 = ~w533 & pi240;
assign w3773 = w531 & w3124;
assign w3774 = w533 & pi119;
assign w3775 = ~w533 & pi247;
assign w3776 = w531 & w3126;
assign w3777 = w531 & w3128;
assign w3778 = (w2793 & w2792) | (w2793 & w2788) | (w2792 & w2788);
assign w3779 = (w2793 & w2792) | (w2793 & w2787) | (w2792 & w2787);
assign w3780 = w1427 & ~w1357;
assign w3781 = ~w27 & w32;
assign w3782 = w583 & ~w576;
assign w3783 = w583 & ~w3651;
assign w3784 = ~w592 & w595;
assign w3785 = w533 & pi015;
assign w3786 = ~w533 & pi143;
assign w3787 = w3652 | pi016;
assign w3788 = (pi016 & w3652) | (pi016 & ~w531) | (w3652 & ~w531);
assign w3789 = w531 & w3653;
assign w3790 = w3654 | pi018;
assign w3791 = (pi018 & w3654) | (pi018 & ~w531) | (w3654 & ~w531);
assign w3792 = w531 & w3655;
assign w3793 = w3656 | pi017;
assign w3794 = (pi017 & w3656) | (pi017 & ~w531) | (w3656 & ~w531);
assign w3795 = w531 & w3657;
assign w3796 = w3658 | pi019;
assign w3797 = (pi019 & w3658) | (pi019 & ~w531) | (w3658 & ~w531);
assign w3798 = w531 & w3659;
assign w3799 = w3660 | pi021;
assign w3800 = (pi021 & w3660) | (pi021 & ~w531) | (w3660 & ~w531);
assign w3801 = w531 & w3661;
assign w3802 = w533 & pi020;
assign w3803 = ~w533 & pi148;
assign w3804 = w3662 | pi022;
assign w3805 = (pi022 & w3662) | (pi022 & ~w531) | (w3662 & ~w531);
assign w3806 = w531 & w3663;
assign w3807 = w3664 | pi023;
assign w3808 = (pi023 & w3664) | (pi023 & ~w531) | (w3664 & ~w531);
assign w3809 = w531 & w3665;
assign w3810 = w3666 | pi024;
assign w3811 = (pi024 & w3666) | (pi024 & ~w531) | (w3666 & ~w531);
assign w3812 = w531 & w3667;
assign w3813 = w3668 | pi026;
assign w3814 = (pi026 & w3668) | (pi026 & ~w531) | (w3668 & ~w531);
assign w3815 = w531 & w3669;
assign w3816 = w3670 | pi025;
assign w3817 = (pi025 & w3670) | (pi025 & ~w531) | (w3670 & ~w531);
assign w3818 = w531 & w3671;
assign w3819 = w533 & pi027;
assign w3820 = ~w533 & pi155;
assign w3821 = w533 & pi029;
assign w3822 = ~w533 & pi157;
assign w3823 = (pi033 & w3072) | (pi033 & ~w531) | (w3072 & ~w531);
assign w3824 = (pi033 & w3072) | (pi033 & ~w4090) | (w3072 & ~w4090);
assign w3825 = ~w523 & w3672;
assign w3826 = w531 & w3674;
assign w3827 = w531 & w3676;
assign w3828 = w531 & w3678;
assign w3829 = (pi032 & w3074) | (pi032 & ~w531) | (w3074 & ~w531);
assign w3830 = (pi032 & w3074) | (pi032 & ~w4090) | (w3074 & ~w4090);
assign w3831 = ~w523 & w3679;
assign w3832 = (pi031 & w3076) | (pi031 & ~w531) | (w3076 & ~w531);
assign w3833 = (pi031 & w3076) | (pi031 & ~w4090) | (w3076 & ~w4090);
assign w3834 = ~w523 & w3680;
assign w3835 = ~w1530 & w1664;
assign w3836 = ~w1690 & w1581;
assign w3837 = w533 & pi067;
assign w3838 = ~w533 & pi195;
assign w3839 = w531 & w3712;
assign w3840 = w531 & w3714;
assign w3841 = w531 & w3716;
assign w3842 = w1736 & w1729;
assign w3843 = ~w533 & pi203;
assign w3844 = ~w1739 & ~w1743;
assign w3845 = w533 & pi074;
assign w3846 = ~w533 & pi202;
assign w3847 = (pi070 & w3099) | (pi070 & ~w531) | (w3099 & ~w531);
assign w3848 = (pi070 & w3099) | (pi070 & ~w4090) | (w3099 & ~w4090);
assign w3849 = ~w523 & w3717;
assign w3850 = (pi069 & w3101) | (pi069 & ~w531) | (w3101 & ~w531);
assign w3851 = (pi069 & w3101) | (pi069 & ~w4090) | (w3101 & ~w4090);
assign w3852 = ~w523 & w3718;
assign w3853 = (pi068 & w3103) | (pi068 & ~w531) | (w3103 & ~w531);
assign w3854 = (pi068 & w3103) | (pi068 & ~w4090) | (w3103 & ~w4090);
assign w3855 = ~w523 & w3719;
assign w3856 = w3720 | pi073;
assign w3857 = (pi073 & w3720) | (pi073 & ~w531) | (w3720 & ~w531);
assign w3858 = w531 & w3721;
assign w3859 = w3722 | pi072;
assign w3860 = (pi072 & w3722) | (pi072 & ~w531) | (w3722 & ~w531);
assign w3861 = w531 & w3723;
assign w3862 = w3724 | pi071;
assign w3863 = (pi071 & w3724) | (pi071 & ~w531) | (w3724 & ~w531);
assign w3864 = w531 & w3725;
assign w3865 = (pi079 & w3105) | (pi079 & ~w531) | (w3105 & ~w531);
assign w3866 = (pi079 & w3105) | (pi079 & ~w4090) | (w3105 & ~w4090);
assign w3867 = ~w523 & w3726;
assign w3868 = w3727 | pi077;
assign w3869 = (pi077 & w3727) | (pi077 & ~w531) | (w3727 & ~w531);
assign w3870 = w531 & w3728;
assign w3871 = w3729 | pi076;
assign w3872 = (pi076 & w3729) | (pi076 & ~w531) | (w3729 & ~w531);
assign w3873 = w531 & w3730;
assign w3874 = (pi078 & w3107) | (pi078 & ~w531) | (w3107 & ~w531);
assign w3875 = (pi078 & w3107) | (pi078 & ~w4090) | (w3107 & ~w4090);
assign w3876 = ~w523 & w3731;
assign w3877 = ~w523 & w3734;
assign w3878 = w3735 | pi085;
assign w3879 = (pi085 & w3735) | (pi085 & ~w531) | (w3735 & ~w531);
assign w3880 = w531 & w3736;
assign w3881 = w3737 | pi087;
assign w3882 = (pi087 & w3737) | (pi087 & ~w531) | (w3737 & ~w531);
assign w3883 = w531 & w3738;
assign w3884 = w533 & pi086;
assign w3885 = ~w533 & pi214;
assign w3886 = ~w523 & w3741;
assign w3887 = ~w523 & w3744;
assign w3888 = w3745 | pi083;
assign w3889 = (pi083 & w3745) | (pi083 & ~w531) | (w3745 & ~w531);
assign w3890 = w531 & w3746;
assign w3891 = ~w523 & w3749;
assign w3892 = w3750 | pi091;
assign w3893 = (pi091 & w3750) | (pi091 & ~w531) | (w3750 & ~w531);
assign w3894 = w531 & w3751;
assign w3895 = ~w523 & w3754;
assign w3896 = ~w523 & w3757;
assign w3897 = ~w523 & w3760;
assign w3898 = w533 & pi099;
assign w3899 = ~w533 & pi227;
assign w3900 = w533 & pi098;
assign w3901 = ~w533 & pi226;
assign w3902 = w531 & w3762;
assign w3903 = w531 & w3764;
assign w3904 = w531 & w3766;
assign w3905 = w533 & pi095;
assign w3906 = ~w533 & pi223;
assign w3907 = w533 & pi097;
assign w3908 = ~w533 & pi225;
assign w3909 = w533 & pi103;
assign w3910 = ~w533 & pi231;
assign w3911 = w533 & pi102;
assign w3912 = ~w533 & pi230;
assign w3913 = w533 & pi115;
assign w3914 = ~w533 & pi243;
assign w3915 = w531 & w3768;
assign w3916 = w531 & w3770;
assign w3917 = w531 & w3772;
assign w3918 = (pi116 & w3123) | (pi116 & ~w531) | (w3123 & ~w531);
assign w3919 = (pi116 & w3123) | (pi116 & ~w4090) | (w3123 & ~w4090);
assign w3920 = ~w523 & w3773;
assign w3921 = w3774 | pi119;
assign w3922 = (pi119 & w3774) | (pi119 & ~w531) | (w3774 & ~w531);
assign w3923 = w531 & w3775;
assign w3924 = w533 & pi120;
assign w3925 = ~w533 & pi248;
assign w3926 = (pi118 & w3125) | (pi118 & ~w531) | (w3125 & ~w531);
assign w3927 = (pi118 & w3125) | (pi118 & ~w4090) | (w3125 & ~w4090);
assign w3928 = ~w523 & w3776;
assign w3929 = (pi117 & w3127) | (pi117 & ~w531) | (w3127 & ~w531);
assign w3930 = (pi117 & w3127) | (pi117 & ~w4090) | (w3127 & ~w4090);
assign w3931 = ~w523 & w3777;
assign w3932 = w38 & ~w32;
assign w3933 = w38 & ~w3781;
assign w3934 = ~w539 & ~w595;
assign w3935 = ~w539 & ~w3784;
assign w3936 = ~w599 & w605;
assign w3937 = (pi033 & w3072) | (pi033 & w4207) | (w3072 & w4207);
assign w3938 = (w3824 & w3823) | (w3824 & ~w515) | (w3823 & ~w515);
assign w3939 = w3825 & w3672;
assign w3940 = (w3672 & w3825) | (w3672 & w515) | (w3825 & w515);
assign w3941 = (pi034 & w3673) | (pi034 & ~w531) | (w3673 & ~w531);
assign w3942 = (pi034 & w3673) | (pi034 & ~w4090) | (w3673 & ~w4090);
assign w3943 = ~w523 & w3826;
assign w3944 = w533 & pi037;
assign w3945 = ~w533 & pi165;
assign w3946 = (pi036 & w3675) | (pi036 & ~w531) | (w3675 & ~w531);
assign w3947 = (pi036 & w3675) | (pi036 & ~w4090) | (w3675 & ~w4090);
assign w3948 = ~w523 & w3827;
assign w3949 = (pi035 & w3677) | (pi035 & ~w531) | (w3677 & ~w531);
assign w3950 = (pi035 & w3677) | (pi035 & ~w4090) | (w3677 & ~w4090);
assign w3951 = ~w523 & w3828;
assign w3952 = (pi032 & w3074) | (pi032 & w4207) | (w3074 & w4207);
assign w3953 = (w3830 & w3829) | (w3830 & ~w515) | (w3829 & ~w515);
assign w3954 = w3831 & w3679;
assign w3955 = (w3679 & w3831) | (w3679 & w515) | (w3831 & w515);
assign w3956 = (pi031 & w3076) | (pi031 & w4207) | (w3076 & w4207);
assign w3957 = (w3833 & w3832) | (w3833 & ~w515) | (w3832 & ~w515);
assign w3958 = w3834 & w3680;
assign w3959 = (w3680 & w3834) | (w3680 & w515) | (w3834 & w515);
assign w3960 = w533 & pi047;
assign w3961 = ~w533 & pi175;
assign w3962 = w533 & pi046;
assign w3963 = ~w533 & pi174;
assign w3964 = w533 & pi045;
assign w3965 = ~w533 & pi173;
assign w3966 = w531 & w3684;
assign w3967 = w531 & w3686;
assign w3968 = w531 & w3688;
assign w3969 = w531 & w3690;
assign w3970 = w531 & w3692;
assign w3971 = w533 & pi057;
assign w3972 = ~w533 & pi185;
assign w3973 = w533 & pi059;
assign w3974 = ~w533 & pi187;
assign w3975 = w533 & pi058;
assign w3976 = ~w533 & pi186;
assign w3977 = (w57 & w51) | (w57 & w3998) | (w51 & w3998);
assign w3978 = (w57 & ~w54) | (w57 & w3989) | (~w54 & w3989);
assign w3979 = w612 & ~w605;
assign w3980 = w612 & ~w3936;
assign w3981 = w620 & ~w3979;
assign w3982 = w620 & ~w3980;
assign w3983 = w1 & w60;
assign w3984 = w66 & ~w60;
assign w3985 = w66 & ~w3983;
assign w3986 = w623 & ~w3982;
assign w3987 = w623 & ~w3981;
assign w3988 = w538 & w627;
assign w3989 = w46 & w57;
assign w3990 = (w3985 & w3984) | (w3985 & ~w3978) | (w3984 & ~w3978);
assign w3991 = w66 & w4208;
assign w3992 = ~w80 & w4008;
assign w3993 = w615 & ~w607;
assign w3994 = w633 & ~w627;
assign w3995 = w633 & ~w3988;
assign w3996 = w638 & ~w3995;
assign w3997 = w638 & ~w3994;
assign w3998 = ~w53 & w57;
assign w3999 = w0 & w87;
assign w4000 = w644 & ~w3997;
assign w4001 = w644 & ~w3996;
assign w4002 = ~w682 & ~w679;
assign w4003 = ~pi416 & pi288;
assign w4004 = ~w705 & w657;
assign w4005 = ~w727 & w770;
assign w4006 = ~w733 & w772;
assign w4007 = ~w799 & w819;
assign w4008 = w81 & ~w74;
assign w4009 = (w80 & w4022) | (w80 & w4036) | (w4022 & w4036);
assign w4010 = ~w93 & w98;
assign w4011 = w664 & ~w4001;
assign w4012 = w664 & ~w4000;
assign w4013 = w678 & w691;
assign w4014 = w698 & ~w645;
assign w4015 = w730 & ~w772;
assign w4016 = w730 & ~w4006;
assign w4017 = w759 & w724;
assign w4018 = w853 & ~w819;
assign w4019 = w853 & ~w4007;
assign w4020 = ~w81 & w84;
assign w4021 = w3999 & w87;
assign w4022 = (w87 & w3999) | (w87 & w84) | (w3999 & w84);
assign w4023 = (~w3992 & w4037) | (~w3992 & w4038) | (w4037 & w4038);
assign w4024 = ~w143 & ~w140;
assign w4025 = ~pi160 & pi032;
assign w4026 = ~w167 & w118;
assign w4027 = ~w191 & w235;
assign w4028 = ~w197 & w237;
assign w4029 = w675 & ~w691;
assign w4030 = w675 & ~w4013;
assign w4031 = w707 & w645;
assign w4032 = w707 & ~w4014;
assign w4033 = ~w711 & w749;
assign w4034 = ~w775 & w741;
assign w4035 = ~w873 & w905;
assign w4036 = (w87 & w3999) | (w87 & w4020) | (w3999 & w4020);
assign w4037 = (w98 & w4010) | (w98 & w4022) | (w4010 & w4022);
assign w4038 = (w98 & w4010) | (w98 & w4021) | (w4010 & w4021);
assign w4039 = ~w262 & w282;
assign w4040 = w104 & ~w4023;
assign w4041 = w104 & w4209;
assign w4042 = w139 & w152;
assign w4043 = w160 & ~w106;
assign w4044 = w155 & w172;
assign w4045 = w315 & ~w282;
assign w4046 = (~w241 & w4045) | (~w241 & w4055) | (w4045 & w4055);
assign w4047 = w650 & ~w4032;
assign w4048 = w650 & ~w4031;
assign w4049 = w693 & w709;
assign w4050 = ~w720 & ~w758;
assign w4051 = w925 & ~w905;
assign w4052 = w925 & ~w4035;
assign w4053 = w959 & ~w4051;
assign w4054 = w959 & ~w4052;
assign w4055 = w315 & ~w4039;
assign w4056 = w77 & ~w69;
assign w4057 = w334 & ~w4045;
assign w4058 = w334 & ~w4046;
assign w4059 = ~w368 & w388;
assign w4060 = ~w864 & ~w861;
assign w4061 = w895 & ~w881;
assign w4062 = w978 & ~w4053;
assign w4063 = w978 & ~w4054;
assign w4064 = ~w1012 & w1032;
assign w4065 = w224 & w188;
assign w4066 = ~w245 & ~w242;
assign w4067 = ~w278 & w297;
assign w4068 = (w388 & w4059) | (w388 & w4057) | (w4059 & w4057);
assign w4069 = (w388 & w4059) | (w388 & w4058) | (w4059 & w4058);
assign w4070 = ~w423 & w442;
assign w4071 = ~w887 & ~w884;
assign w4072 = w1049 & ~w1032;
assign w4073 = w1049 & ~w4064;
assign w4074 = w1056 & ~w4073;
assign w4075 = w1056 & ~w4072;
assign w4076 = ~w240 & w205;
assign w4077 = w312 & ~w283;
assign w4078 = w476 & ~w442;
assign w4079 = w496 & ~w4078;
assign w4080 = (w496 & w4070) | (w496 & w4197) | (w4070 & w4197);
assign w4081 = ~w1041 & w1019;
assign w4082 = w1063 & ~w4075;
assign w4083 = w1063 & ~w4074;
assign w4084 = w1073 & pi289;
assign w4085 = ~w1073 & pi417;
assign w4086 = w1073 & pi288;
assign w4087 = ~w1073 & pi416;
assign w4088 = w515 & ~w4079;
assign w4089 = w515 & ~w4080;
assign w4090 = ~w523 & w531;
assign w4091 = ~w969 & ~w966;
assign w4092 = w1002 & ~w987;
assign w4093 = ~w1044 & w1027;
assign w4094 = ~w1073 & w4083;
assign w4095 = ~w1073 & w4082;
assign w4096 = (w3937 & w3938) | (w3937 & w4079) | (w3938 & w4079);
assign w4097 = (w3937 & w3938) | (w3937 & w4080) | (w3938 & w4080);
assign w4098 = (w3939 & w3940) | (w3939 & ~w4079) | (w3940 & ~w4079);
assign w4099 = (w3939 & w3940) | (w3939 & ~w4080) | (w3940 & ~w4080);
assign w4100 = (pi289 & w4084) | (pi289 & ~w4083) | (w4084 & ~w4083);
assign w4101 = (pi289 & w4084) | (pi289 & ~w4082) | (w4084 & ~w4082);
assign w4102 = w4085 & w4083;
assign w4103 = w4085 & w4082;
assign w4104 = (pi288 & w4086) | (pi288 & ~w4083) | (w4086 & ~w4083);
assign w4105 = (pi288 & w4086) | (pi288 & ~w4082) | (w4086 & ~w4082);
assign w4106 = w4087 & w4083;
assign w4107 = w4087 & w4082;
assign w4108 = (w3952 & w3953) | (w3952 & w4079) | (w3953 & w4079);
assign w4109 = (w3952 & w3953) | (w3952 & w4080) | (w3953 & w4080);
assign w4110 = (w3954 & w3955) | (w3954 & ~w4079) | (w3955 & ~w4079);
assign w4111 = (w3954 & w3955) | (w3954 & ~w4080) | (w3955 & ~w4080);
assign w4112 = (w3956 & w3957) | (w3956 & w4079) | (w3957 & w4079);
assign w4113 = (w3956 & w3957) | (w3956 & w4080) | (w3957 & w4080);
assign w4114 = (w3958 & w3959) | (w3958 & ~w4079) | (w3959 & ~w4079);
assign w4115 = (w3958 & w3959) | (w3958 & ~w4080) | (w3959 & ~w4080);
assign w4116 = (pi287 & w3078) | (pi287 & ~w4083) | (w3078 & ~w4083);
assign w4117 = (pi287 & w3078) | (pi287 & ~w4082) | (w3078 & ~w4082);
assign w4118 = w3079 & w4083;
assign w4119 = w3079 & w4082;
assign w4120 = ~w1387 & ~w1448;
assign w4121 = (pi044 & w3683) | (pi044 & ~w531) | (w3683 & ~w531);
assign w4122 = (pi044 & w3683) | (pi044 & ~w4090) | (w3683 & ~w4090);
assign w4123 = ~w523 & w3966;
assign w4124 = (pi043 & w3685) | (pi043 & ~w531) | (w3685 & ~w531);
assign w4125 = (pi043 & w3685) | (pi043 & ~w4090) | (w3685 & ~w4090);
assign w4126 = ~w523 & w3967;
assign w4127 = (pi042 & w3687) | (pi042 & ~w531) | (w3687 & ~w531);
assign w4128 = (pi042 & w3687) | (pi042 & ~w4090) | (w3687 & ~w4090);
assign w4129 = ~w523 & w3968;
assign w4130 = (pi041 & w3689) | (pi041 & ~w531) | (w3689 & ~w531);
assign w4131 = (pi041 & w3689) | (pi041 & ~w4090) | (w3689 & ~w4090);
assign w4132 = ~w523 & w3969;
assign w4133 = (pi040 & w3691) | (pi040 & ~w531) | (w3691 & ~w531);
assign w4134 = (pi040 & w3691) | (pi040 & ~w4090) | (w3691 & ~w4090);
assign w4135 = ~w523 & w3970;
assign w4136 = (pi305 & w3083) | (pi305 & ~w4083) | (w3083 & ~w4083);
assign w4137 = (pi305 & w3083) | (pi305 & ~w4082) | (w3083 & ~w4082);
assign w4138 = (pi306 & w3085) | (pi306 & ~w4083) | (w3085 & ~w4083);
assign w4139 = (pi306 & w3085) | (pi306 & ~w4082) | (w3085 & ~w4082);
assign w4140 = (pi053 & w3088) | (pi053 & ~w531) | (w3088 & ~w531);
assign w4141 = (pi053 & w3088) | (pi053 & ~w4090) | (w3088 & ~w4090);
assign w4142 = ~w523 & w3700;
assign w4143 = (pi052 & w3090) | (pi052 & ~w531) | (w3090 & ~w531);
assign w4144 = (pi052 & w3090) | (pi052 & ~w4090) | (w3090 & ~w4090);
assign w4145 = ~w523 & w3701;
assign w4146 = ~w523 & w3704;
assign w4147 = (pi054 & w3094) | (pi054 & ~w531) | (w3094 & ~w531);
assign w4148 = (pi054 & w3094) | (pi054 & ~w4090) | (w3094 & ~w4090);
assign w4149 = ~w523 & w3705;
assign w4150 = (pi304 & w3096) | (pi304 & ~w4083) | (w3096 & ~w4083);
assign w4151 = (pi304 & w3096) | (pi304 & ~w4082) | (w3096 & ~w4082);
assign w4152 = ~w1671 & ~w1650;
assign w4153 = ~w1671 & ~w2780;
assign w4154 = (pi066 & w3711) | (pi066 & ~w531) | (w3711 & ~w531);
assign w4155 = (pi066 & w3711) | (pi066 & ~w4090) | (w3711 & ~w4090);
assign w4156 = ~w523 & w3839;
assign w4157 = (pi065 & w3713) | (pi065 & ~w531) | (w3713 & ~w531);
assign w4158 = (pi065 & w3713) | (pi065 & ~w4090) | (w3713 & ~w4090);
assign w4159 = ~w523 & w3840;
assign w4160 = (pi064 & w3715) | (pi064 & ~w531) | (w3715 & ~w531);
assign w4161 = (pi064 & w3715) | (pi064 & ~w4090) | (w3715 & ~w4090);
assign w4162 = ~w523 & w3841;
assign w4163 = ~w523 & w3858;
assign w4164 = ~w523 & w3861;
assign w4165 = ~w523 & w3864;
assign w4166 = ~w1822 & w1752;
assign w4167 = ~w523 & w3870;
assign w4168 = ~w523 & w3873;
assign w4169 = ~w523 & w3880;
assign w4170 = ~w523 & w3883;
assign w4171 = ~w523 & w3890;
assign w4172 = ~w523 & w3894;
assign w4173 = ~w1948 & ~w1939;
assign w4174 = ~w1982 & w1896;
assign w4175 = (pi093 & w3761) | (pi093 & ~w531) | (w3761 & ~w531);
assign w4176 = (pi093 & w3761) | (pi093 & ~w4090) | (w3761 & ~w4090);
assign w4177 = ~w523 & w3902;
assign w4178 = (pi094 & w3763) | (pi094 & ~w531) | (w3763 & ~w531);
assign w4179 = (pi094 & w3763) | (pi094 & ~w4090) | (w3763 & ~w4090);
assign w4180 = ~w523 & w3903;
assign w4181 = (pi092 & w3765) | (pi092 & ~w531) | (w3765 & ~w531);
assign w4182 = (pi092 & w3765) | (pi092 & ~w4090) | (w3765 & ~w4090);
assign w4183 = ~w523 & w3904;
assign w4184 = (pi114 & w3767) | (pi114 & ~w531) | (w3767 & ~w531);
assign w4185 = (pi114 & w3767) | (pi114 & ~w4090) | (w3767 & ~w4090);
assign w4186 = ~w523 & w3915;
assign w4187 = (pi113 & w3769) | (pi113 & ~w531) | (w3769 & ~w531);
assign w4188 = (pi113 & w3769) | (pi113 & ~w4090) | (w3769 & ~w4090);
assign w4189 = ~w523 & w3916;
assign w4190 = (pi112 & w3771) | (pi112 & ~w531) | (w3771 & ~w531);
assign w4191 = (pi112 & w3771) | (pi112 & ~w4090) | (w3771 & ~w4090);
assign w4192 = ~w523 & w3917;
assign w4193 = ~w523 & w3923;
assign w4194 = ~w2286 & ~w2310;
assign w4195 = w2054 & ~w1986;
assign w4196 = w2054 & ~w1863;
assign w4197 = ~w476 & w496;
assign w4198 = w523 & ~w4089;
assign w4199 = w523 & ~w4088;
assign w4200 = w533 & pi000;
assign w4201 = ~w533 & pi128;
assign w4202 = (w106 & ~w4043) | (w106 & ~w168) | (~w4043 & ~w168);
assign w4203 = (~w237 & ~w4028) | (~w237 & ~w236) | (~w4028 & ~w236);
assign w4204 = (~w4075 & ~w4074) | (~w4075 & ~w979) | (~w4074 & ~w979);
assign w4205 = (w4083 & w4082) | (w4083 & ~w979) | (w4082 & ~w979);
assign w4206 = w523 & ~w516;
assign w4207 = ~w531 | ~w4090;
assign w4208 = (~w3983 & ~w60) | (~w3983 & ~w3977) | (~w60 & ~w3977);
assign w4209 = (~w98 & ~w4010) | (~w98 & ~w4009) | (~w4010 & ~w4009);
assign one = 1;
assign po000 = ~w2360;// level 29
assign po001 = ~w2363;// level 29
assign po002 = ~w2366;// level 29
assign po003 = ~w2369;// level 29
assign po004 = ~w2372;// level 29
assign po005 = ~w2375;// level 29
assign po006 = ~w2378;// level 29
assign po007 = ~w2381;// level 29
assign po008 = w2384;// level 29
assign po009 = ~w2387;// level 29
assign po010 = ~w2390;// level 29
assign po011 = ~w2393;// level 29
assign po012 = w2396;// level 29
assign po013 = ~w2399;// level 29
assign po014 = ~w2402;// level 29
assign po015 = ~w2405;// level 29
assign po016 = ~w2408;// level 29
assign po017 = ~w2411;// level 29
assign po018 = ~w2414;// level 29
assign po019 = ~w2417;// level 29
assign po020 = ~w2420;// level 29
assign po021 = ~w2423;// level 29
assign po022 = ~w2426;// level 29
assign po023 = ~w2429;// level 29
assign po024 = ~w2432;// level 29
assign po025 = ~w2435;// level 29
assign po026 = ~w2438;// level 29
assign po027 = ~w2441;// level 29
assign po028 = ~w2444;// level 29
assign po029 = ~w2447;// level 29
assign po030 = ~w2450;// level 29
assign po031 = ~w2453;// level 29
assign po032 = w2456;// level 29
assign po033 = ~w2459;// level 29
assign po034 = w2462;// level 29
assign po035 = ~w2465;// level 29
assign po036 = ~w2468;// level 29
assign po037 = ~w2471;// level 29
assign po038 = w2474;// level 29
assign po039 = ~w2477;// level 29
assign po040 = w2480;// level 29
assign po041 = ~w2483;// level 29
assign po042 = ~w2486;// level 29
assign po043 = ~w2489;// level 29
assign po044 = ~w2492;// level 29
assign po045 = ~w2495;// level 29
assign po046 = ~w2498;// level 29
assign po047 = ~w2501;// level 29
assign po048 = w2504;// level 29
assign po049 = ~w2507;// level 29
assign po050 = w2510;// level 29
assign po051 = ~w2513;// level 29
assign po052 = w2516;// level 29
assign po053 = ~w2519;// level 29
assign po054 = w2522;// level 29
assign po055 = w2525;// level 29
assign po056 = w2528;// level 29
assign po057 = ~w2531;// level 29
assign po058 = ~w2534;// level 29
assign po059 = ~w2537;// level 29
assign po060 = ~w2540;// level 29
assign po061 = ~w2543;// level 29
assign po062 = w2546;// level 29
assign po063 = ~w2549;// level 29
assign po064 = w2552;// level 29
assign po065 = ~w2555;// level 29
assign po066 = w2558;// level 29
assign po067 = ~w2561;// level 29
assign po068 = ~w2564;// level 29
assign po069 = ~w2567;// level 29
assign po070 = w2570;// level 29
assign po071 = ~w2573;// level 29
assign po072 = w2576;// level 29
assign po073 = ~w2579;// level 29
assign po074 = w2582;// level 29
assign po075 = ~w2585;// level 29
assign po076 = w2588;// level 29
assign po077 = ~w2591;// level 29
assign po078 = ~w2594;// level 29
assign po079 = ~w2597;// level 29
assign po080 = w2600;// level 29
assign po081 = ~w2603;// level 29
assign po082 = w2606;// level 29
assign po083 = ~w2609;// level 29
assign po084 = ~w2612;// level 29
assign po085 = ~w2615;// level 29
assign po086 = w2618;// level 29
assign po087 = ~w2621;// level 29
assign po088 = w2624;// level 29
assign po089 = ~w2627;// level 29
assign po090 = w2630;// level 29
assign po091 = ~w2633;// level 29
assign po092 = ~w2636;// level 29
assign po093 = ~w2639;// level 29
assign po094 = w2642;// level 29
assign po095 = ~w2645;// level 29
assign po096 = w2648;// level 29
assign po097 = ~w2651;// level 29
assign po098 = w2654;// level 29
assign po099 = ~w2657;// level 29
assign po100 = w2660;// level 29
assign po101 = ~w2663;// level 29
assign po102 = ~w2666;// level 29
assign po103 = ~w2669;// level 29
assign po104 = w2672;// level 29
assign po105 = ~w2675;// level 29
assign po106 = w2678;// level 29
assign po107 = ~w2681;// level 29
assign po108 = ~w2684;// level 29
assign po109 = ~w2687;// level 29
assign po110 = w2690;// level 29
assign po111 = ~w2693;// level 29
assign po112 = w2696;// level 29
assign po113 = ~w2699;// level 29
assign po114 = w2702;// level 29
assign po115 = ~w2705;// level 29
assign po116 = w2708;// level 29
assign po117 = ~w2711;// level 29
assign po118 = w2714;// level 29
assign po119 = ~w2717;// level 29
assign po120 = w2720;// level 29
assign po121 = ~w2723;// level 29
assign po122 = w2726;// level 29
assign po123 = ~w2729;// level 29
assign po124 = ~w2732;// level 29
assign po125 = ~w2735;// level 29
assign po126 = ~w2738;// level 29
assign po127 = w2739;// level 17
assign po128 = ~w2742;// level 29
assign po129 = ~w2357;// level 29
endmodule
