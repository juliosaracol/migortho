module systemcdes ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278, pi279,
    pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288, pi289,
    pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298, pi299,
    pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308, pi309,
    pi310, pi311, pi312, pi313,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287, pi288,
    pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296, pi297, pi298,
    pi299, pi300, pi301, pi302, pi303, pi304, pi305, pi306, pi307, pi308,
    pi309, pi310, pi311, pi312, pi313;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257;
  wire n574, n575, n576, n577, n578, n579, n580, n581, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n639, n640, n641, n642, n643, n644, n645, n646,
    n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n689, n690, n691, n692, n693, n694, n695, n696,
    n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
    n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n739, n740, n741, n742, n743, n744, n745, n746,
    n747, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n829, n830, n831, n832, n833,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n846, n847,
    n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
    n933, n934, n935, n936, n937, n938, n939, n940, n942, n943, n944, n945,
    n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
    n983, n984, n985, n986, n987, n989, n990, n991, n992, n993, n994, n995,
    n996, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
    n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1083, n1084, n1085, n1086, n1087, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1109, n1110,
    n1111, n1112, n1113, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1166, n1167, n1168, n1169, n1170, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
    n1214, n1216, n1217, n1218, n1219, n1220, n1222, n1223, n1224, n1225,
    n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1374, n1375,
    n1376, n1377, n1378, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
    n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
    n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
    n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688, n1690, n1691, n1692, n1693,
    n1694, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
    n1727, n1728, n1729, n1730, n1731, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1773, n1774, n1775, n1776, n1777, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
    n1793, n1794, n1795, n1796, n1797, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
    n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
    n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
    n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
    n1896, n1897, n1898, n1899, n1901, n1902, n1903, n1904, n1905, n1906,
    n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
    n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
    n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
    n2052, n2053, n2054, n2055, n2057, n2058, n2059, n2060, n2061, n2063,
    n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2077, n2078, n2079, n2080, n2081, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116,
    n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
    n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2197, n2198, n2199, n2200,
    n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
    n2222, n2223, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
    n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
    n2336, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2363, n2364, n2365, n2366, n2367, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2383, n2384, n2385, n2386, n2387, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
    n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
    n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
    n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2623, n2624, n2625, n2626, n2627, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
    n2652, n2653, n2654, n2655, n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
    n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2694,
    n2695, n2696, n2697, n2698, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
    n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
    n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
    n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3033, n3034, n3035, n3036, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
    n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
    n3206, n3207, n3208, n3209, n3210, n3211, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
    n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3255, n3256, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
    n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
    n3329, n3330, n3331, n3332, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
    n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
    n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3468, n3469, n3470, n3471, n3472, n3473,
    n3474, n3475, n3476, n3477, n3479, n3480, n3481, n3482, n3483, n3484,
    n3485, n3486, n3487, n3488, n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3545, n3546, n3547, n3548, n3549, n3550,
    n3551, n3553, n3554, n3555, n3556, n3558, n3559, n3560, n3561, n3563,
    n3564, n3565, n3566, n3568, n3569, n3571;
  assign n574 = ~pi066 & ~pi068;
  assign n575 = ~pi069 & ~pi081;
  assign n576 = n574 & n575;
  assign n577 = ~pi020 & ~pi192;
  assign n578 = pi192 & ~pi227;
  assign n579 = ~n577 & ~n578;
  assign n580 = n576 & ~n579;
  assign n581 = ~pi020 & ~n576;
  assign po223 = ~n580 & ~n581;
  assign n583 = pi066 & pi081;
  assign n584 = pi068 & n583;
  assign n585 = pi069 & n584;
  assign n586 = pi069 & ~pi081;
  assign n587 = n574 & n586;
  assign n588 = ~pi069 & pi081;
  assign n589 = n574 & n588;
  assign n590 = ~n576 & ~n589;
  assign n591 = ~n587 & n590;
  assign n592 = ~n585 & n591;
  assign n593 = ~pi047 & ~pi192;
  assign n594 = pi192 & ~pi303;
  assign n595 = ~n593 & ~n594;
  assign n596 = n576 & ~n595;
  assign n597 = ~pi047 & ~n576;
  assign n598 = ~n596 & ~n597;
  assign n599 = n592 & n598;
  assign n600 = pi035 & ~n576;
  assign n601 = pi035 & ~pi192;
  assign n602 = pi192 & pi296;
  assign n603 = ~n601 & ~n602;
  assign n604 = n576 & ~n603;
  assign n605 = ~n600 & ~n604;
  assign n606 = ~n592 & ~n605;
  assign n607 = ~n599 & ~n606;
  assign n608 = ~pi193 & ~n607;
  assign n609 = ~n587 & ~n589;
  assign n610 = ~n585 & n609;
  assign n611 = ~n576 & n610;
  assign n612 = pi077 & ~pi192;
  assign n613 = pi192 & pi302;
  assign n614 = ~n612 & ~n613;
  assign n615 = n576 & ~n614;
  assign n616 = pi077 & ~n576;
  assign n617 = ~n615 & ~n616;
  assign n618 = n611 & ~n617;
  assign n619 = ~n585 & ~n589;
  assign n620 = ~n587 & n619;
  assign n621 = pi058 & ~pi192;
  assign n622 = pi192 & pi309;
  assign n623 = ~n621 & ~n622;
  assign n624 = n576 & ~n623;
  assign n625 = pi058 & ~n576;
  assign n626 = ~n624 & ~n625;
  assign n627 = ~n620 & ~n626;
  assign n628 = ~n618 & ~n627;
  assign n629 = pi040 & ~n576;
  assign n630 = pi040 & ~pi192;
  assign n631 = pi192 & pi289;
  assign n632 = ~n630 & ~n631;
  assign n633 = n576 & ~n632;
  assign n634 = ~n629 & ~n633;
  assign n635 = n576 & ~n634;
  assign n636 = n628 & ~n635;
  assign n637 = pi193 & ~n636;
  assign po108 = n608 | n637;
  assign n639 = po223 & po108;
  assign n640 = ~po223 & ~po108;
  assign n641 = ~n639 & ~n640;
  assign n642 = pi192 & pi203;
  assign n643 = pi026 & ~pi192;
  assign n644 = ~n642 & ~n643;
  assign n645 = n576 & ~n644;
  assign n646 = pi026 & ~n576;
  assign po225 = n645 | n646;
  assign n648 = pi076 & ~n576;
  assign n649 = pi076 & ~pi192;
  assign n650 = pi192 & pi287;
  assign n651 = ~n649 & ~n650;
  assign n652 = n576 & ~n651;
  assign n653 = ~n648 & ~n652;
  assign n654 = n592 & ~n653;
  assign n655 = pi091 & ~n576;
  assign n656 = pi091 & ~pi192;
  assign n657 = pi192 & pi280;
  assign n658 = ~n656 & ~n657;
  assign n659 = n576 & ~n658;
  assign n660 = ~n655 & ~n659;
  assign n661 = ~n592 & ~n660;
  assign n662 = ~n654 & ~n661;
  assign n663 = ~pi193 & ~n662;
  assign n664 = pi041 & ~n576;
  assign n665 = pi192 & pi266;
  assign n666 = pi041 & ~pi192;
  assign n667 = ~n665 & ~n666;
  assign n668 = n576 & ~n667;
  assign n669 = ~n664 & ~n668;
  assign n670 = ~n620 & ~n669;
  assign n671 = pi090 & ~n576;
  assign n672 = pi090 & ~pi192;
  assign n673 = pi192 & pi273;
  assign n674 = ~n672 & ~n673;
  assign n675 = n576 & ~n674;
  assign n676 = ~n671 & ~n675;
  assign n677 = n576 & ~n676;
  assign n678 = ~n670 & ~n677;
  assign n679 = pi074 & ~pi192;
  assign n680 = pi192 & pi259;
  assign n681 = ~n679 & ~n680;
  assign n682 = n576 & n681;
  assign n683 = ~pi074 & ~n576;
  assign n684 = ~n682 & ~n683;
  assign n685 = n611 & n684;
  assign n686 = n678 & ~n685;
  assign n687 = pi193 & ~n686;
  assign po158 = n663 | n687;
  assign n689 = po225 & ~po158;
  assign n690 = ~po225 & po158;
  assign n691 = ~n689 & ~n690;
  assign n692 = pi007 & ~pi192;
  assign n693 = pi192 & pi253;
  assign n694 = ~n692 & ~n693;
  assign n695 = n576 & ~n694;
  assign n696 = pi007 & ~n576;
  assign po210 = n695 | n696;
  assign n698 = pi078 & ~pi192;
  assign n699 = pi192 & pi294;
  assign n700 = ~n698 & ~n699;
  assign n701 = n576 & ~n700;
  assign n702 = pi078 & ~n576;
  assign n703 = ~n701 & ~n702;
  assign n704 = n611 & ~n703;
  assign n705 = pi039 & ~n576;
  assign n706 = pi039 & ~pi192;
  assign n707 = pi192 & pi301;
  assign n708 = ~n706 & ~n707;
  assign n709 = n576 & ~n708;
  assign n710 = ~n705 & ~n709;
  assign n711 = ~n620 & ~n710;
  assign n712 = pi080 & ~pi192;
  assign n713 = pi192 & pi308;
  assign n714 = ~n712 & ~n713;
  assign n715 = n576 & ~n714;
  assign n716 = pi080 & ~n576;
  assign n717 = ~n715 & ~n716;
  assign n718 = n576 & ~n717;
  assign n719 = ~n711 & ~n718;
  assign n720 = ~n704 & n719;
  assign n721 = pi193 & ~n720;
  assign n722 = pi059 & ~pi192;
  assign n723 = pi192 & pi260;
  assign n724 = ~n722 & ~n723;
  assign n725 = n576 & ~n724;
  assign n726 = pi059 & ~n576;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n592 & ~n727;
  assign n729 = pi083 & ~n576;
  assign n730 = pi083 & ~pi192;
  assign n731 = pi192 & pi267;
  assign n732 = ~n730 & ~n731;
  assign n733 = n576 & ~n732;
  assign n734 = ~n729 & ~n733;
  assign n735 = n592 & ~n734;
  assign n736 = ~n728 & ~n735;
  assign n737 = ~pi193 & ~n736;
  assign po148 = n721 | n737;
  assign n739 = ~po210 & ~po148;
  assign n740 = po210 & po148;
  assign n741 = ~n739 & ~n740;
  assign n742 = n691 & ~n741;
  assign n743 = pi192 & pi219;
  assign n744 = pi021 & ~pi192;
  assign n745 = ~n743 & ~n744;
  assign n746 = n576 & n745;
  assign n747 = ~pi021 & ~n576;
  assign po218 = ~n746 & ~n747;
  assign n749 = pi045 & ~n576;
  assign n750 = pi045 & ~pi192;
  assign n751 = pi192 & pi279;
  assign n752 = ~n750 & ~n751;
  assign n753 = n576 & ~n752;
  assign n754 = ~n749 & ~n753;
  assign n755 = n611 & ~n754;
  assign n756 = pi065 & ~n576;
  assign n757 = pi065 & ~pi192;
  assign n758 = pi192 & pi293;
  assign n759 = ~n757 & ~n758;
  assign n760 = n576 & ~n759;
  assign n761 = ~n756 & ~n760;
  assign n762 = n576 & ~n761;
  assign n763 = pi192 & ~pi286;
  assign n764 = ~pi048 & ~pi192;
  assign n765 = ~n763 & ~n764;
  assign n766 = n576 & ~n765;
  assign n767 = ~pi048 & ~n576;
  assign n768 = ~n766 & ~n767;
  assign n769 = ~n620 & n768;
  assign n770 = ~n762 & ~n769;
  assign n771 = ~n755 & n770;
  assign n772 = pi193 & ~n771;
  assign n773 = pi037 & ~n576;
  assign n774 = pi037 & ~pi192;
  assign n775 = pi192 & pi300;
  assign n776 = ~n774 & ~n775;
  assign n777 = n576 & ~n776;
  assign n778 = ~n773 & ~n777;
  assign n779 = ~n592 & ~n778;
  assign n780 = pi064 & ~n576;
  assign n781 = pi064 & ~pi192;
  assign n782 = pi192 & pi307;
  assign n783 = ~n781 & ~n782;
  assign n784 = n576 & ~n783;
  assign n785 = ~n780 & ~n784;
  assign n786 = n592 & ~n785;
  assign n787 = ~n779 & ~n786;
  assign n788 = ~pi193 & ~n787;
  assign po133 = n772 | n788;
  assign n790 = po218 & ~po133;
  assign n791 = ~po218 & po133;
  assign n792 = ~n790 & ~n791;
  assign n793 = pi192 & pi281;
  assign n794 = pi042 & ~pi192;
  assign n795 = ~n793 & ~n794;
  assign n796 = n576 & ~n795;
  assign n797 = pi042 & ~n576;
  assign n798 = ~n796 & ~n797;
  assign n799 = ~n620 & ~n798;
  assign n800 = pi092 & ~n576;
  assign n801 = pi092 & ~pi192;
  assign n802 = pi192 & pi288;
  assign n803 = ~n801 & ~n802;
  assign n804 = n576 & ~n803;
  assign n805 = ~n800 & ~n804;
  assign n806 = n576 & ~n805;
  assign n807 = ~n576 & n620;
  assign n808 = pi054 & ~pi192;
  assign n809 = pi192 & pi274;
  assign n810 = ~n808 & ~n809;
  assign n811 = n576 & ~n810;
  assign n812 = pi054 & ~n576;
  assign n813 = ~n811 & ~n812;
  assign n814 = n807 & ~n813;
  assign n815 = ~n806 & ~n814;
  assign n816 = ~n799 & n815;
  assign n817 = pi193 & ~n816;
  assign n818 = pi072 & ~pi192;
  assign n819 = pi192 & pi295;
  assign n820 = ~n818 & ~n819;
  assign n821 = n576 & ~n820;
  assign n822 = pi072 & ~n576;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~n592 & ~n823;
  assign n825 = n592 & ~n617;
  assign n826 = ~n824 & ~n825;
  assign n827 = ~pi193 & ~n826;
  assign po160 = n817 | n827;
  assign n829 = pi192 & ~pi195;
  assign n830 = ~pi017 & ~pi192;
  assign n831 = ~n829 & ~n830;
  assign n832 = n576 & ~n831;
  assign n833 = ~pi017 & ~n576;
  assign po220 = ~n832 & ~n833;
  assign n835 = po160 & ~po220;
  assign n836 = ~po160 & po220;
  assign n837 = ~n835 & ~n836;
  assign n838 = ~n792 & n837;
  assign n839 = n742 & n838;
  assign n840 = pi192 & pi211;
  assign n841 = pi029 & ~pi192;
  assign n842 = ~n840 & ~n841;
  assign n843 = n576 & n842;
  assign n844 = ~pi029 & ~n576;
  assign po212 = ~n843 & ~n844;
  assign n846 = pi061 & ~n576;
  assign n847 = pi061 & ~pi192;
  assign n848 = pi192 & pi310;
  assign n849 = ~n847 & ~n848;
  assign n850 = n576 & ~n849;
  assign n851 = ~n846 & ~n850;
  assign n852 = n576 & ~n851;
  assign n853 = n598 & ~n620;
  assign n854 = ~n605 & n611;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~n852 & n855;
  assign n857 = pi193 & ~n856;
  assign n858 = pi192 & pi258;
  assign n859 = pi053 & ~pi192;
  assign n860 = ~n858 & ~n859;
  assign n861 = n576 & ~n860;
  assign n862 = pi053 & ~n576;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~n592 & ~n863;
  assign n865 = pi075 & ~n576;
  assign n866 = pi192 & pi265;
  assign n867 = pi075 & ~pi192;
  assign n868 = ~n866 & ~n867;
  assign n869 = n576 & ~n868;
  assign n870 = ~n865 & ~n869;
  assign n871 = n592 & ~n870;
  assign n872 = ~n864 & ~n871;
  assign n873 = ~pi193 & ~n872;
  assign po129 = n857 | n873;
  assign n875 = po212 & ~po129;
  assign n876 = ~po212 & po129;
  assign n877 = ~n875 & ~n876;
  assign n878 = n741 & ~n877;
  assign n879 = ~n691 & n878;
  assign n880 = n742 & ~n877;
  assign n881 = ~n879 & ~n880;
  assign n882 = ~n792 & ~n881;
  assign n883 = n741 & n837;
  assign n884 = ~n691 & n883;
  assign n885 = ~n792 & n884;
  assign n886 = n741 & ~n837;
  assign n887 = n691 & n886;
  assign n888 = n877 & n887;
  assign n889 = ~n885 & ~n888;
  assign n890 = ~n741 & ~n837;
  assign n891 = ~n691 & n890;
  assign n892 = ~n883 & ~n891;
  assign n893 = ~n877 & ~n892;
  assign n894 = ~n741 & n837;
  assign n895 = ~n691 & n894;
  assign n896 = n877 & n895;
  assign n897 = ~n893 & ~n896;
  assign n898 = ~n887 & n897;
  assign n899 = n792 & ~n898;
  assign n900 = n889 & ~n899;
  assign n901 = ~n882 & n900;
  assign n902 = ~n839 & n901;
  assign n903 = ~n641 & ~n902;
  assign n904 = n877 & n891;
  assign n905 = ~n792 & n904;
  assign n906 = n742 & n837;
  assign n907 = ~n877 & n906;
  assign n908 = n691 & n890;
  assign n909 = n877 & n908;
  assign n910 = n792 & n909;
  assign n911 = ~n907 & ~n910;
  assign n912 = ~n905 & n911;
  assign n913 = n641 & ~n792;
  assign n914 = ~n877 & n887;
  assign n915 = ~n877 & n894;
  assign n916 = ~n891 & ~n915;
  assign n917 = ~n914 & n916;
  assign n918 = n913 & ~n917;
  assign n919 = n912 & ~n918;
  assign n920 = ~n877 & n884;
  assign n921 = n691 & n883;
  assign n922 = ~n691 & ~n837;
  assign n923 = ~n890 & ~n922;
  assign n924 = ~n921 & n923;
  assign n925 = n877 & ~n924;
  assign n926 = ~n691 & n886;
  assign n927 = n792 & n926;
  assign n928 = ~n925 & ~n927;
  assign n929 = n641 & ~n928;
  assign n930 = ~n920 & ~n929;
  assign n931 = n919 & n930;
  assign n932 = ~n903 & n931;
  assign n933 = ~pi139 & ~pi192;
  assign n934 = pi192 & pi236;
  assign n935 = ~n933 & ~n934;
  assign n936 = n576 & n935;
  assign n937 = pi139 & ~n576;
  assign n938 = ~n936 & ~n937;
  assign n939 = ~n932 & ~n938;
  assign n940 = n932 & n938;
  assign po068 = n939 | n940;
  assign n942 = ~pi070 & ~pi192;
  assign n943 = pi192 & ~pi304;
  assign n944 = ~n942 & ~n943;
  assign n945 = n576 & ~n944;
  assign n946 = ~pi070 & ~n576;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~n620 & n947;
  assign n949 = pi032 & ~n576;
  assign n950 = pi192 & pi297;
  assign n951 = pi032 & ~pi192;
  assign n952 = ~n950 & ~n951;
  assign n953 = n576 & ~n952;
  assign n954 = ~n949 & ~n953;
  assign n955 = n611 & ~n954;
  assign n956 = pi067 & ~n576;
  assign n957 = pi067 & ~pi192;
  assign n958 = pi192 & pi311;
  assign n959 = ~n957 & ~n958;
  assign n960 = n576 & ~n959;
  assign n961 = ~n956 & ~n960;
  assign n962 = n576 & ~n961;
  assign n963 = ~n955 & ~n962;
  assign n964 = ~n948 & n963;
  assign n965 = pi193 & ~n964;
  assign n966 = pi038 & ~n576;
  assign n967 = pi038 & ~pi192;
  assign n968 = pi192 & pi261;
  assign n969 = ~n967 & ~n968;
  assign n970 = n576 & ~n969;
  assign n971 = ~n966 & ~n970;
  assign n972 = ~n592 & ~n971;
  assign n973 = pi052 & ~n576;
  assign n974 = pi192 & pi268;
  assign n975 = pi052 & ~pi192;
  assign n976 = ~n974 & ~n975;
  assign n977 = n576 & ~n976;
  assign n978 = ~n973 & ~n977;
  assign n979 = n592 & ~n978;
  assign n980 = ~n972 & ~n979;
  assign n981 = ~pi193 & ~n980;
  assign po135 = n965 | n981;
  assign n983 = pi002 & ~n576;
  assign n984 = pi192 & pi217;
  assign n985 = pi002 & ~pi192;
  assign n986 = ~n984 & ~n985;
  assign n987 = n576 & ~n986;
  assign po215 = n983 | n987;
  assign n989 = po135 & po215;
  assign n990 = ~po135 & ~po215;
  assign n991 = ~n989 & ~n990;
  assign n992 = pi192 & pi209;
  assign n993 = pi019 & ~pi192;
  assign n994 = ~n992 & ~n993;
  assign n995 = n576 & n994;
  assign n996 = ~pi019 & ~n576;
  assign po219 = ~n995 & ~n996;
  assign n998 = pi088 & ~pi192;
  assign n999 = pi192 & pi277;
  assign n1000 = ~n998 & ~n999;
  assign n1001 = n576 & ~n1000;
  assign n1002 = pi088 & ~n576;
  assign n1003 = ~n1001 & ~n1002;
  assign n1004 = n576 & ~n1003;
  assign n1005 = pi033 & ~n576;
  assign n1006 = pi033 & ~pi192;
  assign n1007 = pi192 & pi263;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = n576 & ~n1008;
  assign n1010 = ~n1005 & ~n1009;
  assign n1011 = n611 & ~n1010;
  assign n1012 = pi036 & ~n576;
  assign n1013 = pi036 & ~pi192;
  assign n1014 = pi192 & pi270;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = n576 & ~n1015;
  assign n1017 = ~n1012 & ~n1016;
  assign n1018 = ~n620 & ~n1017;
  assign n1019 = ~n1011 & ~n1018;
  assign n1020 = ~n1004 & n1019;
  assign n1021 = pi193 & ~n1020;
  assign n1022 = pi073 & ~n576;
  assign n1023 = pi073 & ~pi192;
  assign n1024 = pi192 & pi284;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = n576 & ~n1025;
  assign n1027 = ~n1022 & ~n1026;
  assign n1028 = ~n807 & ~n1027;
  assign n1029 = pi044 & ~n576;
  assign n1030 = pi044 & ~pi192;
  assign n1031 = pi192 & pi291;
  assign n1032 = ~n1030 & ~n1031;
  assign n1033 = n576 & ~n1032;
  assign n1034 = ~n1029 & ~n1033;
  assign n1035 = n592 & ~n1034;
  assign n1036 = ~n1028 & ~n1035;
  assign n1037 = ~pi193 & ~n1036;
  assign po156 = n1021 | n1037;
  assign n1039 = ~po219 & ~po156;
  assign n1040 = po219 & po156;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = pi192 & pi269;
  assign n1043 = pi034 & ~pi192;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = n576 & ~n1044;
  assign n1046 = pi034 & ~n576;
  assign n1047 = ~n1045 & ~n1046;
  assign n1048 = ~n592 & ~n1047;
  assign n1049 = pi055 & ~pi192;
  assign n1050 = pi192 & pi276;
  assign n1051 = ~n1049 & ~n1050;
  assign n1052 = n576 & ~n1051;
  assign n1053 = pi055 & ~n576;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = n592 & ~n1054;
  assign n1056 = ~n1048 & ~n1055;
  assign n1057 = ~pi193 & ~n1056;
  assign n1058 = pi057 & ~n576;
  assign n1059 = pi057 & ~pi192;
  assign n1060 = pi192 & pi305;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = n576 & ~n1061;
  assign n1063 = ~n1058 & ~n1062;
  assign n1064 = n611 & ~n1063;
  assign n1065 = pi089 & ~pi192;
  assign n1066 = pi192 & pi262;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = n576 & ~n1067;
  assign n1069 = pi089 & ~n576;
  assign n1070 = ~n1068 & ~n1069;
  assign n1071 = n576 & ~n1070;
  assign n1072 = pi079 & ~n576;
  assign n1073 = pi192 & pi312;
  assign n1074 = pi079 & ~pi192;
  assign n1075 = ~n1073 & ~n1074;
  assign n1076 = n576 & ~n1075;
  assign n1077 = ~n1072 & ~n1076;
  assign n1078 = ~n620 & ~n1077;
  assign n1079 = ~n1071 & ~n1078;
  assign n1080 = ~n1064 & n1079;
  assign n1081 = pi193 & ~n1080;
  assign po157 = n1057 | n1081;
  assign n1083 = pi023 & ~n576;
  assign n1084 = pi023 & ~pi192;
  assign n1085 = pi192 & pi201;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = n576 & ~n1086;
  assign po199 = n1083 | n1087;
  assign n1089 = ~po157 & po199;
  assign n1090 = po157 & ~po199;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = pi192 & pi298;
  assign n1093 = pi085 & ~pi192;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = n576 & n1094;
  assign n1096 = ~pi085 & ~n576;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = n576 & n1097;
  assign n1099 = ~n620 & ~n1034;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = n611 & ~n1027;
  assign n1102 = n1100 & ~n1101;
  assign n1103 = pi193 & ~n1102;
  assign n1104 = n592 & ~n1077;
  assign n1105 = ~n592 & ~n1063;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~pi193 & ~n1106;
  assign po153 = n1103 | n1107;
  assign n1109 = pi192 & pi251;
  assign n1110 = pi003 & ~pi192;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = n576 & n1111;
  assign n1113 = ~pi003 & ~n576;
  assign po217 = ~n1112 & ~n1113;
  assign n1115 = po153 & ~po217;
  assign n1116 = ~n1107 & po217;
  assign n1117 = ~n1103 & n1116;
  assign n1118 = ~n1115 & ~n1117;
  assign n1119 = ~n1091 & n1118;
  assign n1120 = ~n1041 & n1119;
  assign n1121 = n1091 & n1118;
  assign n1122 = n1041 & n1121;
  assign n1123 = ~n1120 & ~n1122;
  assign n1124 = ~n991 & ~n1123;
  assign n1125 = pi046 & ~n576;
  assign n1126 = pi046 & ~pi192;
  assign n1127 = pi192 & pi264;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = n576 & ~n1128;
  assign n1130 = ~n1125 & ~n1129;
  assign n1131 = n576 & ~n1130;
  assign n1132 = pi084 & ~n576;
  assign n1133 = pi192 & pi282;
  assign n1134 = pi084 & ~pi192;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = n576 & ~n1135;
  assign n1137 = ~n1132 & ~n1136;
  assign n1138 = ~n620 & ~n1137;
  assign n1139 = pi051 & ~n576;
  assign n1140 = pi192 & pi275;
  assign n1141 = pi051 & ~pi192;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = n576 & ~n1142;
  assign n1144 = ~n1139 & ~n1143;
  assign n1145 = n611 & ~n1144;
  assign n1146 = ~n1138 & ~n1145;
  assign n1147 = ~n1131 & n1146;
  assign n1148 = pi193 & ~n1147;
  assign n1149 = pi086 & ~pi192;
  assign n1150 = pi192 & pi278;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = n576 & ~n1151;
  assign n1153 = pi086 & ~n576;
  assign n1154 = ~n1152 & ~n1153;
  assign n1155 = n592 & ~n1154;
  assign n1156 = pi043 & ~n576;
  assign n1157 = pi192 & pi271;
  assign n1158 = pi043 & ~pi192;
  assign n1159 = ~n1157 & ~n1158;
  assign n1160 = n576 & ~n1159;
  assign n1161 = ~n1156 & ~n1160;
  assign n1162 = ~n592 & ~n1161;
  assign n1163 = ~n1155 & ~n1162;
  assign n1164 = ~pi193 & ~n1163;
  assign po114 = n1148 | n1164;
  assign n1166 = pi028 & ~n576;
  assign n1167 = pi028 & ~pi192;
  assign n1168 = pi192 & pi225;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = n576 & ~n1169;
  assign po194 = n1166 | n1170;
  assign n1172 = po114 & ~po194;
  assign n1173 = ~po114 & po194;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = ~n1091 & ~n1118;
  assign n1176 = ~n991 & n1175;
  assign n1177 = n1041 & n1176;
  assign n1178 = n1174 & n1177;
  assign n1179 = ~n1124 & ~n1178;
  assign n1180 = n991 & ~n1174;
  assign n1181 = pi062 & ~n576;
  assign n1182 = pi062 & ~pi192;
  assign n1183 = pi192 & pi285;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = n576 & ~n1184;
  assign n1186 = ~n1181 & ~n1185;
  assign n1187 = ~n620 & ~n1186;
  assign n1188 = pi049 & ~n576;
  assign n1189 = pi049 & ~pi192;
  assign n1190 = pi192 & pi292;
  assign n1191 = ~n1189 & ~n1190;
  assign n1192 = n576 & ~n1191;
  assign n1193 = ~n1188 & ~n1192;
  assign n1194 = n576 & ~n1193;
  assign n1195 = n611 & ~n1154;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = ~n1187 & n1196;
  assign n1198 = pi193 & ~n1197;
  assign n1199 = pi192 & pi299;
  assign n1200 = pi063 & ~pi192;
  assign n1201 = ~n1199 & ~n1200;
  assign n1202 = n576 & ~n1201;
  assign n1203 = pi063 & ~n576;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~n592 & ~n1204;
  assign n1206 = pi087 & ~n576;
  assign n1207 = pi192 & pi306;
  assign n1208 = pi087 & ~pi192;
  assign n1209 = ~n1207 & ~n1208;
  assign n1210 = n576 & ~n1209;
  assign n1211 = ~n1206 & ~n1210;
  assign n1212 = n592 & ~n1211;
  assign n1213 = ~n1205 & ~n1212;
  assign n1214 = ~pi193 & ~n1213;
  assign po117 = n1198 | n1214;
  assign n1216 = ~pi030 & ~pi192;
  assign n1217 = pi192 & ~pi233;
  assign n1218 = ~n1216 & ~n1217;
  assign n1219 = n576 & ~n1218;
  assign n1220 = ~pi030 & ~n576;
  assign po224 = ~n1219 & ~n1220;
  assign n1222 = ~po117 & po224;
  assign n1223 = po117 & ~po224;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = n1041 & n1119;
  assign n1226 = n1224 & n1225;
  assign n1227 = n1180 & n1226;
  assign n1228 = ~n1041 & n1175;
  assign n1229 = n1180 & n1228;
  assign n1230 = n1091 & ~n1118;
  assign n1231 = ~n1041 & n1174;
  assign n1232 = n1230 & n1231;
  assign n1233 = ~n991 & n1232;
  assign n1234 = n991 & n1041;
  assign n1235 = ~n1091 & n1234;
  assign n1236 = ~n1041 & n1118;
  assign n1237 = n1091 & n1236;
  assign n1238 = n991 & n1237;
  assign n1239 = ~n1235 & ~n1238;
  assign n1240 = n1174 & ~n1239;
  assign n1241 = n991 & n1230;
  assign n1242 = ~n1174 & n1241;
  assign n1243 = n991 & ~n1041;
  assign n1244 = ~n1118 & n1243;
  assign n1245 = ~n1091 & n1244;
  assign n1246 = ~n1242 & ~n1245;
  assign n1247 = ~n1240 & n1246;
  assign n1248 = ~n1233 & n1247;
  assign n1249 = ~n1041 & ~n1091;
  assign n1250 = ~n991 & n1121;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = ~n1174 & ~n1251;
  assign n1253 = n1248 & ~n1252;
  assign n1254 = ~n1224 & ~n1253;
  assign n1255 = n1041 & n1230;
  assign n1256 = ~n1174 & n1224;
  assign n1257 = n1255 & n1256;
  assign n1258 = n1174 & n1241;
  assign n1259 = ~n1177 & ~n1258;
  assign n1260 = ~n1122 & ~n1176;
  assign n1261 = ~n1120 & n1260;
  assign n1262 = ~n1250 & n1261;
  assign n1263 = n1174 & ~n1262;
  assign n1264 = n1259 & ~n1263;
  assign n1265 = n1224 & ~n1264;
  assign n1266 = ~n1257 & ~n1265;
  assign n1267 = ~n1254 & n1266;
  assign n1268 = ~n1229 & n1267;
  assign n1269 = ~n1227 & n1268;
  assign n1270 = n1179 & n1269;
  assign n1271 = ~pi145 & ~pi192;
  assign n1272 = pi192 & pi244;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = n576 & n1273;
  assign n1275 = pi145 & ~n576;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = ~n1270 & ~n1276;
  assign n1278 = n1269 & n1276;
  assign n1279 = n1179 & n1278;
  assign po069 = n1277 | n1279;
  assign n1281 = pi192 & pi229;
  assign n1282 = pi024 & ~pi192;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = n576 & n1283;
  assign n1285 = ~pi024 & ~n576;
  assign po208 = ~n1284 & ~n1285;
  assign n1287 = n592 & ~n863;
  assign n1288 = ~n592 & ~n851;
  assign n1289 = ~n1287 & ~n1288;
  assign n1290 = ~pi193 & ~n1289;
  assign n1291 = n611 & ~n634;
  assign n1292 = ~n605 & ~n620;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n576 & n598;
  assign n1295 = n1293 & ~n1294;
  assign n1296 = pi193 & ~n1295;
  assign po115 = n1290 | n1296;
  assign n1298 = po208 & ~po115;
  assign n1299 = ~po208 & po115;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = pi031 & ~n576;
  assign n1302 = pi192 & pi213;
  assign n1303 = pi031 & ~pi192;
  assign n1304 = ~n1302 & ~n1303;
  assign n1305 = n576 & ~n1304;
  assign po221 = n1301 | n1305;
  assign n1307 = n576 & n684;
  assign n1308 = ~n620 & ~n785;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = n611 & ~n778;
  assign n1311 = n1309 & ~n1310;
  assign n1312 = pi193 & ~n1311;
  assign n1313 = n592 & ~n676;
  assign n1314 = ~n592 & ~n669;
  assign n1315 = ~n1313 & ~n1314;
  assign n1316 = ~pi193 & ~n1315;
  assign po142 = n1312 | n1316;
  assign n1318 = po221 & ~po142;
  assign n1319 = ~po221 & po142;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = pi192 & pi255;
  assign n1322 = pi014 & ~pi192;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = n576 & ~n1323;
  assign n1325 = pi014 & ~n576;
  assign po214 = n1324 | n1325;
  assign n1327 = n611 & ~n676;
  assign n1328 = n576 & ~n653;
  assign n1329 = ~n620 & ~n660;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~n1327 & n1330;
  assign n1332 = pi193 & ~n1331;
  assign n1333 = n592 & ~n710;
  assign n1334 = ~n592 & ~n703;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~pi193 & ~n1335;
  assign po144 = n1332 | n1336;
  assign n1338 = po214 & ~po144;
  assign n1339 = ~po214 & po144;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = pi013 & ~n576;
  assign n1342 = pi192 & pi197;
  assign n1343 = pi013 & ~pi192;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = n576 & ~n1344;
  assign po195 = n1341 | n1345;
  assign n1347 = n576 & ~n626;
  assign n1348 = ~n617 & ~n620;
  assign n1349 = ~n1347 & ~n1348;
  assign n1350 = n611 & ~n823;
  assign n1351 = n1349 & ~n1350;
  assign n1352 = pi193 & ~n1351;
  assign n1353 = n592 & ~n605;
  assign n1354 = ~n592 & ~n634;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = ~pi193 & ~n1355;
  assign po126 = n1352 | n1356;
  assign n1358 = po195 & ~po126;
  assign n1359 = ~po195 & po126;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~n1340 & n1360;
  assign n1362 = ~n1320 & n1361;
  assign n1363 = ~n592 & ~n798;
  assign n1364 = n592 & ~n805;
  assign n1365 = ~n1363 & ~n1364;
  assign n1366 = ~pi193 & ~n1365;
  assign n1367 = n576 & ~n813;
  assign n1368 = ~n620 & ~n734;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = n611 & ~n727;
  assign n1371 = n1369 & ~n1370;
  assign n1372 = pi193 & ~n1371;
  assign po122 = n1366 | n1372;
  assign n1374 = pi012 & ~n576;
  assign n1375 = pi012 & ~pi192;
  assign n1376 = pi192 & pi221;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = n576 & ~n1377;
  assign po206 = n1374 | n1378;
  assign n1380 = po122 & ~po206;
  assign n1381 = ~n1372 & po206;
  assign n1382 = ~n1366 & n1381;
  assign n1383 = ~n1380 & ~n1382;
  assign n1384 = ~n1362 & n1383;
  assign n1385 = n1340 & n1360;
  assign n1386 = pi192 & pi205;
  assign n1387 = pi027 & ~pi192;
  assign n1388 = ~n1386 & ~n1387;
  assign n1389 = n576 & n1388;
  assign n1390 = ~pi027 & ~n576;
  assign po211 = ~n1389 & ~n1390;
  assign n1392 = ~n592 & ~n754;
  assign n1393 = n592 & n768;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~pi193 & ~n1394;
  assign n1396 = pi071 & ~pi192;
  assign n1397 = pi192 & pi272;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = n576 & ~n1398;
  assign n1400 = pi071 & ~n576;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = n576 & ~n1401;
  assign n1403 = ~n620 & ~n870;
  assign n1404 = n611 & ~n863;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1402 & n1405;
  assign n1407 = pi193 & ~n1406;
  assign po139 = n1395 | n1407;
  assign n1409 = po211 & ~po139;
  assign n1410 = ~po211 & po139;
  assign n1411 = ~n1409 & ~n1410;
  assign n1412 = n1385 & ~n1411;
  assign n1413 = n1384 & ~n1412;
  assign n1414 = n1300 & ~n1413;
  assign n1415 = n1340 & ~n1360;
  assign n1416 = ~n1320 & n1415;
  assign n1417 = ~n1360 & n1411;
  assign n1418 = n1320 & ~n1411;
  assign n1419 = ~n1340 & n1418;
  assign n1420 = ~n1417 & ~n1419;
  assign n1421 = ~n1320 & n1411;
  assign n1422 = n1420 & ~n1421;
  assign n1423 = ~n1416 & n1422;
  assign n1424 = ~n1383 & n1423;
  assign n1425 = n1414 & ~n1424;
  assign n1426 = ~n1340 & ~n1360;
  assign n1427 = n1411 & n1426;
  assign n1428 = n1320 & n1427;
  assign n1429 = n1300 & n1428;
  assign n1430 = ~n1425 & ~n1429;
  assign n1431 = ~po208 & ~po115;
  assign n1432 = po208 & po115;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1320 & n1412;
  assign n1435 = ~n1340 & ~n1383;
  assign n1436 = ~n1320 & n1435;
  assign n1437 = n1320 & n1361;
  assign n1438 = n1411 & n1415;
  assign n1439 = ~n1437 & ~n1438;
  assign n1440 = n1383 & ~n1439;
  assign n1441 = n1320 & n1385;
  assign n1442 = ~n1383 & n1441;
  assign n1443 = ~n1440 & ~n1442;
  assign n1444 = ~n1436 & n1443;
  assign n1445 = ~n1434 & n1444;
  assign n1446 = ~n1360 & n1418;
  assign n1447 = n1340 & n1446;
  assign n1448 = ~n1320 & n1426;
  assign n1449 = ~n1411 & n1448;
  assign n1450 = ~n1447 & ~n1449;
  assign n1451 = n1445 & n1450;
  assign n1452 = n1433 & ~n1451;
  assign n1453 = n1415 & n1421;
  assign n1454 = ~n1447 & ~n1453;
  assign n1455 = n1383 & ~n1454;
  assign n1456 = ~n1452 & ~n1455;
  assign n1457 = n1430 & n1456;
  assign n1458 = ~n1383 & n1427;
  assign n1459 = n1457 & ~n1458;
  assign n1460 = ~pi147 & ~pi192;
  assign n1461 = pi192 & pi216;
  assign n1462 = ~n1460 & ~n1461;
  assign n1463 = n576 & n1462;
  assign n1464 = pi147 & ~n576;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~n1459 & ~n1465;
  assign n1467 = ~n1458 & n1465;
  assign n1468 = n1457 & n1467;
  assign po070 = n1466 | n1468;
  assign n1470 = ~pi149 & ~pi192;
  assign n1471 = pi192 & pi250;
  assign n1472 = ~n1470 & ~n1471;
  assign n1473 = n576 & n1472;
  assign n1474 = pi149 & ~n576;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = n691 & n878;
  assign n1477 = ~n904 & ~n1476;
  assign n1478 = ~n792 & ~n1477;
  assign n1479 = ~n877 & n921;
  assign n1480 = ~n895 & ~n921;
  assign n1481 = ~n792 & ~n1480;
  assign n1482 = n691 & ~n837;
  assign n1483 = ~n886 & ~n1482;
  assign n1484 = ~n792 & ~n877;
  assign n1485 = ~n1483 & n1484;
  assign n1486 = n877 & n886;
  assign n1487 = n742 & n877;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n906 & n1488;
  assign n1490 = n792 & ~n1489;
  assign n1491 = n792 & ~n892;
  assign n1492 = ~n877 & n1491;
  assign n1493 = ~n1490 & ~n1492;
  assign n1494 = ~n1485 & n1493;
  assign n1495 = ~n1481 & n1494;
  assign n1496 = n641 & ~n1495;
  assign n1497 = ~n1479 & ~n1496;
  assign n1498 = ~n877 & n895;
  assign n1499 = n837 & n1484;
  assign n1500 = ~n888 & ~n1499;
  assign n1501 = n837 & n877;
  assign n1502 = ~n691 & n1501;
  assign n1503 = ~n877 & n926;
  assign n1504 = n691 & ~n877;
  assign n1505 = ~n837 & n1504;
  assign n1506 = ~n741 & n1505;
  assign n1507 = ~n1503 & ~n1506;
  assign n1508 = ~n1502 & n1507;
  assign n1509 = n792 & ~n1508;
  assign n1510 = n877 & n890;
  assign n1511 = ~n792 & n1510;
  assign n1512 = ~n839 & ~n1511;
  assign n1513 = ~n1509 & n1512;
  assign n1514 = n1500 & n1513;
  assign n1515 = ~n1498 & n1514;
  assign n1516 = ~n641 & ~n1515;
  assign n1517 = n1497 & ~n1516;
  assign n1518 = ~n1478 & n1517;
  assign n1519 = ~n1475 & ~n1518;
  assign n1520 = n1475 & n1518;
  assign po071 = n1519 | n1520;
  assign n1522 = ~pi129 & ~pi192;
  assign n1523 = pi192 & pi248;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = n576 & n1524;
  assign n1526 = pi129 & ~n576;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = ~n792 & n888;
  assign n1529 = ~n691 & ~n877;
  assign n1530 = n886 & n1529;
  assign n1531 = n792 & n1530;
  assign n1532 = ~n908 & ~n921;
  assign n1533 = ~n877 & ~n1532;
  assign n1534 = n792 & n1533;
  assign n1535 = ~n1531 & ~n1534;
  assign n1536 = ~n1528 & n1535;
  assign n1537 = ~n691 & ~n741;
  assign n1538 = n1484 & n1537;
  assign n1539 = ~n691 & n741;
  assign n1540 = ~n906 & ~n1539;
  assign n1541 = ~n792 & n877;
  assign n1542 = ~n1540 & n1541;
  assign n1543 = ~n1538 & ~n1542;
  assign n1544 = ~n1533 & n1543;
  assign n1545 = n792 & ~n877;
  assign n1546 = n883 & n1545;
  assign n1547 = n792 & n877;
  assign n1548 = n1537 & n1547;
  assign n1549 = n792 & ~n1532;
  assign n1550 = ~n1548 & ~n1549;
  assign n1551 = ~n1546 & n1550;
  assign n1552 = n1544 & n1551;
  assign n1553 = ~n641 & ~n1552;
  assign n1554 = n1536 & ~n1553;
  assign n1555 = n837 & n1545;
  assign n1556 = ~n741 & n1555;
  assign n1557 = n883 & n1484;
  assign n1558 = ~n691 & n1557;
  assign n1559 = ~n792 & n887;
  assign n1560 = n691 & n741;
  assign n1561 = ~n1537 & ~n1560;
  assign n1562 = ~n890 & n1561;
  assign n1563 = n1541 & ~n1562;
  assign n1564 = ~n1559 & ~n1563;
  assign n1565 = ~n1558 & n1564;
  assign n1566 = ~n1556 & n1565;
  assign n1567 = n877 & n884;
  assign n1568 = ~n906 & ~n1567;
  assign n1569 = n792 & ~n1568;
  assign n1570 = n1566 & ~n1569;
  assign n1571 = ~n888 & ~n907;
  assign n1572 = n1570 & n1571;
  assign n1573 = n641 & ~n1572;
  assign n1574 = n1554 & ~n1573;
  assign n1575 = ~n1527 & ~n1574;
  assign n1576 = ~n1553 & ~n1573;
  assign n1577 = n1535 & n1576;
  assign n1578 = ~n1528 & n1577;
  assign n1579 = n1527 & n1578;
  assign po072 = n1575 | n1579;
  assign n1581 = ~n1383 & n1418;
  assign n1582 = n1361 & n1581;
  assign n1583 = ~n1320 & ~n1433;
  assign n1584 = n1427 & n1583;
  assign n1585 = ~n1320 & n1383;
  assign n1586 = n1385 & n1585;
  assign n1587 = n1411 & n1586;
  assign n1588 = n1361 & ~n1411;
  assign n1589 = n1585 & n1588;
  assign n1590 = n1383 & ~n1411;
  assign n1591 = ~n1360 & n1590;
  assign n1592 = n1340 & n1591;
  assign n1593 = n1320 & n1411;
  assign n1594 = ~n1340 & n1593;
  assign n1595 = n1320 & n1426;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = n1383 & ~n1596;
  assign n1598 = ~n1592 & ~n1597;
  assign n1599 = ~n1589 & n1598;
  assign n1600 = ~n1587 & n1599;
  assign n1601 = ~n1433 & ~n1600;
  assign n1602 = n1385 & n1418;
  assign n1603 = n1383 & n1602;
  assign n1604 = n1383 & n1427;
  assign n1605 = n1320 & n1604;
  assign n1606 = ~n1603 & ~n1605;
  assign n1607 = n1340 & n1593;
  assign n1608 = ~n1438 & ~n1607;
  assign n1609 = ~n1434 & n1608;
  assign n1610 = ~n1448 & n1609;
  assign n1611 = ~n1383 & ~n1610;
  assign n1612 = ~n1433 & n1611;
  assign n1613 = n1606 & ~n1612;
  assign n1614 = ~n1601 & n1613;
  assign n1615 = ~n1584 & n1614;
  assign n1616 = ~n1582 & n1615;
  assign n1617 = ~n1588 & ~n1595;
  assign n1618 = ~n1383 & ~n1617;
  assign n1619 = n1361 & n1421;
  assign n1620 = n1360 & n1421;
  assign n1621 = ~n1320 & ~n1411;
  assign n1622 = ~n1360 & n1621;
  assign n1623 = n1340 & n1622;
  assign n1624 = ~n1620 & ~n1623;
  assign n1625 = ~n1383 & ~n1624;
  assign n1626 = ~n1619 & ~n1625;
  assign n1627 = ~n1438 & ~n1441;
  assign n1628 = ~n1412 & ~n1449;
  assign n1629 = n1627 & n1628;
  assign n1630 = n1383 & ~n1629;
  assign n1631 = ~n1602 & ~n1630;
  assign n1632 = n1626 & n1631;
  assign n1633 = ~n1618 & n1632;
  assign n1634 = ~n1300 & ~n1633;
  assign n1635 = n1616 & ~n1634;
  assign n1636 = ~pi136 & ~pi192;
  assign n1637 = pi192 & pi238;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = n576 & n1638;
  assign n1640 = pi136 & ~n576;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = ~n1635 & ~n1641;
  assign n1643 = ~n1582 & n1641;
  assign n1644 = n1615 & ~n1634;
  assign n1645 = n1643 & n1644;
  assign po073 = n1642 | n1645;
  assign n1647 = ~pi121 & ~pi192;
  assign n1648 = pi192 & pi256;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = n576 & n1649;
  assign n1651 = pi121 & ~n576;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = ~n1453 & ~n1588;
  assign n1654 = ~n1428 & n1653;
  assign n1655 = ~n1383 & ~n1654;
  assign n1656 = n1385 & n1411;
  assign n1657 = ~n1447 & ~n1656;
  assign n1658 = ~n1383 & ~n1657;
  assign n1659 = n1360 & n1593;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = ~n1453 & n1660;
  assign n1662 = ~n1411 & n1595;
  assign n1663 = n1361 & n1411;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = n1383 & ~n1664;
  assign n1666 = ~n1458 & ~n1665;
  assign n1667 = n1661 & n1666;
  assign n1668 = ~n1300 & ~n1667;
  assign n1669 = ~n1340 & ~n1411;
  assign n1670 = ~n1320 & n1669;
  assign n1671 = ~n1362 & ~n1670;
  assign n1672 = ~n1383 & ~n1671;
  assign n1673 = n1320 & n1415;
  assign n1674 = n1383 & n1673;
  assign n1675 = ~n1604 & ~n1674;
  assign n1676 = ~n1442 & n1675;
  assign n1677 = ~n1623 & n1676;
  assign n1678 = ~n1672 & n1677;
  assign n1679 = n1361 & n1418;
  assign n1680 = n1678 & ~n1679;
  assign n1681 = ~n1433 & ~n1680;
  assign n1682 = n1340 & ~n1411;
  assign n1683 = n1585 & n1682;
  assign n1684 = ~n1681 & ~n1683;
  assign n1685 = ~n1668 & n1684;
  assign n1686 = ~n1655 & n1685;
  assign n1687 = ~n1652 & ~n1686;
  assign n1688 = n1652 & n1686;
  assign po074 = n1687 | n1688;
  assign n1690 = ~pi010 & ~pi192;
  assign n1691 = pi192 & ~pi231;
  assign n1692 = ~n1690 & ~n1691;
  assign n1693 = n576 & ~n1692;
  assign n1694 = ~pi010 & ~n576;
  assign po216 = ~n1693 & ~n1694;
  assign n1696 = pi050 & ~n576;
  assign n1697 = pi050 & ~pi192;
  assign n1698 = pi192 & pi313;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = n576 & ~n1699;
  assign n1701 = ~n1696 & ~n1700;
  assign n1702 = n576 & ~n1701;
  assign n1703 = n611 & ~n1204;
  assign n1704 = ~n620 & ~n1211;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = ~n1702 & n1705;
  assign n1707 = pi193 & ~n1706;
  assign n1708 = n592 & ~n1017;
  assign n1709 = ~n592 & ~n1010;
  assign n1710 = ~n1708 & ~n1709;
  assign n1711 = ~pi193 & ~n1710;
  assign po118 = n1707 | n1711;
  assign n1713 = ~po216 & ~po118;
  assign n1714 = po216 & po118;
  assign n1715 = ~n1713 & ~n1714;
  assign n1716 = n592 & ~n1204;
  assign n1717 = ~n592 & ~n1193;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = ~pi193 & ~n1718;
  assign n1720 = ~n620 & ~n1154;
  assign n1721 = n611 & ~n1161;
  assign n1722 = n576 & ~n1186;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = ~n1720 & n1723;
  assign n1725 = pi193 & ~n1724;
  assign po130 = n1719 | n1725;
  assign n1727 = pi011 & ~n576;
  assign n1728 = pi011 & ~pi192;
  assign n1729 = pi192 & pi215;
  assign n1730 = ~n1728 & ~n1729;
  assign n1731 = n576 & ~n1730;
  assign po191 = n1727 | n1731;
  assign n1733 = ~po130 & po191;
  assign n1734 = po130 & ~po191;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = pi192 & pi223;
  assign n1737 = pi025 & ~pi192;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = n576 & n1738;
  assign n1740 = ~pi025 & ~n576;
  assign po209 = ~n1739 & ~n1740;
  assign n1742 = ~n592 & ~n1144;
  assign n1743 = n592 & ~n1137;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = ~pi193 & ~n1744;
  assign n1746 = n611 & ~n961;
  assign n1747 = n576 & ~n978;
  assign n1748 = ~n620 & ~n971;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~n1746 & n1749;
  assign n1751 = pi193 & ~n1750;
  assign po120 = n1745 | n1751;
  assign n1753 = po209 & ~po120;
  assign n1754 = ~po209 & po120;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = n576 & n947;
  assign n1757 = ~n620 & ~n954;
  assign n1758 = ~n1756 & ~n1757;
  assign n1759 = pi056 & ~n576;
  assign n1760 = pi056 & ~pi192;
  assign n1761 = pi192 & pi290;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = n576 & ~n1762;
  assign n1764 = ~n1759 & ~n1763;
  assign n1765 = n611 & ~n1764;
  assign n1766 = n1758 & ~n1765;
  assign n1767 = pi193 & ~n1766;
  assign n1768 = ~n592 & ~n961;
  assign n1769 = n592 & ~n971;
  assign n1770 = ~n1768 & ~n1769;
  assign n1771 = ~pi193 & ~n1770;
  assign po138 = n1767 | n1771;
  assign n1773 = pi006 & ~n576;
  assign n1774 = pi006 & ~pi192;
  assign n1775 = pi192 & pi257;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = n576 & ~n1776;
  assign po189 = n1773 | n1777;
  assign n1779 = po138 & ~po189;
  assign n1780 = ~po138 & po189;
  assign n1781 = ~n1779 & ~n1780;
  assign n1782 = ~n592 & ~n1034;
  assign n1783 = n592 & n1097;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~pi193 & ~n1784;
  assign n1786 = ~n620 & ~n1003;
  assign n1787 = n576 & ~n1027;
  assign n1788 = ~n1786 & ~n1787;
  assign n1789 = n611 & ~n1017;
  assign n1790 = n1788 & ~n1789;
  assign n1791 = pi193 & ~n1790;
  assign po141 = n1785 | n1791;
  assign n1793 = pi016 & ~n576;
  assign n1794 = pi016 & ~pi192;
  assign n1795 = pi192 & pi207;
  assign n1796 = ~n1794 & ~n1795;
  assign n1797 = n576 & ~n1796;
  assign po203 = n1793 | n1797;
  assign n1799 = ~po141 & po203;
  assign n1800 = po141 & ~po203;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = ~n1781 & ~n1801;
  assign n1803 = ~n1755 & n1802;
  assign n1804 = n1735 & n1803;
  assign n1805 = pi192 & pi199;
  assign n1806 = pi008 & ~pi192;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = n576 & n1807;
  assign n1809 = ~pi008 & ~n576;
  assign po222 = ~n1808 & ~n1809;
  assign n1811 = n576 & ~n1054;
  assign n1812 = ~n620 & ~n1047;
  assign n1813 = n611 & ~n1070;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = ~n1811 & n1814;
  assign n1816 = pi193 & ~n1815;
  assign n1817 = n592 & ~n1764;
  assign n1818 = pi060 & ~pi192;
  assign n1819 = pi192 & pi283;
  assign n1820 = ~n1818 & ~n1819;
  assign n1821 = n576 & ~n1820;
  assign n1822 = pi060 & ~n576;
  assign n1823 = ~n1821 & ~n1822;
  assign n1824 = ~n592 & ~n1823;
  assign n1825 = ~n1817 & ~n1824;
  assign n1826 = ~pi193 & ~n1825;
  assign po123 = n1816 | n1826;
  assign n1828 = po222 & ~po123;
  assign n1829 = ~po222 & po123;
  assign n1830 = ~n1828 & ~n1829;
  assign n1831 = n1781 & ~n1830;
  assign n1832 = ~n1801 & n1831;
  assign n1833 = ~n1735 & n1832;
  assign n1834 = ~n1735 & n1801;
  assign n1835 = ~n1781 & n1834;
  assign n1836 = ~n1833 & ~n1835;
  assign n1837 = ~n1755 & ~n1836;
  assign n1838 = ~n1804 & ~n1837;
  assign n1839 = ~n1715 & ~n1838;
  assign n1840 = n1735 & n1801;
  assign n1841 = ~n1781 & n1840;
  assign n1842 = n1755 & n1841;
  assign n1843 = n1735 & n1830;
  assign n1844 = ~n1781 & n1843;
  assign n1845 = ~n1801 & n1844;
  assign n1846 = ~n1842 & ~n1845;
  assign n1847 = ~n1735 & n1755;
  assign n1848 = n1781 & n1801;
  assign n1849 = ~n1781 & ~n1830;
  assign n1850 = ~n1801 & n1849;
  assign n1851 = ~n1848 & ~n1850;
  assign n1852 = n1781 & n1830;
  assign n1853 = n1851 & ~n1852;
  assign n1854 = n1847 & ~n1853;
  assign n1855 = n1846 & ~n1854;
  assign n1856 = ~n1715 & ~n1855;
  assign n1857 = ~n1839 & ~n1856;
  assign n1858 = n1781 & n1840;
  assign n1859 = ~n1830 & n1858;
  assign n1860 = n1781 & n1834;
  assign n1861 = n1830 & n1860;
  assign n1862 = ~n1859 & ~n1861;
  assign n1863 = ~n1845 & n1862;
  assign n1864 = ~n1755 & ~n1863;
  assign n1865 = n1715 & n1755;
  assign n1866 = ~n1781 & n1830;
  assign n1867 = ~n1735 & n1866;
  assign n1868 = n1735 & ~n1830;
  assign n1869 = ~n1801 & n1868;
  assign n1870 = ~n1867 & ~n1869;
  assign n1871 = ~n1832 & n1870;
  assign n1872 = ~n1835 & n1871;
  assign n1873 = n1865 & ~n1872;
  assign n1874 = ~n1735 & n1852;
  assign n1875 = ~n1735 & n1850;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = n1801 & n1831;
  assign n1878 = ~n1841 & ~n1877;
  assign n1879 = n1876 & n1878;
  assign n1880 = ~n1755 & ~n1879;
  assign n1881 = n1735 & n1832;
  assign n1882 = ~n1880 & ~n1881;
  assign n1883 = n1715 & ~n1882;
  assign n1884 = n1840 & n1852;
  assign n1885 = ~n1881 & ~n1884;
  assign n1886 = n1755 & ~n1885;
  assign n1887 = ~n1883 & ~n1886;
  assign n1888 = ~n1873 & n1887;
  assign n1889 = ~n1864 & n1888;
  assign n1890 = n1857 & n1889;
  assign n1891 = ~pi142 & ~pi192;
  assign n1892 = pi192 & pi252;
  assign n1893 = ~n1891 & ~n1892;
  assign n1894 = n576 & n1893;
  assign n1895 = pi142 & ~n576;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = ~n1890 & ~n1896;
  assign n1898 = n1889 & n1896;
  assign n1899 = n1857 & n1898;
  assign po075 = n1897 | n1899;
  assign n1901 = ~pi154 & ~pi192;
  assign n1902 = pi192 & pi198;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = n576 & n1903;
  assign n1905 = pi154 & ~n576;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = ~n1122 & ~n1241;
  assign n1908 = ~n991 & ~n1091;
  assign n1909 = n1907 & ~n1908;
  assign n1910 = n1256 & ~n1909;
  assign n1911 = n991 & n1174;
  assign n1912 = n1121 & n1911;
  assign n1913 = n1041 & n1912;
  assign n1914 = n991 & n1232;
  assign n1915 = ~n1913 & ~n1914;
  assign n1916 = ~n1910 & n1915;
  assign n1917 = ~n991 & n1230;
  assign n1918 = ~n1041 & n1917;
  assign n1919 = ~n991 & n1041;
  assign n1920 = n1174 & n1919;
  assign n1921 = ~n1180 & ~n1920;
  assign n1922 = ~n1091 & ~n1921;
  assign n1923 = ~n1123 & n1174;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = ~n1918 & n1924;
  assign n1926 = ~n991 & ~n1041;
  assign n1927 = n1091 & n1926;
  assign n1928 = ~n1917 & ~n1927;
  assign n1929 = ~n1174 & ~n1928;
  assign n1930 = n1925 & ~n1929;
  assign n1931 = ~n1224 & ~n1930;
  assign n1932 = ~n991 & n1228;
  assign n1933 = n991 & n1249;
  assign n1934 = n1118 & n1933;
  assign n1935 = ~n1932 & ~n1934;
  assign n1936 = ~n1174 & ~n1935;
  assign n1937 = ~n1931 & ~n1936;
  assign n1938 = n1174 & n1228;
  assign n1939 = ~n1041 & n1091;
  assign n1940 = n1118 & n1939;
  assign n1941 = ~n991 & n1255;
  assign n1942 = ~n1940 & ~n1941;
  assign n1943 = n1174 & ~n1942;
  assign n1944 = ~n1938 & ~n1943;
  assign n1945 = n1224 & ~n1944;
  assign n1946 = n1937 & ~n1945;
  assign n1947 = n1916 & n1946;
  assign n1948 = ~n1906 & ~n1947;
  assign n1949 = n1916 & n1937;
  assign n1950 = n1906 & n1949;
  assign n1951 = ~n1945 & n1950;
  assign po076 = n1948 | n1951;
  assign n1953 = ~n1118 & n1919;
  assign n1954 = ~n1908 & ~n1953;
  assign n1955 = ~n1175 & n1954;
  assign n1956 = n1174 & ~n1955;
  assign n1957 = n1118 & n1919;
  assign n1958 = ~n1225 & ~n1957;
  assign n1959 = ~n1918 & n1958;
  assign n1960 = ~n1174 & ~n1959;
  assign n1961 = ~n1238 & ~n1245;
  assign n1962 = ~n1960 & n1961;
  assign n1963 = ~n1956 & n1962;
  assign n1964 = n1224 & ~n1963;
  assign n1965 = ~n991 & n1225;
  assign n1966 = n1180 & n1255;
  assign n1967 = ~n1938 & ~n1966;
  assign n1968 = ~n1965 & n1967;
  assign n1969 = ~n1912 & n1968;
  assign n1970 = ~n1118 & n1234;
  assign n1971 = ~n991 & n1940;
  assign n1972 = ~n1970 & ~n1971;
  assign n1973 = ~n1255 & ~n1934;
  assign n1974 = n1972 & n1973;
  assign n1975 = ~n1174 & ~n1974;
  assign n1976 = ~n1118 & n1174;
  assign n1977 = n1926 & n1976;
  assign n1978 = ~n1975 & ~n1977;
  assign n1979 = ~n1932 & n1978;
  assign n1980 = n1091 & n1234;
  assign n1981 = n1174 & n1225;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = n1979 & n1982;
  assign n1984 = ~n1224 & ~n1983;
  assign n1985 = n1969 & ~n1984;
  assign n1986 = ~n1964 & n1985;
  assign n1987 = ~pi130 & ~pi192;
  assign n1988 = pi192 & pi242;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = n576 & n1989;
  assign n1991 = pi130 & ~n576;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = ~n1986 & ~n1992;
  assign n1994 = n1969 & n1992;
  assign n1995 = ~n1964 & n1994;
  assign n1996 = ~n1984 & n1995;
  assign po077 = n1993 | n1996;
  assign n1998 = ~pi148 & ~pi192;
  assign n1999 = pi192 & pi230;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = n576 & n2000;
  assign n2002 = pi148 & ~n576;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = n592 & ~n1027;
  assign n2005 = ~n592 & ~n1003;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = ~pi193 & n2006;
  assign n2008 = n611 & ~n1701;
  assign n2009 = ~n620 & ~n1010;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = n576 & ~n1017;
  assign n2012 = n2010 & ~n2011;
  assign n2013 = pi193 & n2012;
  assign po104 = ~n2007 & ~n2013;
  assign n2015 = ~po222 & po104;
  assign n2016 = po222 & ~po104;
  assign n2017 = ~n2015 & ~n2016;
  assign n2018 = n592 & n947;
  assign n2019 = ~n592 & ~n954;
  assign n2020 = ~n2018 & ~n2019;
  assign n2021 = ~pi193 & ~n2020;
  assign n2022 = ~n620 & ~n1823;
  assign n2023 = n576 & ~n1764;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = n611 & ~n1054;
  assign n2026 = n2024 & ~n2025;
  assign n2027 = pi193 & ~n2026;
  assign po124 = n2021 | n2027;
  assign n2029 = ~po189 & po124;
  assign n2030 = po189 & ~po124;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = ~n620 & ~n1161;
  assign n2033 = n611 & ~n1130;
  assign n2034 = n576 & ~n1154;
  assign n2035 = ~n2033 & ~n2034;
  assign n2036 = ~n2032 & n2035;
  assign n2037 = pi193 & ~n2036;
  assign n2038 = ~n592 & ~n1186;
  assign n2039 = n592 & ~n1193;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~pi193 & ~n2040;
  assign po154 = n2037 | n2041;
  assign n2043 = po194 & ~po154;
  assign n2044 = ~po194 & po154;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = n592 & ~n1701;
  assign n2047 = ~n592 & ~n1211;
  assign n2048 = ~n2046 & ~n2047;
  assign n2049 = ~pi193 & ~n2048;
  assign n2050 = n611 & ~n1186;
  assign n2051 = n576 & ~n1204;
  assign n2052 = ~n620 & ~n1193;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n2050 & n2053;
  assign n2055 = pi193 & ~n2054;
  assign po131 = n2049 | n2055;
  assign n2057 = pi004 & ~n576;
  assign n2058 = pi004 & ~pi192;
  assign n2059 = pi192 & pi249;
  assign n2060 = ~n2058 & ~n2059;
  assign n2061 = n576 & ~n2060;
  assign po197 = n2057 | n2061;
  assign n2063 = po131 & ~po197;
  assign n2064 = ~po131 & po197;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = n592 & ~n1070;
  assign n2067 = ~n592 & ~n1077;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = ~pi193 & ~n2068;
  assign n2070 = n611 & ~n1034;
  assign n2071 = n576 & ~n1063;
  assign n2072 = ~n620 & n1097;
  assign n2073 = ~n2071 & ~n2072;
  assign n2074 = ~n2070 & n2073;
  assign n2075 = pi193 & ~n2074;
  assign po125 = n2069 | n2075;
  assign n2077 = pi192 & pi241;
  assign n2078 = pi022 & ~pi192;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = n576 & n2079;
  assign n2081 = ~pi022 & ~n576;
  assign po205 = ~n2080 & ~n2081;
  assign n2083 = ~po125 & po205;
  assign n2084 = po125 & ~po205;
  assign n2085 = ~n2083 & ~n2084;
  assign n2086 = n2065 & n2085;
  assign n2087 = ~n2045 & n2086;
  assign n2088 = n576 & ~n1137;
  assign n2089 = ~n620 & ~n1144;
  assign n2090 = n611 & ~n978;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2088 & n2091;
  assign n2093 = pi193 & ~n2092;
  assign n2094 = ~n592 & ~n1130;
  assign n2095 = n592 & ~n1161;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~pi193 & ~n2096;
  assign po152 = n2093 | n2097;
  assign n2099 = ~po224 & ~po152;
  assign n2100 = po224 & po152;
  assign n2101 = ~n2099 & ~n2100;
  assign n2102 = ~n2085 & n2101;
  assign n2103 = ~n2065 & n2102;
  assign n2104 = ~n2087 & ~n2103;
  assign n2105 = n2045 & ~n2101;
  assign n2106 = ~n2085 & n2105;
  assign n2107 = ~n2045 & ~n2101;
  assign n2108 = n2085 & n2107;
  assign n2109 = ~n2106 & ~n2108;
  assign n2110 = n2104 & n2109;
  assign n2111 = n2031 & ~n2110;
  assign n2112 = ~n2065 & n2106;
  assign n2113 = ~n2111 & ~n2112;
  assign n2114 = ~n2085 & n2107;
  assign n2115 = n2045 & n2086;
  assign n2116 = ~n2114 & ~n2115;
  assign n2117 = n2045 & n2101;
  assign n2118 = n2065 & n2117;
  assign n2119 = n2116 & ~n2118;
  assign n2120 = ~n2045 & n2085;
  assign n2121 = ~n2065 & n2120;
  assign n2122 = n2101 & n2121;
  assign n2123 = n2119 & ~n2122;
  assign n2124 = ~n2031 & ~n2123;
  assign n2125 = n2113 & ~n2124;
  assign n2126 = n2017 & ~n2125;
  assign n2127 = ~n2065 & n2107;
  assign n2128 = ~n2045 & n2101;
  assign n2129 = n2065 & n2128;
  assign n2130 = ~n2127 & ~n2129;
  assign n2131 = ~n2085 & n2117;
  assign n2132 = ~n2065 & n2131;
  assign n2133 = n2065 & ~n2085;
  assign n2134 = n2045 & n2133;
  assign n2135 = ~n2101 & n2134;
  assign n2136 = ~n2132 & ~n2135;
  assign n2137 = n2130 & n2136;
  assign n2138 = ~n2031 & ~n2137;
  assign n2139 = n2085 & n2105;
  assign n2140 = ~n2114 & ~n2139;
  assign n2141 = n2065 & n2102;
  assign n2142 = ~n2065 & n2085;
  assign n2143 = n2101 & n2142;
  assign n2144 = ~n2141 & ~n2143;
  assign n2145 = n2140 & n2144;
  assign n2146 = n2031 & ~n2145;
  assign n2147 = n2105 & n2142;
  assign n2148 = ~n2146 & ~n2147;
  assign n2149 = ~n2138 & n2148;
  assign n2150 = ~n2017 & ~n2149;
  assign n2151 = n2031 & ~n2065;
  assign n2152 = n2085 & n2151;
  assign n2153 = n2117 & n2152;
  assign n2154 = ~n2085 & n2128;
  assign n2155 = ~n2031 & n2154;
  assign n2156 = n2085 & n2117;
  assign n2157 = ~n2031 & n2156;
  assign n2158 = ~n2155 & ~n2157;
  assign n2159 = n2065 & ~n2158;
  assign n2160 = ~n2153 & ~n2159;
  assign n2161 = ~n2150 & n2160;
  assign n2162 = ~n2126 & n2161;
  assign n2163 = n2003 & ~n2162;
  assign n2164 = ~n2003 & n2162;
  assign po078 = n2163 | n2164;
  assign n2166 = ~n592 & ~n761;
  assign n2167 = n592 & ~n778;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~pi193 & ~n2168;
  assign n2170 = ~n620 & ~n754;
  assign n2171 = n576 & n768;
  assign n2172 = n611 & ~n1401;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = ~n2170 & n2173;
  assign n2175 = pi193 & ~n2174;
  assign po116 = n2169 | n2175;
  assign n2177 = po210 & ~po116;
  assign n2178 = ~po210 & po116;
  assign n2179 = ~n2177 & ~n2178;
  assign n2180 = pi192 & pi237;
  assign n2181 = pi000 & ~pi192;
  assign n2182 = ~n2180 & ~n2181;
  assign n2183 = n576 & n2182;
  assign n2184 = ~pi000 & ~n576;
  assign po207 = ~n2183 & ~n2184;
  assign n2186 = n576 & ~n617;
  assign n2187 = ~n620 & ~n823;
  assign n2188 = n611 & ~n805;
  assign n2189 = ~n2187 & ~n2188;
  assign n2190 = ~n2186 & n2189;
  assign n2191 = pi193 & ~n2190;
  assign n2192 = n592 & ~n634;
  assign n2193 = ~n592 & ~n626;
  assign n2194 = ~n2192 & ~n2193;
  assign n2195 = ~pi193 & ~n2194;
  assign po145 = n2191 | n2195;
  assign n2197 = ~po207 & ~po145;
  assign n2198 = po207 & po145;
  assign n2199 = ~n2197 & ~n2198;
  assign n2200 = n611 & ~n669;
  assign n2201 = ~n620 & ~n676;
  assign n2202 = n576 & ~n660;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = ~n2200 & n2203;
  assign n2205 = pi193 & ~n2204;
  assign n2206 = ~n592 & ~n653;
  assign n2207 = n592 & ~n703;
  assign n2208 = ~n2206 & ~n2207;
  assign n2209 = ~pi193 & ~n2208;
  assign po159 = n2205 | n2209;
  assign n2211 = ~po208 & po159;
  assign n2212 = po208 & ~po159;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = ~n592 & ~n1401;
  assign n2215 = n592 & ~n754;
  assign n2216 = ~n2214 & ~n2215;
  assign n2217 = ~pi193 & ~n2216;
  assign n2218 = n611 & ~n851;
  assign n2219 = ~n620 & ~n863;
  assign n2220 = n576 & ~n870;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = ~n2218 & n2221;
  assign n2223 = pi193 & ~n2222;
  assign po143 = n2217 | n2223;
  assign n2225 = ~po206 & ~po143;
  assign n2226 = po206 & po143;
  assign n2227 = ~n2225 & ~n2226;
  assign n2228 = n2213 & ~n2227;
  assign n2229 = n2199 & n2228;
  assign n2230 = pi192 & pi245;
  assign n2231 = pi001 & ~pi192;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = n576 & ~n2232;
  assign n2234 = pi001 & ~n576;
  assign po213 = n2233 | n2234;
  assign n2236 = ~n592 & ~n734;
  assign n2237 = n592 & ~n813;
  assign n2238 = ~n2236 & ~n2237;
  assign n2239 = ~pi193 & ~n2238;
  assign n2240 = n611 & ~n710;
  assign n2241 = ~n620 & ~n717;
  assign n2242 = n576 & ~n727;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = ~n2240 & n2243;
  assign n2245 = pi193 & ~n2244;
  assign po127 = n2239 | n2245;
  assign n2247 = ~po213 & ~po127;
  assign n2248 = po213 & po127;
  assign n2249 = ~n2247 & ~n2248;
  assign n2250 = n2199 & ~n2227;
  assign n2251 = n2249 & n2250;
  assign n2252 = ~n2229 & ~n2251;
  assign n2253 = ~n2179 & ~n2252;
  assign n2254 = n2199 & ~n2249;
  assign n2255 = ~n2213 & n2254;
  assign n2256 = ~n2227 & n2255;
  assign n2257 = ~n2199 & ~n2227;
  assign n2258 = n2249 & n2257;
  assign n2259 = ~n2256 & ~n2258;
  assign n2260 = n2179 & ~n2259;
  assign n2261 = n2229 & n2249;
  assign n2262 = n2213 & n2227;
  assign n2263 = ~n2249 & n2262;
  assign n2264 = n2199 & n2263;
  assign n2265 = n2199 & ~n2213;
  assign n2266 = n2227 & n2265;
  assign n2267 = n2249 & n2266;
  assign n2268 = ~n2264 & ~n2267;
  assign n2269 = ~n2261 & n2268;
  assign n2270 = ~n2260 & n2269;
  assign n2271 = ~n2253 & n2270;
  assign n2272 = n592 & ~n823;
  assign n2273 = ~n592 & ~n805;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~pi193 & ~n2274;
  assign n2276 = ~n620 & ~n813;
  assign n2277 = n576 & ~n798;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = n611 & ~n734;
  assign n2280 = n2278 & ~n2279;
  assign n2281 = pi193 & ~n2280;
  assign po110 = n2275 | n2281;
  assign n2283 = po220 & ~po110;
  assign n2284 = ~po220 & po110;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = ~n2271 & ~n2285;
  assign n2287 = ~n2199 & n2249;
  assign n2288 = n2213 & n2287;
  assign n2289 = n2227 & n2288;
  assign n2290 = ~n2261 & ~n2289;
  assign n2291 = ~n2213 & ~n2227;
  assign n2292 = ~n2199 & n2291;
  assign n2293 = n2199 & n2227;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = ~n2249 & ~n2294;
  assign n2296 = n2290 & ~n2295;
  assign n2297 = ~n2179 & ~n2296;
  assign n2298 = ~n2286 & ~n2297;
  assign n2299 = ~n2249 & n2257;
  assign n2300 = n2199 & n2291;
  assign n2301 = n2249 & n2300;
  assign n2302 = n2249 & n2262;
  assign n2303 = n2199 & n2302;
  assign n2304 = ~n2301 & ~n2303;
  assign n2305 = n2228 & ~n2249;
  assign n2306 = n2304 & ~n2305;
  assign n2307 = n2179 & ~n2306;
  assign n2308 = ~n2299 & ~n2307;
  assign n2309 = ~n2249 & n2266;
  assign n2310 = n2308 & ~n2309;
  assign n2311 = n2285 & ~n2310;
  assign n2312 = ~n2213 & n2227;
  assign n2313 = ~n2249 & n2312;
  assign n2314 = ~n2292 & ~n2313;
  assign n2315 = ~n2179 & n2285;
  assign n2316 = ~n2314 & n2315;
  assign n2317 = ~n2311 & ~n2316;
  assign n2318 = ~n2199 & n2227;
  assign n2319 = ~n2213 & n2318;
  assign n2320 = n2249 & n2319;
  assign n2321 = ~n2199 & n2262;
  assign n2322 = ~n2249 & n2321;
  assign n2323 = ~n2320 & ~n2322;
  assign n2324 = n2179 & ~n2323;
  assign n2325 = n2317 & ~n2324;
  assign n2326 = n2298 & n2325;
  assign n2327 = ~pi123 & ~pi192;
  assign n2328 = pi192 & pi214;
  assign n2329 = ~n2327 & ~n2328;
  assign n2330 = n576 & n2329;
  assign n2331 = pi123 & ~n576;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = ~n2326 & n2332;
  assign n2334 = n2298 & ~n2332;
  assign n2335 = n2317 & n2334;
  assign n2336 = ~n2324 & n2335;
  assign po079 = n2333 | n2336;
  assign n2338 = ~n592 & n1097;
  assign n2339 = n592 & ~n1063;
  assign n2340 = ~n2338 & ~n2339;
  assign n2341 = ~pi193 & ~n2340;
  assign n2342 = n611 & ~n1003;
  assign n2343 = ~n620 & ~n1027;
  assign n2344 = n576 & ~n1034;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2342 & n2345;
  assign n2347 = pi193 & ~n2346;
  assign po112 = n2341 | n2347;
  assign n2349 = po214 & ~po112;
  assign n2350 = ~po214 & po112;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n620 & ~n1054;
  assign n2353 = n611 & ~n1047;
  assign n2354 = ~n2352 & ~n2353;
  assign n2355 = n576 & ~n1823;
  assign n2356 = n2354 & ~n2355;
  assign n2357 = pi193 & ~n2356;
  assign n2358 = ~n592 & ~n1764;
  assign n2359 = n592 & ~n954;
  assign n2360 = ~n2358 & ~n2359;
  assign n2361 = ~pi193 & ~n2360;
  assign po128 = n2357 | n2361;
  assign n2363 = pi192 & pi247;
  assign n2364 = pi015 & ~pi192;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = n576 & n2365;
  assign n2367 = ~pi015 & ~n576;
  assign po193 = ~n2366 & ~n2367;
  assign n2369 = ~po128 & po193;
  assign n2370 = po128 & ~po193;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = ~n592 & ~n1137;
  assign n2373 = n592 & ~n1130;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = ~pi193 & ~n2374;
  assign n2376 = n611 & ~n971;
  assign n2377 = n576 & ~n1144;
  assign n2378 = ~n620 & ~n978;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = ~n2376 & n2379;
  assign n2381 = pi193 & ~n2380;
  assign po119 = n2375 | n2381;
  assign n2383 = pi192 & pi239;
  assign n2384 = pi005 & ~pi192;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = n576 & n2385;
  assign n2387 = ~pi005 & ~n576;
  assign po204 = ~n2386 & ~n2387;
  assign n2389 = po119 & ~po204;
  assign n2390 = ~n2381 & po204;
  assign n2391 = ~n2375 & n2390;
  assign n2392 = ~n2389 & ~n2391;
  assign n2393 = ~n592 & ~n1701;
  assign n2394 = n592 & ~n1010;
  assign n2395 = ~n2393 & ~n2394;
  assign n2396 = ~pi193 & ~n2395;
  assign n2397 = n576 & ~n1211;
  assign n2398 = ~n620 & ~n1204;
  assign n2399 = n611 & ~n1193;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = ~n2397 & n2400;
  assign n2402 = pi193 & ~n2401;
  assign po155 = n2396 | n2402;
  assign n2404 = po216 & ~po155;
  assign n2405 = ~po216 & po155;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = ~n592 & ~n1070;
  assign n2408 = n592 & ~n1047;
  assign n2409 = ~n2407 & ~n2408;
  assign n2410 = ~pi193 & ~n2409;
  assign n2411 = n611 & n1097;
  assign n2412 = n576 & ~n1077;
  assign n2413 = ~n620 & ~n1063;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = ~n2411 & n2414;
  assign n2416 = pi193 & ~n2415;
  assign po147 = n2410 | n2416;
  assign n2418 = ~po209 & po147;
  assign n2419 = po209 & ~n2410;
  assign n2420 = ~n2416 & n2419;
  assign n2421 = ~n2418 & ~n2420;
  assign n2422 = ~n2406 & n2421;
  assign n2423 = n2392 & n2422;
  assign n2424 = ~n2371 & n2423;
  assign n2425 = ~n2406 & ~n2421;
  assign n2426 = ~n2392 & n2425;
  assign n2427 = ~n2371 & n2426;
  assign n2428 = ~n2424 & ~n2427;
  assign n2429 = n2351 & ~n2428;
  assign n2430 = n2406 & ~n2421;
  assign n2431 = n2392 & n2430;
  assign n2432 = n2371 & n2422;
  assign n2433 = ~n2392 & n2432;
  assign n2434 = ~n2431 & ~n2433;
  assign n2435 = n2351 & ~n2434;
  assign n2436 = ~n2429 & ~n2435;
  assign n2437 = ~n2371 & n2431;
  assign n2438 = n2371 & n2392;
  assign n2439 = n2421 & n2438;
  assign n2440 = ~n2406 & n2439;
  assign n2441 = ~n2437 & ~n2440;
  assign n2442 = ~n2371 & n2425;
  assign n2443 = n2351 & n2442;
  assign n2444 = n2406 & n2421;
  assign n2445 = ~n2392 & n2444;
  assign n2446 = n2351 & n2445;
  assign n2447 = ~n2371 & n2444;
  assign n2448 = n2371 & ~n2406;
  assign n2449 = ~n2421 & n2448;
  assign n2450 = ~n2447 & ~n2449;
  assign n2451 = ~n2351 & ~n2450;
  assign n2452 = ~n2446 & ~n2451;
  assign n2453 = ~n2443 & n2452;
  assign n2454 = n2441 & n2453;
  assign n2455 = n592 & ~n1186;
  assign n2456 = ~n592 & ~n1154;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~pi193 & ~n2457;
  assign n2459 = n611 & ~n1137;
  assign n2460 = ~n620 & ~n1130;
  assign n2461 = ~n2459 & ~n2460;
  assign n2462 = n576 & ~n1161;
  assign n2463 = n2461 & ~n2462;
  assign n2464 = pi193 & ~n2463;
  assign po111 = n2458 | n2464;
  assign n2466 = po195 & po111;
  assign n2467 = ~po195 & ~po111;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = ~n2454 & ~n2468;
  assign n2470 = n2436 & ~n2469;
  assign n2471 = ~n2351 & n2392;
  assign n2472 = n2442 & n2471;
  assign n2473 = n2438 & n2444;
  assign n2474 = ~n2422 & ~n2430;
  assign n2475 = ~n2392 & ~n2474;
  assign n2476 = ~n2473 & ~n2475;
  assign n2477 = ~n2351 & ~n2476;
  assign n2478 = n2371 & n2430;
  assign n2479 = ~n2392 & n2478;
  assign n2480 = ~n2477 & ~n2479;
  assign n2481 = ~n2472 & n2480;
  assign n2482 = n2392 & ~n2421;
  assign n2483 = n2371 & n2482;
  assign n2484 = ~n2447 & ~n2483;
  assign n2485 = n2351 & ~n2484;
  assign n2486 = n2481 & ~n2485;
  assign n2487 = n2468 & ~n2486;
  assign n2488 = ~n2351 & n2478;
  assign n2489 = ~n2392 & n2488;
  assign n2490 = ~n2371 & n2445;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = ~n2487 & n2491;
  assign n2493 = n2470 & n2492;
  assign n2494 = ~pi138 & ~pi192;
  assign n2495 = pi192 & pi220;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = n576 & n2496;
  assign n2498 = pi138 & ~n576;
  assign n2499 = ~n2497 & ~n2498;
  assign n2500 = ~n2493 & n2499;
  assign n2501 = ~n2489 & ~n2499;
  assign n2502 = ~n2490 & n2501;
  assign n2503 = n2470 & ~n2487;
  assign n2504 = n2502 & n2503;
  assign po080 = n2500 | n2504;
  assign n2506 = ~pi127 & ~pi192;
  assign n2507 = pi192 & pi196;
  assign n2508 = ~n2506 & ~n2507;
  assign n2509 = n576 & n2508;
  assign n2510 = pi127 & ~n576;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = ~n991 & ~n1174;
  assign n2513 = n1940 & n2512;
  assign n2514 = n991 & n1119;
  assign n2515 = ~n1250 & ~n2514;
  assign n2516 = n1256 & ~n2515;
  assign n2517 = ~n1932 & ~n1941;
  assign n2518 = ~n1939 & ~n1965;
  assign n2519 = n1174 & ~n2518;
  assign n2520 = n2517 & ~n2519;
  assign n2521 = n1224 & ~n2520;
  assign n2522 = n1122 & n1174;
  assign n2523 = ~n991 & n1119;
  assign n2524 = ~n1970 & ~n2523;
  assign n2525 = ~n1174 & ~n2524;
  assign n2526 = ~n2522 & ~n2525;
  assign n2527 = ~n1238 & ~n1918;
  assign n2528 = n2526 & n2527;
  assign n2529 = ~n1224 & ~n2528;
  assign n2530 = ~n2521 & ~n2529;
  assign n2531 = ~n2516 & n2530;
  assign n2532 = ~n2513 & n2531;
  assign n2533 = ~n1229 & ~n1977;
  assign n2534 = ~n1041 & ~n1118;
  assign n2535 = n1041 & ~n1175;
  assign n2536 = n1911 & ~n2535;
  assign n2537 = ~n2534 & n2536;
  assign n2538 = n1174 & n1917;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = n2533 & n2539;
  assign n2541 = n2532 & n2540;
  assign n2542 = ~n2511 & ~n2541;
  assign n2543 = ~n2516 & n2539;
  assign n2544 = ~n2521 & n2543;
  assign n2545 = ~n2529 & n2544;
  assign n2546 = ~n1229 & ~n2513;
  assign n2547 = ~n1977 & n2546;
  assign n2548 = n2511 & n2547;
  assign n2549 = n2545 & n2548;
  assign po081 = n2542 | n2549;
  assign n2551 = ~n1849 & ~n1852;
  assign n2552 = n1755 & ~n2551;
  assign n2553 = ~n1801 & n2552;
  assign n2554 = n1801 & n1866;
  assign n2555 = n1735 & n2554;
  assign n2556 = ~n2553 & ~n2555;
  assign n2557 = ~n1735 & ~n1755;
  assign n2558 = ~n2551 & n2557;
  assign n2559 = ~n1831 & ~n1866;
  assign n2560 = ~n1755 & ~n2559;
  assign n2561 = n1735 & n2560;
  assign n2562 = ~n2558 & ~n2561;
  assign n2563 = n2556 & n2562;
  assign n2564 = ~n1715 & ~n2563;
  assign n2565 = n1735 & n1852;
  assign n2566 = ~n1735 & n1802;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = ~n1850 & n2567;
  assign n2569 = n1715 & ~n1755;
  assign n2570 = ~n2568 & n2569;
  assign n2571 = n1801 & n1849;
  assign n2572 = ~n1832 & ~n1845;
  assign n2573 = ~n2571 & n2572;
  assign n2574 = n1755 & ~n2573;
  assign n2575 = n1801 & ~n2551;
  assign n2576 = n1735 & n2575;
  assign n2577 = ~n2574 & ~n2576;
  assign n2578 = n1715 & ~n2577;
  assign n2579 = ~n2570 & ~n2578;
  assign n2580 = ~n2564 & n2579;
  assign n2581 = ~n1801 & n1852;
  assign n2582 = ~n2554 & ~n2581;
  assign n2583 = n1847 & ~n2582;
  assign n2584 = ~n1735 & n1877;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = n2580 & n2585;
  assign n2587 = ~pi146 & ~pi192;
  assign n2588 = pi192 & pi254;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = n576 & n2589;
  assign n2591 = pi146 & ~n576;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = ~n2586 & ~n2592;
  assign n2594 = n2585 & n2592;
  assign n2595 = n2579 & n2594;
  assign n2596 = ~n2564 & n2595;
  assign po082 = n2593 | n2596;
  assign n2598 = ~n592 & ~n870;
  assign n2599 = n592 & ~n1401;
  assign n2600 = ~n2598 & ~n2599;
  assign n2601 = ~pi193 & ~n2600;
  assign n2602 = n598 & n611;
  assign n2603 = n576 & ~n863;
  assign n2604 = ~n620 & ~n851;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = ~n2602 & n2605;
  assign n2607 = pi193 & ~n2606;
  assign po121 = n2601 | n2607;
  assign n2609 = ~po217 & po121;
  assign n2610 = po217 & ~po121;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = ~n592 & n684;
  assign n2613 = n592 & ~n669;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = ~pi193 & ~n2614;
  assign n2616 = n576 & ~n785;
  assign n2617 = ~n620 & ~n778;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = n611 & ~n761;
  assign n2620 = n2618 & ~n2619;
  assign n2621 = pi193 & ~n2620;
  assign po132 = n2615 | n2621;
  assign n2623 = pi009 & ~n576;
  assign n2624 = pi009 & ~pi192;
  assign n2625 = pi192 & pi243;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = n576 & ~n2626;
  assign po198 = n2623 | n2627;
  assign n2629 = po132 & ~po198;
  assign n2630 = ~po132 & po198;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = n592 & ~n798;
  assign n2633 = ~n592 & ~n813;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = ~pi193 & ~n2634;
  assign n2636 = n576 & ~n734;
  assign n2637 = ~n620 & ~n727;
  assign n2638 = n611 & ~n717;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~n2636 & n2639;
  assign n2641 = pi193 & ~n2640;
  assign po151 = n2635 | n2641;
  assign n2643 = ~po218 & ~po151;
  assign n2644 = po218 & po151;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = n611 & ~n660;
  assign n2647 = n576 & ~n703;
  assign n2648 = ~n620 & ~n653;
  assign n2649 = ~n2647 & ~n2648;
  assign n2650 = ~n2646 & n2649;
  assign n2651 = pi193 & ~n2650;
  assign n2652 = ~n592 & ~n710;
  assign n2653 = n592 & ~n717;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = ~pi193 & ~n2654;
  assign po146 = n2651 | n2655;
  assign n2657 = po223 & ~po146;
  assign n2658 = ~po223 & po146;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = ~n2645 & ~n2659;
  assign n2661 = ~n2631 & n2660;
  assign n2662 = ~n2645 & n2659;
  assign n2663 = n2631 & n2662;
  assign n2664 = ~n2661 & ~n2663;
  assign n2665 = ~n2611 & ~n2664;
  assign n2666 = n576 & ~n754;
  assign n2667 = ~n620 & ~n1401;
  assign n2668 = n611 & ~n870;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = ~n2666 & n2669;
  assign n2671 = pi193 & ~n2670;
  assign n2672 = n592 & ~n761;
  assign n2673 = ~n592 & n768;
  assign n2674 = ~n2672 & ~n2673;
  assign n2675 = ~pi193 & ~n2674;
  assign po113 = n2671 | n2675;
  assign n2677 = ~po199 & ~po113;
  assign n2678 = po199 & po113;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = n2645 & ~n2659;
  assign n2681 = ~n2611 & n2631;
  assign n2682 = n2680 & n2681;
  assign n2683 = n576 & ~n823;
  assign n2684 = n611 & ~n798;
  assign n2685 = ~n620 & ~n805;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = ~n2683 & n2686;
  assign n2688 = pi193 & ~n2687;
  assign n2689 = n592 & ~n626;
  assign n2690 = ~n592 & ~n617;
  assign n2691 = ~n2689 & ~n2690;
  assign n2692 = ~pi193 & ~n2691;
  assign po140 = n2688 | n2692;
  assign n2694 = pi018 & ~n576;
  assign n2695 = pi018 & ~pi192;
  assign n2696 = pi192 & pi235;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = n576 & ~n2697;
  assign po196 = n2694 | n2698;
  assign n2700 = ~po140 & po196;
  assign n2701 = po140 & ~po196;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = n2645 & n2659;
  assign n2704 = n2702 & n2703;
  assign n2705 = n2631 & n2704;
  assign n2706 = ~n2631 & n2702;
  assign n2707 = ~n2659 & n2706;
  assign n2708 = ~n2645 & n2702;
  assign n2709 = ~n2659 & n2708;
  assign n2710 = ~n2707 & ~n2709;
  assign n2711 = n2611 & ~n2710;
  assign n2712 = ~n2631 & ~n2702;
  assign n2713 = n2703 & n2712;
  assign n2714 = ~n2711 & ~n2713;
  assign n2715 = ~n2705 & n2714;
  assign n2716 = ~n2682 & n2715;
  assign n2717 = ~n2679 & ~n2716;
  assign n2718 = n2659 & ~n2702;
  assign n2719 = n2631 & n2718;
  assign n2720 = n2660 & ~n2702;
  assign n2721 = ~n2719 & ~n2720;
  assign n2722 = ~n2611 & ~n2721;
  assign n2723 = n2645 & n2706;
  assign n2724 = n2659 & n2723;
  assign n2725 = ~n2659 & ~n2702;
  assign n2726 = n2645 & n2725;
  assign n2727 = ~n2631 & n2726;
  assign n2728 = ~n2724 & ~n2727;
  assign n2729 = n2611 & n2680;
  assign n2730 = n2631 & n2729;
  assign n2731 = n2728 & ~n2730;
  assign n2732 = ~n2722 & n2731;
  assign n2733 = n2679 & ~n2732;
  assign n2734 = ~n2717 & ~n2733;
  assign n2735 = ~n2665 & n2734;
  assign n2736 = n2631 & n2726;
  assign n2737 = ~n2705 & ~n2736;
  assign n2738 = n2662 & ~n2702;
  assign n2739 = n2737 & ~n2738;
  assign n2740 = n2611 & ~n2739;
  assign n2741 = ~n2645 & n2706;
  assign n2742 = ~n2659 & n2741;
  assign n2743 = ~n2740 & ~n2742;
  assign n2744 = n2735 & n2743;
  assign n2745 = ~pi125 & ~pi192;
  assign n2746 = pi192 & pi246;
  assign n2747 = ~n2745 & ~n2746;
  assign n2748 = n576 & n2747;
  assign n2749 = pi125 & ~n576;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = ~n2744 & ~n2750;
  assign n2752 = n2743 & n2750;
  assign n2753 = n2734 & n2752;
  assign n2754 = ~n2665 & n2753;
  assign po083 = n2751 | n2754;
  assign n2756 = ~pi135 & ~pi192;
  assign n2757 = pi192 & pi206;
  assign n2758 = ~n2756 & ~n2757;
  assign n2759 = n576 & n2758;
  assign n2760 = pi135 & ~n576;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = ~n2351 & ~n2468;
  assign n2763 = ~n2371 & n2421;
  assign n2764 = ~n2392 & n2763;
  assign n2765 = ~n2478 & ~n2764;
  assign n2766 = n2762 & ~n2765;
  assign n2767 = ~n2371 & n2430;
  assign n2768 = ~n2392 & n2767;
  assign n2769 = ~n2433 & ~n2768;
  assign n2770 = ~n2425 & ~n2444;
  assign n2771 = n2392 & ~n2770;
  assign n2772 = n2769 & ~n2771;
  assign n2773 = n2351 & ~n2772;
  assign n2774 = ~n2371 & n2392;
  assign n2775 = n2421 & n2774;
  assign n2776 = n2406 & n2775;
  assign n2777 = ~n2773 & ~n2776;
  assign n2778 = ~n2468 & ~n2777;
  assign n2779 = ~n2766 & ~n2778;
  assign n2780 = n2371 & n2426;
  assign n2781 = ~n2440 & ~n2780;
  assign n2782 = ~n2445 & n2781;
  assign n2783 = ~n2351 & ~n2782;
  assign n2784 = ~n2351 & n2432;
  assign n2785 = ~n2427 & ~n2784;
  assign n2786 = ~n2351 & n2431;
  assign n2787 = ~n2371 & n2422;
  assign n2788 = ~n2478 & ~n2787;
  assign n2789 = n2351 & ~n2788;
  assign n2790 = ~n2786 & ~n2789;
  assign n2791 = n2371 & n2445;
  assign n2792 = n2790 & ~n2791;
  assign n2793 = n2785 & n2792;
  assign n2794 = n2468 & ~n2793;
  assign n2795 = ~n2783 & ~n2794;
  assign n2796 = n2351 & n2392;
  assign n2797 = n2447 & n2796;
  assign n2798 = n2371 & n2431;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = ~n2472 & n2799;
  assign n2801 = n2795 & n2800;
  assign n2802 = n2779 & n2801;
  assign n2803 = ~n2761 & ~n2802;
  assign n2804 = n2779 & n2795;
  assign n2805 = n2800 & n2804;
  assign n2806 = n2761 & n2805;
  assign po084 = n2803 | n2806;
  assign n2808 = ~n1449 & ~n1619;
  assign n2809 = ~n1383 & ~n2808;
  assign n2810 = n1360 & n1418;
  assign n2811 = ~n1416 & ~n2810;
  assign n2812 = n1433 & ~n2811;
  assign n2813 = ~n1383 & n2812;
  assign n2814 = ~n1453 & ~n1589;
  assign n2815 = n1320 & n1383;
  assign n2816 = ~n1360 & ~n1411;
  assign n2817 = ~n1340 & n1411;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = n2815 & ~n2818;
  assign n2820 = ~n1320 & ~n1383;
  assign n2821 = n1656 & ~n2820;
  assign n2822 = ~n2819 & ~n2821;
  assign n2823 = ~n1428 & n2822;
  assign n2824 = n1433 & ~n2823;
  assign n2825 = n1385 & n1593;
  assign n2826 = ~n1595 & ~n2825;
  assign n2827 = n1383 & ~n2826;
  assign n2828 = ~n2824 & ~n2827;
  assign n2829 = n2814 & n2828;
  assign n2830 = ~n2813 & n2829;
  assign n2831 = ~n2809 & n2830;
  assign n2832 = n1360 & ~n1411;
  assign n2833 = ~n1416 & ~n2832;
  assign n2834 = n1383 & ~n2833;
  assign n2835 = ~n1412 & ~n1662;
  assign n2836 = ~n1383 & n1663;
  assign n2837 = n2835 & ~n2836;
  assign n2838 = ~n2834 & n2837;
  assign n2839 = n1300 & ~n2838;
  assign n2840 = n2831 & ~n2839;
  assign n2841 = ~pi152 & ~pi192;
  assign n2842 = pi192 & pi194;
  assign n2843 = ~n2841 & ~n2842;
  assign n2844 = n576 & n2843;
  assign n2845 = pi152 & ~n576;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = ~n2840 & ~n2846;
  assign n2848 = ~n2839 & n2846;
  assign n2849 = n2830 & n2848;
  assign n2850 = ~n2809 & n2849;
  assign po085 = n2847 | n2850;
  assign n2852 = ~pi128 & ~pi192;
  assign n2853 = pi192 & pi234;
  assign n2854 = ~n2852 & ~n2853;
  assign n2855 = n576 & n2854;
  assign n2856 = pi128 & ~n576;
  assign n2857 = ~n2855 & ~n2856;
  assign n2858 = ~n1735 & ~n1801;
  assign n2859 = ~n2571 & ~n2858;
  assign n2860 = n1781 & ~n1801;
  assign n2861 = ~n2565 & ~n2860;
  assign n2862 = n2859 & n2861;
  assign n2863 = n1755 & ~n2862;
  assign n2864 = n1735 & n2581;
  assign n2865 = ~n2863 & ~n2864;
  assign n2866 = n1735 & n1866;
  assign n2867 = ~n1860 & ~n2866;
  assign n2868 = ~n1850 & n2867;
  assign n2869 = ~n1755 & ~n2868;
  assign n2870 = n2865 & ~n2869;
  assign n2871 = ~n1715 & ~n2870;
  assign n2872 = ~n1881 & ~n2571;
  assign n2873 = n1830 & n1840;
  assign n2874 = ~n1735 & n1830;
  assign n2875 = ~n1801 & n2874;
  assign n2876 = ~n2873 & ~n2875;
  assign n2877 = n2872 & n2876;
  assign n2878 = n2569 & ~n2877;
  assign n2879 = n1735 & n1865;
  assign n2880 = ~n1802 & ~n1877;
  assign n2881 = n2879 & ~n2880;
  assign n2882 = ~n2878 & ~n2881;
  assign n2883 = ~n2871 & n2882;
  assign n2884 = ~n1849 & ~n2860;
  assign n2885 = ~n1735 & ~n2884;
  assign n2886 = ~n2581 & ~n2885;
  assign n2887 = n1755 & ~n2886;
  assign n2888 = ~n1755 & n2584;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = n2883 & n2889;
  assign n2891 = ~n2857 & ~n2890;
  assign n2892 = n2857 & n2889;
  assign n2893 = n2882 & n2892;
  assign n2894 = ~n2871 & n2893;
  assign po086 = n2891 | n2894;
  assign n2896 = ~pi151 & ~pi192;
  assign n2897 = pi192 & pi208;
  assign n2898 = ~n2896 & ~n2897;
  assign n2899 = n576 & n2898;
  assign n2900 = pi151 & ~n576;
  assign n2901 = ~n2899 & ~n2900;
  assign n2902 = ~n2065 & ~n2085;
  assign n2903 = ~n2045 & n2902;
  assign n2904 = n2101 & n2903;
  assign n2905 = ~n2101 & n2133;
  assign n2906 = n2107 & n2142;
  assign n2907 = n2065 & n2105;
  assign n2908 = ~n2906 & ~n2907;
  assign n2909 = ~n2905 & n2908;
  assign n2910 = ~n2904 & n2909;
  assign n2911 = n2031 & ~n2910;
  assign n2912 = n2031 & n2106;
  assign n2913 = ~n2153 & ~n2912;
  assign n2914 = n2017 & ~n2913;
  assign n2915 = n2065 & n2156;
  assign n2916 = ~n2065 & n2128;
  assign n2917 = ~n2108 & ~n2916;
  assign n2918 = ~n2154 & n2917;
  assign n2919 = ~n2915 & n2918;
  assign n2920 = n2017 & ~n2919;
  assign n2921 = n2017 & n2103;
  assign n2922 = ~n2147 & ~n2921;
  assign n2923 = ~n2920 & n2922;
  assign n2924 = ~n2031 & ~n2923;
  assign n2925 = ~n2914 & ~n2924;
  assign n2926 = n2086 & n2128;
  assign n2927 = n2085 & n2128;
  assign n2928 = ~n2131 & ~n2927;
  assign n2929 = n2031 & ~n2928;
  assign n2930 = ~n2926 & ~n2929;
  assign n2931 = ~n2017 & ~n2930;
  assign n2932 = ~n2017 & ~n2031;
  assign n2933 = ~n2085 & ~n2101;
  assign n2934 = n2045 & n2142;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n2932 & ~n2935;
  assign n2937 = ~n2931 & ~n2936;
  assign n2938 = ~n2135 & n2937;
  assign n2939 = n2925 & n2938;
  assign n2940 = ~n2911 & n2939;
  assign n2941 = ~n2901 & ~n2940;
  assign n2942 = n2901 & ~n2911;
  assign n2943 = n2925 & n2942;
  assign n2944 = n2938 & n2943;
  assign po087 = n2941 | n2944;
  assign n2946 = n2179 & ~n2268;
  assign n2947 = n2199 & n2213;
  assign n2948 = ~n2249 & n2947;
  assign n2949 = ~n2258 & ~n2292;
  assign n2950 = ~n2263 & ~n2266;
  assign n2951 = n2949 & n2950;
  assign n2952 = n2179 & ~n2951;
  assign n2953 = ~n2948 & ~n2952;
  assign n2954 = n2285 & ~n2953;
  assign n2955 = ~n2305 & ~n2947;
  assign n2956 = ~n2319 & n2955;
  assign n2957 = n2315 & ~n2956;
  assign n2958 = ~n2954 & ~n2957;
  assign n2959 = ~n2946 & n2958;
  assign n2960 = ~n2249 & ~n2291;
  assign n2961 = ~n2321 & n2960;
  assign n2962 = ~n2265 & n2961;
  assign n2963 = ~n2199 & n2228;
  assign n2964 = n2249 & ~n2963;
  assign n2965 = ~n2179 & ~n2964;
  assign n2966 = ~n2962 & n2965;
  assign n2967 = ~n2199 & ~n2249;
  assign n2968 = n2213 & n2967;
  assign n2969 = ~n2227 & n2968;
  assign n2970 = ~n2319 & ~n2969;
  assign n2971 = n2179 & ~n2970;
  assign n2972 = n2227 & n2287;
  assign n2973 = ~n2251 & ~n2972;
  assign n2974 = n2179 & ~n2973;
  assign n2975 = ~n2971 & ~n2974;
  assign n2976 = ~n2966 & n2975;
  assign n2977 = ~n2300 & n2976;
  assign n2978 = ~n2285 & ~n2977;
  assign n2979 = ~n2179 & ~n2304;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = n2959 & n2980;
  assign n2982 = ~pi155 & ~pi192;
  assign n2983 = pi192 & pi226;
  assign n2984 = ~n2982 & ~n2983;
  assign n2985 = n576 & n2984;
  assign n2986 = pi155 & ~n576;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = ~n2981 & n2987;
  assign n2989 = n2959 & ~n2987;
  assign n2990 = n2980 & n2989;
  assign po088 = n2988 | n2990;
  assign n2992 = ~n2065 & n2105;
  assign n2993 = n2065 & n2114;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~n2031 & ~n2994;
  assign n2996 = ~n2127 & ~n2907;
  assign n2997 = n2928 & n2996;
  assign n2998 = n2017 & ~n2997;
  assign n2999 = n2031 & n2998;
  assign n3000 = ~n2065 & n2114;
  assign n3001 = ~n2134 & ~n3000;
  assign n3002 = n2031 & ~n3001;
  assign n3003 = ~n2031 & ~n2065;
  assign n3004 = n2128 & n3003;
  assign n3005 = ~n2031 & n2065;
  assign n3006 = n2107 & n3005;
  assign n3007 = ~n3004 & ~n3006;
  assign n3008 = ~n2157 & n3007;
  assign n3009 = n2017 & ~n3008;
  assign n3010 = ~n3002 & ~n3009;
  assign n3011 = ~n2999 & n3010;
  assign n3012 = ~n2122 & n3011;
  assign n3013 = ~n2995 & n3012;
  assign n3014 = n2128 & n2151;
  assign n3015 = ~n2108 & ~n2117;
  assign n3016 = n2065 & ~n3015;
  assign n3017 = n2031 & n3016;
  assign n3018 = ~n2129 & ~n2139;
  assign n3019 = n2045 & n2902;
  assign n3020 = n3018 & ~n3019;
  assign n3021 = ~n2031 & ~n3020;
  assign n3022 = ~n2147 & ~n3021;
  assign n3023 = ~n3017 & n3022;
  assign n3024 = ~n3014 & n3023;
  assign n3025 = ~n2017 & ~n3024;
  assign n3026 = n3013 & ~n3025;
  assign n3027 = ~pi150 & ~pi192;
  assign n3028 = pi192 & pi218;
  assign n3029 = ~n3027 & ~n3028;
  assign n3030 = n576 & n3029;
  assign n3031 = pi150 & ~n576;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = ~n3026 & ~n3032;
  assign n3034 = ~n3025 & n3032;
  assign n3035 = n3012 & n3034;
  assign n3036 = ~n2995 & n3035;
  assign po089 = n3033 | n3036;
  assign n3038 = ~pi137 & ~pi192;
  assign n3039 = pi192 & pi240;
  assign n3040 = ~n3038 & ~n3039;
  assign n3041 = n576 & n3040;
  assign n3042 = pi137 & ~n576;
  assign n3043 = ~n3041 & ~n3042;
  assign n3044 = n1735 & n2571;
  assign n3045 = ~n1845 & ~n3044;
  assign n3046 = ~n1755 & ~n3045;
  assign n3047 = ~n1801 & n1866;
  assign n3048 = ~n1832 & ~n2575;
  assign n3049 = ~n3047 & n3048;
  assign n3050 = n2569 & ~n3049;
  assign n3051 = ~n1735 & n1831;
  assign n3052 = ~n2565 & ~n3051;
  assign n3053 = ~n2554 & n3052;
  assign n3054 = n1755 & ~n3053;
  assign n3055 = n1735 & n1850;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = n1715 & ~n3056;
  assign n3058 = ~n3050 & ~n3057;
  assign n3059 = ~n3046 & n3058;
  assign n3060 = ~n1877 & ~n2581;
  assign n3061 = ~n1755 & ~n3060;
  assign n3062 = ~n1850 & ~n2554;
  assign n3063 = ~n1755 & ~n3062;
  assign n3064 = ~n1735 & n3063;
  assign n3065 = ~n3061 & ~n3064;
  assign n3066 = ~n1715 & ~n3065;
  assign n3067 = n1735 & n1755;
  assign n3068 = n2554 & n3067;
  assign n3069 = ~n1715 & n1755;
  assign n3070 = ~n1868 & ~n2875;
  assign n3071 = ~n1874 & n3070;
  assign n3072 = n3069 & ~n3071;
  assign n3073 = ~n3068 & ~n3072;
  assign n3074 = ~n3066 & n3073;
  assign n3075 = n3059 & n3074;
  assign n3076 = ~n3043 & ~n3075;
  assign n3077 = n3058 & n3074;
  assign n3078 = n3043 & n3077;
  assign n3079 = ~n3046 & n3078;
  assign po090 = n3076 | n3079;
  assign n3081 = ~pi131 & ~pi192;
  assign n3082 = pi192 & pi200;
  assign n3083 = ~n3081 & ~n3082;
  assign n3084 = n576 & n3083;
  assign n3085 = pi131 & ~n576;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = n2371 & n2406;
  assign n3088 = ~n2392 & n3087;
  assign n3089 = ~n2787 & ~n3088;
  assign n3090 = n2351 & ~n3089;
  assign n3091 = ~n2427 & ~n3090;
  assign n3092 = ~n2433 & ~n2437;
  assign n3093 = ~n2351 & ~n3092;
  assign n3094 = n3091 & ~n3093;
  assign n3095 = n2351 & n2421;
  assign n3096 = ~n2371 & n3095;
  assign n3097 = n2392 & n3096;
  assign n3098 = ~n2798 & ~n3097;
  assign n3099 = ~n2426 & ~n2445;
  assign n3100 = ~n2442 & n3099;
  assign n3101 = ~n2351 & ~n3100;
  assign n3102 = n3098 & ~n3101;
  assign n3103 = ~n2784 & n3102;
  assign n3104 = ~n2468 & ~n3103;
  assign n3105 = n3094 & ~n3104;
  assign n3106 = ~n2423 & n3099;
  assign n3107 = n2351 & ~n3106;
  assign n3108 = n2371 & n2771;
  assign n3109 = ~n2767 & ~n3108;
  assign n3110 = ~n2351 & ~n3109;
  assign n3111 = ~n2423 & ~n2431;
  assign n3112 = ~n2371 & ~n3111;
  assign n3113 = ~n3110 & ~n3112;
  assign n3114 = ~n3107 & n3113;
  assign n3115 = n2468 & ~n3114;
  assign n3116 = n3105 & ~n3115;
  assign n3117 = n3086 & ~n3116;
  assign n3118 = n3094 & ~n3115;
  assign n3119 = ~n3086 & n3118;
  assign n3120 = ~n3104 & n3119;
  assign po091 = n3117 | n3120;
  assign n3122 = n2631 & n2709;
  assign n3123 = n2631 & n2738;
  assign n3124 = ~n3122 & ~n3123;
  assign n3125 = ~n2704 & n3124;
  assign n3126 = ~n2611 & ~n3125;
  assign n3127 = ~n2709 & ~n2726;
  assign n3128 = ~n2611 & ~n3127;
  assign n3129 = ~n2611 & ~n2631;
  assign n3130 = n2703 & n3129;
  assign n3131 = ~n3128 & ~n3130;
  assign n3132 = n2679 & ~n3131;
  assign n3133 = n2631 & n2702;
  assign n3134 = n2662 & n3133;
  assign n3135 = ~n2631 & ~n2645;
  assign n3136 = ~n2702 & n3135;
  assign n3137 = n2659 & n3136;
  assign n3138 = ~n3134 & ~n3137;
  assign n3139 = n2611 & ~n3138;
  assign n3140 = n2663 & n2679;
  assign n3141 = n2702 & n3140;
  assign n3142 = ~n2736 & ~n3141;
  assign n3143 = ~n3139 & n3142;
  assign n3144 = ~n3132 & n3143;
  assign n3145 = ~n3126 & n3144;
  assign n3146 = ~n2645 & ~n2702;
  assign n3147 = n2611 & n3146;
  assign n3148 = ~n2631 & n3147;
  assign n3149 = ~n2662 & ~n2680;
  assign n3150 = n2611 & ~n3149;
  assign n3151 = n2702 & n3150;
  assign n3152 = ~n3148 & ~n3151;
  assign n3153 = n2679 & ~n3152;
  assign n3154 = ~n2631 & n3146;
  assign n3155 = ~n2723 & ~n3154;
  assign n3156 = ~n2611 & ~n2679;
  assign n3157 = ~n3155 & n3156;
  assign n3158 = n2631 & n2725;
  assign n3159 = n2631 & n2703;
  assign n3160 = ~n3158 & ~n3159;
  assign n3161 = ~n2742 & n3160;
  assign n3162 = ~n2726 & n3161;
  assign n3163 = n2611 & ~n3162;
  assign n3164 = ~n2679 & n3163;
  assign n3165 = ~n3157 & ~n3164;
  assign n3166 = ~n3153 & n3165;
  assign n3167 = n3145 & n3166;
  assign n3168 = ~pi140 & ~pi192;
  assign n3169 = pi192 & pi228;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = n576 & n3170;
  assign n3172 = pi140 & ~n576;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3167 & ~n3173;
  assign n3175 = n3145 & n3173;
  assign n3176 = n3166 & n3175;
  assign po092 = n3174 | n3176;
  assign n3178 = ~pi141 & ~pi192;
  assign n3179 = pi192 & pi222;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = n576 & n3180;
  assign n3182 = pi141 & ~n576;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = n792 & n894;
  assign n3185 = n877 & n3184;
  assign n3186 = ~n837 & ~n877;
  assign n3187 = ~n891 & ~n3186;
  assign n3188 = ~n792 & ~n3187;
  assign n3189 = ~n885 & ~n3188;
  assign n3190 = n641 & ~n3189;
  assign n3191 = ~n3185 & ~n3190;
  assign n3192 = n886 & n1547;
  assign n3193 = ~n691 & n3192;
  assign n3194 = ~n1549 & ~n3193;
  assign n3195 = n641 & ~n3194;
  assign n3196 = n3191 & ~n3195;
  assign n3197 = ~n1486 & n1532;
  assign n3198 = ~n792 & ~n3197;
  assign n3199 = ~n1499 & ~n3198;
  assign n3200 = ~n641 & ~n3199;
  assign n3201 = ~n884 & ~n891;
  assign n3202 = ~n914 & n3201;
  assign n3203 = n792 & ~n3202;
  assign n3204 = ~n641 & n3203;
  assign n3205 = ~n792 & n880;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = ~n3200 & n3206;
  assign n3208 = ~n1528 & n3207;
  assign n3209 = n3196 & n3208;
  assign n3210 = ~n3183 & ~n3209;
  assign n3211 = n3183 & n3209;
  assign po093 = n3210 | n3211;
  assign n3213 = ~pi157 & ~pi192;
  assign n3214 = pi192 & pi202;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = n576 & n3215;
  assign n3217 = pi157 & ~n576;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = ~n2426 & n3111;
  assign n3220 = ~n2351 & ~n3219;
  assign n3221 = n2371 & n2444;
  assign n3222 = ~n2371 & n2475;
  assign n3223 = ~n3221 & ~n3222;
  assign n3224 = n2351 & ~n3223;
  assign n3225 = n2371 & ~n3099;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = ~n3220 & n3226;
  assign n3228 = ~n2468 & ~n3227;
  assign n3229 = ~n2371 & n2406;
  assign n3230 = n2392 & n3229;
  assign n3231 = ~n2449 & ~n3230;
  assign n3232 = ~n2351 & ~n3231;
  assign n3233 = n2371 & ~n2421;
  assign n3234 = ~n2351 & n3233;
  assign n3235 = ~n2392 & n3234;
  assign n3236 = ~n2490 & ~n3235;
  assign n3237 = ~n2432 & ~n2442;
  assign n3238 = n3111 & n3237;
  assign n3239 = n2351 & ~n3238;
  assign n3240 = n3236 & ~n3239;
  assign n3241 = n2468 & ~n3240;
  assign n3242 = ~n3232 & ~n3241;
  assign n3243 = n2442 & n2796;
  assign n3244 = n2351 & n2371;
  assign n3245 = n2445 & n3244;
  assign n3246 = ~n3243 & ~n3245;
  assign n3247 = ~n2440 & n3246;
  assign n3248 = n3242 & n3247;
  assign n3249 = ~n3228 & n3248;
  assign n3250 = n3218 & ~n3249;
  assign n3251 = ~n3228 & n3247;
  assign n3252 = n3242 & n3251;
  assign n3253 = ~n3218 & n3252;
  assign po094 = n3250 | n3253;
  assign n3255 = ~n2065 & n2117;
  assign n3256 = n2031 & n3255;
  assign n3257 = ~n2102 & ~n2139;
  assign n3258 = ~n2031 & ~n3257;
  assign n3259 = n2065 & ~n2101;
  assign n3260 = ~n2927 & ~n3259;
  assign n3261 = n2031 & ~n3260;
  assign n3262 = ~n2993 & ~n3261;
  assign n3263 = ~n3258 & n3262;
  assign n3264 = ~n3256 & n3263;
  assign n3265 = ~n2017 & ~n3264;
  assign n3266 = ~n2154 & ~n2906;
  assign n3267 = ~n2031 & ~n3266;
  assign n3268 = n2065 & n2927;
  assign n3269 = n2031 & n3268;
  assign n3270 = ~n3267 & ~n3269;
  assign n3271 = n2065 & n2154;
  assign n3272 = n2031 & n3019;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = ~n2031 & n2907;
  assign n3275 = ~n2127 & ~n3274;
  assign n3276 = ~n2157 & n3275;
  assign n3277 = ~n2115 & n3276;
  assign n3278 = n3273 & n3277;
  assign n3279 = n2017 & ~n3278;
  assign n3280 = n3270 & ~n3279;
  assign n3281 = ~n3265 & n3280;
  assign n3282 = ~pi143 & ~pi192;
  assign n3283 = pi192 & pi204;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = n576 & n3284;
  assign n3286 = pi143 & ~n576;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n3281 & ~n3287;
  assign n3289 = n3281 & n3287;
  assign po095 = n3288 | n3289;
  assign n3291 = ~n2179 & n2301;
  assign n3292 = n2228 & n2249;
  assign n3293 = ~n2295 & ~n3292;
  assign n3294 = ~n2320 & n3293;
  assign n3295 = n2315 & ~n3294;
  assign n3296 = ~n2199 & n2213;
  assign n3297 = ~n2249 & n2250;
  assign n3298 = ~n3296 & ~n3297;
  assign n3299 = n2179 & ~n3298;
  assign n3300 = ~n2322 & ~n3299;
  assign n3301 = n2285 & ~n3300;
  assign n3302 = ~n3295 & ~n3301;
  assign n3303 = ~n3291 & n3302;
  assign n3304 = n2249 & ~n2294;
  assign n3305 = ~n2302 & ~n2305;
  assign n3306 = ~n2300 & n3305;
  assign n3307 = ~n2179 & ~n3306;
  assign n3308 = ~n2249 & n2319;
  assign n3309 = n2249 & n2947;
  assign n3310 = n2199 & n2262;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = n2179 & ~n3311;
  assign n3313 = ~n3308 & ~n3312;
  assign n3314 = ~n3307 & n3313;
  assign n3315 = ~n3304 & n3314;
  assign n3316 = ~n2285 & ~n3315;
  assign n3317 = n2199 & n2249;
  assign n3318 = n2227 & n3317;
  assign n3319 = ~n2969 & ~n3318;
  assign n3320 = n2179 & ~n3319;
  assign n3321 = ~n3316 & ~n3320;
  assign n3322 = n3303 & n3321;
  assign n3323 = ~pi126 & ~pi192;
  assign n3324 = pi192 & pi224;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = n576 & n3325;
  assign n3327 = pi126 & ~n576;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = ~n3322 & ~n3328;
  assign n3330 = n3302 & n3321;
  assign n3331 = n3328 & n3330;
  assign n3332 = ~n3291 & n3331;
  assign po096 = n3329 | n3332;
  assign n3334 = ~pi144 & ~pi192;
  assign n3335 = pi192 & pi210;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = n576 & n3336;
  assign n3338 = pi144 & ~n576;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = n2611 & ~n2728;
  assign n3341 = ~n2680 & ~n3135;
  assign n3342 = n2702 & ~n3341;
  assign n3343 = ~n2719 & ~n3342;
  assign n3344 = n3156 & ~n3343;
  assign n3345 = ~n2704 & ~n2725;
  assign n3346 = ~n2631 & n2703;
  assign n3347 = ~n2663 & ~n3346;
  assign n3348 = n3345 & n3347;
  assign n3349 = n2611 & ~n3348;
  assign n3350 = ~n2631 & n2720;
  assign n3351 = ~n3349 & ~n3350;
  assign n3352 = ~n2679 & ~n3351;
  assign n3353 = ~n3344 & ~n3352;
  assign n3354 = ~n2702 & n3159;
  assign n3355 = ~n2709 & ~n3354;
  assign n3356 = n2611 & ~n3355;
  assign n3357 = n2611 & ~n2631;
  assign n3358 = n2662 & n3357;
  assign n3359 = n2659 & ~n2708;
  assign n3360 = n2631 & ~n3359;
  assign n3361 = ~n2611 & n3360;
  assign n3362 = ~n3130 & ~n3361;
  assign n3363 = ~n2659 & n3133;
  assign n3364 = ~n3137 & ~n3363;
  assign n3365 = n3362 & n3364;
  assign n3366 = ~n3358 & n3365;
  assign n3367 = ~n3356 & n3366;
  assign n3368 = n2679 & ~n3367;
  assign n3369 = n3353 & ~n3368;
  assign n3370 = ~n3340 & n3369;
  assign n3371 = ~n3339 & ~n3370;
  assign n3372 = n3339 & ~n3340;
  assign n3373 = ~n3368 & n3372;
  assign n3374 = n3353 & n3373;
  assign po097 = n3371 | n3374;
  assign n3376 = ~pi156 & ~pi192;
  assign n3377 = pi192 & pi232;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = n576 & n3378;
  assign n3380 = pi156 & ~n576;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = ~n2736 & ~n3154;
  assign n3383 = ~n2611 & ~n3382;
  assign n3384 = n2631 & ~n2702;
  assign n3385 = ~n2645 & n3384;
  assign n3386 = ~n2659 & n3385;
  assign n3387 = ~n2742 & ~n3386;
  assign n3388 = ~n2705 & ~n2727;
  assign n3389 = n3387 & n3388;
  assign n3390 = n2611 & ~n3389;
  assign n3391 = n2659 & n3133;
  assign n3392 = ~n3159 & ~n3391;
  assign n3393 = n2611 & ~n3392;
  assign n3394 = ~n2723 & ~n2738;
  assign n3395 = ~n3122 & n3394;
  assign n3396 = ~n2611 & ~n3395;
  assign n3397 = ~n3393 & ~n3396;
  assign n3398 = n2737 & ~n3137;
  assign n3399 = n3397 & n3398;
  assign n3400 = n2679 & ~n3399;
  assign n3401 = n2680 & n3133;
  assign n3402 = ~n2724 & ~n3401;
  assign n3403 = ~n3386 & n3402;
  assign n3404 = n2611 & n2631;
  assign n3405 = n3146 & n3404;
  assign n3406 = ~n2631 & n2659;
  assign n3407 = n2662 & n2702;
  assign n3408 = ~n3406 & ~n3407;
  assign n3409 = ~n2611 & ~n3408;
  assign n3410 = ~n3405 & ~n3409;
  assign n3411 = n3403 & n3410;
  assign n3412 = ~n2679 & ~n3411;
  assign n3413 = ~n3400 & ~n3412;
  assign n3414 = ~n3390 & n3413;
  assign n3415 = ~n3383 & n3414;
  assign n3416 = ~n3381 & n3415;
  assign n3417 = n3381 & ~n3415;
  assign po098 = n3416 | n3417;
  assign n3419 = ~pi153 & ~pi192;
  assign n3420 = pi192 & pi212;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = n576 & n3421;
  assign n3423 = pi153 & ~n576;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~n2257 & ~n2291;
  assign n3426 = ~n2249 & ~n3425;
  assign n3427 = ~n2179 & n3426;
  assign n3428 = n2179 & n2291;
  assign n3429 = n2249 & n3428;
  assign n3430 = n2229 & ~n2249;
  assign n3431 = ~n3308 & ~n3430;
  assign n3432 = n2179 & ~n3431;
  assign n3433 = ~n3429 & ~n3432;
  assign n3434 = n2179 & n2947;
  assign n3435 = n2249 & n2312;
  assign n3436 = ~n2263 & ~n3435;
  assign n3437 = ~n2179 & ~n3436;
  assign n3438 = ~n3434 & ~n3437;
  assign n3439 = ~n2229 & ~n2319;
  assign n3440 = n2249 & ~n3439;
  assign n3441 = n3438 & ~n3440;
  assign n3442 = ~n2285 & ~n3441;
  assign n3443 = ~n2266 & ~n2321;
  assign n3444 = n2179 & ~n3443;
  assign n3445 = ~n2302 & ~n2963;
  assign n3446 = ~n2179 & ~n3445;
  assign n3447 = ~n3444 & ~n3446;
  assign n3448 = ~n2301 & ~n2309;
  assign n3449 = n3447 & n3448;
  assign n3450 = n2285 & ~n3449;
  assign n3451 = ~n3442 & ~n3450;
  assign n3452 = n3433 & n3451;
  assign n3453 = ~n3427 & n3452;
  assign n3454 = n3424 & n3453;
  assign n3455 = ~n3424 & ~n3453;
  assign po099 = n3454 | n3455;
  assign n3457 = n576 & ~n954;
  assign n3458 = ~n620 & ~n1764;
  assign n3459 = ~n3457 & ~n3458;
  assign n3460 = n611 & ~n1823;
  assign n3461 = n3459 & ~n3460;
  assign n3462 = pi193 & ~n3461;
  assign n3463 = n592 & ~n961;
  assign n3464 = ~n592 & n947;
  assign n3465 = ~n3463 & ~n3464;
  assign n3466 = ~pi193 & ~n3465;
  assign po100 = n3462 | n3466;
  assign n3468 = n611 & ~n1211;
  assign n3469 = ~n620 & ~n1701;
  assign n3470 = ~n3468 & ~n3469;
  assign n3471 = n576 & ~n1010;
  assign n3472 = n3470 & ~n3471;
  assign n3473 = pi193 & ~n3472;
  assign n3474 = n592 & ~n1003;
  assign n3475 = ~n592 & ~n1017;
  assign n3476 = ~n3474 & ~n3475;
  assign n3477 = ~pi193 & ~n3476;
  assign po101 = n3473 | n3477;
  assign n3479 = n611 & ~n1077;
  assign n3480 = ~n620 & ~n1070;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = n576 & ~n1047;
  assign n3483 = n3481 & ~n3482;
  assign n3484 = pi193 & ~n3483;
  assign n3485 = n592 & ~n1823;
  assign n3486 = ~n592 & ~n1054;
  assign n3487 = ~n3485 & ~n3486;
  assign n3488 = ~pi193 & ~n3487;
  assign po102 = n3484 | n3488;
  assign n3490 = n576 & ~n605;
  assign n3491 = n611 & ~n626;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = ~n620 & ~n634;
  assign n3494 = n3492 & ~n3493;
  assign n3495 = pi193 & ~n3494;
  assign n3496 = n592 & ~n851;
  assign n3497 = ~n592 & n598;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = ~pi193 & ~n3498;
  assign po103 = n3495 | n3499;
  assign n3501 = n576 & ~n778;
  assign n3502 = n611 & n768;
  assign n3503 = ~n3501 & ~n3502;
  assign n3504 = ~n620 & ~n761;
  assign n3505 = n3503 & ~n3504;
  assign n3506 = pi193 & ~n3505;
  assign n3507 = n592 & ~n684;
  assign n3508 = ~n592 & n785;
  assign n3509 = ~n3507 & ~n3508;
  assign n3510 = ~pi193 & n3509;
  assign po105 = n3506 | n3510;
  assign n3512 = n576 & ~n971;
  assign n3513 = n611 & n947;
  assign n3514 = ~n3512 & ~n3513;
  assign n3515 = ~n620 & ~n961;
  assign n3516 = n3514 & ~n3515;
  assign n3517 = pi193 & ~n3516;
  assign n3518 = n592 & ~n1144;
  assign n3519 = ~n592 & ~n978;
  assign n3520 = ~n3518 & ~n3519;
  assign n3521 = ~pi193 & ~n3520;
  assign po106 = n3517 | n3521;
  assign n3523 = n611 & ~n653;
  assign n3524 = ~n620 & ~n703;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = n576 & ~n710;
  assign n3527 = n3525 & ~n3526;
  assign n3528 = pi193 & ~n3527;
  assign n3529 = n592 & ~n727;
  assign n3530 = ~n592 & ~n717;
  assign n3531 = ~n3529 & ~n3530;
  assign n3532 = ~pi193 & ~n3531;
  assign po107 = n3528 | n3532;
  assign n3534 = n576 & ~n669;
  assign n3535 = ~n620 & n684;
  assign n3536 = ~n3534 & ~n3535;
  assign n3537 = n611 & ~n785;
  assign n3538 = n3536 & ~n3537;
  assign n3539 = pi193 & ~n3538;
  assign n3540 = n592 & ~n660;
  assign n3541 = ~n592 & ~n676;
  assign n3542 = ~n3540 & ~n3541;
  assign n3543 = ~pi193 & ~n3542;
  assign po109 = n3539 | n3543;
  assign n3545 = pi082 & ~pi192;
  assign n3546 = n576 & n3545;
  assign n3547 = pi066 & n3546;
  assign n3548 = ~pi066 & ~pi081;
  assign n3549 = ~n583 & ~n3548;
  assign n3550 = ~n576 & ~n585;
  assign n3551 = n3549 & n3550;
  assign po134 = n3547 | n3551;
  assign n3553 = pi068 & n3546;
  assign n3554 = ~pi068 & ~n583;
  assign n3555 = ~n584 & ~n3554;
  assign n3556 = n3550 & n3555;
  assign po136 = n3553 | n3556;
  assign n3558 = pi069 & n3546;
  assign n3559 = ~pi069 & ~n584;
  assign n3560 = ~n585 & ~n3559;
  assign n3561 = n3550 & n3560;
  assign po137 = n3558 | n3561;
  assign n3563 = pi081 & pi082;
  assign n3564 = ~pi192 & ~n3563;
  assign n3565 = n576 & ~n3564;
  assign n3566 = ~pi081 & n3550;
  assign po149 = n3565 | n3566;
  assign n3568 = pi082 & ~n576;
  assign n3569 = ~pi192 & n576;
  assign po150 = n3568 | n3569;
  assign n3571 = ~pi082 & ~pi192;
  assign po161 = n576 & n3571;
  assign po066 = 1'b1;
  assign po162 = ~pi130;
  assign po163 = ~pi126;
  assign po164 = ~pi131;
  assign po165 = ~pi129;
  assign po166 = ~pi127;
  assign po167 = ~pi121;
  assign po168 = ~pi125;
  assign po169 = ~pi128;
  assign po170 = ~pi123;
  assign po171 = ~pi141;
  assign po172 = ~pi139;
  assign po173 = ~pi144;
  assign po174 = ~pi143;
  assign po175 = ~pi140;
  assign po176 = ~pi142;
  assign po177 = ~pi137;
  assign po178 = ~pi138;
  assign po179 = ~pi136;
  assign po180 = ~pi135;
  assign po181 = ~pi145;
  assign po182 = ~pi146;
  assign po183 = ~pi155;
  assign po184 = ~pi148;
  assign po185 = ~pi147;
  assign po186 = ~pi149;
  assign po187 = ~pi152;
  assign po188 = ~pi154;
  assign po190 = ~pi153;
  assign po192 = ~pi150;
  assign po200 = ~pi156;
  assign po201 = ~pi151;
  assign po202 = ~pi157;
  assign po000 = pi170;
  assign po001 = pi119;
  assign po002 = pi186;
  assign po003 = pi098;
  assign po004 = pi165;
  assign po005 = pi120;
  assign po006 = pi184;
  assign po007 = pi096;
  assign po008 = pi174;
  assign po009 = pi134;
  assign po010 = pi162;
  assign po011 = pi106;
  assign po012 = pi183;
  assign po013 = pi112;
  assign po014 = pi163;
  assign po015 = pi133;
  assign po016 = pi168;
  assign po017 = pi105;
  assign po018 = pi158;
  assign po019 = pi122;
  assign po020 = pi181;
  assign po021 = pi102;
  assign po022 = pi173;
  assign po023 = pi117;
  assign po024 = pi175;
  assign po025 = pi124;
  assign po026 = pi189;
  assign po027 = pi110;
  assign po028 = pi160;
  assign po029 = pi103;
  assign po030 = pi188;
  assign po031 = pi095;
  assign po032 = pi172;
  assign po033 = pi115;
  assign po034 = pi171;
  assign po035 = pi107;
  assign po036 = pi166;
  assign po037 = pi116;
  assign po038 = pi169;
  assign po039 = pi132;
  assign po040 = pi182;
  assign po041 = pi101;
  assign po042 = pi159;
  assign po043 = pi104;
  assign po044 = pi161;
  assign po045 = pi111;
  assign po046 = pi167;
  assign po047 = pi109;
  assign po048 = pi179;
  assign po049 = pi094;
  assign po050 = pi164;
  assign po051 = pi113;
  assign po052 = pi176;
  assign po053 = pi100;
  assign po054 = pi185;
  assign po055 = pi097;
  assign po056 = pi178;
  assign po057 = pi118;
  assign po058 = pi187;
  assign po059 = pi108;
  assign po060 = pi177;
  assign po061 = pi114;
  assign po062 = pi180;
  assign po063 = pi099;
  assign po064 = pi093;
  assign po065 = pi191;
  assign po067 = pi190;
  assign po226 = pi031;
  assign po227 = pi000;
  assign po228 = pi025;
  assign po229 = pi005;
  assign po230 = pi027;
  assign po231 = pi019;
  assign po232 = pi001;
  assign po233 = pi008;
  assign po234 = pi010;
  assign po235 = pi022;
  assign po236 = pi029;
  assign po237 = pi030;
  assign po238 = pi017;
  assign po239 = pi024;
  assign po240 = pi020;
  assign po241 = pi002;
  assign po242 = pi026;
  assign po243 = pi021;
  assign po244 = pi015;
  assign po245 = pi014;
  assign po246 = pi003;
  assign po247 = pi009;
  assign po248 = pi006;
  assign po249 = pi011;
  assign po250 = pi018;
  assign po251 = pi016;
  assign po252 = pi023;
  assign po253 = pi004;
  assign po254 = pi013;
  assign po255 = pi007;
  assign po256 = pi028;
  assign po257 = pi012;
endmodule


