module top (
            pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197, 
            po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224);
input pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196, pi1197;
output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223, po1224;
wire one, w0, w1, w2, w3, w4, w5, w6, w7, w8, w9, w10, w11, w12, w13, w14, w15, w16, w17, w18, w19, w20, w21, w22, w23, w24, w25, w26, w27, w28, w29, w30, w31, w32, w33, w34, w35, w36, w37, w38, w39, w40, w41, w42, w43, w44, w45, w46, w47, w48, w49, w50, w51, w52, w53, w54, w55, w56, w57, w58, w59, w60, w61, w62, w63, w64, w65, w66, w67, w68, w69, w70, w71, w72, w73, w74, w75, w76, w77, w78, w79, w80, w81, w82, w83, w84, w85, w86, w87, w88, w89, w90, w91, w92, w93, w94, w95, w96, w97, w98, w99, w100, w101, w102, w103, w104, w105, w106, w107, w108, w109, w110, w111, w112, w113, w114, w115, w116, w117, w118, w119, w120, w121, w122, w123, w124, w125, w126, w127, w128, w129, w130, w131, w132, w133, w134, w135, w136, w137, w138, w139, w140, w141, w142, w143, w144, w145, w146, w147, w148, w149, w150, w151, w152, w153, w154, w155, w156, w157, w158, w159, w160, w161, w162, w163, w164, w165, w166, w167, w168, w169, w170, w171, w172, w173, w174, w175, w176, w177, w178, w179, w180, w181, w182, w183, w184, w185, w186, w187, w188, w189, w190, w191, w192, w193, w194, w195, w196, w197, w198, w199, w200, w201, w202, w203, w204, w205, w206, w207, w208, w209, w210, w211, w212, w213, w214, w215, w216, w217, w218, w219, w220, w221, w222, w223, w224, w225, w226, w227, w228, w229, w230, w231, w232, w233, w234, w235, w236, w237, w238, w239, w240, w241, w242, w243, w244, w245, w246, w247, w248, w249, w250, w251, w252, w253, w254, w255, w256, w257, w258, w259, w260, w261, w262, w263, w264, w265, w266, w267, w268, w269, w270, w271, w272, w273, w274, w275, w276, w277, w278, w279, w280, w281, w282, w283, w284, w285, w286, w287, w288, w289, w290, w291, w292, w293, w294, w295, w296, w297, w298, w299, w300, w301, w302, w303, w304, w305, w306, w307, w308, w309, w310, w311, w312, w313, w314, w315, w316, w317, w318, w319, w320, w321, w322, w323, w324, w325, w326, w327, w328, w329, w330, w331, w332, w333, w334, w335, w336, w337, w338, w339, w340, w341, w342, w343, w344, w345, w346, w347, w348, w349, w350, w351, w352, w353, w354, w355, w356, w357, w358, w359, w360, w361, w362, w363, w364, w365, w366, w367, w368, w369, w370, w371, w372, w373, w374, w375, w376, w377, w378, w379, w380, w381, w382, w383, w384, w385, w386, w387, w388, w389, w390, w391, w392, w393, w394, w395, w396, w397, w398, w399, w400, w401, w402, w403, w404, w405, w406, w407, w408, w409, w410, w411, w412, w413, w414, w415, w416, w417, w418, w419, w420, w421, w422, w423, w424, w425, w426, w427, w428, w429, w430, w431, w432, w433, w434, w435, w436, w437, w438, w439, w440, w441, w442, w443, w444, w445, w446, w447, w448, w449, w450, w451, w452, w453, w454, w455, w456, w457, w458, w459, w460, w461, w462, w463, w464, w465, w466, w467, w468, w469, w470, w471, w472, w473, w474, w475, w476, w477, w478, w479, w480, w481, w482, w483, w484, w485, w486, w487, w488, w489, w490, w491, w492, w493, w494, w495, w496, w497, w498, w499, w500, w501, w502, w503, w504, w505, w506, w507, w508, w509, w510, w511, w512, w513, w514, w515, w516, w517, w518, w519, w520, w521, w522, w523, w524, w525, w526, w527, w528, w529, w530, w531, w532, w533, w534, w535, w536, w537, w538, w539, w540, w541, w542, w543, w544, w545, w546, w547, w548, w549, w550, w551, w552, w553, w554, w555, w556, w557, w558, w559, w560, w561, w562, w563, w564, w565, w566, w567, w568, w569, w570, w571, w572, w573, w574, w575, w576, w577, w578, w579, w580, w581, w582, w583, w584, w585, w586, w587, w588, w589, w590, w591, w592, w593, w594, w595, w596, w597, w598, w599, w600, w601, w602, w603, w604, w605, w606, w607, w608, w609, w610, w611, w612, w613, w614, w615, w616, w617, w618, w619, w620, w621, w622, w623, w624, w625, w626, w627, w628, w629, w630, w631, w632, w633, w634, w635, w636, w637, w638, w639, w640, w641, w642, w643, w644, w645, w646, w647, w648, w649, w650, w651, w652, w653, w654, w655, w656, w657, w658, w659, w660, w661, w662, w663, w664, w665, w666, w667, w668, w669, w670, w671, w672, w673, w674, w675, w676, w677, w678, w679, w680, w681, w682, w683, w684, w685, w686, w687, w688, w689, w690, w691, w692, w693, w694, w695, w696, w697, w698, w699, w700, w701, w702, w703, w704, w705, w706, w707, w708, w709, w710, w711, w712, w713, w714, w715, w716, w717, w718, w719, w720, w721, w722, w723, w724, w725, w726, w727, w728, w729, w730, w731, w732, w733, w734, w735, w736, w737, w738, w739, w740, w741, w742, w743, w744, w745, w746, w747, w748, w749, w750, w751, w752, w753, w754, w755, w756, w757, w758, w759, w760, w761, w762, w763, w764, w765, w766, w767, w768, w769, w770, w771, w772, w773, w774, w775, w776, w777, w778, w779, w780, w781, w782, w783, w784, w785, w786, w787, w788, w789, w790, w791, w792, w793, w794, w795, w796, w797, w798, w799, w800, w801, w802, w803, w804, w805, w806, w807, w808, w809, w810, w811, w812, w813, w814, w815, w816, w817, w818, w819, w820, w821, w822, w823, w824, w825, w826, w827, w828, w829, w830, w831, w832, w833, w834, w835, w836, w837, w838, w839, w840, w841, w842, w843, w844, w845, w846, w847, w848, w849, w850, w851, w852, w853, w854, w855, w856, w857, w858, w859, w860, w861, w862, w863, w864, w865, w866, w867, w868, w869, w870, w871, w872, w873, w874, w875, w876, w877, w878, w879, w880, w881, w882, w883, w884, w885, w886, w887, w888, w889, w890, w891, w892, w893, w894, w895, w896, w897, w898, w899, w900, w901, w902, w903, w904, w905, w906, w907, w908, w909, w910, w911, w912, w913, w914, w915, w916, w917, w918, w919, w920, w921, w922, w923, w924, w925, w926, w927, w928, w929, w930, w931, w932, w933, w934, w935, w936, w937, w938, w939, w940, w941, w942, w943, w944, w945, w946, w947, w948, w949, w950, w951, w952, w953, w954, w955, w956, w957, w958, w959, w960, w961, w962, w963, w964, w965, w966, w967, w968, w969, w970, w971, w972, w973, w974, w975, w976, w977, w978, w979, w980, w981, w982, w983, w984, w985, w986, w987, w988, w989, w990, w991, w992, w993, w994, w995, w996, w997, w998, w999, w1000, w1001, w1002, w1003, w1004, w1005, w1006, w1007, w1008, w1009, w1010, w1011, w1012, w1013, w1014, w1015, w1016, w1017, w1018, w1019, w1020, w1021, w1022, w1023, w1024, w1025, w1026, w1027, w1028, w1029, w1030, w1031, w1032, w1033, w1034, w1035, w1036, w1037, w1038, w1039, w1040, w1041, w1042, w1043, w1044, w1045, w1046, w1047, w1048, w1049, w1050, w1051, w1052, w1053, w1054, w1055, w1056, w1057, w1058, w1059, w1060, w1061, w1062, w1063, w1064, w1065, w1066, w1067, w1068, w1069, w1070, w1071, w1072, w1073, w1074, w1075, w1076, w1077, w1078, w1079, w1080, w1081, w1082, w1083, w1084, w1085, w1086, w1087, w1088, w1089, w1090, w1091, w1092, w1093, w1094, w1095, w1096, w1097, w1098, w1099, w1100, w1101, w1102, w1103, w1104, w1105, w1106, w1107, w1108, w1109, w1110, w1111, w1112, w1113, w1114, w1115, w1116, w1117, w1118, w1119, w1120, w1121, w1122, w1123, w1124, w1125, w1126, w1127, w1128, w1129, w1130, w1131, w1132, w1133, w1134, w1135, w1136, w1137, w1138, w1139, w1140, w1141, w1142, w1143, w1144, w1145, w1146, w1147, w1148, w1149, w1150, w1151, w1152, w1153, w1154, w1155, w1156, w1157, w1158, w1159, w1160, w1161, w1162, w1163, w1164, w1165, w1166, w1167, w1168, w1169, w1170, w1171, w1172, w1173, w1174, w1175, w1176, w1177, w1178, w1179, w1180, w1181, w1182, w1183, w1184, w1185, w1186, w1187, w1188, w1189, w1190, w1191, w1192, w1193, w1194, w1195, w1196, w1197, w1198, w1199, w1200, w1201, w1202, w1203, w1204, w1205, w1206, w1207, w1208, w1209, w1210, w1211, w1212, w1213, w1214, w1215, w1216, w1217, w1218, w1219, w1220, w1221, w1222, w1223, w1224, w1225, w1226, w1227, w1228, w1229, w1230, w1231, w1232, w1233, w1234, w1235, w1236, w1237, w1238, w1239, w1240, w1241, w1242, w1243, w1244, w1245, w1246, w1247, w1248, w1249, w1250, w1251, w1252, w1253, w1254, w1255, w1256, w1257, w1258, w1259, w1260, w1261, w1262, w1263, w1264, w1265, w1266, w1267, w1268, w1269, w1270, w1271, w1272, w1273, w1274, w1275, w1276, w1277, w1278, w1279, w1280, w1281, w1282, w1283, w1284, w1285, w1286, w1287, w1288, w1289, w1290, w1291, w1292, w1293, w1294, w1295, w1296, w1297, w1298, w1299, w1300, w1301, w1302, w1303, w1304, w1305, w1306, w1307, w1308, w1309, w1310, w1311, w1312, w1313, w1314, w1315, w1316, w1317, w1318, w1319, w1320, w1321, w1322, w1323, w1324, w1325, w1326, w1327, w1328, w1329, w1330, w1331, w1332, w1333, w1334, w1335, w1336, w1337, w1338, w1339, w1340, w1341, w1342, w1343, w1344, w1345, w1346, w1347, w1348, w1349, w1350, w1351, w1352, w1353, w1354, w1355, w1356, w1357, w1358, w1359, w1360, w1361, w1362, w1363, w1364, w1365, w1366, w1367, w1368, w1369, w1370, w1371, w1372, w1373, w1374, w1375, w1376, w1377, w1378, w1379, w1380, w1381, w1382, w1383, w1384, w1385, w1386, w1387, w1388, w1389, w1390, w1391, w1392, w1393, w1394, w1395, w1396, w1397, w1398, w1399, w1400, w1401, w1402, w1403, w1404, w1405, w1406, w1407, w1408, w1409, w1410, w1411, w1412, w1413, w1414, w1415, w1416, w1417, w1418, w1419, w1420, w1421, w1422, w1423, w1424, w1425, w1426, w1427, w1428, w1429, w1430, w1431, w1432, w1433, w1434, w1435, w1436, w1437, w1438, w1439, w1440, w1441, w1442, w1443, w1444, w1445, w1446, w1447, w1448, w1449, w1450, w1451, w1452, w1453, w1454, w1455, w1456, w1457, w1458, w1459, w1460, w1461, w1462, w1463, w1464, w1465, w1466, w1467, w1468, w1469, w1470, w1471, w1472, w1473, w1474, w1475, w1476, w1477, w1478, w1479, w1480, w1481, w1482, w1483, w1484, w1485, w1486, w1487, w1488, w1489, w1490, w1491, w1492, w1493, w1494, w1495, w1496, w1497, w1498, w1499, w1500, w1501, w1502, w1503, w1504, w1505, w1506, w1507, w1508, w1509, w1510, w1511, w1512, w1513, w1514, w1515, w1516, w1517, w1518, w1519, w1520, w1521, w1522, w1523, w1524, w1525, w1526, w1527, w1528, w1529, w1530, w1531, w1532, w1533, w1534, w1535, w1536, w1537, w1538, w1539, w1540, w1541, w1542, w1543, w1544, w1545, w1546, w1547, w1548, w1549, w1550, w1551, w1552, w1553, w1554, w1555, w1556, w1557, w1558, w1559, w1560, w1561, w1562, w1563, w1564, w1565, w1566, w1567, w1568, w1569, w1570, w1571, w1572, w1573, w1574, w1575, w1576, w1577, w1578, w1579, w1580, w1581, w1582, w1583, w1584, w1585, w1586, w1587, w1588, w1589, w1590, w1591, w1592, w1593, w1594, w1595, w1596, w1597, w1598, w1599, w1600, w1601, w1602, w1603, w1604, w1605, w1606, w1607, w1608, w1609, w1610, w1611, w1612, w1613, w1614, w1615, w1616, w1617, w1618, w1619, w1620, w1621, w1622, w1623, w1624, w1625, w1626, w1627, w1628, w1629, w1630, w1631, w1632, w1633, w1634, w1635, w1636, w1637, w1638, w1639, w1640, w1641, w1642, w1643, w1644, w1645, w1646, w1647, w1648, w1649, w1650, w1651, w1652, w1653, w1654, w1655, w1656, w1657, w1658, w1659, w1660, w1661, w1662, w1663, w1664, w1665, w1666, w1667, w1668, w1669, w1670, w1671, w1672, w1673, w1674, w1675, w1676, w1677, w1678, w1679, w1680, w1681, w1682, w1683, w1684, w1685, w1686, w1687, w1688, w1689, w1690, w1691, w1692, w1693, w1694, w1695, w1696, w1697, w1698, w1699, w1700, w1701, w1702, w1703, w1704, w1705, w1706, w1707, w1708, w1709, w1710, w1711, w1712, w1713, w1714, w1715, w1716, w1717, w1718, w1719, w1720, w1721, w1722, w1723, w1724, w1725, w1726, w1727, w1728, w1729, w1730, w1731, w1732, w1733, w1734, w1735, w1736, w1737, w1738, w1739, w1740, w1741, w1742, w1743, w1744, w1745, w1746, w1747, w1748, w1749, w1750, w1751, w1752, w1753, w1754, w1755, w1756, w1757, w1758, w1759, w1760, w1761, w1762, w1763, w1764, w1765, w1766, w1767, w1768, w1769, w1770, w1771, w1772, w1773, w1774, w1775, w1776, w1777, w1778, w1779, w1780, w1781, w1782, w1783, w1784, w1785, w1786, w1787, w1788, w1789, w1790, w1791, w1792, w1793, w1794, w1795, w1796, w1797, w1798, w1799, w1800, w1801, w1802, w1803, w1804, w1805, w1806, w1807, w1808, w1809, w1810, w1811, w1812, w1813, w1814, w1815, w1816, w1817, w1818, w1819, w1820, w1821, w1822, w1823, w1824, w1825, w1826, w1827, w1828, w1829, w1830, w1831, w1832, w1833, w1834, w1835, w1836, w1837, w1838, w1839, w1840, w1841, w1842, w1843, w1844, w1845, w1846, w1847, w1848, w1849, w1850, w1851, w1852, w1853, w1854, w1855, w1856, w1857, w1858, w1859, w1860, w1861, w1862, w1863, w1864, w1865, w1866, w1867, w1868, w1869, w1870, w1871, w1872, w1873, w1874, w1875, w1876, w1877, w1878, w1879, w1880, w1881, w1882, w1883, w1884, w1885, w1886, w1887, w1888, w1889, w1890, w1891, w1892, w1893, w1894, w1895, w1896, w1897, w1898, w1899, w1900, w1901, w1902, w1903, w1904, w1905, w1906, w1907, w1908, w1909, w1910, w1911, w1912, w1913, w1914, w1915, w1916, w1917, w1918, w1919, w1920, w1921, w1922, w1923, w1924, w1925, w1926, w1927, w1928, w1929, w1930, w1931, w1932, w1933, w1934, w1935, w1936, w1937, w1938, w1939, w1940, w1941, w1942, w1943, w1944, w1945, w1946, w1947, w1948, w1949, w1950, w1951, w1952, w1953, w1954, w1955, w1956, w1957, w1958, w1959, w1960, w1961, w1962, w1963, w1964, w1965, w1966, w1967, w1968, w1969, w1970, w1971, w1972, w1973, w1974, w1975, w1976, w1977, w1978, w1979, w1980, w1981, w1982, w1983, w1984, w1985, w1986, w1987, w1988, w1989, w1990, w1991, w1992, w1993, w1994, w1995, w1996, w1997, w1998, w1999, w2000, w2001, w2002, w2003, w2004, w2005, w2006, w2007, w2008, w2009, w2010, w2011, w2012, w2013, w2014, w2015, w2016, w2017, w2018, w2019, w2020, w2021, w2022, w2023, w2024, w2025, w2026, w2027, w2028, w2029, w2030, w2031, w2032, w2033, w2034, w2035, w2036, w2037, w2038, w2039, w2040, w2041, w2042, w2043, w2044, w2045, w2046, w2047, w2048, w2049, w2050, w2051, w2052, w2053, w2054, w2055, w2056, w2057, w2058, w2059, w2060, w2061, w2062, w2063, w2064, w2065, w2066, w2067, w2068, w2069, w2070, w2071, w2072, w2073, w2074, w2075, w2076, w2077, w2078, w2079, w2080, w2081, w2082, w2083, w2084, w2085, w2086, w2087, w2088, w2089, w2090, w2091, w2092, w2093, w2094, w2095, w2096, w2097, w2098, w2099, w2100, w2101, w2102, w2103, w2104, w2105, w2106, w2107, w2108, w2109, w2110, w2111, w2112, w2113, w2114, w2115, w2116, w2117, w2118, w2119, w2120, w2121, w2122, w2123, w2124, w2125, w2126, w2127, w2128, w2129, w2130, w2131, w2132, w2133, w2134, w2135, w2136, w2137, w2138, w2139, w2140, w2141, w2142, w2143, w2144, w2145, w2146, w2147, w2148, w2149, w2150, w2151, w2152, w2153, w2154, w2155, w2156, w2157, w2158, w2159, w2160, w2161, w2162, w2163, w2164, w2165, w2166, w2167, w2168, w2169, w2170, w2171, w2172, w2173, w2174, w2175, w2176, w2177, w2178, w2179, w2180, w2181, w2182, w2183, w2184, w2185, w2186, w2187, w2188, w2189, w2190, w2191, w2192, w2193, w2194, w2195, w2196, w2197, w2198, w2199, w2200, w2201, w2202, w2203, w2204, w2205, w2206, w2207, w2208, w2209, w2210, w2211, w2212, w2213, w2214, w2215, w2216, w2217, w2218, w2219, w2220, w2221, w2222, w2223, w2224, w2225, w2226, w2227, w2228, w2229, w2230, w2231, w2232, w2233, w2234, w2235, w2236, w2237, w2238, w2239, w2240, w2241, w2242, w2243, w2244, w2245, w2246, w2247, w2248, w2249, w2250, w2251, w2252, w2253, w2254, w2255, w2256, w2257, w2258, w2259, w2260, w2261, w2262, w2263, w2264, w2265, w2266, w2267, w2268, w2269, w2270, w2271, w2272, w2273, w2274, w2275, w2276, w2277, w2278, w2279, w2280, w2281, w2282, w2283, w2284, w2285, w2286, w2287, w2288, w2289, w2290, w2291, w2292, w2293, w2294, w2295, w2296, w2297, w2298, w2299, w2300, w2301, w2302, w2303, w2304, w2305, w2306, w2307, w2308, w2309, w2310, w2311, w2312, w2313, w2314, w2315, w2316, w2317, w2318, w2319, w2320, w2321, w2322, w2323, w2324, w2325, w2326, w2327, w2328, w2329, w2330, w2331, w2332, w2333, w2334, w2335, w2336, w2337, w2338, w2339, w2340, w2341, w2342, w2343, w2344, w2345, w2346, w2347, w2348, w2349, w2350, w2351, w2352, w2353, w2354, w2355, w2356, w2357, w2358, w2359, w2360, w2361, w2362, w2363, w2364, w2365, w2366, w2367, w2368, w2369, w2370, w2371, w2372, w2373, w2374, w2375, w2376, w2377, w2378, w2379, w2380, w2381, w2382, w2383, w2384, w2385, w2386, w2387, w2388, w2389, w2390, w2391, w2392, w2393, w2394, w2395, w2396, w2397, w2398, w2399, w2400, w2401, w2402, w2403, w2404, w2405, w2406, w2407, w2408, w2409, w2410, w2411, w2412, w2413, w2414, w2415, w2416, w2417, w2418, w2419, w2420, w2421, w2422, w2423, w2424, w2425, w2426, w2427, w2428, w2429, w2430, w2431, w2432, w2433, w2434, w2435, w2436, w2437, w2438, w2439, w2440, w2441, w2442, w2443, w2444, w2445, w2446, w2447, w2448, w2449, w2450, w2451, w2452, w2453, w2454, w2455, w2456, w2457, w2458, w2459, w2460, w2461, w2462, w2463, w2464, w2465, w2466, w2467, w2468, w2469, w2470, w2471, w2472, w2473, w2474, w2475, w2476, w2477, w2478, w2479, w2480, w2481, w2482, w2483, w2484, w2485, w2486, w2487, w2488, w2489, w2490, w2491, w2492, w2493, w2494, w2495, w2496, w2497, w2498, w2499, w2500, w2501, w2502, w2503, w2504, w2505, w2506, w2507, w2508, w2509, w2510, w2511, w2512, w2513, w2514, w2515, w2516, w2517, w2518, w2519, w2520, w2521, w2522, w2523, w2524, w2525, w2526, w2527, w2528, w2529, w2530, w2531, w2532, w2533, w2534, w2535, w2536, w2537, w2538, w2539, w2540, w2541, w2542, w2543, w2544, w2545, w2546, w2547, w2548, w2549, w2550, w2551, w2552, w2553, w2554, w2555, w2556, w2557, w2558, w2559, w2560, w2561, w2562, w2563, w2564, w2565, w2566, w2567, w2568, w2569, w2570, w2571, w2572, w2573, w2574, w2575, w2576, w2577, w2578, w2579, w2580, w2581, w2582, w2583, w2584, w2585, w2586, w2587, w2588, w2589, w2590, w2591, w2592, w2593, w2594, w2595, w2596, w2597, w2598, w2599, w2600, w2601, w2602, w2603, w2604, w2605, w2606, w2607, w2608, w2609, w2610, w2611, w2612, w2613, w2614, w2615, w2616, w2617, w2618, w2619, w2620, w2621, w2622, w2623, w2624, w2625, w2626, w2627, w2628, w2629, w2630, w2631, w2632, w2633, w2634, w2635, w2636, w2637, w2638, w2639, w2640, w2641, w2642, w2643, w2644, w2645, w2646, w2647, w2648, w2649, w2650, w2651, w2652, w2653, w2654, w2655, w2656, w2657, w2658, w2659, w2660, w2661, w2662, w2663, w2664, w2665, w2666, w2667, w2668, w2669, w2670, w2671, w2672, w2673, w2674, w2675, w2676, w2677, w2678, w2679, w2680, w2681, w2682, w2683, w2684, w2685, w2686, w2687, w2688, w2689, w2690, w2691, w2692, w2693, w2694, w2695, w2696, w2697, w2698, w2699, w2700, w2701, w2702, w2703, w2704, w2705, w2706, w2707, w2708, w2709, w2710, w2711, w2712, w2713, w2714, w2715, w2716, w2717, w2718, w2719, w2720, w2721, w2722, w2723, w2724, w2725, w2726, w2727, w2728, w2729, w2730, w2731, w2732, w2733, w2734, w2735, w2736, w2737, w2738, w2739, w2740, w2741, w2742, w2743, w2744, w2745, w2746, w2747, w2748, w2749, w2750, w2751, w2752, w2753, w2754, w2755, w2756, w2757, w2758, w2759, w2760, w2761, w2762, w2763, w2764, w2765, w2766, w2767, w2768, w2769, w2770, w2771, w2772, w2773, w2774, w2775, w2776, w2777, w2778, w2779, w2780, w2781, w2782, w2783, w2784, w2785, w2786, w2787, w2788, w2789, w2790, w2791, w2792, w2793, w2794, w2795, w2796, w2797, w2798, w2799, w2800, w2801, w2802, w2803, w2804, w2805, w2806, w2807, w2808, w2809, w2810, w2811, w2812, w2813, w2814, w2815, w2816, w2817, w2818, w2819, w2820, w2821, w2822, w2823, w2824, w2825, w2826, w2827, w2828, w2829, w2830, w2831, w2832, w2833, w2834, w2835, w2836, w2837, w2838, w2839, w2840, w2841, w2842, w2843, w2844, w2845, w2846, w2847, w2848, w2849, w2850, w2851, w2852, w2853, w2854, w2855, w2856, w2857, w2858, w2859, w2860, w2861, w2862, w2863, w2864, w2865, w2866, w2867, w2868, w2869, w2870, w2871, w2872, w2873, w2874, w2875, w2876, w2877, w2878, w2879, w2880, w2881, w2882, w2883, w2884, w2885, w2886, w2887, w2888, w2889, w2890, w2891, w2892, w2893, w2894, w2895, w2896, w2897, w2898, w2899, w2900, w2901, w2902, w2903, w2904, w2905, w2906, w2907, w2908, w2909, w2910, w2911, w2912, w2913, w2914, w2915, w2916, w2917, w2918, w2919, w2920, w2921, w2922, w2923, w2924, w2925, w2926, w2927, w2928, w2929, w2930, w2931, w2932, w2933, w2934, w2935, w2936, w2937, w2938, w2939, w2940, w2941, w2942, w2943, w2944, w2945, w2946, w2947, w2948, w2949, w2950, w2951, w2952, w2953, w2954, w2955, w2956, w2957, w2958, w2959, w2960, w2961, w2962, w2963, w2964, w2965, w2966, w2967, w2968, w2969, w2970, w2971, w2972, w2973, w2974, w2975, w2976, w2977, w2978, w2979, w2980, w2981, w2982, w2983, w2984, w2985, w2986, w2987, w2988, w2989, w2990, w2991, w2992, w2993, w2994, w2995, w2996, w2997, w2998, w2999, w3000, w3001, w3002, w3003, w3004, w3005, w3006, w3007, w3008, w3009, w3010, w3011, w3012, w3013, w3014, w3015, w3016, w3017, w3018, w3019, w3020, w3021, w3022, w3023, w3024, w3025, w3026, w3027, w3028, w3029, w3030, w3031, w3032, w3033, w3034, w3035, w3036, w3037, w3038, w3039, w3040, w3041, w3042, w3043, w3044, w3045, w3046, w3047, w3048, w3049, w3050, w3051, w3052, w3053, w3054, w3055, w3056, w3057, w3058, w3059, w3060, w3061, w3062, w3063, w3064, w3065, w3066, w3067, w3068, w3069, w3070, w3071, w3072, w3073, w3074, w3075, w3076, w3077, w3078, w3079, w3080, w3081, w3082, w3083, w3084, w3085, w3086, w3087, w3088, w3089, w3090, w3091, w3092, w3093, w3094, w3095, w3096, w3097, w3098, w3099, w3100, w3101, w3102, w3103, w3104, w3105, w3106, w3107, w3108, w3109, w3110, w3111, w3112, w3113, w3114, w3115, w3116, w3117, w3118, w3119, w3120, w3121, w3122, w3123, w3124, w3125, w3126, w3127, w3128, w3129, w3130, w3131, w3132, w3133, w3134, w3135, w3136, w3137, w3138, w3139, w3140, w3141, w3142, w3143, w3144, w3145, w3146, w3147, w3148, w3149, w3150, w3151, w3152, w3153, w3154, w3155, w3156, w3157, w3158, w3159, w3160, w3161, w3162, w3163, w3164, w3165, w3166, w3167, w3168, w3169, w3170, w3171, w3172, w3173, w3174, w3175, w3176, w3177, w3178, w3179, w3180, w3181, w3182, w3183, w3184, w3185, w3186, w3187, w3188, w3189, w3190, w3191, w3192, w3193, w3194, w3195, w3196, w3197, w3198, w3199, w3200, w3201, w3202, w3203, w3204, w3205, w3206, w3207, w3208, w3209, w3210, w3211, w3212, w3213, w3214, w3215, w3216, w3217, w3218, w3219, w3220, w3221, w3222, w3223, w3224, w3225, w3226, w3227, w3228, w3229, w3230, w3231, w3232, w3233, w3234, w3235, w3236, w3237, w3238, w3239, w3240, w3241, w3242, w3243, w3244, w3245, w3246, w3247, w3248, w3249, w3250, w3251, w3252, w3253, w3254, w3255, w3256, w3257, w3258, w3259, w3260, w3261, w3262, w3263, w3264, w3265, w3266, w3267, w3268, w3269, w3270, w3271, w3272, w3273, w3274, w3275, w3276, w3277, w3278, w3279, w3280, w3281, w3282, w3283, w3284, w3285, w3286, w3287, w3288, w3289, w3290, w3291, w3292, w3293, w3294, w3295, w3296, w3297, w3298, w3299, w3300, w3301, w3302, w3303, w3304, w3305, w3306, w3307, w3308, w3309, w3310, w3311, w3312, w3313, w3314, w3315, w3316, w3317, w3318, w3319, w3320, w3321, w3322, w3323, w3324, w3325, w3326, w3327, w3328, w3329, w3330, w3331, w3332, w3333, w3334, w3335, w3336, w3337, w3338, w3339, w3340, w3341, w3342, w3343, w3344, w3345, w3346, w3347, w3348, w3349, w3350, w3351, w3352, w3353, w3354, w3355, w3356, w3357, w3358, w3359, w3360, w3361, w3362, w3363, w3364, w3365, w3366, w3367, w3368, w3369, w3370, w3371, w3372, w3373, w3374, w3375, w3376, w3377, w3378, w3379, w3380, w3381, w3382, w3383, w3384, w3385, w3386, w3387, w3388, w3389, w3390, w3391, w3392, w3393, w3394, w3395, w3396, w3397, w3398, w3399, w3400, w3401, w3402, w3403, w3404, w3405, w3406, w3407, w3408, w3409, w3410, w3411, w3412, w3413, w3414, w3415, w3416, w3417, w3418, w3419, w3420, w3421, w3422, w3423, w3424, w3425, w3426, w3427, w3428, w3429, w3430, w3431, w3432, w3433, w3434, w3435, w3436, w3437, w3438, w3439, w3440, w3441, w3442, w3443, w3444, w3445, w3446, w3447, w3448, w3449, w3450, w3451, w3452, w3453, w3454, w3455, w3456, w3457, w3458, w3459, w3460, w3461, w3462, w3463, w3464, w3465, w3466, w3467, w3468, w3469, w3470, w3471, w3472, w3473, w3474, w3475, w3476, w3477, w3478, w3479, w3480, w3481, w3482, w3483, w3484, w3485, w3486, w3487, w3488, w3489, w3490, w3491, w3492, w3493, w3494, w3495, w3496, w3497, w3498, w3499, w3500, w3501, w3502, w3503, w3504, w3505, w3506, w3507, w3508, w3509, w3510, w3511, w3512, w3513, w3514, w3515, w3516, w3517, w3518, w3519, w3520, w3521, w3522, w3523, w3524, w3525, w3526, w3527, w3528, w3529, w3530, w3531, w3532, w3533, w3534, w3535, w3536, w3537, w3538, w3539, w3540, w3541, w3542, w3543, w3544, w3545, w3546, w3547, w3548, w3549, w3550, w3551, w3552, w3553, w3554, w3555, w3556, w3557, w3558, w3559, w3560, w3561, w3562, w3563, w3564, w3565, w3566, w3567, w3568, w3569, w3570, w3571, w3572, w3573, w3574, w3575, w3576, w3577, w3578, w3579, w3580, w3581, w3582, w3583, w3584, w3585, w3586, w3587, w3588, w3589, w3590, w3591, w3592, w3593, w3594, w3595, w3596, w3597, w3598, w3599, w3600, w3601, w3602, w3603, w3604, w3605, w3606, w3607, w3608, w3609, w3610, w3611, w3612, w3613, w3614, w3615, w3616, w3617, w3618, w3619, w3620, w3621, w3622, w3623, w3624, w3625, w3626, w3627, w3628, w3629, w3630, w3631, w3632, w3633, w3634, w3635, w3636, w3637, w3638, w3639, w3640, w3641, w3642, w3643, w3644, w3645, w3646, w3647, w3648, w3649, w3650, w3651, w3652, w3653, w3654, w3655, w3656, w3657, w3658, w3659, w3660, w3661, w3662, w3663, w3664, w3665, w3666, w3667, w3668, w3669, w3670, w3671, w3672, w3673, w3674, w3675, w3676, w3677, w3678, w3679, w3680, w3681, w3682, w3683, w3684, w3685, w3686, w3687, w3688, w3689, w3690, w3691, w3692, w3693, w3694, w3695, w3696, w3697, w3698, w3699, w3700, w3701, w3702, w3703, w3704, w3705, w3706, w3707, w3708, w3709, w3710, w3711, w3712, w3713, w3714, w3715, w3716, w3717, w3718, w3719, w3720, w3721, w3722, w3723, w3724, w3725, w3726, w3727, w3728, w3729, w3730, w3731, w3732, w3733, w3734, w3735, w3736, w3737, w3738, w3739, w3740, w3741, w3742, w3743, w3744, w3745, w3746, w3747, w3748, w3749, w3750, w3751, w3752, w3753, w3754, w3755, w3756, w3757, w3758, w3759, w3760, w3761, w3762, w3763, w3764, w3765, w3766, w3767, w3768, w3769, w3770, w3771, w3772, w3773, w3774, w3775, w3776, w3777, w3778, w3779, w3780, w3781, w3782, w3783, w3784, w3785, w3786, w3787, w3788, w3789, w3790, w3791, w3792, w3793, w3794, w3795, w3796, w3797, w3798, w3799, w3800, w3801, w3802, w3803, w3804, w3805, w3806, w3807, w3808, w3809, w3810, w3811, w3812, w3813, w3814, w3815, w3816, w3817, w3818, w3819, w3820, w3821, w3822, w3823, w3824, w3825, w3826, w3827, w3828, w3829, w3830, w3831, w3832, w3833, w3834, w3835, w3836, w3837, w3838, w3839, w3840, w3841, w3842, w3843, w3844, w3845, w3846, w3847, w3848, w3849, w3850, w3851, w3852, w3853, w3854, w3855, w3856, w3857, w3858, w3859, w3860, w3861, w3862, w3863, w3864, w3865, w3866, w3867, w3868, w3869, w3870, w3871, w3872, w3873, w3874, w3875, w3876, w3877, w3878, w3879, w3880, w3881, w3882, w3883, w3884, w3885, w3886, w3887, w3888, w3889, w3890, w3891, w3892, w3893, w3894, w3895, w3896, w3897, w3898, w3899, w3900, w3901, w3902, w3903, w3904, w3905, w3906, w3907, w3908, w3909, w3910, w3911, w3912, w3913, w3914, w3915, w3916, w3917, w3918, w3919, w3920, w3921, w3922, w3923, w3924, w3925, w3926, w3927, w3928, w3929, w3930, w3931, w3932, w3933, w3934, w3935, w3936, w3937, w3938, w3939, w3940, w3941, w3942, w3943, w3944, w3945, w3946, w3947, w3948, w3949, w3950, w3951, w3952, w3953, w3954, w3955, w3956, w3957, w3958, w3959, w3960, w3961, w3962, w3963, w3964, w3965, w3966, w3967, w3968, w3969, w3970, w3971, w3972, w3973, w3974, w3975, w3976, w3977, w3978, w3979, w3980, w3981, w3982, w3983, w3984, w3985, w3986, w3987, w3988, w3989, w3990, w3991, w3992, w3993, w3994, w3995, w3996, w3997, w3998, w3999, w4000, w4001, w4002, w4003, w4004, w4005, w4006, w4007, w4008, w4009, w4010, w4011, w4012, w4013, w4014, w4015, w4016, w4017, w4018, w4019, w4020, w4021, w4022, w4023, w4024, w4025, w4026, w4027, w4028, w4029, w4030, w4031, w4032, w4033, w4034, w4035, w4036, w4037, w4038, w4039, w4040, w4041, w4042, w4043, w4044, w4045, w4046, w4047, w4048, w4049, w4050, w4051, w4052, w4053, w4054, w4055, w4056, w4057, w4058, w4059, w4060, w4061, w4062, w4063, w4064, w4065, w4066, w4067, w4068, w4069, w4070, w4071, w4072, w4073, w4074, w4075, w4076, w4077, w4078, w4079, w4080, w4081, w4082, w4083, w4084, w4085, w4086, w4087, w4088, w4089, w4090, w4091, w4092, w4093, w4094, w4095, w4096, w4097, w4098, w4099, w4100, w4101, w4102, w4103, w4104, w4105, w4106, w4107, w4108, w4109, w4110, w4111, w4112, w4113, w4114, w4115, w4116, w4117, w4118, w4119, w4120, w4121, w4122, w4123, w4124, w4125, w4126, w4127, w4128, w4129, w4130, w4131, w4132, w4133, w4134, w4135, w4136, w4137, w4138, w4139, w4140, w4141, w4142, w4143, w4144, w4145, w4146, w4147, w4148, w4149, w4150, w4151, w4152, w4153, w4154, w4155, w4156, w4157, w4158, w4159, w4160, w4161, w4162, w4163, w4164, w4165, w4166, w4167, w4168, w4169, w4170, w4171, w4172, w4173, w4174, w4175, w4176, w4177, w4178, w4179, w4180, w4181, w4182, w4183, w4184, w4185, w4186, w4187, w4188, w4189, w4190, w4191, w4192, w4193, w4194, w4195, w4196, w4197, w4198, w4199, w4200, w4201, w4202, w4203, w4204, w4205, w4206, w4207, w4208, w4209, w4210, w4211, w4212, w4213, w4214, w4215, w4216, w4217, w4218, w4219, w4220, w4221, w4222, w4223, w4224, w4225, w4226, w4227, w4228, w4229, w4230, w4231, w4232, w4233, w4234, w4235, w4236, w4237, w4238, w4239, w4240, w4241, w4242, w4243, w4244, w4245, w4246, w4247, w4248, w4249, w4250, w4251, w4252, w4253, w4254, w4255, w4256, w4257, w4258, w4259, w4260, w4261, w4262, w4263, w4264, w4265, w4266, w4267, w4268, w4269, w4270, w4271, w4272, w4273, w4274, w4275, w4276, w4277, w4278, w4279, w4280, w4281, w4282, w4283, w4284, w4285, w4286, w4287, w4288, w4289, w4290, w4291, w4292, w4293, w4294, w4295, w4296, w4297, w4298, w4299, w4300, w4301, w4302, w4303, w4304, w4305, w4306, w4307, w4308, w4309, w4310, w4311, w4312, w4313, w4314, w4315, w4316, w4317, w4318, w4319, w4320, w4321, w4322, w4323, w4324, w4325, w4326, w4327, w4328, w4329, w4330, w4331, w4332, w4333, w4334, w4335, w4336, w4337, w4338, w4339, w4340, w4341, w4342, w4343, w4344, w4345, w4346, w4347, w4348, w4349, w4350, w4351, w4352, w4353, w4354, w4355, w4356, w4357, w4358, w4359, w4360, w4361, w4362, w4363, w4364, w4365, w4366, w4367, w4368, w4369, w4370, w4371, w4372, w4373, w4374, w4375, w4376, w4377, w4378, w4379, w4380, w4381, w4382, w4383, w4384, w4385, w4386, w4387, w4388, w4389, w4390, w4391, w4392, w4393, w4394, w4395, w4396, w4397, w4398, w4399, w4400, w4401, w4402, w4403, w4404, w4405, w4406, w4407, w4408, w4409, w4410, w4411, w4412, w4413, w4414, w4415, w4416, w4417, w4418, w4419, w4420, w4421, w4422, w4423, w4424, w4425, w4426, w4427, w4428, w4429, w4430, w4431, w4432, w4433, w4434, w4435, w4436, w4437, w4438, w4439, w4440, w4441, w4442, w4443, w4444, w4445, w4446, w4447, w4448, w4449, w4450, w4451, w4452, w4453, w4454, w4455, w4456, w4457, w4458, w4459, w4460, w4461, w4462, w4463, w4464, w4465, w4466, w4467, w4468, w4469, w4470, w4471, w4472, w4473, w4474, w4475, w4476, w4477, w4478, w4479, w4480, w4481, w4482, w4483, w4484, w4485, w4486, w4487, w4488, w4489, w4490, w4491, w4492, w4493, w4494, w4495, w4496, w4497, w4498, w4499, w4500, w4501, w4502, w4503, w4504, w4505, w4506, w4507, w4508, w4509, w4510, w4511, w4512, w4513, w4514, w4515, w4516, w4517, w4518, w4519, w4520, w4521, w4522, w4523, w4524, w4525, w4526, w4527, w4528, w4529, w4530, w4531, w4532, w4533, w4534, w4535, w4536, w4537, w4538, w4539, w4540, w4541, w4542, w4543, w4544, w4545, w4546, w4547, w4548, w4549, w4550, w4551, w4552, w4553, w4554, w4555, w4556, w4557, w4558, w4559, w4560, w4561, w4562, w4563, w4564, w4565, w4566, w4567, w4568, w4569, w4570, w4571, w4572, w4573, w4574, w4575, w4576, w4577, w4578, w4579, w4580, w4581, w4582, w4583, w4584, w4585, w4586, w4587, w4588, w4589, w4590, w4591, w4592, w4593, w4594, w4595, w4596, w4597, w4598, w4599, w4600, w4601, w4602, w4603, w4604, w4605, w4606, w4607, w4608, w4609, w4610, w4611, w4612, w4613, w4614, w4615, w4616, w4617, w4618, w4619, w4620, w4621, w4622, w4623, w4624, w4625, w4626, w4627, w4628, w4629, w4630, w4631, w4632, w4633, w4634, w4635, w4636, w4637, w4638, w4639, w4640, w4641, w4642, w4643, w4644, w4645, w4646, w4647, w4648, w4649, w4650, w4651, w4652, w4653, w4654, w4655, w4656, w4657, w4658, w4659, w4660, w4661, w4662, w4663, w4664, w4665, w4666, w4667, w4668, w4669, w4670, w4671, w4672, w4673, w4674, w4675, w4676, w4677, w4678, w4679, w4680, w4681, w4682, w4683, w4684, w4685, w4686, w4687, w4688, w4689, w4690, w4691, w4692, w4693, w4694, w4695, w4696, w4697, w4698, w4699, w4700, w4701, w4702, w4703, w4704, w4705, w4706, w4707, w4708, w4709, w4710, w4711, w4712, w4713, w4714, w4715, w4716, w4717, w4718, w4719, w4720, w4721, w4722, w4723, w4724, w4725, w4726, w4727, w4728, w4729, w4730, w4731, w4732, w4733, w4734, w4735, w4736, w4737, w4738, w4739, w4740, w4741, w4742, w4743, w4744, w4745, w4746, w4747, w4748, w4749, w4750, w4751, w4752, w4753, w4754, w4755, w4756, w4757, w4758, w4759, w4760, w4761, w4762, w4763, w4764, w4765, w4766, w4767, w4768, w4769, w4770, w4771, w4772, w4773, w4774, w4775, w4776, w4777, w4778, w4779, w4780, w4781, w4782, w4783, w4784, w4785, w4786, w4787, w4788, w4789, w4790, w4791, w4792, w4793, w4794, w4795, w4796, w4797, w4798, w4799, w4800, w4801, w4802, w4803, w4804, w4805, w4806, w4807, w4808, w4809, w4810, w4811, w4812, w4813, w4814, w4815, w4816, w4817, w4818, w4819, w4820, w4821, w4822, w4823, w4824, w4825, w4826, w4827, w4828, w4829, w4830, w4831, w4832, w4833, w4834, w4835, w4836, w4837, w4838, w4839, w4840, w4841, w4842, w4843, w4844, w4845, w4846, w4847, w4848, w4849, w4850, w4851, w4852, w4853, w4854, w4855, w4856, w4857, w4858, w4859, w4860, w4861, w4862, w4863, w4864, w4865, w4866, w4867, w4868, w4869, w4870, w4871, w4872, w4873, w4874, w4875, w4876, w4877, w4878, w4879, w4880, w4881, w4882, w4883, w4884, w4885, w4886, w4887, w4888, w4889, w4890, w4891, w4892, w4893, w4894, w4895, w4896, w4897, w4898, w4899, w4900, w4901, w4902, w4903, w4904, w4905, w4906, w4907, w4908, w4909, w4910, w4911, w4912, w4913, w4914, w4915, w4916, w4917, w4918, w4919, w4920, w4921, w4922, w4923, w4924, w4925, w4926, w4927, w4928, w4929, w4930, w4931, w4932, w4933, w4934, w4935, w4936, w4937, w4938, w4939, w4940, w4941, w4942, w4943, w4944, w4945, w4946, w4947, w4948, w4949, w4950, w4951, w4952, w4953, w4954, w4955, w4956, w4957, w4958, w4959, w4960, w4961, w4962, w4963, w4964, w4965, w4966, w4967, w4968, w4969, w4970, w4971, w4972, w4973, w4974, w4975, w4976, w4977, w4978, w4979, w4980, w4981, w4982, w4983, w4984, w4985, w4986, w4987, w4988, w4989, w4990, w4991, w4992, w4993, w4994, w4995, w4996, w4997, w4998, w4999, w5000, w5001, w5002, w5003, w5004, w5005, w5006, w5007, w5008, w5009, w5010, w5011, w5012, w5013, w5014, w5015, w5016, w5017, w5018, w5019, w5020, w5021, w5022, w5023, w5024, w5025, w5026, w5027, w5028, w5029, w5030, w5031, w5032, w5033, w5034, w5035, w5036, w5037, w5038, w5039, w5040, w5041, w5042, w5043, w5044, w5045, w5046, w5047, w5048, w5049, w5050, w5051, w5052, w5053, w5054, w5055, w5056, w5057, w5058, w5059, w5060, w5061, w5062, w5063, w5064, w5065, w5066, w5067, w5068, w5069, w5070, w5071, w5072, w5073, w5074, w5075, w5076, w5077, w5078, w5079, w5080, w5081, w5082, w5083, w5084, w5085, w5086, w5087, w5088, w5089, w5090, w5091, w5092, w5093, w5094, w5095, w5096, w5097, w5098, w5099, w5100, w5101, w5102, w5103, w5104, w5105, w5106, w5107, w5108, w5109, w5110, w5111, w5112, w5113, w5114, w5115, w5116, w5117, w5118, w5119, w5120, w5121, w5122, w5123, w5124, w5125, w5126, w5127, w5128, w5129, w5130, w5131, w5132, w5133, w5134, w5135, w5136, w5137, w5138, w5139, w5140, w5141, w5142, w5143, w5144, w5145, w5146, w5147, w5148, w5149, w5150, w5151, w5152, w5153, w5154, w5155, w5156, w5157, w5158, w5159, w5160, w5161, w5162, w5163, w5164, w5165, w5166, w5167, w5168, w5169, w5170, w5171, w5172, w5173, w5174, w5175, w5176, w5177, w5178, w5179, w5180, w5181, w5182, w5183, w5184, w5185, w5186, w5187, w5188, w5189, w5190, w5191, w5192, w5193, w5194, w5195, w5196, w5197, w5198, w5199, w5200, w5201, w5202, w5203, w5204, w5205, w5206, w5207, w5208, w5209, w5210, w5211, w5212, w5213, w5214, w5215, w5216, w5217, w5218, w5219, w5220, w5221, w5222, w5223, w5224, w5225, w5226, w5227, w5228, w5229, w5230, w5231, w5232, w5233, w5234, w5235, w5236, w5237, w5238, w5239, w5240, w5241, w5242, w5243, w5244, w5245, w5246, w5247, w5248, w5249, w5250, w5251, w5252, w5253, w5254, w5255, w5256, w5257, w5258, w5259, w5260, w5261, w5262, w5263, w5264, w5265, w5266, w5267, w5268, w5269, w5270, w5271, w5272, w5273, w5274, w5275, w5276, w5277, w5278, w5279, w5280, w5281, w5282, w5283, w5284, w5285, w5286, w5287, w5288, w5289, w5290, w5291, w5292, w5293, w5294, w5295, w5296, w5297, w5298, w5299, w5300, w5301, w5302, w5303, w5304, w5305, w5306, w5307, w5308, w5309, w5310, w5311, w5312, w5313, w5314, w5315, w5316, w5317, w5318, w5319, w5320, w5321, w5322, w5323, w5324, w5325, w5326, w5327, w5328, w5329, w5330, w5331, w5332, w5333, w5334, w5335, w5336, w5337, w5338, w5339, w5340, w5341, w5342, w5343, w5344, w5345, w5346, w5347, w5348, w5349, w5350, w5351, w5352, w5353, w5354, w5355, w5356, w5357, w5358, w5359, w5360, w5361, w5362, w5363, w5364, w5365, w5366, w5367, w5368, w5369, w5370, w5371, w5372, w5373, w5374, w5375, w5376, w5377, w5378, w5379, w5380, w5381, w5382, w5383, w5384, w5385, w5386, w5387, w5388, w5389, w5390, w5391, w5392, w5393, w5394, w5395, w5396, w5397, w5398, w5399, w5400, w5401, w5402, w5403, w5404, w5405, w5406, w5407, w5408, w5409, w5410, w5411, w5412, w5413, w5414, w5415, w5416, w5417, w5418, w5419, w5420, w5421, w5422, w5423, w5424, w5425, w5426, w5427, w5428, w5429, w5430, w5431, w5432, w5433, w5434, w5435, w5436, w5437, w5438, w5439, w5440, w5441, w5442, w5443, w5444, w5445, w5446, w5447, w5448, w5449, w5450, w5451, w5452, w5453, w5454, w5455, w5456, w5457, w5458, w5459, w5460, w5461, w5462, w5463, w5464, w5465, w5466, w5467, w5468, w5469, w5470, w5471, w5472, w5473, w5474, w5475, w5476, w5477, w5478, w5479, w5480, w5481, w5482, w5483, w5484, w5485, w5486, w5487, w5488, w5489, w5490, w5491, w5492, w5493, w5494, w5495, w5496, w5497, w5498, w5499, w5500, w5501, w5502, w5503, w5504, w5505, w5506, w5507, w5508, w5509, w5510, w5511, w5512, w5513, w5514, w5515, w5516, w5517, w5518, w5519, w5520, w5521, w5522, w5523, w5524, w5525, w5526, w5527, w5528, w5529, w5530, w5531, w5532, w5533, w5534, w5535, w5536, w5537, w5538, w5539, w5540, w5541, w5542, w5543, w5544, w5545, w5546, w5547, w5548, w5549, w5550, w5551, w5552, w5553, w5554, w5555, w5556, w5557, w5558, w5559, w5560, w5561, w5562, w5563, w5564, w5565, w5566, w5567, w5568, w5569, w5570, w5571, w5572, w5573, w5574, w5575, w5576, w5577, w5578, w5579, w5580, w5581, w5582, w5583, w5584, w5585, w5586, w5587, w5588, w5589, w5590, w5591, w5592, w5593, w5594, w5595, w5596, w5597, w5598, w5599, w5600, w5601, w5602, w5603, w5604, w5605, w5606, w5607, w5608, w5609, w5610, w5611, w5612, w5613, w5614, w5615, w5616, w5617, w5618, w5619, w5620, w5621, w5622, w5623, w5624, w5625, w5626, w5627, w5628, w5629, w5630, w5631, w5632, w5633, w5634, w5635, w5636, w5637, w5638, w5639, w5640, w5641, w5642, w5643, w5644, w5645, w5646, w5647, w5648, w5649, w5650, w5651, w5652, w5653, w5654, w5655, w5656, w5657, w5658, w5659, w5660, w5661, w5662, w5663, w5664, w5665, w5666, w5667, w5668, w5669, w5670, w5671, w5672, w5673, w5674, w5675, w5676, w5677, w5678, w5679, w5680, w5681, w5682, w5683, w5684, w5685, w5686, w5687, w5688, w5689, w5690, w5691, w5692, w5693, w5694, w5695, w5696, w5697, w5698, w5699, w5700, w5701, w5702, w5703, w5704, w5705, w5706, w5707, w5708, w5709, w5710, w5711, w5712, w5713, w5714, w5715, w5716, w5717, w5718, w5719, w5720, w5721, w5722, w5723, w5724, w5725, w5726, w5727, w5728, w5729, w5730, w5731, w5732, w5733, w5734, w5735, w5736, w5737, w5738, w5739, w5740, w5741, w5742, w5743, w5744, w5745, w5746, w5747, w5748, w5749, w5750, w5751, w5752, w5753, w5754, w5755, w5756, w5757, w5758, w5759, w5760, w5761, w5762, w5763, w5764, w5765, w5766, w5767, w5768, w5769, w5770, w5771, w5772, w5773, w5774, w5775, w5776, w5777, w5778, w5779, w5780, w5781, w5782, w5783, w5784, w5785, w5786, w5787, w5788, w5789, w5790, w5791, w5792, w5793, w5794, w5795, w5796, w5797, w5798, w5799, w5800, w5801, w5802, w5803, w5804, w5805, w5806, w5807, w5808, w5809, w5810, w5811, w5812, w5813, w5814, w5815, w5816, w5817, w5818, w5819, w5820, w5821, w5822, w5823, w5824, w5825, w5826, w5827, w5828, w5829, w5830, w5831, w5832, w5833, w5834, w5835, w5836, w5837, w5838, w5839, w5840, w5841, w5842, w5843, w5844, w5845, w5846, w5847, w5848, w5849, w5850, w5851, w5852, w5853, w5854, w5855, w5856, w5857, w5858, w5859, w5860, w5861, w5862, w5863, w5864, w5865, w5866, w5867, w5868, w5869, w5870, w5871, w5872, w5873, w5874, w5875, w5876, w5877, w5878, w5879, w5880, w5881, w5882, w5883, w5884, w5885, w5886, w5887, w5888, w5889, w5890, w5891, w5892, w5893, w5894, w5895, w5896, w5897, w5898, w5899, w5900, w5901, w5902, w5903, w5904, w5905, w5906, w5907, w5908, w5909, w5910, w5911, w5912, w5913, w5914, w5915, w5916, w5917, w5918, w5919, w5920, w5921, w5922, w5923, w5924, w5925, w5926, w5927, w5928, w5929, w5930, w5931, w5932, w5933, w5934, w5935, w5936, w5937, w5938, w5939, w5940, w5941, w5942, w5943, w5944, w5945, w5946, w5947, w5948, w5949, w5950, w5951, w5952, w5953, w5954, w5955, w5956, w5957, w5958, w5959, w5960, w5961, w5962, w5963, w5964, w5965, w5966, w5967, w5968, w5969, w5970, w5971, w5972, w5973, w5974, w5975, w5976, w5977, w5978, w5979, w5980, w5981, w5982, w5983, w5984, w5985, w5986, w5987, w5988, w5989, w5990, w5991, w5992, w5993, w5994, w5995, w5996, w5997, w5998, w5999, w6000, w6001, w6002, w6003, w6004, w6005, w6006, w6007, w6008, w6009, w6010, w6011, w6012, w6013, w6014, w6015, w6016, w6017, w6018, w6019, w6020, w6021, w6022, w6023, w6024, w6025, w6026, w6027, w6028, w6029, w6030, w6031, w6032, w6033, w6034, w6035, w6036, w6037, w6038, w6039, w6040, w6041, w6042, w6043, w6044, w6045, w6046, w6047, w6048, w6049, w6050, w6051, w6052, w6053, w6054, w6055, w6056, w6057, w6058, w6059, w6060, w6061, w6062, w6063, w6064, w6065, w6066, w6067, w6068, w6069, w6070, w6071, w6072, w6073, w6074, w6075, w6076, w6077, w6078, w6079, w6080, w6081, w6082, w6083, w6084, w6085, w6086, w6087, w6088, w6089, w6090, w6091, w6092, w6093, w6094, w6095, w6096, w6097, w6098, w6099, w6100, w6101, w6102, w6103, w6104, w6105, w6106, w6107, w6108, w6109, w6110, w6111, w6112, w6113, w6114, w6115, w6116, w6117, w6118, w6119, w6120, w6121, w6122, w6123, w6124, w6125, w6126, w6127, w6128, w6129, w6130, w6131, w6132, w6133, w6134, w6135, w6136, w6137, w6138, w6139, w6140, w6141, w6142, w6143, w6144, w6145, w6146, w6147, w6148, w6149, w6150, w6151, w6152, w6153, w6154, w6155, w6156, w6157, w6158, w6159, w6160, w6161, w6162, w6163, w6164, w6165, w6166, w6167, w6168, w6169, w6170, w6171, w6172, w6173, w6174, w6175, w6176, w6177, w6178, w6179, w6180, w6181, w6182, w6183, w6184, w6185, w6186, w6187, w6188, w6189, w6190, w6191, w6192, w6193, w6194, w6195, w6196, w6197, w6198, w6199, w6200, w6201, w6202, w6203, w6204, w6205, w6206, w6207, w6208, w6209, w6210, w6211, w6212, w6213, w6214, w6215, w6216, w6217, w6218, w6219, w6220, w6221, w6222, w6223, w6224, w6225, w6226, w6227, w6228, w6229, w6230, w6231, w6232, w6233, w6234, w6235, w6236, w6237, w6238, w6239, w6240, w6241, w6242, w6243, w6244, w6245, w6246, w6247, w6248, w6249, w6250, w6251, w6252, w6253, w6254, w6255, w6256, w6257, w6258, w6259, w6260, w6261, w6262, w6263, w6264, w6265, w6266, w6267, w6268, w6269, w6270, w6271, w6272, w6273, w6274, w6275, w6276, w6277, w6278, w6279, w6280, w6281, w6282, w6283, w6284, w6285, w6286, w6287, w6288, w6289, w6290, w6291, w6292, w6293, w6294, w6295, w6296, w6297, w6298, w6299, w6300, w6301, w6302, w6303, w6304, w6305, w6306, w6307, w6308, w6309, w6310, w6311, w6312, w6313, w6314, w6315, w6316, w6317, w6318, w6319, w6320, w6321, w6322, w6323, w6324, w6325, w6326, w6327, w6328, w6329, w6330, w6331, w6332, w6333, w6334, w6335, w6336, w6337, w6338, w6339, w6340, w6341, w6342, w6343, w6344, w6345, w6346, w6347, w6348, w6349, w6350, w6351, w6352, w6353, w6354, w6355, w6356, w6357, w6358, w6359, w6360, w6361, w6362, w6363, w6364, w6365, w6366, w6367, w6368, w6369, w6370, w6371, w6372, w6373, w6374, w6375, w6376, w6377, w6378, w6379, w6380, w6381, w6382, w6383, w6384, w6385, w6386, w6387, w6388, w6389, w6390, w6391, w6392, w6393, w6394, w6395, w6396, w6397, w6398, w6399, w6400, w6401, w6402, w6403, w6404, w6405, w6406, w6407, w6408, w6409, w6410, w6411, w6412, w6413, w6414, w6415, w6416, w6417, w6418, w6419, w6420, w6421, w6422, w6423, w6424, w6425, w6426, w6427, w6428, w6429, w6430, w6431, w6432, w6433, w6434, w6435, w6436, w6437, w6438, w6439, w6440, w6441, w6442, w6443, w6444, w6445, w6446, w6447, w6448, w6449, w6450, w6451, w6452, w6453, w6454, w6455, w6456, w6457, w6458, w6459, w6460, w6461, w6462, w6463, w6464, w6465, w6466, w6467, w6468, w6469, w6470, w6471, w6472, w6473, w6474, w6475, w6476, w6477, w6478, w6479, w6480, w6481, w6482, w6483, w6484, w6485, w6486, w6487, w6488, w6489, w6490, w6491, w6492, w6493, w6494, w6495, w6496, w6497, w6498, w6499, w6500, w6501, w6502, w6503, w6504, w6505, w6506, w6507, w6508, w6509, w6510, w6511, w6512, w6513, w6514, w6515, w6516, w6517, w6518, w6519, w6520, w6521, w6522, w6523, w6524, w6525, w6526, w6527, w6528, w6529, w6530, w6531, w6532, w6533, w6534, w6535, w6536, w6537, w6538, w6539, w6540, w6541, w6542, w6543, w6544, w6545, w6546, w6547, w6548, w6549, w6550, w6551, w6552, w6553, w6554, w6555, w6556, w6557, w6558, w6559, w6560, w6561, w6562, w6563, w6564, w6565, w6566, w6567, w6568, w6569, w6570, w6571, w6572, w6573, w6574, w6575, w6576, w6577, w6578, w6579, w6580, w6581, w6582, w6583, w6584, w6585, w6586, w6587, w6588, w6589, w6590, w6591, w6592, w6593, w6594, w6595, w6596, w6597, w6598, w6599, w6600, w6601, w6602, w6603, w6604, w6605, w6606, w6607, w6608, w6609, w6610, w6611, w6612, w6613, w6614, w6615, w6616, w6617, w6618, w6619, w6620, w6621, w6622, w6623, w6624, w6625, w6626, w6627, w6628, w6629, w6630, w6631, w6632, w6633, w6634, w6635, w6636, w6637, w6638, w6639, w6640, w6641, w6642, w6643, w6644, w6645, w6646, w6647, w6648, w6649, w6650, w6651, w6652, w6653, w6654, w6655, w6656, w6657, w6658, w6659, w6660, w6661, w6662, w6663, w6664, w6665, w6666, w6667, w6668, w6669, w6670, w6671, w6672, w6673, w6674, w6675, w6676, w6677, w6678, w6679, w6680, w6681, w6682, w6683, w6684, w6685, w6686, w6687, w6688, w6689, w6690, w6691, w6692, w6693, w6694, w6695, w6696, w6697, w6698, w6699, w6700, w6701, w6702, w6703, w6704, w6705, w6706, w6707, w6708, w6709, w6710, w6711, w6712, w6713, w6714, w6715, w6716, w6717, w6718, w6719, w6720, w6721, w6722, w6723, w6724, w6725, w6726, w6727, w6728, w6729, w6730, w6731, w6732, w6733, w6734, w6735, w6736, w6737, w6738, w6739, w6740, w6741, w6742, w6743, w6744, w6745, w6746, w6747, w6748, w6749, w6750, w6751, w6752, w6753, w6754, w6755, w6756, w6757, w6758, w6759, w6760, w6761, w6762, w6763, w6764, w6765, w6766, w6767, w6768, w6769, w6770, w6771, w6772, w6773, w6774, w6775, w6776, w6777, w6778, w6779, w6780, w6781, w6782, w6783, w6784, w6785, w6786, w6787, w6788, w6789, w6790, w6791, w6792, w6793, w6794, w6795, w6796, w6797, w6798, w6799, w6800, w6801, w6802, w6803, w6804, w6805, w6806, w6807, w6808, w6809, w6810, w6811, w6812, w6813, w6814, w6815, w6816, w6817, w6818, w6819, w6820, w6821, w6822, w6823, w6824, w6825, w6826, w6827, w6828, w6829, w6830, w6831, w6832, w6833, w6834, w6835, w6836, w6837, w6838, w6839, w6840, w6841, w6842, w6843, w6844, w6845, w6846, w6847, w6848, w6849, w6850, w6851, w6852, w6853, w6854, w6855, w6856, w6857, w6858, w6859, w6860, w6861, w6862, w6863, w6864, w6865, w6866, w6867, w6868, w6869, w6870, w6871, w6872, w6873, w6874, w6875, w6876, w6877, w6878, w6879, w6880, w6881, w6882, w6883, w6884, w6885, w6886, w6887, w6888, w6889, w6890, w6891, w6892, w6893, w6894, w6895, w6896, w6897, w6898, w6899, w6900, w6901, w6902, w6903, w6904, w6905, w6906, w6907, w6908, w6909, w6910, w6911, w6912, w6913, w6914, w6915, w6916, w6917, w6918, w6919, w6920, w6921, w6922, w6923, w6924, w6925, w6926, w6927, w6928, w6929, w6930, w6931, w6932, w6933, w6934, w6935, w6936, w6937, w6938, w6939, w6940, w6941, w6942, w6943, w6944, w6945, w6946, w6947, w6948, w6949, w6950, w6951, w6952, w6953, w6954, w6955, w6956, w6957, w6958, w6959, w6960, w6961, w6962, w6963, w6964, w6965, w6966, w6967, w6968, w6969, w6970, w6971, w6972, w6973, w6974, w6975, w6976, w6977, w6978, w6979, w6980, w6981, w6982, w6983, w6984, w6985, w6986, w6987, w6988, w6989, w6990, w6991, w6992, w6993, w6994, w6995, w6996, w6997, w6998, w6999, w7000, w7001, w7002, w7003, w7004, w7005, w7006, w7007, w7008, w7009, w7010, w7011, w7012, w7013, w7014, w7015, w7016, w7017, w7018, w7019, w7020, w7021, w7022, w7023, w7024, w7025, w7026, w7027, w7028, w7029, w7030, w7031, w7032, w7033, w7034, w7035, w7036, w7037, w7038, w7039, w7040, w7041, w7042, w7043, w7044, w7045, w7046, w7047, w7048, w7049, w7050, w7051, w7052, w7053, w7054, w7055, w7056, w7057, w7058, w7059, w7060, w7061, w7062, w7063, w7064, w7065, w7066, w7067, w7068, w7069, w7070, w7071, w7072, w7073, w7074, w7075, w7076, w7077, w7078, w7079, w7080, w7081, w7082, w7083, w7084, w7085, w7086, w7087, w7088, w7089, w7090, w7091, w7092, w7093, w7094, w7095, w7096, w7097, w7098, w7099, w7100, w7101, w7102, w7103, w7104, w7105, w7106, w7107, w7108, w7109, w7110, w7111, w7112, w7113, w7114, w7115, w7116, w7117, w7118, w7119, w7120, w7121, w7122, w7123, w7124, w7125, w7126, w7127, w7128, w7129, w7130, w7131, w7132, w7133, w7134, w7135, w7136, w7137, w7138, w7139, w7140, w7141, w7142;
assign w0 = ~pi0055 & ~pi0057;
assign w1 = ~pi0056 & ~pi0062;
assign w2 = w0 & w1;
assign w3 = ~pi0059 & ~pi0299;
assign w4 = w2 & w3;
assign w5 = (pi0221 & ~w2) | (pi0221 & w6515) | (~w2 & w6515);
assign w6 = w2 & w6516;
assign w7 = ~w5 & ~w6;
assign w8 = (pi0215 & ~w2) | (pi0215 & w6517) | (~w2 & w6517);
assign w9 = w2 & w6518;
assign w10 = ~w8 & ~w9;
assign w11 = w7 & w10;
assign w12 = (pi0216 & ~w2) | (pi0216 & w6519) | (~w2 & w6519);
assign w13 = w2 & w6520;
assign w14 = ~w12 & ~w13;
assign w15 = w11 & w14;
assign w16 = pi0105 & pi0228;
assign w17 = (~w16 & ~w2) | (~w16 & w6521) | (~w2 & w6521);
assign w18 = pi0228 & w17;
assign w19 = ~pi0035 & ~pi0070;
assign w20 = ~pi0095 & w19;
assign w21 = ~pi0089 & ~pi0108;
assign w22 = w20 & w21;
assign w23 = ~pi0039 & ~pi0048;
assign w24 = w20 & w6329;
assign w25 = ~pi0075 & ~pi0100;
assign w26 = ~pi0094 & w25;
assign w27 = ~pi0074 & ~pi0096;
assign w28 = ~pi0097 & w27;
assign w29 = w26 & w28;
assign w30 = ~pi0032 & ~pi0038;
assign w31 = ~pi0050 & w30;
assign w32 = ~pi0049 & ~pi0076;
assign w33 = w31 & w32;
assign w34 = w29 & w33;
assign w35 = w24 & w34;
assign w36 = ~pi0053 & ~pi0054;
assign w37 = ~pi0045 & ~pi0106;
assign w38 = w36 & w37;
assign w39 = w2 & w38;
assign w40 = ~pi0063 & ~pi0107;
assign w41 = ~pi0064 & w40;
assign w42 = ~pi0046 & ~pi0059;
assign w43 = ~pi0060 & ~pi0061;
assign w44 = w42 & w43;
assign w45 = w41 & w44;
assign w46 = w39 & w45;
assign w47 = ~pi0065 & ~pi0102;
assign w48 = ~pi0068 & ~pi0081;
assign w49 = ~pi0040 & w48;
assign w50 = w47 & w49;
assign w51 = w46 & w50;
assign w52 = w35 & w51;
assign w53 = ~pi0088 & ~pi0110;
assign w54 = ~pi0047 & ~pi0104;
assign w55 = w53 & w54;
assign w56 = ~pi0036 & ~pi0091;
assign w57 = w55 & w56;
assign w58 = ~pi0092 & ~pi0098;
assign w59 = ~pi0058 & ~pi0093;
assign w60 = w58 & w59;
assign w61 = ~pi0073 & ~pi0090;
assign w62 = w60 & w61;
assign w63 = w57 & w62;
assign w64 = ~pi0077 & ~pi0086;
assign w65 = ~pi0072 & ~pi0111;
assign w66 = ~pi0087 & ~pi0103;
assign w67 = w65 & w66;
assign w68 = w64 & w67;
assign w69 = ~pi0067 & ~pi0069;
assign w70 = ~pi0109 & w69;
assign w71 = ~pi0071 & ~pi0085;
assign w72 = w70 & w71;
assign w73 = w68 & w72;
assign w74 = w63 & w73;
assign w75 = ~pi0066 & ~pi0084;
assign w76 = ~pi0083 & w75;
assign w77 = pi0051 & ~pi0082;
assign w78 = w76 & w77;
assign w79 = w74 & w78;
assign w80 = w52 & w79;
assign w81 = ~pi0051 & ~pi0082;
assign w82 = w75 & w81;
assign w83 = ~pi0040 & ~pi0083;
assign w84 = w48 & w83;
assign w85 = w82 & w84;
assign w86 = w71 & w85;
assign w87 = w64 & w70;
assign w88 = w67 & w87;
assign w89 = w86 & w88;
assign w90 = w55 & w6330;
assign w91 = w46 & w47;
assign w92 = w35 & w91;
assign w93 = ~pi0092 & pi0098;
assign w94 = w59 & w93;
assign w95 = w90 & w94;
assign w96 = w89 & w95;
assign w97 = w92 & w96;
assign w98 = ~w80 & ~w97;
assign w99 = w47 & w85;
assign w100 = w74 & w99;
assign w101 = w39 & w41;
assign w102 = ~pi0060 & pi0061;
assign w103 = w42 & w102;
assign w104 = w39 & w6331;
assign w105 = w35 & w104;
assign w106 = w100 & w105;
assign w107 = w63 & w67;
assign w108 = pi0109 & w64;
assign w109 = w69 & w108;
assign w110 = w86 & w109;
assign w111 = w107 & w110;
assign w112 = w92 & w111;
assign w113 = w63 & w87;
assign w114 = ~pi0087 & pi0103;
assign w115 = w65 & w114;
assign w116 = w85 & w6332;
assign w117 = w113 & w116;
assign w118 = w92 & w117;
assign w119 = w24 & w46;
assign w120 = pi0049 & ~pi0076;
assign w121 = w29 & w6333;
assign w122 = w119 & w121;
assign w123 = w100 & w122;
assign w124 = ~pi0064 & w44;
assign w125 = w39 & w124;
assign w126 = ~pi0063 & pi0107;
assign w127 = w125 & w126;
assign w128 = w35 & w127;
assign w129 = w100 & w128;
assign w130 = ~pi0045 & pi0106;
assign w131 = w36 & w130;
assign w132 = w45 & w6334;
assign w133 = w35 & w132;
assign w134 = w100 & w133;
assign w135 = ~pi0072 & w66;
assign w136 = w66 & w6522;
assign w137 = w85 & w6523;
assign w138 = w92 & w6335;
assign w139 = w60 & w6330;
assign w140 = ~pi0088 & pi0110;
assign w141 = w54 & w140;
assign w142 = w139 & w141;
assign w143 = w92 & w6336;
assign w144 = ~w138 & ~w143;
assign w145 = w92 & w6337;
assign w146 = ~pi0047 & pi0104;
assign w147 = w53 & w146;
assign w148 = pi0088 & ~pi0110;
assign w149 = w54 & w148;
assign w150 = ~w147 & ~w149;
assign w151 = pi0047 & ~pi0104;
assign w152 = w53 & w151;
assign w153 = w150 & ~w152;
assign w154 = w145 & ~w153;
assign w155 = (w82 & w74) | (w82 & w6338) | (w74 & w6338);
assign w156 = pi0071 & ~pi0085;
assign w157 = ~pi0071 & pi0085;
assign w158 = ~w156 & ~w157;
assign w159 = w67 & ~w158;
assign w160 = w87 & w159;
assign w161 = w63 & w160;
assign w162 = ~pi0083 & ~w161;
assign w163 = w52 & ~w162;
assign w164 = w155 & w163;
assign w165 = pi0073 & ~pi0090;
assign w166 = w57 & w6339;
assign w167 = w89 & w166;
assign w168 = w92 & w167;
assign w169 = w67 & w6340;
assign w170 = w63 & w169;
assign w171 = pi0067 & ~pi0069;
assign w172 = w85 & w6341;
assign w173 = w170 & w172;
assign w174 = w92 & w173;
assign w175 = pi0068 & pi0081;
assign w176 = w83 & ~w175;
assign w177 = w82 & w176;
assign w178 = w74 & w177;
assign w179 = w92 & w178;
assign w180 = pi0068 & w179;
assign w181 = ~pi0083 & w74;
assign w182 = ~pi0066 & pi0084;
assign w183 = w81 & w182;
assign w184 = pi0066 & ~pi0084;
assign w185 = w81 & w184;
assign w186 = ~w183 & ~w185;
assign w187 = w74 & w6342;
assign w188 = w52 & w187;
assign w189 = ~w168 & ~w174;
assign w190 = ~w164 & w189;
assign w191 = ~w180 & ~w188;
assign w192 = w190 & w191;
assign w193 = pi0081 & w179;
assign w194 = w35 & w100;
assign w195 = pi0045 & ~pi0106;
assign w196 = w36 & w195;
assign w197 = w45 & w6524;
assign w198 = w100 & w6343;
assign w199 = pi0097 & w27;
assign w200 = w33 & w6344;
assign w201 = w119 & w200;
assign w202 = w100 & w201;
assign w203 = ~pi0074 & pi0096;
assign w204 = ~pi0097 & w203;
assign w205 = w33 & w6345;
assign w206 = w119 & w205;
assign w207 = w100 & w206;
assign w208 = ~w202 & ~w207;
assign w209 = pi0058 & ~pi0093;
assign w210 = w58 & w209;
assign w211 = w90 & w210;
assign w212 = w92 & w6346;
assign w213 = ~w106 & ~w112;
assign w214 = ~w118 & ~w123;
assign w215 = ~w129 & ~w134;
assign w216 = w214 & w215;
assign w217 = w98 & w213;
assign w218 = ~w193 & ~w198;
assign w219 = w208 & ~w212;
assign w220 = w218 & w219;
assign w221 = w216 & w217;
assign w222 = w144 & ~w154;
assign w223 = w221 & w222;
assign w224 = w192 & w220;
assign w225 = w223 & w224;
assign w226 = (pi0166 & ~w2) | (pi0166 & w6347) | (~w2 & w6347);
assign w227 = w2 & w6348;
assign w228 = ~w226 & ~w227;
assign w229 = (pi0161 & ~w2) | (pi0161 & w6349) | (~w2 & w6349);
assign w230 = w2 & w6350;
assign w231 = ~w229 & ~w230;
assign w232 = w228 & w231;
assign w233 = (pi0152 & ~w2) | (pi0152 & w6351) | (~w2 & w6351);
assign w234 = w2 & w6352;
assign w235 = ~w233 & ~w234;
assign w236 = pi0252 & w235;
assign w237 = w232 & w236;
assign w238 = (pi0146 & ~w2) | (pi0146 & w6525) | (~w2 & w6525);
assign w239 = w2 & w6526;
assign w240 = ~w238 & ~w239;
assign w241 = pi0252 & ~w240;
assign w242 = ~w237 & ~w241;
assign w243 = w100 & w119;
assign w244 = w33 & w6527;
assign w245 = ~pi0075 & pi0100;
assign w246 = w244 & w245;
assign w247 = w100 & w6528;
assign w248 = w242 & w247;
assign w249 = w232 & w235;
assign w250 = ~pi0250 & w240;
assign w251 = ~w249 & w250;
assign w252 = (pi0129 & w249) | (pi0129 & w6529) | (w249 & w6529);
assign w253 = pi1085 & pi1087;
assign w254 = pi0957 & pi1086;
assign w255 = ~pi0833 & w253;
assign w256 = w254 & w255;
assign w257 = (pi0950 & ~w255) | (pi0950 & w6530) | (~w255 & w6530);
assign w258 = pi0824 & pi1086;
assign w259 = w257 & w258;
assign w260 = ~pi1085 & pi1087;
assign w261 = pi0829 & pi1086;
assign w262 = ~w260 & w261;
assign w263 = w257 & w262;
assign w264 = ~w259 & ~w263;
assign w265 = ~pi1087 & ~w264;
assign w266 = w251 & ~w265;
assign w267 = ~w252 & ~w266;
assign w268 = w248 & w267;
assign w269 = w38 & w45;
assign w270 = w35 & w269;
assign w271 = w100 & w270;
assign w272 = pi0056 & ~pi0062;
assign w273 = w0 & w272;
assign w274 = w271 & w273;
assign w275 = pi0064 & w40;
assign w276 = w44 & w275;
assign w277 = w39 & w276;
assign w278 = w100 & w6353;
assign w279 = ~w274 & ~w278;
assign w280 = w23 & w46;
assign w281 = w20 & w34;
assign w282 = w280 & w281;
assign w283 = w100 & w282;
assign w284 = ~pi0089 & pi0108;
assign w285 = w283 & w284;
assign w286 = w22 & w39;
assign w287 = w34 & w286;
assign w288 = ~pi0039 & pi0048;
assign w289 = w45 & w288;
assign w290 = w287 & w289;
assign w291 = w100 & w290;
assign w292 = ~w285 & ~w291;
assign w293 = w279 & w292;
assign w294 = ~pi0111 & w66;
assign w295 = w66 & w6531;
assign w296 = w85 & w6532;
assign w297 = w113 & w296;
assign w298 = w92 & w297;
assign w299 = pi0036 & ~pi0091;
assign w300 = w62 & w6533;
assign w301 = w92 & w6354;
assign w302 = ~w298 & ~w301;
assign w303 = w293 & w302;
assign w304 = ~w268 & w303;
assign w305 = w225 & w304;
assign w306 = pi0094 & w25;
assign w307 = w33 & w6355;
assign w308 = w119 & w307;
assign w309 = w100 & w308;
assign w310 = ~pi0056 & pi0062;
assign w311 = w0 & w310;
assign w312 = w45 & w6356;
assign w313 = w35 & w312;
assign w314 = w100 & w313;
assign w315 = ~pi0049 & pi0076;
assign w316 = w29 & w6534;
assign w317 = w100 & w6357;
assign w318 = ~w309 & ~w314;
assign w319 = ~w317 & w318;
assign w320 = pi0087 & ~pi0103;
assign w321 = w65 & w320;
assign w322 = w85 & w6358;
assign w323 = w113 & w322;
assign w324 = w92 & w323;
assign w325 = pi0040 & ~pi0083;
assign w326 = w48 & w325;
assign w327 = w82 & w326;
assign w328 = w74 & w327;
assign w329 = w92 & w328;
assign w330 = ~w324 & ~w329;
assign w331 = ~pi0067 & pi0069;
assign w332 = w85 & w6359;
assign w333 = w170 & w332;
assign w334 = w92 & w333;
assign w335 = w49 & w82;
assign w336 = pi0065 & pi0102;
assign w337 = ~w47 & ~w336;
assign w338 = w335 & w337;
assign w339 = w46 & w338;
assign w340 = w35 & w339;
assign w341 = w181 & w340;
assign w342 = ~w334 & ~w341;
assign w343 = w330 & w342;
assign w344 = w319 & w343;
assign w345 = pi0089 & ~pi0108;
assign w346 = w283 & w345;
assign w347 = pi0039 & ~pi0048;
assign w348 = w45 & w347;
assign w349 = w287 & w348;
assign w350 = w100 & w349;
assign w351 = ~w346 & ~w350;
assign w352 = pi0063 & ~pi0107;
assign w353 = w125 & w352;
assign w354 = w35 & w353;
assign w355 = w100 & w354;
assign w356 = pi0050 & w30;
assign w357 = w29 & w6360;
assign w358 = w119 & w357;
assign w359 = w100 & w358;
assign w360 = ~w355 & ~w359;
assign w361 = ~pi0036 & pi0091;
assign w362 = w62 & w6361;
assign w363 = w89 & w362;
assign w364 = w92 & w363;
assign w365 = w360 & ~w364;
assign w366 = w351 & w365;
assign w367 = w344 & w366;
assign w368 = w63 & w6362;
assign w369 = ~pi0077 & pi0086;
assign w370 = pi0077 & ~pi0086;
assign w371 = ~w369 & ~w370;
assign w372 = w85 & w6535;
assign w373 = w92 & w6363;
assign w374 = pi0092 & ~pi0098;
assign w375 = w59 & w374;
assign w376 = w90 & w375;
assign w377 = w92 & w6364;
assign w378 = ~w373 & ~w377;
assign w379 = ~pi0051 & pi0082;
assign w380 = w76 & w379;
assign w381 = w74 & w380;
assign w382 = w52 & w381;
assign w383 = w21 & w34;
assign w384 = w280 & w383;
assign w385 = pi0095 & w19;
assign w386 = w85 & w6365;
assign w387 = w74 & w386;
assign w388 = w384 & w387;
assign w389 = ~w382 & ~w388;
assign w390 = pi0032 & ~pi0038;
assign w391 = w29 & w6537;
assign w392 = w100 & w6538;
assign w393 = pi0053 & pi0054;
assign w394 = w37 & ~w393;
assign w395 = w2 & w394;
assign w396 = pi0053 & w45;
assign w397 = w395 & w396;
assign w398 = w35 & w397;
assign w399 = w100 & w398;
assign w400 = pi0055 & ~pi0057;
assign w401 = w1 & w400;
assign w402 = w45 & w6366;
assign w403 = w35 & w402;
assign w404 = w100 & w403;
assign w405 = ~w399 & ~w404;
assign w406 = ~pi0035 & pi0070;
assign w407 = ~pi0095 & w406;
assign w408 = w85 & w6367;
assign w409 = w74 & w408;
assign w410 = w384 & w409;
assign w411 = pi0060 & ~pi0061;
assign w412 = w42 & w411;
assign w413 = w39 & w6368;
assign w414 = w35 & w413;
assign w415 = w100 & w414;
assign w416 = ~w410 & ~w415;
assign w417 = w405 & w416;
assign w418 = w389 & ~w392;
assign w419 = ~w248 & w418;
assign w420 = w378 & w417;
assign w421 = w419 & w420;
assign w422 = w367 & w421;
assign w423 = ~pi0073 & pi0090;
assign w424 = w57 & w6369;
assign w425 = w89 & w424;
assign w426 = w92 & w425;
assign w427 = ~pi0058 & pi0093;
assign w428 = w58 & w427;
assign w429 = w90 & w428;
assign w430 = w89 & w429;
assign w431 = w92 & w430;
assign w432 = ~w426 & ~w431;
assign w433 = w100 & w384;
assign w434 = pi0035 & ~pi0070;
assign w435 = ~pi0095 & w434;
assign w436 = w433 & w435;
assign w437 = w432 & ~w436;
assign w438 = w17 & w437;
assign w439 = w422 & w438;
assign w440 = w305 & w439;
assign w441 = pi0095 & ~pi0479;
assign w442 = ~w207 & ~w441;
assign w443 = ~w440 & w6370;
assign w444 = w92 & w6371;
assign w445 = w370 & w444;
assign w446 = pi0074 & ~pi0096;
assign w447 = ~pi0097 & w446;
assign w448 = w33 & w6539;
assign w449 = w243 & w448;
assign w450 = ~w445 & ~w449;
assign w451 = w225 & w450;
assign w452 = pi0075 & ~pi0100;
assign w453 = w244 & w452;
assign w454 = w100 & w6540;
assign w455 = ~w247 & ~w454;
assign w456 = ~w301 & ~w377;
assign w457 = w455 & w456;
assign w458 = w293 & w457;
assign w459 = w369 & w444;
assign w460 = ~pi0032 & pi0038;
assign w461 = w29 & w6541;
assign w462 = w243 & w461;
assign w463 = ~w459 & ~w462;
assign w464 = ~pi0055 & pi0057;
assign w465 = w1 & w464;
assign w466 = w271 & w465;
assign w467 = w389 & ~w466;
assign w468 = ~w298 & ~w364;
assign w469 = w35 & w101;
assign w470 = w100 & w469;
assign w471 = ~pi0046 & pi0059;
assign w472 = w43 & w471;
assign w473 = w470 & w472;
assign w474 = w468 & ~w473;
assign w475 = w467 & w474;
assign w476 = w463 & w475;
assign w477 = w458 & w476;
assign w478 = ~w36 & w45;
assign w479 = w395 & w478;
assign w480 = ~w132 & ~w479;
assign w481 = w194 & ~w480;
assign w482 = w194 & w6372;
assign w483 = pi0046 & ~pi0059;
assign w484 = w43 & w483;
assign w485 = w470 & w484;
assign w486 = w360 & w432;
assign w487 = ~w485 & w486;
assign w488 = w351 & ~w482;
assign w489 = w487 & w488;
assign w490 = w344 & w489;
assign w491 = w477 & w490;
assign w492 = w451 & w491;
assign w493 = (pi0210 & ~w2) | (pi0210 & w6542) | (~w2 & w6542);
assign w494 = w2 & w6543;
assign w495 = ~w493 & ~w494;
assign w496 = ~pi0841 & w495;
assign w497 = w392 & ~w496;
assign w498 = ~w436 & ~w497;
assign w499 = pi0225 & ~w498;
assign w500 = w406 & w6544;
assign w501 = w433 & w500;
assign w502 = (w240 & ~w232) | (w240 & w6545) | (~w232 & w6545);
assign w503 = w257 & w6546;
assign w504 = w202 & w503;
assign w505 = w257 & w6547;
assign w506 = w207 & w505;
assign w507 = ~w504 & ~w506;
assign w508 = w495 & ~w502;
assign w509 = (w508 & ~w507) | (w508 & w6548) | (~w507 & w6548);
assign w510 = w405 & ~w415;
assign w511 = ~w501 & w510;
assign w512 = ~w499 & w511;
assign w513 = ~w509 & w512;
assign w514 = (w513 & w492) | (w513 & w6373) | (w492 & w6373);
assign w515 = w443 & ~w514;
assign w516 = (pi0234 & w207) | (pi0234 & w6549) | (w207 & w6549);
assign w517 = ~w440 & w6374;
assign w518 = (~pi0153 & w440) | (~pi0153 & w6375) | (w440 & w6375);
assign w519 = ~w517 & ~w518;
assign w520 = ~w515 & w519;
assign w521 = w15 & ~w520;
assign w522 = w11 & ~w14;
assign w523 = w11 & w6550;
assign w524 = ~w7 & w10;
assign w525 = w14 & w524;
assign w526 = w524 & w6551;
assign w527 = ~w11 & ~w526;
assign w528 = ~w526 & w6552;
assign w529 = pi0929 & w526;
assign w530 = ~pi0332 & ~w523;
assign w531 = ~w529 & w530;
assign w532 = ~w528 & w531;
assign w533 = ~w521 & w532;
assign w534 = ~w440 & w6440;
assign w535 = (~pi0154 & w440) | (~pi0154 & w6441) | (w440 & w6441);
assign w536 = ~w534 & ~w535;
assign w537 = w15 & ~w536;
assign w538 = w11 & w6553;
assign w539 = ~w526 & w6554;
assign w540 = pi0939 & w526;
assign w541 = ~w538 & ~w540;
assign w542 = ~w539 & w541;
assign w543 = ~w537 & w542;
assign w544 = ~w440 & w6442;
assign w545 = (~pi0151 & w440) | (~pi0151 & w6443) | (w440 & w6443);
assign w546 = ~w544 & ~w545;
assign w547 = w15 & ~w546;
assign w548 = w11 & w6555;
assign w549 = ~w526 & w6556;
assign w550 = pi0927 & w526;
assign w551 = ~w548 & ~w550;
assign w552 = ~w549 & w551;
assign w553 = ~w547 & w552;
assign w554 = ~w440 & w6444;
assign w555 = ~w440 & w6557;
assign w556 = (~w440 & w6445) | (~w440 & w6446) | (w6445 & w6446);
assign w557 = ~w554 & w556;
assign w558 = ~w555 & w557;
assign w559 = w11 & w6558;
assign w560 = ~w526 & w6559;
assign w561 = pi0944 & w526;
assign w562 = ~w559 & ~w561;
assign w563 = ~w560 & w562;
assign w564 = ~w558 & w563;
assign w565 = ~w440 & w6447;
assign w566 = ~w440 & w6560;
assign w567 = (~w440 & w6448) | (~w440 & w6449) | (w6448 & w6449);
assign w568 = ~w565 & w567;
assign w569 = ~w566 & w568;
assign w570 = w11 & w6561;
assign w571 = ~w526 & w6562;
assign w572 = pi0932 & w526;
assign w573 = ~w570 & ~w572;
assign w574 = ~w571 & w573;
assign w575 = ~w569 & w574;
assign w576 = ~w440 & w6450;
assign w577 = ~w440 & w6563;
assign w578 = (~w440 & w6451) | (~w440 & w6452) | (w6451 & w6452);
assign w579 = ~w576 & w578;
assign w580 = ~w577 & w579;
assign w581 = w11 & w6564;
assign w582 = ~w526 & w6565;
assign w583 = pi0935 & w526;
assign w584 = ~w581 & ~w583;
assign w585 = ~w582 & w584;
assign w586 = ~w580 & w585;
assign w587 = ~w440 & w6453;
assign w588 = ~w440 & w6566;
assign w589 = (~w440 & w6454) | (~w440 & w6455) | (w6454 & w6455);
assign w590 = ~w587 & w589;
assign w591 = ~w588 & w590;
assign w592 = w11 & w6567;
assign w593 = ~w526 & w6568;
assign w594 = pi0921 & w526;
assign w595 = ~w592 & ~w594;
assign w596 = ~w593 & w595;
assign w597 = ~w591 & w596;
assign w598 = ~w440 & w6456;
assign w599 = ~w440 & w6569;
assign w600 = (~w440 & w6457) | (~w440 & w6458) | (w6457 & w6458);
assign w601 = ~w598 & w600;
assign w602 = ~w599 & w601;
assign w603 = w11 & w6570;
assign w604 = ~w526 & w6571;
assign w605 = pi0920 & w526;
assign w606 = ~w603 & ~w605;
assign w607 = ~w604 & w606;
assign w608 = ~w602 & w607;
assign w609 = ~w440 & w6459;
assign w610 = ~w440 & w6572;
assign w611 = (~w440 & w6460) | (~w440 & w6461) | (w6460 & w6461);
assign w612 = ~w609 & w611;
assign w613 = ~w610 & w612;
assign w614 = w11 & w6573;
assign w615 = ~w526 & w6574;
assign w616 = pi0940 & w526;
assign w617 = ~w614 & ~w616;
assign w618 = ~w615 & w617;
assign w619 = ~w613 & w618;
assign w620 = ~w440 & w6462;
assign w621 = ~w440 & w6575;
assign w622 = (~w440 & w6463) | (~w440 & w6464) | (w6463 & w6464);
assign w623 = ~w620 & w622;
assign w624 = ~w621 & w623;
assign w625 = w11 & w6576;
assign w626 = ~w526 & w6577;
assign w627 = pi0933 & w526;
assign w628 = ~w625 & ~w627;
assign w629 = ~w626 & w628;
assign w630 = ~w624 & w629;
assign w631 = ~w440 & w6465;
assign w632 = ~w440 & w6578;
assign w633 = (~w440 & w6466) | (~w440 & w6467) | (w6466 & w6467);
assign w634 = ~w631 & w633;
assign w635 = ~w632 & w634;
assign w636 = w11 & w6579;
assign w637 = ~w526 & w6580;
assign w638 = pi0928 & w526;
assign w639 = ~w636 & ~w638;
assign w640 = ~w637 & w639;
assign w641 = ~w635 & w640;
assign w642 = ~w440 & w6468;
assign w643 = ~w440 & w6581;
assign w644 = (~w440 & w6469) | (~w440 & w6470) | (w6469 & w6470);
assign w645 = ~w642 & w644;
assign w646 = ~w643 & w645;
assign w647 = w11 & w6582;
assign w648 = ~w526 & w6583;
assign w649 = pi0938 & w526;
assign w650 = ~w647 & ~w649;
assign w651 = ~w648 & w650;
assign w652 = ~w646 & w651;
assign w653 = ~w440 & w6471;
assign w654 = ~w440 & w6584;
assign w655 = (~w440 & w6472) | (~w440 & w6473) | (w6472 & w6473);
assign w656 = ~w653 & w655;
assign w657 = ~w654 & w656;
assign w658 = w11 & w6585;
assign w659 = ~w526 & w6586;
assign w660 = pi0930 & w526;
assign w661 = ~w658 & ~w660;
assign w662 = ~w659 & w661;
assign w663 = ~w657 & w662;
assign w664 = ~pi0252 & ~pi0995;
assign w665 = pi0835 & pi0984;
assign w666 = ~pi0287 & ~pi0979;
assign w667 = ~w665 & w666;
assign w668 = ~w664 & w667;
assign w669 = w350 & ~w668;
assign w670 = ~w346 & ~w355;
assign w671 = ~w669 & w670;
assign w672 = w319 & w467;
assign w673 = w671 & w672;
assign w674 = ~pi0841 & w431;
assign w675 = ~w426 & ~w449;
assign w676 = ~w334 & ~w485;
assign w677 = w350 & w524;
assign w678 = w350 & w6587;
assign w679 = w350 & w6588;
assign w680 = ~pi0332 & ~pi0468;
assign w681 = w2 & w6387;
assign w682 = ~pi0961 & ~pi0969;
assign w683 = ~pi0971 & ~pi0974;
assign w684 = ~pi0977 & w683;
assign w685 = w682 & w684;
assign w686 = w681 & w685;
assign w687 = (~pi0970 & ~w2) | (~pi0970 & w6474) | (~w2 & w6474);
assign w688 = ~pi0960 & ~pi0963;
assign w689 = ~pi0972 & ~pi0975;
assign w690 = ~pi0978 & w689;
assign w691 = w688 & w690;
assign w692 = w687 & w691;
assign w693 = w680 & ~w686;
assign w694 = ~w692 & w693;
assign w695 = (pi0947 & ~w2) | (pi0947 & w6388) | (~w2 & w6388);
assign w696 = w2 & w6389;
assign w697 = ~w695 & ~w696;
assign w698 = ~pi0614 & ~pi0616;
assign w699 = ~pi0642 & w698;
assign w700 = w698 & w6589;
assign w701 = ~w680 & w700;
assign w702 = (~w701 & w697) | (~w701 & w6590) | (w697 & w6590);
assign w703 = (pi0907 & ~w2) | (pi0907 & w6475) | (~w2 & w6475);
assign w704 = w2 & w6476;
assign w705 = ~w703 & ~w704;
assign w706 = ~pi0661 & ~pi0662;
assign w707 = ~pi0681 & w706;
assign w708 = w706 & w6591;
assign w709 = ~w680 & w708;
assign w710 = (~w709 & w705) | (~w709 & w6592) | (w705 & w6592);
assign w711 = ~w694 & w6593;
assign w712 = pi0835 & ~w264;
assign w713 = ~w711 & w712;
assign w714 = ~w11 & ~w525;
assign w715 = (w350 & ~w713) | (w350 & w6594) | (~w713 & w6594);
assign w716 = ~pi0041 & ~pi0044;
assign w717 = ~pi0101 & w716;
assign w718 = w716 & w6595;
assign w719 = ~pi0113 & ~pi0116;
assign w720 = w718 & w719;
assign w721 = ~pi0114 & ~pi0115;
assign w722 = w718 & w6596;
assign w723 = ~pi0042 & w722;
assign w724 = ~pi0043 & ~pi0052;
assign w725 = w722 & w6597;
assign w726 = w502 & ~w725;
assign w727 = w502 & w6598;
assign w728 = w248 & ~w727;
assign w729 = w330 & ~w341;
assign w730 = ~w462 & ~w674;
assign w731 = w729 & w730;
assign w732 = w675 & w676;
assign w733 = w731 & w732;
assign w734 = w498 & ~w679;
assign w735 = w733 & w734;
assign w736 = w673 & ~w728;
assign w737 = w735 & w736;
assign w738 = ~w715 & w737;
assign w739 = w305 & w738;
assign w740 = pi0232 & w680;
assign w741 = pi0332 & w345;
assign w742 = w283 & w741;
assign w743 = pi0287 & w350;
assign w744 = ~w485 & ~w501;
assign w745 = ~w742 & ~w743;
assign w746 = w744 & w745;
assign w747 = ~w4 & w740;
assign w748 = (w747 & ~w243) | (w747 & w6599) | (~w243 & w6599);
assign w749 = w746 & w6390;
assign w750 = w4 & w740;
assign w751 = (w750 & ~w243) | (w750 & w6600) | (~w243 & w6600);
assign w752 = w746 & w751;
assign w753 = w746 & w6391;
assign w754 = ~w749 & ~w753;
assign w755 = (pi0197 & ~w2) | (pi0197 & w6601) | (~w2 & w6601);
assign w756 = w2 & w6602;
assign w757 = ~w755 & ~w756;
assign w758 = w746 & w6392;
assign w759 = w746 & w6393;
assign w760 = ~w758 & ~w759;
assign w761 = w746 & w6394;
assign w762 = w746 & w6395;
assign w763 = ~w761 & ~w762;
assign w764 = ~w754 & ~w757;
assign w765 = ~w760 & ~w763;
assign w766 = w764 & w765;
assign w767 = w112 & ~w766;
assign w768 = (w378 & w766) | (w378 & w6477) | (w766 & w6477);
assign w769 = ~w711 & w6478;
assign w770 = ~w263 & w769;
assign w771 = w350 & w1854;
assign w772 = w770 & w771;
assign w773 = w417 & w6603;
assign w774 = w474 & w676;
assign w775 = w773 & w774;
assign w776 = ~w454 & ~w466;
assign w777 = w350 & w668;
assign w778 = pi0835 & w503;
assign w779 = w350 & w6604;
assign w780 = ~w711 & w779;
assign w781 = w678 & w780;
assign w782 = ~w242 & w247;
assign w783 = ~pi0252 & ~w502;
assign w784 = (w247 & w266) | (w247 & w6605) | (w266 & w6605);
assign w785 = ~w783 & w784;
assign w786 = w784 & w6606;
assign w787 = pi0841 & w431;
assign w788 = w392 & w496;
assign w789 = ~w462 & ~w788;
assign w790 = ~pi0479 & w388;
assign w791 = ~pi0314 & w118;
assign w792 = ~w193 & ~w382;
assign w793 = ~w787 & ~w790;
assign w794 = ~w791 & w793;
assign w795 = w675 & w792;
assign w796 = w776 & ~w782;
assign w797 = w795 & w796;
assign w798 = w192 & w794;
assign w799 = w789 & w798;
assign w800 = ~w781 & w797;
assign w801 = w799 & w800;
assign w802 = ~w772 & ~w786;
assign w803 = w801 & w6607;
assign w804 = w768 & w803;
assign w805 = w768 & w6608;
assign w806 = ~pi0030 & pi0228;
assign w807 = ~w710 & ~w806;
assign w808 = ~w805 & w807;
assign w809 = ~w702 & ~w806;
assign w810 = ~w805 & w809;
assign w811 = w680 & ~w806;
assign w812 = ~w681 & w811;
assign w813 = ~w687 & w812;
assign w814 = ~w805 & w813;
assign w815 = (~pi0972 & ~w2) | (~pi0972 & w6609) | (~w2 & w6609);
assign w816 = w2 & w6610;
assign w817 = w811 & ~w815;
assign w818 = ~w816 & w817;
assign w819 = ~w805 & w818;
assign w820 = (~pi0960 & ~w2) | (~pi0960 & w6611) | (~w2 & w6611);
assign w821 = w2 & w6612;
assign w822 = w811 & ~w820;
assign w823 = ~w821 & w822;
assign w824 = ~w805 & w823;
assign w825 = (~pi0963 & ~w2) | (~pi0963 & w6613) | (~w2 & w6613);
assign w826 = w2 & w6614;
assign w827 = w811 & ~w825;
assign w828 = ~w826 & w827;
assign w829 = ~w805 & w828;
assign w830 = (~pi0975 & ~w2) | (~pi0975 & w6615) | (~w2 & w6615);
assign w831 = w2 & w6616;
assign w832 = w811 & ~w830;
assign w833 = ~w831 & w832;
assign w834 = ~w805 & w833;
assign w835 = (~pi0978 & ~w2) | (~pi0978 & w6617) | (~w2 & w6617);
assign w836 = w2 & w6618;
assign w837 = w811 & ~w835;
assign w838 = ~w836 & w837;
assign w839 = ~w805 & w838;
assign w840 = (~pi0954 & ~w768) | (~pi0954 & w6619) | (~w768 & w6619);
assign w841 = ~pi0024 & pi0954;
assign w842 = ~w840 & ~w841;
assign w843 = w422 & w437;
assign w844 = w305 & w843;
assign w845 = ~pi0228 & ~w844;
assign w846 = ~w16 & ~w845;
assign w847 = ~pi0228 & pi0252;
assign w848 = (~pi0468 & w847) | (~pi0468 & w6620) | (w847 & w6620);
assign w849 = pi0119 & pi1050;
assign w850 = w848 & ~w849;
assign w851 = pi0119 & pi1071;
assign w852 = w848 & ~w851;
assign w853 = pi0119 & pi1067;
assign w854 = w848 & ~w853;
assign w855 = pi0119 & pi1035;
assign w856 = w848 & ~w855;
assign w857 = ~pi0024 & w364;
assign w858 = ~pi0122 & w503;
assign w859 = w364 & w6621;
assign w860 = w232 & w6622;
assign w861 = (w860 & ~w243) | (w860 & w6623) | (~w243 & w6623);
assign w862 = w746 & w861;
assign w863 = ~pi0024 & pi0252;
assign w864 = w100 & w6624;
assign w865 = w100 & w6625;
assign w866 = ~w864 & ~w865;
assign w867 = ~w725 & w858;
assign w868 = ~w866 & w867;
assign w869 = (~w859 & w862) | (~w859 & w6398) | (w862 & w6398);
assign w870 = w779 & w6479;
assign w871 = ~pi0122 & ~w507;
assign w872 = w98 & ~w324;
assign w873 = ~pi0841 & ~w432;
assign w874 = w872 & ~w873;
assign w875 = ~w871 & w874;
assign w876 = (~pi0122 & w264) | (~pi0122 & w6626) | (w264 & w6626);
assign w877 = ~pi0286 & ~pi0288;
assign w878 = ~pi0285 & ~pi0289;
assign w879 = w877 & w878;
assign w880 = w257 & w6627;
assign w881 = ~w253 & w880;
assign w882 = w876 & w881;
assign w883 = w875 & w6480;
assign w884 = (~w264 & ~w883) | (~w264 & w6399) | (~w883 & w6399);
assign w885 = ~pi1155 & ~pi1156;
assign w886 = ~pi1157 & w885;
assign w887 = (w6399 & w6628) | (w6399 & w6629) | (w6628 & w6629);
assign w888 = ~pi0588 & ~pi0590;
assign w889 = pi0591 & ~pi0592;
assign w890 = w888 & w889;
assign w891 = pi0392 & w890;
assign w892 = ~pi0591 & ~pi0592;
assign w893 = pi0588 & ~pi0590;
assign w894 = w892 & w893;
assign w895 = pi0417 & w894;
assign w896 = ~pi0588 & pi0590;
assign w897 = w892 & w896;
assign w898 = pi0345 & w897;
assign w899 = ~pi0591 & pi0592;
assign w900 = w888 & w899;
assign w901 = pi0367 & w900;
assign w902 = ~w891 & ~w895;
assign w903 = ~w898 & ~w901;
assign w904 = w902 & w903;
assign w905 = pi0335 & w890;
assign w906 = pi0344 & w897;
assign w907 = pi0416 & w894;
assign w908 = pi0366 & w900;
assign w909 = ~w905 & ~w906;
assign w910 = ~w907 & ~w908;
assign w911 = w909 & w910;
assign w912 = ~w904 & ~w911;
assign w913 = w904 & w911;
assign w914 = ~w912 & ~w913;
assign w915 = pi0413 & w890;
assign w916 = pi0389 & w900;
assign w917 = pi0450 & w897;
assign w918 = pi0438 & w894;
assign w919 = ~w915 & ~w916;
assign w920 = ~w917 & ~w918;
assign w921 = w919 & w920;
assign w922 = pi0393 & w890;
assign w923 = pi0346 & w897;
assign w924 = pi0418 & w894;
assign w925 = pi0368 & w900;
assign w926 = ~w922 & ~w923;
assign w927 = ~w924 & ~w925;
assign w928 = w926 & w927;
assign w929 = w921 & ~w928;
assign w930 = ~w921 & w928;
assign w931 = ~w929 & ~w930;
assign w932 = w914 & w931;
assign w933 = ~w914 & ~w931;
assign w934 = ~w932 & ~w933;
assign w935 = pi0336 & w900;
assign w936 = pi0362 & w897;
assign w937 = pi0437 & w894;
assign w938 = pi0463 & w890;
assign w939 = ~w935 & ~w936;
assign w940 = ~w937 & ~w938;
assign w941 = w939 & w940;
assign w942 = pi0391 & w890;
assign w943 = pi0343 & w897;
assign w944 = pi0364 & w900;
assign w945 = pi0415 & w894;
assign w946 = ~w942 & ~w943;
assign w947 = ~w944 & ~w945;
assign w948 = w946 & w947;
assign w949 = w941 & ~w948;
assign w950 = ~w941 & w948;
assign w951 = ~w949 & ~w950;
assign w952 = pi0407 & w890;
assign w953 = pi0358 & w897;
assign w954 = pi0383 & w900;
assign w955 = pi0431 & w894;
assign w956 = ~w952 & ~w953;
assign w957 = ~w954 & ~w955;
assign w958 = w956 & w957;
assign w959 = pi0334 & w890;
assign w960 = pi0323 & w897;
assign w961 = pi0365 & w900;
assign w962 = pi0464 & w894;
assign w963 = ~w959 & ~w960;
assign w964 = ~w961 & ~w962;
assign w965 = w963 & w964;
assign w966 = ~w958 & w965;
assign w967 = w958 & ~w965;
assign w968 = ~w966 & ~w967;
assign w969 = pi0333 & w890;
assign w970 = pi0447 & w900;
assign w971 = pi0453 & w894;
assign w972 = pi0327 & w897;
assign w973 = ~w969 & ~w970;
assign w974 = ~w971 & ~w972;
assign w975 = w973 & w974;
assign w976 = w968 & ~w975;
assign w977 = ~w968 & w975;
assign w978 = ~w976 & ~w977;
assign w979 = w951 & w978;
assign w980 = ~w951 & ~w978;
assign w981 = ~w979 & ~w980;
assign w982 = ~w934 & w981;
assign w983 = (pi1191 & w981) | (pi1191 & w6400) | (w981 & w6400);
assign w984 = ~w982 & w983;
assign w985 = pi0394 & w890;
assign w986 = pi0369 & w900;
assign w987 = pi0419 & w894;
assign w988 = pi0315 & w897;
assign w989 = ~w985 & ~w986;
assign w990 = ~w987 & ~w988;
assign w991 = w989 & w990;
assign w992 = pi0349 & w897;
assign w993 = pi0329 & w890;
assign w994 = pi0454 & w894;
assign w995 = pi0440 & w900;
assign w996 = ~w992 & ~w993;
assign w997 = ~w994 & ~w995;
assign w998 = w996 & w997;
assign w999 = ~w991 & ~w998;
assign w1000 = w991 & w998;
assign w1001 = ~w999 & ~w1000;
assign w1002 = pi0424 & w894;
assign w1003 = pi0399 & w890;
assign w1004 = pi0375 & w900;
assign w1005 = pi0316 & w897;
assign w1006 = ~w1002 & ~w1003;
assign w1007 = ~w1004 & ~w1005;
assign w1008 = w1006 & w1007;
assign w1009 = pi0396 & w890;
assign w1010 = pi0322 & w897;
assign w1011 = pi0421 & w894;
assign w1012 = pi0371 & w900;
assign w1013 = ~w1009 & ~w1010;
assign w1014 = ~w1011 & ~w1012;
assign w1015 = w1013 & w1014;
assign w1016 = w1008 & ~w1015;
assign w1017 = ~w1008 & w1015;
assign w1018 = ~w1016 & ~w1017;
assign w1019 = w1001 & w1018;
assign w1020 = ~w1001 & ~w1018;
assign w1021 = ~w1019 & ~w1020;
assign w1022 = pi0347 & w897;
assign w1023 = pi0420 & w894;
assign w1024 = pi0370 & w900;
assign w1025 = pi0395 & w890;
assign w1026 = ~w1022 & ~w1023;
assign w1027 = ~w1024 & ~w1025;
assign w1028 = w1026 & w1027;
assign w1029 = pi0400 & w890;
assign w1030 = pi0374 & w900;
assign w1031 = pi0350 & w897;
assign w1032 = pi0425 & w894;
assign w1033 = ~w1029 & ~w1030;
assign w1034 = ~w1031 & ~w1032;
assign w1035 = w1033 & w1034;
assign w1036 = w1028 & ~w1035;
assign w1037 = ~w1028 & w1035;
assign w1038 = ~w1036 & ~w1037;
assign w1039 = pi0408 & w890;
assign w1040 = pi0384 & w900;
assign w1041 = pi0359 & w897;
assign w1042 = pi0432 & w894;
assign w1043 = ~w1039 & ~w1040;
assign w1044 = ~w1041 & ~w1042;
assign w1045 = w1043 & w1044;
assign w1046 = pi0398 & w890;
assign w1047 = pi0373 & w900;
assign w1048 = pi0348 & w897;
assign w1049 = pi0423 & w894;
assign w1050 = ~w1046 & ~w1047;
assign w1051 = ~w1048 & ~w1049;
assign w1052 = w1050 & w1051;
assign w1053 = w1045 & ~w1052;
assign w1054 = ~w1045 & w1052;
assign w1055 = ~w1053 & ~w1054;
assign w1056 = pi0459 & w894;
assign w1057 = pi0442 & w900;
assign w1058 = pi0328 & w890;
assign w1059 = pi0321 & w897;
assign w1060 = ~w1056 & ~w1057;
assign w1061 = ~w1058 & ~w1059;
assign w1062 = w1060 & w1061;
assign w1063 = w1055 & ~w1062;
assign w1064 = ~w1055 & w1062;
assign w1065 = ~w1063 & ~w1064;
assign w1066 = w1038 & w1065;
assign w1067 = ~w1038 & ~w1065;
assign w1068 = ~w1066 & ~w1067;
assign w1069 = ~w1021 & w1068;
assign w1070 = (pi1192 & w1068) | (pi1192 & w6401) | (w1068 & w6401);
assign w1071 = ~w1069 & w1070;
assign w1072 = pi0456 & w890;
assign w1073 = pi0443 & w894;
assign w1074 = pi0441 & w897;
assign w1075 = pi0337 & w900;
assign w1076 = ~w1072 & ~w1073;
assign w1077 = ~w1074 & ~w1075;
assign w1078 = w1076 & w1077;
assign w1079 = pi0404 & w890;
assign w1080 = pi0355 & w897;
assign w1081 = pi0429 & w894;
assign w1082 = pi0380 & w900;
assign w1083 = ~w1079 & ~w1080;
assign w1084 = ~w1081 & ~w1082;
assign w1085 = w1083 & w1084;
assign w1086 = w1078 & ~w1085;
assign w1087 = ~w1078 & w1085;
assign w1088 = ~w1086 & ~w1087;
assign w1089 = pi0324 & w890;
assign w1090 = pi0460 & w897;
assign w1091 = pi0339 & w900;
assign w1092 = pi0446 & w894;
assign w1093 = ~w1089 & ~w1090;
assign w1094 = ~w1091 & ~w1092;
assign w1095 = w1093 & w1094;
assign w1096 = pi0319 & w890;
assign w1097 = pi0338 & w900;
assign w1098 = pi0444 & w894;
assign w1099 = pi0458 & w897;
assign w1100 = ~w1096 & ~w1097;
assign w1101 = ~w1098 & ~w1099;
assign w1102 = w1100 & w1101;
assign w1103 = w1095 & ~w1102;
assign w1104 = ~w1095 & w1102;
assign w1105 = ~w1103 & ~w1104;
assign w1106 = pi0390 & w890;
assign w1107 = pi0414 & w894;
assign w1108 = pi0363 & w900;
assign w1109 = pi0342 & w897;
assign w1110 = ~w1106 & ~w1107;
assign w1111 = ~w1108 & ~w1109;
assign w1112 = w1110 & w1111;
assign w1113 = w1105 & ~w1112;
assign w1114 = ~w1105 & w1112;
assign w1115 = ~w1113 & ~w1114;
assign w1116 = w1088 & w1115;
assign w1117 = ~w1088 & ~w1115;
assign w1118 = ~w1116 & ~w1117;
assign w1119 = pi0388 & w900;
assign w1120 = pi0412 & w890;
assign w1121 = pi0436 & w894;
assign w1122 = pi0455 & w897;
assign w1123 = ~w1119 & ~w1120;
assign w1124 = ~w1121 & ~w1122;
assign w1125 = w1123 & w1124;
assign w1126 = pi0422 & w894;
assign w1127 = pi0397 & w890;
assign w1128 = pi0372 & w900;
assign w1129 = pi0320 & w897;
assign w1130 = ~w1126 & ~w1127;
assign w1131 = ~w1128 & ~w1129;
assign w1132 = w1130 & w1131;
assign w1133 = ~w1125 & ~w1132;
assign w1134 = w1125 & w1132;
assign w1135 = ~w1133 & ~w1134;
assign w1136 = pi0411 & w890;
assign w1137 = pi0435 & w894;
assign w1138 = pi0387 & w900;
assign w1139 = pi0452 & w897;
assign w1140 = ~w1136 & ~w1137;
assign w1141 = ~w1138 & ~w1139;
assign w1142 = w1140 & w1141;
assign w1143 = pi0386 & w900;
assign w1144 = pi0410 & w890;
assign w1145 = pi0361 & w897;
assign w1146 = pi0434 & w894;
assign w1147 = ~w1143 & ~w1144;
assign w1148 = ~w1145 & ~w1146;
assign w1149 = w1147 & w1148;
assign w1150 = w1142 & ~w1149;
assign w1151 = ~w1142 & w1149;
assign w1152 = ~w1150 & ~w1151;
assign w1153 = w1135 & w1152;
assign w1154 = ~w1135 & ~w1152;
assign w1155 = ~w1153 & ~w1154;
assign w1156 = ~w1118 & w1155;
assign w1157 = (pi1190 & ~w1118) | (pi1190 & w6402) | (~w1118 & w6402);
assign w1158 = ~w1156 & w1157;
assign w1159 = pi0405 & w890;
assign w1160 = pi0356 & w897;
assign w1161 = pi0445 & w894;
assign w1162 = pi0381 & w900;
assign w1163 = ~w1159 & ~w1160;
assign w1164 = ~w1161 & ~w1162;
assign w1165 = w1163 & w1164;
assign w1166 = pi0403 & w890;
assign w1167 = pi0428 & w894;
assign w1168 = pi0354 & w897;
assign w1169 = pi0379 & w900;
assign w1170 = ~w1166 & ~w1167;
assign w1171 = ~w1168 & ~w1169;
assign w1172 = w1170 & w1171;
assign w1173 = ~w1165 & ~w1172;
assign w1174 = w1165 & w1172;
assign w1175 = ~w1173 & ~w1174;
assign w1176 = pi0448 & w894;
assign w1177 = pi0462 & w897;
assign w1178 = pi0318 & w890;
assign w1179 = pi0377 & w900;
assign w1180 = ~w1176 & ~w1177;
assign w1181 = ~w1178 & ~w1179;
assign w1182 = w1180 & w1181;
assign w1183 = pi0378 & w900;
assign w1184 = pi0325 & w890;
assign w1185 = pi0451 & w894;
assign w1186 = pi0353 & w897;
assign w1187 = ~w1183 & ~w1184;
assign w1188 = ~w1185 & ~w1186;
assign w1189 = w1187 & w1188;
assign w1190 = w1182 & ~w1189;
assign w1191 = ~w1182 & w1189;
assign w1192 = ~w1190 & ~w1191;
assign w1193 = w1175 & w1192;
assign w1194 = ~w1175 & ~w1192;
assign w1195 = ~w1193 & ~w1194;
assign w1196 = pi0352 & w897;
assign w1197 = pi0427 & w894;
assign w1198 = pi0402 & w890;
assign w1199 = pi0317 & w900;
assign w1200 = ~w1196 & ~w1197;
assign w1201 = ~w1198 & ~w1199;
assign w1202 = w1200 & w1201;
assign w1203 = pi0401 & w890;
assign w1204 = pi0351 & w897;
assign w1205 = pi0426 & w894;
assign w1206 = pi0376 & w900;
assign w1207 = ~w1203 & ~w1204;
assign w1208 = ~w1205 & ~w1206;
assign w1209 = w1207 & w1208;
assign w1210 = w1202 & ~w1209;
assign w1211 = ~w1202 & w1209;
assign w1212 = ~w1210 & ~w1211;
assign w1213 = pi0409 & w890;
assign w1214 = pi0360 & w897;
assign w1215 = pi0385 & w900;
assign w1216 = pi0433 & w894;
assign w1217 = ~w1213 & ~w1214;
assign w1218 = ~w1215 & ~w1216;
assign w1219 = w1217 & w1218;
assign w1220 = pi0449 & w894;
assign w1221 = pi0439 & w900;
assign w1222 = pi0461 & w897;
assign w1223 = pi0326 & w890;
assign w1224 = ~w1220 & ~w1221;
assign w1225 = ~w1222 & ~w1223;
assign w1226 = w1224 & w1225;
assign w1227 = w1219 & ~w1226;
assign w1228 = ~w1219 & w1226;
assign w1229 = ~w1227 & ~w1228;
assign w1230 = pi0430 & w894;
assign w1231 = pi0357 & w897;
assign w1232 = pi0382 & w900;
assign w1233 = pi0406 & w890;
assign w1234 = ~w1230 & ~w1231;
assign w1235 = ~w1232 & ~w1233;
assign w1236 = w1234 & w1235;
assign w1237 = w1229 & ~w1236;
assign w1238 = ~w1229 & w1236;
assign w1239 = ~w1237 & ~w1238;
assign w1240 = w1212 & w1239;
assign w1241 = ~w1212 & ~w1239;
assign w1242 = ~w1240 & ~w1241;
assign w1243 = w1195 & ~w1242;
assign w1244 = (pi1193 & ~w1242) | (pi1193 & w6403) | (~w1242 & w6403);
assign w1245 = ~w1243 & w1244;
assign w1246 = ~w984 & ~w1071;
assign w1247 = ~w1158 & ~w1245;
assign w1248 = w1246 & w1247;
assign w1249 = ~pi0217 & ~pi1085;
assign w1250 = (w6399 & w6481) | (w6399 & w6482) | (w6481 & w6482);
assign w1251 = ~pi0098 & pi0567;
assign w1252 = (w1251 & w1248) | (w1251 & w6483) | (w1248 & w6483);
assign w1253 = w887 & w1252;
assign w1254 = pi1086 & pi1087;
assign w1255 = pi1155 & pi1156;
assign w1256 = ~pi1157 & w1255;
assign w1257 = ~pi0031 & w1254;
assign w1258 = w1256 & w1257;
assign w1259 = (~w1258 & ~w887) | (~w1258 & w6630) | (~w887 & w6630);
assign w1260 = ~w1253 & w1259;
assign w1261 = ~pi0024 & w359;
assign w1262 = (~w725 & ~w746) | (~w725 & w6404) | (~w746 & w6404);
assign w1263 = w785 & ~w1262;
assign w1264 = (w746 & w6631) | (w746 & w6632) | (w6631 & w6632);
assign w1265 = w454 & w6633;
assign w1266 = ~w726 & w1265;
assign w1267 = ~w1264 & w1266;
assign w1268 = ~w1263 & ~w1267;
assign w1269 = ~pi0137 & ~w1268;
assign w1270 = ~pi0137 & w495;
assign w1271 = (~w879 & ~w257) | (~w879 & w6634) | (~w257 & w6634);
assign w1272 = w317 & w6635;
assign w1273 = (~pi0841 & ~w495) | (~pi0841 & w6636) | (~w495 & w6636);
assign w1274 = w392 & ~w1273;
assign w1275 = ~w1261 & ~w1274;
assign w1276 = ~w1272 & w1275;
assign w1277 = ~w1269 & w1276;
assign w1278 = ~pi0841 & w426;
assign w1279 = ~w212 & ~w1278;
assign w1280 = w770 & w6637;
assign w1281 = ~w168 & ~w1280;
assign w1282 = ~w1280 & w6638;
assign w1283 = w25 & w1282;
assign w1284 = w746 & w6484;
assign w1285 = w746 & w6485;
assign w1286 = ~w1284 & ~w1285;
assign w1287 = ~pi0038 & ~pi0054;
assign w1288 = ~pi0057 & ~pi0059;
assign w1289 = w1287 & w1288;
assign w1290 = w417 & w6639;
assign w1291 = ~pi0074 & ~w790;
assign w1292 = ~pi0040 & w1289;
assign w1293 = w1289 & w6640;
assign w1294 = ~pi0033 & ~pi0954;
assign w1295 = ~pi0033 & ~pi0034;
assign w1296 = ~pi0079 & ~pi0118;
assign w1297 = ~pi0138 & ~pi0139;
assign w1298 = ~pi0195 & ~pi0196;
assign w1299 = w1297 & w1298;
assign w1300 = w1295 & w1296;
assign w1301 = w1299 & w1300;
assign w1302 = w1294 & ~w1301;
assign w1303 = pi0033 & pi0954;
assign w1304 = w1293 & ~w1303;
assign w1305 = ~w1302 & w1304;
assign w1306 = w1290 & w6641;
assign w1307 = (w1306 & w1286) | (w1306 & w6642) | (w1286 & w6642);
assign w1308 = w746 & w6405;
assign w1309 = w746 & w6406;
assign w1310 = ~w1308 & ~w1309;
assign w1311 = pi0074 & w1310;
assign w1312 = w760 & w790;
assign w1313 = ~w462 & w746;
assign w1314 = (pi0149 & ~w2) | (pi0149 & w6643) | (~w2 & w6643);
assign w1315 = w2 & w6644;
assign w1316 = ~w1314 & ~w1315;
assign w1317 = w746 & w6645;
assign w1318 = ~w1290 & ~w1317;
assign w1319 = ~w1311 & ~w1312;
assign w1320 = w1319 & w6646;
assign w1321 = w1283 & ~w1320;
assign w1322 = (~w377 & ~w780) | (~w377 & w6486) | (~w780 & w6486);
assign w1323 = w746 & w6647;
assign w1324 = ~w1281 & ~w1323;
assign w1325 = w746 & w6648;
assign w1326 = w746 & w6649;
assign w1327 = ~w1325 & ~w1326;
assign w1328 = ~w1279 & w1327;
assign w1329 = (pi0157 & ~w2) | (pi0157 & w6650) | (~w2 & w6650);
assign w1330 = w2 & w6651;
assign w1331 = ~w1329 & ~w1330;
assign w1332 = ~w1316 & ~w1331;
assign w1333 = w1316 & w1331;
assign w1334 = ~w25 & ~w1332;
assign w1335 = ~w1333 & w1334;
assign w1336 = w746 & w6652;
assign w1337 = w1322 & ~w1336;
assign w1338 = ~w1328 & w6653;
assign w1339 = ~w1321 & w1338;
assign w1340 = w746 & w6654;
assign w1341 = w746 & w6655;
assign w1342 = ~w1340 & ~w1341;
assign w1343 = ~w1322 & ~w1342;
assign w1344 = ~w1339 & ~w1343;
assign w1345 = ~w1301 & w6656;
assign w1346 = pi0034 & ~w1294;
assign w1347 = w1293 & ~w1346;
assign w1348 = ~w1345 & w1347;
assign w1349 = w746 & w6487;
assign w1350 = w746 & w6488;
assign w1351 = ~w1349 & ~w1350;
assign w1352 = w1290 & w6657;
assign w1353 = (w1352 & w1351) | (w1352 & w6658) | (w1351 & w6658);
assign w1354 = pi0162 & ~w4;
assign w1355 = w2 & w6659;
assign w1356 = ~w1354 & ~w1355;
assign w1357 = w746 & w6489;
assign w1358 = ~w1290 & ~w1357;
assign w1359 = w763 & w790;
assign w1360 = w746 & w6490;
assign w1361 = w746 & w6491;
assign w1362 = ~w1360 & ~w1361;
assign w1363 = pi0074 & w1362;
assign w1364 = ~w1358 & ~w1359;
assign w1365 = w1364 & w6660;
assign w1366 = w1283 & ~w1365;
assign w1367 = w746 & w6661;
assign w1368 = w746 & w6662;
assign w1369 = ~w1367 & ~w1368;
assign w1370 = ~w1322 & w1369;
assign w1371 = w746 & w6663;
assign w1372 = ~w1281 & ~w1371;
assign w1373 = ~w1370 & ~w1372;
assign w1374 = w757 & w1356;
assign w1375 = ~w757 & ~w1356;
assign w1376 = ~w1374 & ~w1375;
assign w1377 = w1333 & w1376;
assign w1378 = ~w1333 & ~w1376;
assign w1379 = ~w1377 & ~w1378;
assign w1380 = w746 & w6664;
assign w1381 = ~w25 & ~w1380;
assign w1382 = w746 & w6665;
assign w1383 = ~w1279 & ~w1382;
assign w1384 = ~w1381 & ~w1383;
assign w1385 = w1373 & w1384;
assign w1386 = ~w1366 & w1385;
assign w1387 = ~w1370 & w6666;
assign w1388 = ~w1386 & ~w1387;
assign w1389 = w1265 & w6667;
assign w1390 = ~w726 & w784;
assign w1391 = (~w864 & ~w784) | (~w864 & w6668) | (~w784 & w6668);
assign w1392 = ~w1262 & ~w1391;
assign w1393 = (~w746 & w6492) | (~w746 & w6493) | (w6492 & w6493);
assign w1394 = pi0683 & w1393;
assign w1395 = w1393 & w6669;
assign w1396 = w317 & w6670;
assign w1397 = w876 & w1396;
assign w1398 = pi1076 & w329;
assign w1399 = w433 & w6671;
assign w1400 = w783 & w784;
assign w1401 = ~w473 & ~w482;
assign w1402 = w789 & w1401;
assign w1403 = ~pi0024 & ~w1402;
assign w1404 = ~w212 & ~w674;
assign w1405 = w1404 & w6672;
assign w1406 = w1405 & w6673;
assign w1407 = ~w1400 & ~w1403;
assign w1408 = w1406 & w1407;
assign w1409 = ~w1392 & w1408;
assign w1410 = ~w1395 & w1409;
assign w1411 = ~w301 & ~w857;
assign w1412 = w265 & ~w1411;
assign w1413 = (~pi0841 & w742) | (~pi0841 & w6674) | (w742 & w6674);
assign w1414 = pi0024 & w462;
assign w1415 = ~w1413 & ~w1414;
assign w1416 = w145 & w152;
assign w1417 = pi0314 & w285;
assign w1418 = w285 & w1729;
assign w1419 = pi0786 & ~pi1076;
assign w1420 = (w1419 & w711) | (w1419 & w6678) | (w711 & w6678);
assign w1421 = w350 & ~w1420;
assign w1422 = ~w711 & w6679;
assign w1423 = w668 & ~w769;
assign w1424 = ~w1422 & w1423;
assign w1425 = w1421 & w1424;
assign w1426 = w392 & ~w495;
assign w1427 = ~w291 & ~w436;
assign w1428 = (~pi0841 & ~w1427) | (~pi0841 & w6680) | (~w1427 & w6680);
assign w1429 = ~w1416 & ~w1418;
assign w1430 = ~w1428 & w1429;
assign w1431 = ~w1425 & w1430;
assign w1432 = pi0102 & w341;
assign w1433 = ~pi1076 & w329;
assign w1434 = ~w1432 & ~w1433;
assign w1435 = w875 & w6494;
assign w1436 = ~pi0480 & pi0949;
assign w1437 = w143 & w1436;
assign w1438 = ~pi0250 & pi0252;
assign w1439 = pi0901 & ~pi0959;
assign w1440 = w1438 & w1439;
assign w1441 = w309 & w1440;
assign w1442 = ~w1437 & ~w1441;
assign w1443 = ~pi0228 & w1442;
assign w1444 = (w6408 & w6495) | (w6408 & w6496) | (w6495 & w6496);
assign w1445 = ~pi0101 & w1444;
assign w1446 = (pi0041 & ~w1444) | (pi0041 & w6681) | (~w1444 & w6681);
assign w1447 = ~pi0039 & ~pi0072;
assign w1448 = (w6408 & w6497) | (w6408 & w6498) | (w6497 & w6498);
assign w1449 = w1447 & ~w1448;
assign w1450 = ~w1446 & w1449;
assign w1451 = pi0039 & ~pi0072;
assign w1452 = w746 & w6682;
assign w1453 = (w1451 & ~w1452) | (w1451 & w6684) | (~w1452 & w6684);
assign w1454 = ~w1450 & ~w1453;
assign w1455 = (pi0219 & ~w2) | (pi0219 & w6409) | (~w2 & w6409);
assign w1456 = w2 & w6410;
assign w1457 = ~w1455 & ~w1456;
assign w1458 = (pi0214 & ~w2) | (pi0214 & w6685) | (~w2 & w6685);
assign w1459 = w2 & w6686;
assign w1460 = ~w1458 & ~w1459;
assign w1461 = (pi0212 & ~w2) | (pi0212 & w6687) | (~w2 & w6687);
assign w1462 = w2 & w6688;
assign w1463 = ~w1461 & ~w1462;
assign w1464 = ~w1460 & ~w1463;
assign w1465 = (pi0211 & ~w2) | (pi0211 & w6689) | (~w2 & w6689);
assign w1466 = w2 & w6690;
assign w1467 = ~w1465 & ~w1466;
assign w1468 = w1457 & ~w1467;
assign w1469 = w1464 & w1468;
assign w1470 = w1457 & ~w1469;
assign w1471 = ~w1452 & w6691;
assign w1472 = (w6408 & w6499) | (w6408 & w6500) | (w6499 & w6500);
assign w1473 = (w6408 & w6501) | (w6408 & w6502) | (w6501 & w6502);
assign w1474 = pi0042 & ~w1473;
assign w1475 = (w1447 & w1474) | (w1447 & w6692) | (w1474 & w6692);
assign w1476 = ~w1471 & ~w1475;
assign w1477 = w1457 & w1467;
assign w1478 = ~w1464 & w1477;
assign w1479 = w1460 & w1463;
assign w1480 = ~w1469 & w6693;
assign w1481 = ~w1464 & ~w1467;
assign w1482 = (~w1481 & ~w1480) | (~w1481 & w6694) | (~w1480 & w6694);
assign w1483 = ~w1452 & w6695;
assign w1484 = pi0043 & ~w1472;
assign w1485 = ~pi0043 & w1472;
assign w1486 = ~w1484 & ~w1485;
assign w1487 = w1447 & ~w1486;
assign w1488 = ~w1483 & ~w1487;
assign w1489 = w746 & w6696;
assign w1490 = (~w6408 & w6697) | (~w6408 & w6698) | (w6697 & w6698);
assign w1491 = ~w1444 & ~w1490;
assign w1492 = w1447 & ~w1491;
assign w1493 = ~w1489 & ~w1492;
assign w1494 = ~pi0287 & pi0979;
assign w1495 = w350 & w1494;
assign w1496 = w470 & w6699;
assign w1497 = ~pi0841 & w106;
assign w1498 = ~w1496 & ~w1497;
assign w1499 = (~w263 & w264) | (~w263 & w6700) | (w264 & w6700);
assign w1500 = (w1499 & w857) | (w1499 & w2689) | (w857 & w2689);
assign w1501 = ~w150 & ~w259;
assign w1502 = w145 & w1501;
assign w1503 = ~w1500 & ~w1502;
assign w1504 = w317 & w6701;
assign w1505 = ~w274 & w6702;
assign w1506 = w437 & w1505;
assign w1507 = (~w1504 & w1506) | (~w1504 & w6703) | (w1506 & w6703);
assign w1508 = pi0048 & ~w1507;
assign w1509 = pi0841 & w123;
assign w1510 = w243 & w6704;
assign w1511 = ~w1509 & ~w1510;
assign w1512 = pi0024 & w359;
assign w1513 = w257 & w6705;
assign w1514 = (~w746 & w6706) | (~w746 & w6707) | (w6706 & w6707);
assign w1515 = (w309 & w1514) | (w309 & w6708) | (w1514 & w6708);
assign w1516 = w726 & w1265;
assign w1517 = ~w1512 & ~w1516;
assign w1518 = ~w786 & w1517;
assign w1519 = ~w1515 & w1518;
assign w1520 = ~w1452 & w6709;
assign w1521 = w725 & w1447;
assign w1522 = (w6408 & w6710) | (w6408 & w6711) | (w6710 & w6711);
assign w1523 = pi0052 & w1447;
assign w1524 = (w1523 & ~w1472) | (w1523 & w6712) | (~w1472 & w6712);
assign w1525 = ~w1520 & ~w1522;
assign w1526 = ~w1524 & w1525;
assign w1527 = pi0024 & w399;
assign w1528 = w665 & w666;
assign w1529 = w350 & w1528;
assign w1530 = ~w1527 & ~w1529;
assign w1531 = pi0024 & w482;
assign w1532 = ~pi0841 & w134;
assign w1533 = ~w1531 & ~w1532;
assign w1534 = pi0024 & w404;
assign w1535 = ~w198 & ~w1534;
assign w1536 = ~pi0024 & w404;
assign w1537 = (~w1506 & w6713) | (~w1506 & w6714) | (w6713 & w6714);
assign w1538 = ~w1536 & ~w1537;
assign w1539 = (pi0024 & w466) | (pi0024 & w6715) | (w466 & w6715);
assign w1540 = pi0057 & w1539;
assign w1541 = ~pi0924 & w314;
assign w1542 = ~w274 & ~w1541;
assign w1543 = ~pi0841 & ~w1542;
assign w1544 = ~w1540 & ~w1543;
assign w1545 = w470 & w6716;
assign w1546 = ~pi0841 & pi0924;
assign w1547 = w314 & w1546;
assign w1548 = ~w1545 & ~w1547;
assign w1549 = pi0024 & w415;
assign w1550 = w350 & w6717;
assign w1551 = ~w1549 & ~w1550;
assign w1552 = ~pi0024 & w415;
assign w1553 = ~w106 & ~w207;
assign w1554 = ~w346 & w1553;
assign w1555 = pi0841 & ~w1554;
assign w1556 = ~w1554 & w6718;
assign w1557 = ~w1552 & ~w1556;
assign w1558 = w271 & w6719;
assign w1559 = pi0841 & w314;
assign w1560 = ~w1558 & ~w1559;
assign w1561 = pi0993 & w355;
assign w1562 = w470 & w6720;
assign w1563 = ~w1561 & ~w1562;
assign w1564 = (~w1506 & w6721) | (~w1506 & w6722) | (w6721 & w6722);
assign w1565 = ~w129 & ~w1564;
assign w1566 = w777 & w1420;
assign w1567 = w179 & w6723;
assign w1568 = ~w1457 & w1567;
assign w1569 = pi0083 & w335;
assign w1570 = w74 & w1569;
assign w1571 = w92 & w1570;
assign w1572 = pi0314 & w1571;
assign w1573 = w350 & w6724;
assign w1574 = w770 & w1573;
assign w1575 = ~pi0314 & w334;
assign w1576 = w67 & w85;
assign w1577 = w92 & w6725;
assign w1578 = w156 & w1577;
assign w1579 = ~w1575 & ~w1578;
assign w1580 = pi0024 & w410;
assign w1581 = pi0589 & ~w495;
assign w1582 = w15 & w769;
assign w1583 = ~pi0979 & ~w664;
assign w1584 = ~w665 & w1583;
assign w1585 = w1583 & w6726;
assign w1586 = ~w495 & w6727;
assign w1587 = (~pi0287 & ~w769) | (~pi0287 & w6729) | (~w769 & w6729);
assign w1588 = w350 & ~w1587;
assign w1589 = ~w1580 & ~w1588;
assign w1590 = w157 & w1577;
assign w1591 = w179 & w6730;
assign w1592 = ~w1590 & ~w1591;
assign w1593 = pi0314 & ~w1592;
assign w1594 = w257 & w6731;
assign w1595 = w145 & w6732;
assign w1596 = w770 & w6733;
assign w1597 = pi0024 & w298;
assign w1598 = ~w1595 & ~w1597;
assign w1599 = ~w1596 & w1598;
assign w1600 = ~pi0314 & pi1044;
assign w1601 = ~w1280 & ~w1600;
assign w1602 = ~w1281 & ~w1601;
assign w1603 = w243 & w6734;
assign w1604 = (~pi0841 & ~w257) | (~pi0841 & w6735) | (~w257 & w6735);
assign w1605 = w207 & w6736;
assign w1606 = pi0479 & ~w495;
assign w1607 = w202 & w6737;
assign w1608 = ~w1603 & ~w1605;
assign w1609 = ~w1607 & w1608;
assign w1610 = w784 & w6738;
assign w1611 = w1262 & w1610;
assign w1612 = ~w1394 & w1611;
assign w1613 = w143 & w1393;
assign w1614 = w309 & ~w1513;
assign w1615 = (~w746 & w6739) | (~w746 & w6740) | (w6739 & w6740);
assign w1616 = w1614 & w1615;
assign w1617 = ~w1425 & ~w1613;
assign w1618 = ~w1616 & w1617;
assign w1619 = w1618 & w6741;
assign w1620 = pi0075 & ~w1619;
assign w1621 = w507 & ~w1620;
assign w1622 = w317 & w1271;
assign w1623 = (w746 & w6742) | (w746 & w6743) | (w6742 & w6743);
assign w1624 = ~w1504 & ~w1622;
assign w1625 = ~w1623 & w1624;
assign w1626 = (~pi0314 & w445) | (~pi0314 & w6744) | (w445 & w6744);
assign w1627 = (pi0077 & w1626) | (pi0077 & w6745) | (w1626 & w6745);
assign w1628 = ~w459 & ~w1627;
assign w1629 = pi0119 & pi0232;
assign w1630 = ~pi0468 & w1629;
assign w1631 = w746 & w6746;
assign w1632 = w746 & w6747;
assign w1633 = ~w1631 & ~w1632;
assign w1634 = ~w1322 & ~w1633;
assign w1635 = ~w1281 & ~w1452;
assign w1636 = w746 & w6503;
assign w1637 = w746 & w6504;
assign w1638 = ~w1636 & ~w1637;
assign w1639 = (w1322 & ~w1638) | (w1322 & w6748) | (~w1638 & w6748);
assign w1640 = ~w1635 & w1639;
assign w1641 = w1639 & w6749;
assign w1642 = w746 & w6411;
assign w1643 = w746 & w6412;
assign w1644 = ~w1642 & ~w1643;
assign w1645 = (~w1374 & ~w1376) | (~w1374 & w6750) | (~w1376 & w6750);
assign w1646 = w746 & w6505;
assign w1647 = w1644 & ~w1646;
assign w1648 = (~w25 & ~w1644) | (~w25 & w6506) | (~w1644 & w6506);
assign w1649 = ~w1644 & w1646;
assign w1650 = w1648 & ~w1649;
assign w1651 = w1290 & w6751;
assign w1652 = (pi0079 & w1301) | (pi0079 & w6752) | (w1301 & w6752);
assign w1653 = (w40 & ~w1345) | (w40 & w6753) | (~w1345 & w6753);
assign w1654 = (w1292 & ~w1653) | (w1292 & w6754) | (~w1653 & w6754);
assign w1655 = w746 & w6755;
assign w1656 = (~w1289 & ~w746) | (~w1289 & w6756) | (~w746 & w6756);
assign w1657 = ~w1655 & w1656;
assign w1658 = (w1651 & w1657) | (w1651 & w6757) | (w1657 & w6757);
assign w1659 = w754 & w790;
assign w1660 = ~w1290 & w1644;
assign w1661 = ~w1659 & ~w1660;
assign w1662 = ~w1650 & w1661;
assign w1663 = w1662 & w6758;
assign w1664 = ~w1634 & ~w1641;
assign w1665 = ~w1663 & w1664;
assign w1666 = w886 & w1254;
assign w1667 = w886 & w6759;
assign w1668 = ~w1252 & w1667;
assign w1669 = w179 & w6760;
assign w1670 = ~w180 & ~w1669;
assign w1671 = w52 & w181;
assign w1672 = w185 & w1671;
assign w1673 = pi0314 & w334;
assign w1674 = ~w1672 & ~w1673;
assign w1675 = w183 & w1671;
assign w1676 = ~pi0314 & w1571;
assign w1677 = ~w1675 & ~w1676;
assign w1678 = w1477 & w1567;
assign w1679 = w1577 & w6761;
assign w1680 = ~w174 & ~w1679;
assign w1681 = w522 & w780;
assign w1682 = pi0314 & w118;
assign w1683 = w145 & w6762;
assign w1684 = w145 & w6763;
assign w1685 = ~w1683 & ~w1684;
assign w1686 = w259 & ~w1685;
assign w1687 = ~pi0024 & w410;
assign w1688 = ~w1554 & w6764;
assign w1689 = ~w1687 & ~w1688;
assign w1690 = (~w1506 & w6765) | (~w1506 & w6766) | (w6765 & w6766);
assign w1691 = ~pi1044 & w168;
assign w1692 = ~w1690 & ~w1691;
assign w1693 = w301 & w503;
assign w1694 = ~w364 & ~w1693;
assign w1695 = ~pi0024 & ~w503;
assign w1696 = (~w1695 & w1693) | (~w1695 & w6767) | (w1693 & w6767);
assign w1697 = ~w870 & ~w1696;
assign w1698 = (~w1600 & ~w780) | (~w1600 & w6768) | (~w780 & w6768);
assign w1699 = ~w1322 & ~w1698;
assign w1700 = ~pi1044 & w377;
assign w1701 = ~w787 & ~w1700;
assign w1702 = ~pi0841 & w123;
assign w1703 = ~w1616 & ~w1702;
assign w1704 = w1582 & w6769;
assign w1705 = pi0024 & w388;
assign w1706 = ~pi0332 & ~pi0841;
assign w1707 = w283 & w6770;
assign w1708 = ~w1705 & ~w1707;
assign w1709 = ~w1704 & w1708;
assign w1710 = ~pi0024 & w388;
assign w1711 = w207 & w6771;
assign w1712 = (pi0096 & w1555) | (pi0096 & w6772) | (w1555 & w6772);
assign w1713 = ~w1710 & ~w1712;
assign w1714 = ~w263 & w1606;
assign w1715 = ~w265 & ~w1714;
assign w1716 = w202 & ~w1715;
assign w1717 = ~w495 & w6773;
assign w1718 = w1582 & w6774;
assign w1719 = ~w1716 & ~w1718;
assign w1720 = ~w168 & ~w377;
assign w1721 = pi0314 & pi1044;
assign w1722 = ~w1720 & w1721;
assign w1723 = pi0099 & ~w1448;
assign w1724 = (w6408 & w6508) | (w6408 & w6509) | (w6508 & w6509);
assign w1725 = (w1447 & w1723) | (w1447 & w6775) | (w1723 & w6775);
assign w1726 = ~w235 & w1451;
assign w1727 = w1452 & w6776;
assign w1728 = ~w1725 & ~w1727;
assign w1729 = (w264 & w6777) | (w264 & w6778) | (w6777 & w6778);
assign w1730 = w285 & ~w1729;
assign w1731 = ~w266 & w6779;
assign w1732 = ~w1730 & ~w1731;
assign w1733 = w1618 & w6780;
assign w1734 = pi0100 & ~w1733;
assign w1735 = w454 & w6781;
assign w1736 = ~w1264 & w1735;
assign w1737 = ~w1734 & ~w1736;
assign w1738 = pi0101 & ~w1444;
assign w1739 = ~w1445 & ~w1738;
assign w1740 = w1447 & ~w1739;
assign w1741 = w231 & w1726;
assign w1742 = w1452 & w1741;
assign w1743 = ~w1740 & ~w1742;
assign w1744 = pi0065 & w341;
assign w1745 = ~w112 & ~w791;
assign w1746 = w143 & ~w1393;
assign w1747 = w145 & w6782;
assign w1748 = ~w1746 & ~w1747;
assign w1749 = pi0841 & w134;
assign w1750 = ~pi0024 & w399;
assign w1751 = ~w1749 & ~w1750;
assign w1752 = ~pi0993 & w355;
assign w1753 = w872 & ~w1730;
assign w1754 = w444 & w6783;
assign w1755 = pi0314 & w138;
assign w1756 = ~w1613 & ~w1755;
assign w1757 = pi0111 & w1626;
assign w1758 = ~pi0024 & w298;
assign w1759 = ~w1757 & ~w1758;
assign w1760 = pi0124 & ~pi0468;
assign w1761 = pi0113 & ~w1724;
assign w1762 = ~pi0113 & w1724;
assign w1763 = ~w1761 & ~w1762;
assign w1764 = w1447 & ~w1763;
assign w1765 = (w6408 & w6510) | (w6408 & w6511) | (w6510 & w6511);
assign w1766 = ~pi0115 & w1765;
assign w1767 = (pi0114 & ~w1765) | (pi0114 & w6784) | (~w1765 & w6784);
assign w1768 = ~w1473 & ~w1767;
assign w1769 = w1447 & ~w1768;
assign w1770 = pi0115 & ~w1765;
assign w1771 = ~w1766 & ~w1770;
assign w1772 = w1447 & ~w1771;
assign w1773 = (pi0116 & ~w1724) | (pi0116 & w6785) | (~w1724 & w6785);
assign w1774 = ~w1765 & ~w1773;
assign w1775 = w1447 & ~w1774;
assign w1776 = (pi0118 & ~w1345) | (pi0118 & w6786) | (~w1345 & w6786);
assign w1777 = w1345 & w1296;
assign w1778 = ~w1776 & ~w1777;
assign w1779 = w1293 & w1322;
assign w1780 = w1651 & w1779;
assign w1781 = w1780 & w6787;
assign w1782 = w746 & w6413;
assign w1783 = w746 & w6414;
assign w1784 = ~w1782 & ~w1783;
assign w1785 = (w1784 & w1648) | (w1784 & w6788) | (w1648 & w6788);
assign w1786 = ~w25 & ~w1784;
assign w1787 = w1647 & w1786;
assign w1788 = w746 & w6789;
assign w1789 = (~w1289 & ~w746) | (~w1289 & w6790) | (~w746 & w6790);
assign w1790 = ~w1788 & w1789;
assign w1791 = w1651 & w1790;
assign w1792 = w746 & w6791;
assign w1793 = w746 & w6792;
assign w1794 = ~w1792 & ~w1793;
assign w1795 = ~w1281 & w1794;
assign w1796 = w746 & w6513;
assign w1797 = ~w1322 & ~w1796;
assign w1798 = w746 & w6415;
assign w1799 = w746 & w6416;
assign w1800 = ~w1798 & ~w1799;
assign w1801 = ~w1279 & w1800;
assign w1802 = ~w1797 & ~w1801;
assign w1803 = ~w1787 & w1802;
assign w1804 = w1803 & w6793;
assign w1805 = ~w1781 & w1804;
assign w1806 = pi0128 & pi0228;
assign w1807 = ~w522 & ~w524;
assign w1808 = w779 & w6794;
assign w1809 = ~w431 & ~w504;
assign w1810 = w455 & w1809;
assign w1811 = w1810 & w6795;
assign w1812 = ~w767 & w6417;
assign w1813 = (~pi0228 & w767) | (~pi0228 & w6796) | (w767 & w6796);
assign w1814 = ~w1806 & ~w1813;
assign w1815 = ~pi0031 & ~pi0080;
assign w1816 = pi0818 & w1815;
assign w1817 = pi0951 & pi0982;
assign w1818 = w886 & w6797;
assign w1819 = ~w1816 & ~w1818;
assign w1820 = (pi1087 & w1818) | (pi1087 & w6798) | (w1818 & w6798);
assign w1821 = ~pi0120 & ~w1820;
assign w1822 = ~w884 & ~w1821;
assign w1823 = (~pi0024 & ~w444) | (~pi0024 & w6799) | (~w444 & w6799);
assign w1824 = w373 & ~w1823;
assign w1825 = ~w1754 & ~w1824;
assign w1826 = pi0051 & ~w1382;
assign w1827 = ~pi0067 & ~pi0068;
assign w1828 = ~pi0071 & ~pi0084;
assign w1829 = w1827 & w1828;
assign w1830 = ~pi0125 & ~pi0133;
assign w1831 = ~pi0121 & w1830;
assign w1832 = w1830 & w6800;
assign w1833 = w1832 & w6801;
assign w1834 = w1832 & w6802;
assign w1835 = w1834 & w6803;
assign w1836 = pi0121 & ~w1830;
assign w1837 = ~w1831 & ~w1836;
assign w1838 = (w1829 & w1835) | (w1829 & w6804) | (w1835 & w6804);
assign w1839 = ~pi0051 & ~w1838;
assign w1840 = (w1839 & ~w1371) | (w1839 & w6805) | (~w1371 & w6805);
assign w1841 = ~pi0087 & ~w1826;
assign w1842 = ~w1840 & w1841;
assign w1843 = (w1825 & w1644) | (w1825 & w6806) | (w1644 & w6806);
assign w1844 = ~w1842 & w1843;
assign w1845 = w1754 & w1823;
assign w1846 = w760 & w1845;
assign w1847 = ~w298 & ~w677;
assign w1848 = (w1847 & ~w1633) | (w1847 & w6807) | (~w1633 & w6807);
assign w1849 = ~w1846 & w1848;
assign w1850 = ~w1844 & w1849;
assign w1851 = w678 & ~w763;
assign w1852 = ~w1850 & ~w1851;
assign w1853 = pi0110 & ~w1393;
assign w1854 = w524 & w668;
assign w1855 = (pi0039 & ~w769) | (pi0039 & w6809) | (~w769 & w6809);
assign w1856 = ~w52 & ~w179;
assign w1857 = ~w171 & ~w331;
assign w1858 = w63 & w6810;
assign w1859 = ~w135 & ~w294;
assign w1860 = w63 & w6811;
assign w1861 = ~w88 & ~w1860;
assign w1862 = w65 & ~w166;
assign w1863 = ~w424 & w1862;
assign w1864 = ~w1861 & ~w1863;
assign w1865 = (w71 & w1864) | (w71 & w6812) | (w1864 & w6812);
assign w1866 = w48 & ~w187;
assign w1867 = (~w1865 & w6814) | (~w1865 & w6815) | (w6814 & w6815);
assign w1868 = pi0039 & ~pi0110;
assign w1869 = ~pi0039 & pi0110;
assign w1870 = ~w1868 & ~w1869;
assign w1871 = (w1870 & w1867) | (w1870 & w6816) | (w1867 & w6816);
assign w1872 = ~w1853 & ~w1855;
assign w1873 = ~w1871 & w1872;
assign w1874 = w746 & w6817;
assign w1875 = w1845 & ~w1874;
assign w1876 = ~pi0051 & ~pi0087;
assign w1877 = ~w1829 & w1876;
assign w1878 = ~w1323 & w1877;
assign w1879 = pi0087 & ~w1357;
assign w1880 = pi0051 & ~pi0087;
assign w1881 = w1327 & w1880;
assign w1882 = w678 & w760;
assign w1883 = w1369 & w1824;
assign w1884 = w1829 & w1876;
assign w1885 = w1825 & w6818;
assign w1886 = pi0125 & pi0133;
assign w1887 = ~w1830 & ~w1886;
assign w1888 = w1885 & w6819;
assign w1889 = ~w1875 & ~w1878;
assign w1890 = ~w1879 & ~w1881;
assign w1891 = ~w1882 & ~w1883;
assign w1892 = w1890 & w1891;
assign w1893 = w1889 & w1892;
assign w1894 = ~w1888 & w1893;
assign w1895 = pi0087 & ~w1784;
assign w1896 = w678 & ~w754;
assign w1897 = ~w1638 & w1880;
assign w1898 = ~w1796 & w1824;
assign w1899 = w1452 & w1877;
assign w1900 = (w1832 & ~w1834) | (w1832 & w6820) | (~w1834 & w6820);
assign w1901 = (pi0126 & ~w1830) | (pi0126 & w6821) | (~w1830 & w6821);
assign w1902 = w1884 & ~w1901;
assign w1903 = ~w1900 & w1902;
assign w1904 = w1825 & w6822;
assign w1905 = ~w1899 & w1904;
assign w1906 = (~w678 & ~w763) | (~w678 & w6823) | (~w763 & w6823);
assign w1907 = ~w1898 & w1906;
assign w1908 = ~w1905 & w1907;
assign w1909 = ~w1895 & ~w1896;
assign w1910 = ~w1897 & w1909;
assign w1911 = ~w1908 & w1910;
assign w1912 = w225 & w6824;
assign w1913 = ~w346 & w6825;
assign w1914 = w344 & w1913;
assign w1915 = w773 & w1914;
assign w1916 = w477 & w1915;
assign w1917 = w1912 & w1916;
assign w1918 = (pi0127 & ~w1615) | (pi0127 & w6826) | (~w1615 & w6826);
assign w1919 = w1615 & w6827;
assign w1920 = w309 & ~w1918;
assign w1921 = ~w1919 & w1920;
assign w1922 = (pi0129 & ~w1917) | (pi0129 & w6828) | (~w1917 & w6828);
assign w1923 = ~w1921 & w1922;
assign w1924 = (~pi0250 & w1615) | (~pi0250 & w6829) | (w1615 & w6829);
assign w1925 = (w1615 & w6830) | (w1615 & w6831) | (w6830 & w6831);
assign w1926 = (~w455 & w1924) | (~w455 & w6832) | (w1924 & w6832);
assign w1927 = ~w1925 & w1926;
assign w1928 = ~w355 & w455;
assign w1929 = w1917 & w1928;
assign w1930 = ~w1927 & ~w1929;
assign w1931 = w678 & ~w1357;
assign w1932 = pi0087 & w1351;
assign w1933 = (pi0130 & ~w1832) | (pi0130 & w6833) | (~w1832 & w6833);
assign w1934 = ~w1833 & ~w1933;
assign w1935 = w1885 & w6834;
assign w1936 = w1310 & w1877;
assign w1937 = ~w1931 & ~w1932;
assign w1938 = ~w1936 & w1937;
assign w1939 = ~w1935 & w1938;
assign w1940 = w1800 & w1880;
assign w1941 = w1794 & w1877;
assign w1942 = w754 & w1845;
assign w1943 = pi0087 & w1286;
assign w1944 = w678 & ~w1317;
assign w1945 = ~pi0132 & ~w1900;
assign w1946 = pi0132 & w1900;
assign w1947 = ~w1945 & ~w1946;
assign w1948 = w1885 & w1947;
assign w1949 = ~w1940 & ~w1941;
assign w1950 = ~w1942 & ~w1943;
assign w1951 = ~w1944 & w1950;
assign w1952 = ~w1948 & w1949;
assign w1953 = w1951 & w1952;
assign w1954 = w1342 & w1824;
assign w1955 = w678 & ~w1874;
assign w1956 = (~pi0133 & ~w1834) | (~pi0133 & w6835) | (~w1834 & w6835);
assign w1957 = w1884 & ~w1956;
assign w1958 = pi0087 & w1317;
assign w1959 = w1825 & w6836;
assign w1960 = ~w1958 & w1959;
assign w1961 = ~w1954 & ~w1955;
assign w1962 = ~w1960 & w1961;
assign w1963 = w678 & w1286;
assign w1964 = w746 & w6837;
assign w1965 = w746 & w6838;
assign w1966 = ~w1964 & ~w1965;
assign w1967 = w1877 & w1966;
assign w1968 = (pi0134 & ~w1834) | (pi0134 & w6839) | (~w1834 & w6839);
assign w1969 = w1885 & w1968;
assign w1970 = ~w1963 & ~w1967;
assign w1971 = ~w1969 & w1970;
assign w1972 = w678 & w1784;
assign w1973 = w1834 & w6840;
assign w1974 = (w1829 & w1834) | (w1829 & w6841) | (w1834 & w6841);
assign w1975 = ~w1973 & w1974;
assign w1976 = w746 & w6842;
assign w1977 = pi0194 & w752;
assign w1978 = ~w1976 & ~w1977;
assign w1979 = (~w1829 & w1977) | (~w1829 & w6843) | (w1977 & w6843);
assign w1980 = w1876 & ~w1975;
assign w1981 = w1825 & w6844;
assign w1982 = ~w1979 & w1981;
assign w1983 = ~w1972 & ~w1982;
assign w1984 = w1362 & w1877;
assign w1985 = (pi0136 & ~w1832) | (pi0136 & w6845) | (~w1832 & w6845);
assign w1986 = ~w1834 & ~w1985;
assign w1987 = w1885 & w6846;
assign w1988 = w678 & w1644;
assign w1989 = ~w1984 & ~w1988;
assign w1990 = ~w1987 & w1989;
assign w1991 = ~pi0039 & pi0137;
assign w1992 = pi0039 & w495;
assign w1993 = w746 & w6847;
assign w1994 = ~w1991 & ~w1993;
assign w1995 = w1345 & w6848;
assign w1996 = (pi0138 & ~w1345) | (pi0138 & w6849) | (~w1345 & w6849);
assign w1997 = w1345 & w6850;
assign w1998 = ~w1996 & ~w1997;
assign w1999 = w1780 & w6851;
assign w2000 = ~w1281 & w1362;
assign w2001 = ~w1999 & ~w2000;
assign w2002 = (pi0139 & ~w1345) | (pi0139 & w6852) | (~w1345 & w6852);
assign w2003 = ~w1995 & ~w2002;
assign w2004 = w1780 & w6853;
assign w2005 = ~w1281 & w1310;
assign w2006 = ~w2004 & ~w2005;
assign w2007 = (pi0120 & ~w1422) | (pi0120 & w6854) | (~w1422 & w6854);
assign w2008 = w713 & w6418;
assign w2009 = (~pi0287 & w2008) | (~pi0287 & w6855) | (w2008 & w6855);
assign w2010 = (w350 & w2009) | (w350 & w6856) | (w2009 & w6856);
assign w2011 = w433 & w6419;
assign w2012 = (~w265 & w1417) | (~w265 & w6420) | (w1417 & w6420);
assign w2013 = (pi0252 & w2012) | (pi0252 & w6857) | (w2012 & w6857);
assign w2014 = ~pi0841 & pi1087;
assign w2015 = ~w264 & w2014;
assign w2016 = w392 & w6858;
assign w2017 = ~w198 & ~w329;
assign w2018 = ~w462 & ~w1432;
assign w2019 = w2018 & w6859;
assign w2020 = ~w2016 & w2019;
assign w2021 = ~w2013 & w2020;
assign w2022 = w2021 & w6860;
assign w2023 = (~pi0140 & w2022) | (~pi0140 & w6861) | (w2022 & w6861);
assign w2024 = pi0621 & pi1085;
assign w2025 = pi0644 & pi1154;
assign w2026 = ~pi0644 & ~pi1154;
assign w2027 = pi0790 & ~w2025;
assign w2028 = ~pi0629 & ~pi1150;
assign w2029 = pi0629 & pi1150;
assign w2030 = pi0792 & ~w2028;
assign w2031 = ~w2029 & w2030;
assign w2032 = ~pi0626 & pi1152;
assign w2033 = pi0626 & ~pi1152;
assign w2034 = ~w2032 & ~w2033;
assign w2035 = pi0788 & ~w2034;
assign w2036 = ~pi0608 & ~pi1147;
assign w2037 = pi0608 & pi1147;
assign w2038 = pi0778 & ~w2036;
assign w2039 = ~w2037 & w2038;
assign w2040 = ~pi0630 & ~pi1151;
assign w2041 = pi0630 & pi1151;
assign w2042 = pi0787 & ~w2040;
assign w2043 = ~w2041 & w2042;
assign w2044 = ~pi0618 & ~pi1148;
assign w2045 = pi0618 & pi1148;
assign w2046 = pi0781 & ~w2044;
assign w2047 = ~w2045 & w2046;
assign w2048 = ~pi0609 & ~pi1149;
assign w2049 = pi0609 & pi1149;
assign w2050 = pi0785 & ~w2048;
assign w2051 = ~w2049 & w2050;
assign w2052 = ~pi0619 & ~pi1153;
assign w2053 = pi0619 & pi1153;
assign w2054 = pi0789 & ~w2052;
assign w2055 = ~w2053 & w2054;
assign w2056 = (pi0603 & ~w2027) | (pi0603 & w6862) | (~w2027 & w6862);
assign w2057 = ~w2031 & ~w2035;
assign w2058 = ~w2039 & ~w2043;
assign w2059 = ~w2047 & ~w2051;
assign w2060 = ~w2055 & w2059;
assign w2061 = w2057 & w2058;
assign w2062 = w2056 & w2061;
assign w2063 = w2060 & w2062;
assign w2064 = w2062 & w6863;
assign w2065 = ~pi0761 & w1254;
assign w2066 = w2064 & w2065;
assign w2067 = pi0665 & pi1085;
assign w2068 = pi0715 & pi1154;
assign w2069 = ~pi0715 & ~pi1154;
assign w2070 = pi0790 & ~w2068;
assign w2071 = ~pi0647 & ~pi1151;
assign w2072 = pi0647 & pi1151;
assign w2073 = pi0787 & ~w2071;
assign w2074 = ~w2072 & w2073;
assign w2075 = ~pi0641 & pi1152;
assign w2076 = pi0641 & ~pi1152;
assign w2077 = ~w2075 & ~w2076;
assign w2078 = pi0788 & ~w2077;
assign w2079 = ~pi0627 & ~pi1148;
assign w2080 = pi0627 & pi1148;
assign w2081 = pi0781 & ~w2079;
assign w2082 = ~w2080 & w2081;
assign w2083 = ~pi0660 & ~pi1149;
assign w2084 = pi0660 & pi1149;
assign w2085 = pi0785 & ~w2083;
assign w2086 = ~w2084 & w2085;
assign w2087 = ~pi0625 & ~pi1147;
assign w2088 = pi0625 & pi1147;
assign w2089 = pi0778 & ~w2087;
assign w2090 = ~w2088 & w2089;
assign w2091 = ~pi0628 & ~pi1150;
assign w2092 = pi0628 & pi1150;
assign w2093 = pi0792 & ~w2091;
assign w2094 = ~w2092 & w2093;
assign w2095 = ~pi0648 & ~pi1153;
assign w2096 = pi0648 & pi1153;
assign w2097 = pi0789 & ~w2095;
assign w2098 = ~w2096 & w2097;
assign w2099 = (pi0680 & ~w2070) | (pi0680 & w6864) | (~w2070 & w6864);
assign w2100 = ~w2074 & ~w2078;
assign w2101 = ~w2082 & ~w2086;
assign w2102 = ~w2090 & ~w2094;
assign w2103 = ~w2098 & w2102;
assign w2104 = w2100 & w2101;
assign w2105 = w2099 & w2104;
assign w2106 = w2103 & w2105;
assign w2107 = w2105 & w6865;
assign w2108 = ~w2064 & w2107;
assign w2109 = ~pi0738 & w1254;
assign w2110 = w2108 & w2109;
assign w2111 = ~w2066 & ~w2110;
assign w2112 = ~w2022 & ~w2111;
assign w2113 = ~w2023 & ~w2112;
assign w2114 = (~pi0141 & w2022) | (~pi0141 & w6866) | (w2022 & w6866);
assign w2115 = pi0749 & w1254;
assign w2116 = w2064 & w2115;
assign w2117 = pi0706 & w1254;
assign w2118 = w2108 & w2117;
assign w2119 = ~w2116 & ~w2118;
assign w2120 = ~w2022 & ~w2119;
assign w2121 = ~w2114 & ~w2120;
assign w2122 = (pi0142 & w2022) | (pi0142 & w6867) | (w2022 & w6867);
assign w2123 = pi0743 & w1254;
assign w2124 = w2064 & w2123;
assign w2125 = pi0735 & w1254;
assign w2126 = w2108 & w2125;
assign w2127 = ~w2124 & ~w2126;
assign w2128 = ~w2022 & ~w2127;
assign w2129 = ~w2122 & ~w2128;
assign w2130 = (~pi0143 & w2022) | (~pi0143 & w6868) | (w2022 & w6868);
assign w2131 = ~pi0774 & w1254;
assign w2132 = w2064 & w2131;
assign w2133 = pi0687 & w1254;
assign w2134 = w2108 & w2133;
assign w2135 = ~w2132 & ~w2134;
assign w2136 = ~w2022 & ~w2135;
assign w2137 = ~w2130 & ~w2136;
assign w2138 = (pi0144 & w2022) | (pi0144 & w6869) | (w2022 & w6869);
assign w2139 = pi0758 & w1254;
assign w2140 = w2064 & w2139;
assign w2141 = pi0736 & w1254;
assign w2142 = w2108 & w2141;
assign w2143 = ~w2140 & ~w2142;
assign w2144 = ~w2022 & ~w2143;
assign w2145 = ~w2138 & ~w2144;
assign w2146 = (~pi0145 & w2022) | (~pi0145 & w6870) | (w2022 & w6870);
assign w2147 = ~pi0767 & w1254;
assign w2148 = w2064 & w2147;
assign w2149 = ~pi0698 & w1254;
assign w2150 = w2108 & w2149;
assign w2151 = ~w2148 & ~w2150;
assign w2152 = ~w2022 & ~w2151;
assign w2153 = ~w2146 & ~w2152;
assign w2154 = (pi0146 & w2022) | (pi0146 & w6871) | (w2022 & w6871);
assign w2155 = w1254 & w6872;
assign w2156 = pi0907 & ~pi0947;
assign w2157 = w1254 & w2156;
assign w2158 = pi0735 & w2157;
assign w2159 = ~w2155 & ~w2158;
assign w2160 = ~w2022 & ~w2159;
assign w2161 = ~w2154 & ~w2160;
assign w2162 = (~pi0147 & w2022) | (~pi0147 & w6873) | (w2022 & w6873);
assign w2163 = ~pi0770 & w1254;
assign w2164 = w1254 & w6874;
assign w2165 = pi0726 & w2157;
assign w2166 = ~w2164 & ~w2165;
assign w2167 = ~w2022 & ~w2166;
assign w2168 = ~w2162 & ~w2167;
assign w2169 = (~pi0148 & w2022) | (~pi0148 & w6875) | (w2022 & w6875);
assign w2170 = w1254 & w6876;
assign w2171 = pi0706 & w2157;
assign w2172 = ~w2170 & ~w2171;
assign w2173 = ~w2022 & ~w2172;
assign w2174 = ~w2169 & ~w2173;
assign w2175 = (~pi0149 & w2022) | (~pi0149 & w6877) | (w2022 & w6877);
assign w2176 = ~pi0755 & w1254;
assign w2177 = w1254 & w6878;
assign w2178 = ~pi0725 & w2157;
assign w2179 = ~w2177 & ~w2178;
assign w2180 = ~w2022 & ~w2179;
assign w2181 = ~w2175 & ~w2180;
assign w2182 = (~pi0150 & w2022) | (~pi0150 & w6879) | (w2022 & w6879);
assign w2183 = ~pi0751 & w1254;
assign w2184 = w1254 & w6880;
assign w2185 = ~pi0701 & w2157;
assign w2186 = ~w2184 & ~w2185;
assign w2187 = ~w2022 & ~w2186;
assign w2188 = ~w2182 & ~w2187;
assign w2189 = (~pi0151 & w2022) | (~pi0151 & w6881) | (w2022 & w6881);
assign w2190 = ~pi0745 & w1254;
assign w2191 = w1254 & w6882;
assign w2192 = ~pi0723 & w2157;
assign w2193 = ~w2191 & ~w2192;
assign w2194 = ~w2022 & ~w2193;
assign w2195 = ~w2189 & ~w2194;
assign w2196 = (pi0152 & w2022) | (pi0152 & w6883) | (w2022 & w6883);
assign w2197 = pi0759 & w1254;
assign w2198 = w1254 & w6884;
assign w2199 = pi0696 & w2157;
assign w2200 = ~w2198 & ~w2199;
assign w2201 = ~w2022 & ~w2200;
assign w2202 = ~w2196 & ~w2201;
assign w2203 = (~pi0153 & w2022) | (~pi0153 & w6885) | (w2022 & w6885);
assign w2204 = pi0766 & w1254;
assign w2205 = w1254 & w6886;
assign w2206 = pi0700 & w2157;
assign w2207 = ~w2205 & ~w2206;
assign w2208 = ~w2022 & ~w2207;
assign w2209 = ~w2203 & ~w2208;
assign w2210 = (~pi0154 & w2022) | (~pi0154 & w6887) | (w2022 & w6887);
assign w2211 = ~pi0742 & w1254;
assign w2212 = w1254 & w6888;
assign w2213 = ~pi0704 & w2157;
assign w2214 = ~w2212 & ~w2213;
assign w2215 = ~w2022 & ~w2214;
assign w2216 = ~w2210 & ~w2215;
assign w2217 = (~pi0155 & w2022) | (~pi0155 & w6889) | (w2022 & w6889);
assign w2218 = ~pi0757 & w1254;
assign w2219 = w1254 & w6890;
assign w2220 = ~pi0686 & w2157;
assign w2221 = ~w2219 & ~w2220;
assign w2222 = ~w2022 & ~w2221;
assign w2223 = ~w2217 & ~w2222;
assign w2224 = (~pi0156 & w2022) | (~pi0156 & w6891) | (w2022 & w6891);
assign w2225 = ~pi0741 & w1254;
assign w2226 = w1254 & w6892;
assign w2227 = ~pi0724 & w2157;
assign w2228 = ~w2226 & ~w2227;
assign w2229 = ~w2022 & ~w2228;
assign w2230 = ~w2224 & ~w2229;
assign w2231 = (~pi0157 & w2022) | (~pi0157 & w6893) | (w2022 & w6893);
assign w2232 = ~pi0760 & w1254;
assign w2233 = w1254 & w6894;
assign w2234 = ~pi0688 & w2157;
assign w2235 = ~w2233 & ~w2234;
assign w2236 = ~w2022 & ~w2235;
assign w2237 = ~w2231 & ~w2236;
assign w2238 = (~pi0158 & w2022) | (~pi0158 & w6895) | (w2022 & w6895);
assign w2239 = ~pi0753 & w1254;
assign w2240 = w1254 & w6896;
assign w2241 = ~pi0702 & w2157;
assign w2242 = ~w2240 & ~w2241;
assign w2243 = ~w2022 & ~w2242;
assign w2244 = ~w2238 & ~w2243;
assign w2245 = (~pi0159 & w2022) | (~pi0159 & w6897) | (w2022 & w6897);
assign w2246 = ~pi0754 & w1254;
assign w2247 = w1254 & w6898;
assign w2248 = ~pi0709 & w2157;
assign w2249 = ~w2247 & ~w2248;
assign w2250 = ~w2022 & ~w2249;
assign w2251 = ~w2245 & ~w2250;
assign w2252 = (~pi0160 & w2022) | (~pi0160 & w6899) | (w2022 & w6899);
assign w2253 = ~pi0756 & w1254;
assign w2254 = w1254 & w6900;
assign w2255 = ~pi0734 & w2157;
assign w2256 = ~w2254 & ~w2255;
assign w2257 = ~w2022 & ~w2256;
assign w2258 = ~w2252 & ~w2257;
assign w2259 = (pi0161 & w2022) | (pi0161 & w6901) | (w2022 & w6901);
assign w2260 = w1254 & w6902;
assign w2261 = pi0736 & w2157;
assign w2262 = ~w2260 & ~w2261;
assign w2263 = ~w2022 & ~w2262;
assign w2264 = ~w2259 & ~w2263;
assign w2265 = (~pi0162 & w2022) | (~pi0162 & w6903) | (w2022 & w6903);
assign w2266 = w1254 & w6904;
assign w2267 = ~pi0738 & w2157;
assign w2268 = ~w2266 & ~w2267;
assign w2269 = ~w2022 & ~w2268;
assign w2270 = ~w2265 & ~w2269;
assign w2271 = (~pi0163 & w2022) | (~pi0163 & w6905) | (w2022 & w6905);
assign w2272 = ~pi0777 & w1254;
assign w2273 = w1254 & w6906;
assign w2274 = ~pi0737 & w2157;
assign w2275 = ~w2273 & ~w2274;
assign w2276 = ~w2022 & ~w2275;
assign w2277 = ~w2271 & ~w2276;
assign w2278 = (~pi0164 & w2022) | (~pi0164 & w6907) | (w2022 & w6907);
assign w2279 = ~pi0752 & w1254;
assign w2280 = w1254 & w6908;
assign w2281 = pi0703 & w2157;
assign w2282 = ~w2280 & ~w2281;
assign w2283 = ~w2022 & ~w2282;
assign w2284 = ~w2278 & ~w2283;
assign w2285 = (~pi0165 & w2022) | (~pi0165 & w6909) | (w2022 & w6909);
assign w2286 = w1254 & w6910;
assign w2287 = pi0687 & w2157;
assign w2288 = ~w2286 & ~w2287;
assign w2289 = ~w2022 & ~w2288;
assign w2290 = ~w2285 & ~w2289;
assign w2291 = (pi0166 & w2022) | (pi0166 & w6911) | (w2022 & w6911);
assign w2292 = pi0772 & w1254;
assign w2293 = w1254 & w6912;
assign w2294 = pi0727 & w2157;
assign w2295 = ~w2293 & ~w2294;
assign w2296 = ~w2022 & ~w2295;
assign w2297 = ~w2291 & ~w2296;
assign w2298 = (~pi0167 & w2022) | (~pi0167 & w6913) | (w2022 & w6913);
assign w2299 = ~pi0768 & w1254;
assign w2300 = w1254 & w6914;
assign w2301 = pi0705 & w2157;
assign w2302 = ~w2300 & ~w2301;
assign w2303 = ~w2022 & ~w2302;
assign w2304 = ~w2298 & ~w2303;
assign w2305 = (~pi0168 & w2022) | (~pi0168 & w6915) | (w2022 & w6915);
assign w2306 = pi0763 & w1254;
assign w2307 = w1254 & w6916;
assign w2308 = pi0699 & w2157;
assign w2309 = ~w2307 & ~w2308;
assign w2310 = ~w2022 & ~w2309;
assign w2311 = ~w2305 & ~w2310;
assign w2312 = (~pi0169 & w2022) | (~pi0169 & w6917) | (w2022 & w6917);
assign w2313 = pi0746 & w1254;
assign w2314 = w1254 & w6918;
assign w2315 = pi0729 & w2157;
assign w2316 = ~w2314 & ~w2315;
assign w2317 = ~w2022 & ~w2316;
assign w2318 = ~w2312 & ~w2317;
assign w2319 = (~pi0170 & w2022) | (~pi0170 & w6919) | (w2022 & w6919);
assign w2320 = pi0748 & w1254;
assign w2321 = w1254 & w6920;
assign w2322 = pi0730 & w2157;
assign w2323 = ~w2321 & ~w2322;
assign w2324 = ~w2022 & ~w2323;
assign w2325 = ~w2319 & ~w2324;
assign w2326 = (~pi0171 & w2022) | (~pi0171 & w6921) | (w2022 & w6921);
assign w2327 = pi0764 & w1254;
assign w2328 = w1254 & w6922;
assign w2329 = pi0691 & w2157;
assign w2330 = ~w2328 & ~w2329;
assign w2331 = ~w2022 & ~w2330;
assign w2332 = ~w2326 & ~w2331;
assign w2333 = (~pi0172 & w2022) | (~pi0172 & w6923) | (w2022 & w6923);
assign w2334 = pi0739 & w1254;
assign w2335 = w1254 & w6924;
assign w2336 = pi0690 & w2157;
assign w2337 = ~w2335 & ~w2336;
assign w2338 = ~w2022 & ~w2337;
assign w2339 = ~w2333 & ~w2338;
assign w2340 = (~pi0173 & w2022) | (~pi0173 & w6925) | (w2022 & w6925);
assign w2341 = w2064 & w2190;
assign w2342 = ~pi0723 & w1254;
assign w2343 = w2108 & w2342;
assign w2344 = ~w2341 & ~w2343;
assign w2345 = ~w2022 & ~w2344;
assign w2346 = ~w2340 & ~w2345;
assign w2347 = (pi0174 & w2022) | (pi0174 & w6926) | (w2022 & w6926);
assign w2348 = w2064 & w2197;
assign w2349 = pi0696 & w1254;
assign w2350 = w2108 & w2349;
assign w2351 = ~w2348 & ~w2350;
assign w2352 = ~w2022 & ~w2351;
assign w2353 = ~w2347 & ~w2352;
assign w2354 = (~pi0175 & w2022) | (~pi0175 & w6927) | (w2022 & w6927);
assign w2355 = w2064 & w2204;
assign w2356 = pi0700 & w1254;
assign w2357 = w2108 & w2356;
assign w2358 = ~w2355 & ~w2357;
assign w2359 = ~w2022 & ~w2358;
assign w2360 = ~w2354 & ~w2359;
assign w2361 = (~pi0176 & w2022) | (~pi0176 & w6928) | (w2022 & w6928);
assign w2362 = w2064 & w2211;
assign w2363 = ~pi0704 & w1254;
assign w2364 = w2108 & w2363;
assign w2365 = ~w2362 & ~w2364;
assign w2366 = ~w2022 & ~w2365;
assign w2367 = ~w2361 & ~w2366;
assign w2368 = (~pi0177 & w2022) | (~pi0177 & w6929) | (w2022 & w6929);
assign w2369 = w2064 & w2218;
assign w2370 = ~pi0686 & w1254;
assign w2371 = w2108 & w2370;
assign w2372 = ~w2369 & ~w2371;
assign w2373 = ~w2022 & ~w2372;
assign w2374 = ~w2368 & ~w2373;
assign w2375 = (~pi0178 & w2022) | (~pi0178 & w6930) | (w2022 & w6930);
assign w2376 = w2064 & w2232;
assign w2377 = ~pi0688 & w1254;
assign w2378 = w2108 & w2377;
assign w2379 = ~w2376 & ~w2378;
assign w2380 = ~w2022 & ~w2379;
assign w2381 = ~w2375 & ~w2380;
assign w2382 = (~pi0179 & w2022) | (~pi0179 & w6931) | (w2022 & w6931);
assign w2383 = w2064 & w2225;
assign w2384 = ~pi0724 & w1254;
assign w2385 = w2108 & w2384;
assign w2386 = ~w2383 & ~w2385;
assign w2387 = ~w2022 & ~w2386;
assign w2388 = ~w2382 & ~w2387;
assign w2389 = (~pi0180 & w2022) | (~pi0180 & w6932) | (w2022 & w6932);
assign w2390 = w2064 & w2239;
assign w2391 = ~pi0702 & w1254;
assign w2392 = w2108 & w2391;
assign w2393 = ~w2390 & ~w2392;
assign w2394 = ~w2022 & ~w2393;
assign w2395 = ~w2389 & ~w2394;
assign w2396 = (~pi0181 & w2022) | (~pi0181 & w6933) | (w2022 & w6933);
assign w2397 = w2064 & w2246;
assign w2398 = ~pi0709 & w1254;
assign w2399 = w2108 & w2398;
assign w2400 = ~w2397 & ~w2399;
assign w2401 = ~w2022 & ~w2400;
assign w2402 = ~w2396 & ~w2401;
assign w2403 = (~pi0182 & w2022) | (~pi0182 & w6934) | (w2022 & w6934);
assign w2404 = w2064 & w2253;
assign w2405 = ~pi0734 & w1254;
assign w2406 = w2108 & w2405;
assign w2407 = ~w2404 & ~w2406;
assign w2408 = ~w2022 & ~w2407;
assign w2409 = ~w2403 & ~w2408;
assign w2410 = (~pi0183 & w2022) | (~pi0183 & w6935) | (w2022 & w6935);
assign w2411 = w2064 & w2176;
assign w2412 = ~pi0725 & w1254;
assign w2413 = w2108 & w2412;
assign w2414 = ~w2411 & ~w2413;
assign w2415 = ~w2022 & ~w2414;
assign w2416 = ~w2410 & ~w2415;
assign w2417 = (~pi0184 & w2022) | (~pi0184 & w6936) | (w2022 & w6936);
assign w2418 = w2064 & w2272;
assign w2419 = ~pi0737 & w1254;
assign w2420 = w2108 & w2419;
assign w2421 = ~w2418 & ~w2420;
assign w2422 = ~w2022 & ~w2421;
assign w2423 = ~w2417 & ~w2422;
assign w2424 = (~pi0185 & w2022) | (~pi0185 & w6937) | (w2022 & w6937);
assign w2425 = w2064 & w2183;
assign w2426 = ~pi0701 & w1254;
assign w2427 = w2108 & w2426;
assign w2428 = ~w2425 & ~w2427;
assign w2429 = ~w2022 & ~w2428;
assign w2430 = ~w2424 & ~w2429;
assign w2431 = (~pi0186 & w2022) | (~pi0186 & w6938) | (w2022 & w6938);
assign w2432 = w2064 & w2279;
assign w2433 = pi0703 & w1254;
assign w2434 = w2108 & w2433;
assign w2435 = ~w2432 & ~w2434;
assign w2436 = ~w2022 & ~w2435;
assign w2437 = ~w2431 & ~w2436;
assign w2438 = (~pi0187 & w2022) | (~pi0187 & w6939) | (w2022 & w6939);
assign w2439 = w2064 & w2163;
assign w2440 = pi0726 & w1254;
assign w2441 = w2108 & w2440;
assign w2442 = ~w2439 & ~w2441;
assign w2443 = ~w2022 & ~w2442;
assign w2444 = ~w2438 & ~w2443;
assign w2445 = (~pi0188 & w2022) | (~pi0188 & w6940) | (w2022 & w6940);
assign w2446 = w2064 & w2299;
assign w2447 = pi0705 & w1254;
assign w2448 = w2108 & w2447;
assign w2449 = ~w2446 & ~w2448;
assign w2450 = ~w2022 & ~w2449;
assign w2451 = ~w2445 & ~w2450;
assign w2452 = (pi0189 & w2022) | (pi0189 & w6941) | (w2022 & w6941);
assign w2453 = w2064 & w2292;
assign w2454 = pi0727 & w1254;
assign w2455 = w2108 & w2454;
assign w2456 = ~w2453 & ~w2455;
assign w2457 = ~w2022 & ~w2456;
assign w2458 = ~w2452 & ~w2457;
assign w2459 = (~pi0190 & w2022) | (~pi0190 & w6942) | (w2022 & w6942);
assign w2460 = w2064 & w2306;
assign w2461 = pi0699 & w1254;
assign w2462 = w2108 & w2461;
assign w2463 = ~w2460 & ~w2462;
assign w2464 = ~w2022 & ~w2463;
assign w2465 = ~w2459 & ~w2464;
assign w2466 = (~pi0191 & w2022) | (~pi0191 & w6943) | (w2022 & w6943);
assign w2467 = w2064 & w2313;
assign w2468 = pi0729 & w1254;
assign w2469 = w2108 & w2468;
assign w2470 = ~w2467 & ~w2469;
assign w2471 = ~w2022 & ~w2470;
assign w2472 = ~w2466 & ~w2471;
assign w2473 = (~pi0192 & w2022) | (~pi0192 & w6944) | (w2022 & w6944);
assign w2474 = w2064 & w2327;
assign w2475 = pi0691 & w1254;
assign w2476 = w2108 & w2475;
assign w2477 = ~w2474 & ~w2476;
assign w2478 = ~w2022 & ~w2477;
assign w2479 = ~w2473 & ~w2478;
assign w2480 = (~pi0193 & w2022) | (~pi0193 & w6945) | (w2022 & w6945);
assign w2481 = w2064 & w2334;
assign w2482 = pi0690 & w1254;
assign w2483 = w2108 & w2482;
assign w2484 = ~w2481 & ~w2483;
assign w2485 = ~w2022 & ~w2484;
assign w2486 = ~w2480 & ~w2485;
assign w2487 = (~pi0194 & w2022) | (~pi0194 & w6946) | (w2022 & w6946);
assign w2488 = w2064 & w2320;
assign w2489 = pi0730 & w1254;
assign w2490 = w2108 & w2489;
assign w2491 = ~w2488 & ~w2490;
assign w2492 = ~w2022 & ~w2491;
assign w2493 = ~w2487 & ~w2492;
assign w2494 = ~w1281 & w1966;
assign w2495 = w1345 & w6947;
assign w2496 = pi0195 & ~w2495;
assign w2497 = w1780 & w6948;
assign w2498 = ~w2494 & ~w2497;
assign w2499 = (pi0196 & ~w1345) | (pi0196 & w6949) | (~w1345 & w6949);
assign w2500 = ~w2495 & ~w2499;
assign w2501 = w1780 & w6950;
assign w2502 = ~w1281 & w1978;
assign w2503 = ~w2501 & ~w2502;
assign w2504 = (~pi0197 & w2022) | (~pi0197 & w6951) | (w2022 & w6951);
assign w2505 = pi0947 & w2147;
assign w2506 = ~pi0698 & w2157;
assign w2507 = ~w2505 & ~w2506;
assign w2508 = ~w2022 & ~w2507;
assign w2509 = ~w2504 & ~w2508;
assign w2510 = ~w2010 & w2021;
assign w2511 = (w1254 & ~w2021) | (w1254 & w6952) | (~w2021 & w6952);
assign w2512 = pi0634 & w2108;
assign w2513 = pi0633 & w2064;
assign w2514 = ~w2512 & ~w2513;
assign w2515 = w2511 & ~w2514;
assign w2516 = pi0198 & ~w2511;
assign w2517 = ~w2515 & ~w2516;
assign w2518 = pi0637 & w2108;
assign w2519 = pi0617 & w2064;
assign w2520 = ~w2518 & ~w2519;
assign w2521 = w2511 & ~w2520;
assign w2522 = pi0199 & ~w2511;
assign w2523 = ~w2521 & ~w2522;
assign w2524 = pi0643 & w2108;
assign w2525 = pi0606 & w2064;
assign w2526 = ~w2524 & ~w2525;
assign w2527 = w2511 & ~w2526;
assign w2528 = pi0200 & ~w2511;
assign w2529 = ~w2527 & ~w2528;
assign w2530 = pi0233 & pi0237;
assign w2531 = pi0096 & ~w495;
assign w2532 = ~w702 & w2531;
assign w2533 = w2530 & w2532;
assign w2534 = ~w45 & ~w101;
assign w2535 = w36 & ~w412;
assign w2536 = ~w472 & w2535;
assign w2537 = w395 & ~w2536;
assign w2538 = ~w2534 & w2537;
assign w2539 = ~w402 & ~w2538;
assign w2540 = w194 & ~w2539;
assign w2541 = ~pi0032 & pi0070;
assign w2542 = pi0032 & ~pi0070;
assign w2543 = (~w2541 & ~w495) | (~w2541 & w6955) | (~w495 & w6955);
assign w2544 = ~w702 & ~w2543;
assign w2545 = w2530 & w2544;
assign w2546 = (~w2540 & w6958) | (~w2540 & w6959) | (w6958 & w6959);
assign w2547 = ~w2533 & ~w2546;
assign w2548 = ~pi0233 & pi0237;
assign w2549 = w2532 & w2548;
assign w2550 = w2544 & w2548;
assign w2551 = (~w2540 & w6962) | (~w2540 & w6963) | (w6962 & w6963);
assign w2552 = ~w2549 & ~w2551;
assign w2553 = ~pi0233 & ~pi0237;
assign w2554 = w2532 & w2553;
assign w2555 = w2544 & w2553;
assign w2556 = (~w2540 & w6966) | (~w2540 & w6967) | (w6966 & w6967);
assign w2557 = ~w2554 & ~w2556;
assign w2558 = ~w710 & w2531;
assign w2559 = w2530 & w2558;
assign w2560 = ~w710 & ~w2543;
assign w2561 = w2530 & w2560;
assign w2562 = (~w2540 & w6971) | (~w2540 & w6972) | (w6971 & w6972);
assign w2563 = ~w2559 & ~w2562;
assign w2564 = w2548 & w2558;
assign w2565 = w2548 & w2560;
assign w2566 = (~w2540 & w6975) | (~w2540 & w6976) | (w6975 & w6976);
assign w2567 = ~w2564 & ~w2566;
assign w2568 = pi0233 & ~pi0237;
assign w2569 = w2558 & w2568;
assign w2570 = w2560 & w2568;
assign w2571 = (~w2540 & w6979) | (~w2540 & w6980) | (w6979 & w6980);
assign w2572 = ~w2569 & ~w2571;
assign w2573 = pi0710 & w2108;
assign w2574 = pi0623 & w2064;
assign w2575 = ~w2573 & ~w2574;
assign w2576 = w2511 & ~w2575;
assign w2577 = ~pi0207 & ~w2511;
assign w2578 = ~w2576 & ~w2577;
assign w2579 = pi0638 & w2108;
assign w2580 = pi0607 & w2064;
assign w2581 = ~w2579 & ~w2580;
assign w2582 = w2511 & ~w2581;
assign w2583 = ~pi0208 & ~w2511;
assign w2584 = ~w2582 & ~w2583;
assign w2585 = pi0639 & w2108;
assign w2586 = pi0622 & w2064;
assign w2587 = ~w2585 & ~w2586;
assign w2588 = w2511 & ~w2587;
assign w2589 = ~pi0209 & ~w2511;
assign w2590 = ~w2588 & ~w2589;
assign w2591 = pi0633 & pi0947;
assign w2592 = pi0634 & w2156;
assign w2593 = ~w2591 & ~w2592;
assign w2594 = w2511 & ~w2593;
assign w2595 = pi0210 & ~w2511;
assign w2596 = ~w2594 & ~w2595;
assign w2597 = pi0606 & pi0947;
assign w2598 = pi0643 & w2156;
assign w2599 = ~w2597 & ~w2598;
assign w2600 = w2511 & ~w2599;
assign w2601 = pi0211 & ~w2511;
assign w2602 = ~w2600 & ~w2601;
assign w2603 = pi0212 & ~w2511;
assign w2604 = pi0607 & pi0947;
assign w2605 = pi0638 & w2156;
assign w2606 = ~w2604 & ~w2605;
assign w2607 = w2511 & w2606;
assign w2608 = ~w2603 & ~w2607;
assign w2609 = pi0213 & ~w2511;
assign w2610 = pi0622 & pi0947;
assign w2611 = pi0639 & w2156;
assign w2612 = ~w2610 & ~w2611;
assign w2613 = w2511 & w2612;
assign w2614 = ~w2609 & ~w2613;
assign w2615 = pi0214 & ~w2511;
assign w2616 = pi0623 & pi0947;
assign w2617 = pi0710 & w2156;
assign w2618 = ~w2616 & ~w2617;
assign w2619 = w2511 & w2618;
assign w2620 = ~w2615 & ~w2619;
assign w2621 = pi0642 & pi0947;
assign w2622 = pi0681 & w2156;
assign w2623 = ~w2621 & ~w2622;
assign w2624 = w2511 & ~w2623;
assign w2625 = pi0215 & ~w2511;
assign w2626 = ~w2624 & ~w2625;
assign w2627 = pi0614 & pi0947;
assign w2628 = pi0662 & w2156;
assign w2629 = ~w2627 & ~w2628;
assign w2630 = w2511 & ~w2629;
assign w2631 = pi0216 & ~w2511;
assign w2632 = ~w2630 & ~w2631;
assign w2633 = ~pi0695 & w2108;
assign w2634 = pi0612 & w2064;
assign w2635 = ~w2633 & ~w2634;
assign w2636 = w2511 & ~w2635;
assign w2637 = ~pi0217 & ~w2511;
assign w2638 = ~w2636 & ~w2637;
assign w2639 = w2553 & w2558;
assign w2640 = w2553 & w2560;
assign w2641 = (~w2540 & w6981) | (~w2540 & w6982) | (w6981 & w6982);
assign w2642 = ~w2640 & w2641;
assign w2643 = ~w2639 & ~w2642;
assign w2644 = pi0617 & pi0947;
assign w2645 = pi0637 & w2156;
assign w2646 = ~w2644 & ~w2645;
assign w2647 = w2511 & ~w2646;
assign w2648 = pi0219 & ~w2511;
assign w2649 = ~w2647 & ~w2648;
assign w2650 = w2532 & w2568;
assign w2651 = w2544 & w2568;
assign w2652 = (~w2540 & w6983) | (~w2540 & w6984) | (w6983 & w6984);
assign w2653 = ~w2651 & w2652;
assign w2654 = ~w2650 & ~w2653;
assign w2655 = pi0616 & pi0947;
assign w2656 = pi0661 & w2156;
assign w2657 = ~w2655 & ~w2656;
assign w2658 = w2511 & ~w2657;
assign w2659 = pi0221 & ~w2511;
assign w2660 = ~w2658 & ~w2659;
assign w2661 = pi0661 & w2108;
assign w2662 = pi0616 & w2064;
assign w2663 = ~w2661 & ~w2662;
assign w2664 = w2511 & ~w2663;
assign w2665 = pi0222 & ~w2511;
assign w2666 = ~w2664 & ~w2665;
assign w2667 = pi0681 & w2108;
assign w2668 = pi0642 & w2064;
assign w2669 = ~w2667 & ~w2668;
assign w2670 = w2511 & ~w2669;
assign w2671 = pi0223 & ~w2511;
assign w2672 = ~w2670 & ~w2671;
assign w2673 = pi0662 & w2108;
assign w2674 = pi0614 & w2064;
assign w2675 = ~w2673 & ~w2674;
assign w2676 = w2511 & ~w2675;
assign w2677 = pi0224 & ~w2511;
assign w2678 = ~w2676 & ~w2677;
assign w2679 = pi0228 & pi0231;
assign w2680 = pi0479 & w388;
assign w2681 = w225 & w6985;
assign w2682 = ~w298 & ~w382;
assign w2683 = ~w2680 & w2682;
assign w2684 = w2683 & w6986;
assign w2685 = w367 & w2684;
assign w2686 = w2681 & w2685;
assign w2687 = (~pi0228 & ~w2681) | (~pi0228 & w6987) | (~w2681 & w6987);
assign w2688 = ~w2679 & ~w2687;
assign w2689 = w301 & w1499;
assign w2690 = w468 & ~w1416;
assign w2691 = ~w1502 & ~w2689;
assign w2692 = w2690 & w2691;
assign w2693 = ~w1596 & w2692;
assign w2694 = ~pi0039 & pi0228;
assign w2695 = (~w253 & ~w257) | (~w253 & w6988) | (~w257 & w6988);
assign w2696 = (w208 & ~w1582) | (w208 & w6989) | (~w1582 & w6989);
assign w2697 = ~w2695 & ~w2696;
assign w2698 = ~w2694 & ~w2697;
assign w2699 = ~w324 & ~w392;
assign w2700 = ~w1433 & w2699;
assign w2701 = w463 & w2700;
assign w2702 = w673 & w2701;
assign w2703 = w2702 & w6990;
assign w2704 = w2681 & w2703;
assign w2705 = ~pi0230 & pi0233;
assign w2706 = (pi0213 & ~w2) | (pi0213 & w6991) | (~w2 & w6991);
assign w2707 = w2 & w6992;
assign w2708 = ~w2706 & ~w2707;
assign w2709 = pi0230 & ~w2708;
assign w2710 = pi1138 & w1477;
assign w2711 = w1460 & ~w1463;
assign w2712 = ~w1460 & w1463;
assign w2713 = ~w2711 & ~w2712;
assign w2714 = w2710 & ~w2713;
assign w2715 = ~w1457 & w1467;
assign w2716 = ~w1479 & w2715;
assign w2717 = ~w1469 & ~w2716;
assign w2718 = pi1136 & ~w2717;
assign w2719 = w1480 & w6993;
assign w2720 = ~w2714 & ~w2718;
assign w2721 = w2720 & w6994;
assign w2722 = pi1149 & w1477;
assign w2723 = pi1148 & w1468;
assign w2724 = ~w2722 & ~w2723;
assign w2725 = w1464 & ~w2724;
assign w2726 = pi1149 & w1468;
assign w2727 = pi1150 & w1477;
assign w2728 = ~w2726 & ~w2727;
assign w2729 = w2711 & ~w2728;
assign w2730 = ~w2725 & ~w2729;
assign w2731 = pi1148 & w2715;
assign w2732 = pi1150 & w1468;
assign w2733 = pi1151 & w1477;
assign w2734 = pi1149 & w2715;
assign w2735 = ~w2732 & ~w2733;
assign w2736 = (w2712 & ~w2735) | (w2712 & w6995) | (~w2735 & w6995);
assign w2737 = pi0230 & w2708;
assign w2738 = pi1147 & w2715;
assign w2739 = w1464 & w2738;
assign w2740 = (w2737 & ~w2731) | (w2737 & w6996) | (~w2731 & w6996);
assign w2741 = ~w2739 & w2740;
assign w2742 = w2730 & w6997;
assign w2743 = ~w2705 & ~w2742;
assign w2744 = ~w2721 & w2743;
assign w2745 = ~pi0230 & pi0234;
assign w2746 = (~w2731 & w2728) | (~w2731 & w6998) | (w2728 & w6998);
assign w2747 = ~w1479 & ~w2746;
assign w2748 = w2730 & ~w2747;
assign w2749 = pi1148 & w1477;
assign w2750 = ~w2713 & w2749;
assign w2751 = pi1146 & ~w2717;
assign w2752 = w1480 & w6999;
assign w2753 = ~w2750 & ~w2751;
assign w2754 = ~w2752 & w2753;
assign w2755 = (w2737 & ~w2753) | (w2737 & w7000) | (~w2753 & w7000);
assign w2756 = (~w2745 & w2748) | (~w2745 & w7001) | (w2748 & w7001);
assign w2757 = ~w2755 & w2756;
assign w2758 = ~pi0230 & ~pi0235;
assign w2759 = pi1147 & w1469;
assign w2760 = ~w2722 & ~w2738;
assign w2761 = ~w2713 & ~w2760;
assign w2762 = w1480 & w7002;
assign w2763 = ~w2759 & ~w2761;
assign w2764 = w2763 & w7003;
assign w2765 = w1464 & ~w2728;
assign w2766 = (w2711 & ~w2735) | (w2711 & w7004) | (~w2735 & w7004);
assign w2767 = ~w2765 & ~w2766;
assign w2768 = w2709 & ~w2736;
assign w2769 = w2767 & w2768;
assign w2770 = ~w2758 & ~w2769;
assign w2771 = ~w2764 & w2770;
assign w2772 = ~pi0230 & pi0237;
assign w2773 = pi1139 & w1477;
assign w2774 = ~w2713 & w2773;
assign w2775 = pi1137 & ~w2717;
assign w2776 = w1480 & w7005;
assign w2777 = ~w2774 & ~w2775;
assign w2778 = ~w2776 & w2777;
assign w2779 = w2777 & w7006;
assign w2780 = pi1152 & w1477;
assign w2781 = pi1150 & w2715;
assign w2782 = pi1151 & w1468;
assign w2783 = ~w2780 & ~w2781;
assign w2784 = (w2712 & ~w2783) | (w2712 & w7007) | (~w2783 & w7007);
assign w2785 = (w2737 & ~w2731) | (w2737 & w7008) | (~w2731 & w7008);
assign w2786 = ~w2784 & w2785;
assign w2787 = w2767 & w2786;
assign w2788 = ~w2772 & ~w2787;
assign w2789 = ~w2779 & w2788;
assign w2790 = ~pi0230 & pi0238;
assign w2791 = w2763 & w7009;
assign w2792 = w2709 & ~w2791;
assign w2793 = pi1147 & w1477;
assign w2794 = ~w2713 & w2793;
assign w2795 = pi1145 & ~w2717;
assign w2796 = w1480 & w7010;
assign w2797 = ~w2794 & ~w2795;
assign w2798 = (w2737 & ~w2797) | (w2737 & w7011) | (~w2797 & w7011);
assign w2799 = ~w2790 & ~w2798;
assign w2800 = ~w2792 & w2799;
assign w2801 = ~pi0230 & pi0239;
assign w2802 = w2712 & w2737;
assign w2803 = ~w2746 & w2802;
assign w2804 = (~w2801 & ~w2784) | (~w2801 & w7012) | (~w2784 & w7012);
assign w2805 = ~w2803 & w2804;
assign w2806 = pi1141 & w1477;
assign w2807 = ~w2713 & w2806;
assign w2808 = pi1139 & ~w2717;
assign w2809 = w1480 & w7013;
assign w2810 = ~w2807 & ~w2808;
assign w2811 = (w2737 & ~w2810) | (w2737 & w7014) | (~w2810 & w7014);
assign w2812 = pi1143 & w1477;
assign w2813 = ~w2713 & w2812;
assign w2814 = pi1141 & ~w2717;
assign w2815 = w1480 & w7015;
assign w2816 = ~w2813 & ~w2814;
assign w2817 = (w2709 & ~w2816) | (w2709 & w7016) | (~w2816 & w7016);
assign w2818 = ~pi0230 & pi0240;
assign w2819 = ~w2811 & ~w2818;
assign w2820 = ~w2817 & w2819;
assign w2821 = (w2709 & ~w2797) | (w2709 & w7017) | (~w2797 & w7017);
assign w2822 = pi1145 & w1477;
assign w2823 = ~w2713 & w2822;
assign w2824 = pi1143 & ~w2717;
assign w2825 = w1480 & w7018;
assign w2826 = ~w2823 & ~w2824;
assign w2827 = ~w2825 & w2826;
assign w2828 = (w2737 & ~w2826) | (w2737 & w7019) | (~w2826 & w7019);
assign w2829 = ~pi0230 & pi0241;
assign w2830 = ~w2821 & ~w2829;
assign w2831 = ~w2828 & w2830;
assign w2832 = pi1140 & w1477;
assign w2833 = ~w2713 & w2832;
assign w2834 = pi1138 & ~w2717;
assign w2835 = w1480 & w7020;
assign w2836 = ~w2833 & ~w2834;
assign w2837 = (w2709 & ~w2836) | (w2709 & w7021) | (~w2836 & w7021);
assign w2838 = (w2737 & ~w2720) | (w2737 & w7022) | (~w2720 & w7022);
assign w2839 = ~pi0230 & pi0242;
assign w2840 = ~w2837 & ~w2839;
assign w2841 = ~w2838 & w2840;
assign w2842 = ~pi0083 & ~pi0085;
assign w2843 = (w1457 & w7023) | (w1457 & w7024) | (w7023 & w7024);
assign w2844 = w2843 & w7025;
assign w2845 = w2843 & w7026;
assign w2846 = w2843 & w7028;
assign w2847 = w2843 & w7029;
assign w2848 = pi0275 & w2847;
assign w2849 = w2847 & w7030;
assign w2850 = pi0253 & pi0254;
assign w2851 = pi0267 & w2850;
assign w2852 = w2850 & w7031;
assign w2853 = ~pi0230 & ~pi1085;
assign w2854 = (w2853 & ~w2847) | (w2853 & w7033) | (~w2847 & w7033);
assign w2855 = (~w2847 & w7034) | (~w2847 & w7035) | (w7034 & w7035);
assign w2856 = ~pi0243 & w2853;
assign w2857 = w2847 & w7036;
assign w2858 = pi1151 & w2715;
assign w2859 = (~w2853 & ~w1477) | (~w2853 & w7037) | (~w1477 & w7037);
assign w2860 = ~w2732 & ~w2858;
assign w2861 = w2859 & w2860;
assign w2862 = ~w2857 & ~w2861;
assign w2863 = ~w2855 & w2862;
assign w2864 = (w2709 & ~w2810) | (w2709 & w7038) | (~w2810 & w7038);
assign w2865 = w2737 & ~w2778;
assign w2866 = ~pi0230 & pi0244;
assign w2867 = ~w2864 & ~w2866;
assign w2868 = ~w2865 & w2867;
assign w2869 = (w2737 & ~w2836) | (w2737 & w7039) | (~w2836 & w7039);
assign w2870 = pi1142 & w1477;
assign w2871 = ~w2713 & w2870;
assign w2872 = pi1140 & ~w2717;
assign w2873 = w1480 & w7040;
assign w2874 = ~w2871 & ~w2872;
assign w2875 = (w2709 & ~w2874) | (w2709 & w7041) | (~w2874 & w7041);
assign w2876 = ~pi0230 & pi0245;
assign w2877 = ~w2869 & ~w2876;
assign w2878 = ~w2875 & w2877;
assign w2879 = pi1144 & w1477;
assign w2880 = ~w2713 & w2879;
assign w2881 = pi1142 & ~w2717;
assign w2882 = w1480 & w7042;
assign w2883 = ~w2880 & ~w2881;
assign w2884 = (w2709 & ~w2883) | (w2709 & w7043) | (~w2883 & w7043);
assign w2885 = (w2737 & ~w2874) | (w2737 & w7044) | (~w2874 & w7044);
assign w2886 = ~pi0230 & pi0246;
assign w2887 = ~w2884 & ~w2886;
assign w2888 = ~w2885 & w2887;
assign w2889 = (w2737 & ~w2816) | (w2737 & w7045) | (~w2816 & w7045);
assign w2890 = w2709 & ~w2827;
assign w2891 = ~pi0230 & pi0247;
assign w2892 = ~w2889 & ~w2891;
assign w2893 = ~w2890 & w2892;
assign w2894 = (w2737 & ~w2883) | (w2737 & w7046) | (~w2883 & w7046);
assign w2895 = pi1146 & w1477;
assign w2896 = ~w2713 & w2895;
assign w2897 = pi1144 & ~w2717;
assign w2898 = w1480 & w7047;
assign w2899 = ~w2896 & ~w2897;
assign w2900 = (w2709 & ~w2899) | (w2709 & w7048) | (~w2899 & w7048);
assign w2901 = ~pi0230 & pi0248;
assign w2902 = ~w2894 & ~w2901;
assign w2903 = ~w2900 & w2902;
assign w2904 = (w2737 & ~w2899) | (w2737 & w7049) | (~w2899 & w7049);
assign w2905 = w2709 & ~w2754;
assign w2906 = ~pi0230 & pi0249;
assign w2907 = ~w2904 & ~w2906;
assign w2908 = ~w2905 & w2907;
assign w2909 = ~w309 & w455;
assign w2910 = ~pi0250 & ~w2909;
assign w2911 = ~pi0199 & pi0200;
assign w2912 = ~pi0476 & w2911;
assign w2913 = w2911 & w7050;
assign w2914 = ~pi0199 & ~pi0200;
assign w2915 = pi0897 & w2914;
assign w2916 = w2914 & w7051;
assign w2917 = ~w2912 & ~w2915;
assign w2918 = pi0251 & w2917;
assign w2919 = ~w2913 & ~w2916;
assign w2920 = ~w2918 & w2919;
assign w2921 = w713 & w777;
assign w2922 = (pi1087 & ~w885) | (pi1087 & w7052) | (~w885 & w7052);
assign w2923 = pi0252 & pi1086;
assign w2924 = ~w2922 & w2923;
assign w2925 = ~w2921 & ~w2924;
assign w2926 = w2847 & w7053;
assign w2927 = (~pi0253 & ~w2847) | (~pi0253 & w7054) | (~w2847 & w7054);
assign w2928 = ~w2926 & ~w2927;
assign w2929 = w2853 & ~w2928;
assign w2930 = pi1146 & w1468;
assign w2931 = (~w2853 & ~w2715) | (~w2853 & w7055) | (~w2715 & w7055);
assign w2932 = ~w2822 & ~w2930;
assign w2933 = w2931 & w2932;
assign w2934 = ~w2929 & ~w2933;
assign w2935 = (~pi0254 & ~w2847) | (~pi0254 & w7056) | (~w2847 & w7056);
assign w2936 = (w2853 & ~w2847) | (w2853 & w7058) | (~w2847 & w7058);
assign w2937 = ~w2935 & w2936;
assign w2938 = pi1147 & w1468;
assign w2939 = ~w2731 & ~w2895;
assign w2940 = (~w2853 & ~w2939) | (~w2853 & w7059) | (~w2939 & w7059);
assign w2941 = ~w2937 & ~w2940;
assign w2942 = w2914 & w7060;
assign w2943 = w2911 & w7061;
assign w2944 = pi0255 & w2917;
assign w2945 = ~w2942 & ~w2943;
assign w2946 = ~w2944 & w2945;
assign w2947 = w2914 & w7062;
assign w2948 = w2911 & w7063;
assign w2949 = pi0256 & w2917;
assign w2950 = ~w2947 & ~w2948;
assign w2951 = ~w2949 & w2950;
assign w2952 = w2911 & w7064;
assign w2953 = w2914 & w7065;
assign w2954 = pi0257 & w2917;
assign w2955 = ~w2952 & ~w2953;
assign w2956 = ~w2954 & w2955;
assign w2957 = w2911 & w7066;
assign w2958 = w2914 & w7067;
assign w2959 = pi0258 & w2917;
assign w2960 = ~w2957 & ~w2958;
assign w2961 = ~w2959 & w2960;
assign w2962 = w2911 & w7068;
assign w2963 = w2914 & w7069;
assign w2964 = pi0259 & w2917;
assign w2965 = ~w2962 & ~w2963;
assign w2966 = ~w2964 & w2965;
assign w2967 = w2914 & w7070;
assign w2968 = w2911 & w7071;
assign w2969 = pi0260 & w2917;
assign w2970 = ~w2967 & ~w2968;
assign w2971 = ~w2969 & w2970;
assign w2972 = w2911 & w7072;
assign w2973 = w2914 & w7073;
assign w2974 = pi0261 & w2917;
assign w2975 = ~w2972 & ~w2973;
assign w2976 = ~w2974 & w2975;
assign w2977 = ~pi0228 & pi1087;
assign w2978 = ~pi0123 & pi0228;
assign w2979 = ~w2977 & ~w2978;
assign w2980 = ~pi0262 & w2979;
assign w2981 = pi1136 & ~w2979;
assign w2982 = w1480 & w2981;
assign w2983 = ~w2980 & ~w2982;
assign w2984 = w2847 & w7074;
assign w2985 = (pi0263 & ~w2847) | (pi0263 & w7075) | (~w2847 & w7075);
assign w2986 = w2854 & ~w2985;
assign w2987 = ~w2726 & ~w2749;
assign w2988 = (~w2853 & ~w2987) | (~w2853 & w7076) | (~w2987 & w7076);
assign w2989 = ~w2986 & ~w2988;
assign w2990 = (~w1457 & w7077) | (~w1457 & w7078) | (w7077 & w7078);
assign w2991 = pi0264 & w2990;
assign w2992 = (w1457 & w7079) | (w1457 & w7080) | (w7079 & w7080);
assign w2993 = ~pi0796 & w2992;
assign w2994 = pi1136 & w1468;
assign w2995 = pi1135 & w1477;
assign w2996 = (~w2853 & ~w2715) | (~w2853 & w7081) | (~w2715 & w7081);
assign w2997 = ~w2994 & ~w2995;
assign w2998 = (~w2991 & ~w2997) | (~w2991 & w7082) | (~w2997 & w7082);
assign w2999 = ~w2993 & w2998;
assign w3000 = pi0265 & w2990;
assign w3001 = ~pi0819 & w2992;
assign w3002 = pi1137 & w1468;
assign w3003 = pi1136 & w1477;
assign w3004 = (~w2853 & ~w2715) | (~w2853 & w7083) | (~w2715 & w7083);
assign w3005 = ~w3002 & ~w3003;
assign w3006 = (~w3000 & ~w3005) | (~w3000 & w7084) | (~w3005 & w7084);
assign w3007 = ~w3001 & w3006;
assign w3008 = ~pi0266 & w2990;
assign w3009 = ~pi0948 & w2992;
assign w3010 = pi1128 & w1477;
assign w3011 = pi1129 & w1468;
assign w3012 = (~w2853 & ~w2715) | (~w2853 & w7085) | (~w2715 & w7085);
assign w3013 = ~w3010 & ~w3011;
assign w3014 = (~w3008 & ~w3013) | (~w3008 & w7086) | (~w3013 & w7086);
assign w3015 = ~w3009 & w3014;
assign w3016 = (~pi0267 & ~w2847) | (~pi0267 & w7087) | (~w2847 & w7087);
assign w3017 = w2853 & ~w2984;
assign w3018 = ~w3016 & w3017;
assign w3019 = ~w2723 & ~w2734;
assign w3020 = (~w2853 & ~w3019) | (~w2853 & w7088) | (~w3019 & w7088);
assign w3021 = ~w3018 & ~w3020;
assign w3022 = (~pi0268 & ~w2847) | (~pi0268 & w7089) | (~w2847 & w7089);
assign w3023 = ~w2849 & ~w3022;
assign w3024 = w2853 & ~w3023;
assign w3025 = pi1145 & w1468;
assign w3026 = pi1146 & w2715;
assign w3027 = (~w2853 & ~w1477) | (~w2853 & w7090) | (~w1477 & w7090);
assign w3028 = ~w3025 & ~w3026;
assign w3029 = w3027 & w3028;
assign w3030 = ~w3024 & ~w3029;
assign w3031 = pi0269 & w2990;
assign w3032 = ~pi0817 & w2992;
assign w3033 = pi1130 & w1477;
assign w3034 = pi1131 & w1468;
assign w3035 = (~w2853 & ~w2715) | (~w2853 & w7091) | (~w2715 & w7091);
assign w3036 = ~w3033 & ~w3034;
assign w3037 = (~w3031 & ~w3036) | (~w3031 & w7092) | (~w3036 & w7092);
assign w3038 = ~w3032 & w3037;
assign w3039 = pi0270 & w2990;
assign w3040 = ~pi0805 & w2992;
assign w3041 = pi1134 & w1468;
assign w3042 = pi1133 & w1477;
assign w3043 = (~w2853 & ~w2715) | (~w2853 & w7093) | (~w2715 & w7093);
assign w3044 = ~w3041 & ~w3042;
assign w3045 = (~w3039 & ~w3044) | (~w3039 & w7094) | (~w3044 & w7094);
assign w3046 = ~w3040 & w3045;
assign w3047 = (~pi0271 & ~w2843) | (~pi0271 & w7095) | (~w2843 & w7095);
assign w3048 = ~w2845 & ~w3047;
assign w3049 = w2853 & ~w3048;
assign w3050 = pi1140 & w1468;
assign w3051 = pi1141 & w2715;
assign w3052 = (~w2853 & ~w1477) | (~w2853 & w7096) | (~w1477 & w7096);
assign w3053 = ~w3050 & ~w3051;
assign w3054 = w3052 & w3053;
assign w3055 = ~w3049 & ~w3054;
assign w3056 = (~pi0272 & ~w2843) | (~pi0272 & w7097) | (~w2843 & w7097);
assign w3057 = ~w2847 & ~w3056;
assign w3058 = w2853 & ~w3057;
assign w3059 = pi1144 & w2715;
assign w3060 = pi1143 & w1468;
assign w3061 = (~w2853 & ~w1477) | (~w2853 & w7098) | (~w1477 & w7098);
assign w3062 = ~w3059 & ~w3060;
assign w3063 = w3061 & w3062;
assign w3064 = ~w3058 & ~w3063;
assign w3065 = pi1142 & w2715;
assign w3066 = pi1141 & w1468;
assign w3067 = ~w2832 & ~w3065;
assign w3068 = (~w2853 & ~w3067) | (~w2853 & w7099) | (~w3067 & w7099);
assign w3069 = ~pi0273 & ~w2845;
assign w3070 = (w2853 & ~w2843) | (w2853 & w7100) | (~w2843 & w7100);
assign w3071 = ~w3069 & w3070;
assign w3072 = ~w3068 & ~w3071;
assign w3073 = pi0274 & w2990;
assign w3074 = ~pi0659 & w2992;
assign w3075 = pi1137 & w1477;
assign w3076 = pi1138 & w1468;
assign w3077 = pi1139 & w2715;
assign w3078 = (~w2853 & ~w1477) | (~w2853 & w7081) | (~w1477 & w7081);
assign w3079 = ~w3076 & ~w3077;
assign w3080 = (~w3073 & ~w3079) | (~w3073 & w7101) | (~w3079 & w7101);
assign w3081 = ~w3074 & w3080;
assign w3082 = ~pi0275 & ~w2847;
assign w3083 = ~w2848 & ~w3082;
assign w3084 = w2853 & ~w3083;
assign w3085 = pi1144 & w1468;
assign w3086 = pi1145 & w2715;
assign w3087 = (~w2853 & ~w1477) | (~w2853 & w7102) | (~w1477 & w7102);
assign w3088 = ~w3085 & ~w3086;
assign w3089 = w3087 & w3088;
assign w3090 = ~w3084 & ~w3089;
assign w3091 = (~pi0276 & ~w2843) | (~pi0276 & w7103) | (~w2843 & w7103);
assign w3092 = ~w2844 & ~w3091;
assign w3093 = w2853 & ~w3092;
assign w3094 = pi1140 & w2715;
assign w3095 = pi1139 & w1468;
assign w3096 = (~w2853 & ~w1477) | (~w2853 & w7083) | (~w1477 & w7083);
assign w3097 = ~w3094 & ~w3095;
assign w3098 = w3096 & w3097;
assign w3099 = ~w3093 & ~w3098;
assign w3100 = pi0277 & w2990;
assign w3101 = ~pi0820 & w2992;
assign w3102 = pi1135 & w1468;
assign w3103 = pi1134 & w1477;
assign w3104 = (~w2853 & ~w2715) | (~w2853 & w7104) | (~w2715 & w7104);
assign w3105 = ~w3102 & ~w3103;
assign w3106 = (~w3100 & ~w3105) | (~w3100 & w7105) | (~w3105 & w7105);
assign w3107 = ~w3101 & w3106;
assign w3108 = ~pi0278 & w2990;
assign w3109 = ~pi0976 & w2992;
assign w3110 = pi1126 & w1477;
assign w3111 = pi1128 & w2715;
assign w3112 = (~w2853 & ~w1468) | (~w2853 & w7106) | (~w1468 & w7106);
assign w3113 = ~w3110 & ~w3111;
assign w3114 = (~w3108 & ~w3113) | (~w3108 & w7107) | (~w3113 & w7107);
assign w3115 = ~w3109 & w3114;
assign w3116 = ~pi0279 & w2990;
assign w3117 = ~pi0958 & w2992;
assign w3118 = pi1128 & w1468;
assign w3119 = pi1127 & w1477;
assign w3120 = (~w2853 & ~w2715) | (~w2853 & w7108) | (~w2715 & w7108);
assign w3121 = ~w3118 & ~w3119;
assign w3122 = (~w3116 & ~w3121) | (~w3116 & w7109) | (~w3121 & w7109);
assign w3123 = ~w3117 & w3122;
assign w3124 = pi0280 & w2990;
assign w3125 = ~pi0914 & w2992;
assign w3126 = pi1129 & w1477;
assign w3127 = pi1130 & w1468;
assign w3128 = (~w2853 & ~w2715) | (~w2853 & w7110) | (~w2715 & w7110);
assign w3129 = ~w3126 & ~w3127;
assign w3130 = (~w3124 & ~w3129) | (~w3124 & w7111) | (~w3129 & w7111);
assign w3131 = ~w3125 & w3130;
assign w3132 = pi0281 & w2990;
assign w3133 = ~pi0830 & w2992;
assign w3134 = pi1132 & w1468;
assign w3135 = pi1131 & w1477;
assign w3136 = (~w2853 & ~w2715) | (~w2853 & w7112) | (~w2715 & w7112);
assign w3137 = ~w3134 & ~w3135;
assign w3138 = (~w3132 & ~w3137) | (~w3132 & w7113) | (~w3137 & w7113);
assign w3139 = ~w3133 & w3138;
assign w3140 = pi0282 & w2990;
assign w3141 = ~pi0836 & w2992;
assign w3142 = pi1132 & w1477;
assign w3143 = pi1133 & w1468;
assign w3144 = (~w2853 & ~w2715) | (~w2853 & w7114) | (~w2715 & w7114);
assign w3145 = ~w3142 & ~w3143;
assign w3146 = (~w3140 & ~w3145) | (~w3140 & w7115) | (~w3145 & w7115);
assign w3147 = ~w3141 & w3146;
assign w3148 = (~pi0283 & ~w2843) | (~pi0283 & w7116) | (~w2843 & w7116);
assign w3149 = ~w2846 & ~w3148;
assign w3150 = w2853 & ~w3149;
assign w3151 = pi1142 & w1468;
assign w3152 = pi1143 & w2715;
assign w3153 = (~w2853 & ~w1477) | (~w2853 & w7117) | (~w1477 & w7117);
assign w3154 = ~w3151 & ~w3152;
assign w3155 = w3153 & w3154;
assign w3156 = ~w3150 & ~w3155;
assign w3157 = ~pi0284 & w2979;
assign w3158 = ~w2713 & ~w2979;
assign w3159 = w3075 & w3158;
assign w3160 = ~w3157 & ~w3159;
assign w3161 = w882 & w1442;
assign w3162 = w1442 & w7118;
assign w3163 = w1442 & w7119;
assign w3164 = pi0286 & pi0288;
assign w3165 = ~w882 & ~w1442;
assign w3166 = ~w1442 & w7120;
assign w3167 = ~w1442 & w7121;
assign w3168 = pi0285 & w3167;
assign w3169 = ~pi0285 & ~w3167;
assign w3170 = ~pi0793 & ~w3163;
assign w3171 = ~w3168 & w3170;
assign w3172 = ~w3169 & w3171;
assign w3173 = ~w877 & ~w3164;
assign w3174 = ~w3161 & ~w3165;
assign w3175 = ~pi0286 & w3174;
assign w3176 = w1442 & w7123;
assign w3177 = (~pi0793 & w1442) | (~pi0793 & w7124) | (w1442 & w7124);
assign w3178 = ~w3176 & w3177;
assign w3179 = ~w3175 & w3178;
assign w3180 = ~pi0287 & pi0457;
assign w3181 = ~pi0332 & ~w3180;
assign w3182 = ~pi0288 & w3174;
assign w3183 = (~pi0793 & w3174) | (~pi0793 & w7125) | (w3174 & w7125);
assign w3184 = ~w3182 & w3183;
assign w3185 = ~w3162 & ~w3166;
assign w3186 = pi0289 & ~w3185;
assign w3187 = (~pi0793 & ~w3185) | (~pi0793 & w7126) | (~w3185 & w7126);
assign w3188 = ~w3186 & w3187;
assign w3189 = pi0290 & pi0476;
assign w3190 = ~pi0476 & pi1042;
assign w3191 = ~w3189 & ~w3190;
assign w3192 = pi0291 & pi0476;
assign w3193 = ~pi0476 & pi1043;
assign w3194 = ~w3192 & ~w3193;
assign w3195 = pi0292 & pi0476;
assign w3196 = ~pi0476 & pi1078;
assign w3197 = ~w3195 & ~w3196;
assign w3198 = pi0293 & pi0476;
assign w3199 = ~pi0476 & pi1053;
assign w3200 = ~w3198 & ~w3199;
assign w3201 = pi0294 & pi0476;
assign w3202 = ~pi0476 & pi1066;
assign w3203 = ~w3201 & ~w3202;
assign w3204 = pi0295 & pi0476;
assign w3205 = ~pi0476 & pi1047;
assign w3206 = ~w3204 & ~w3205;
assign w3207 = pi0296 & pi0476;
assign w3208 = ~pi0476 & pi1031;
assign w3209 = ~w3207 & ~w3208;
assign w3210 = pi0297 & pi0476;
assign w3211 = ~pi0476 & pi1038;
assign w3212 = ~w3210 & ~w3211;
assign w3213 = pi0298 & pi0478;
assign w3214 = ~pi0478 & pi1038;
assign w3215 = ~w3213 & ~w3214;
assign w3216 = pi0039 & w1528;
assign w3217 = ~w481 & ~w3216;
assign w3218 = w271 & w7127;
assign w3219 = (~pi0055 & ~w271) | (~pi0055 & w7129) | (~w271 & w7129);
assign w3220 = (pi0300 & ~w271) | (pi0300 & w7130) | (~w271 & w7130);
assign w3221 = w3219 & ~w3220;
assign w3222 = (~w271 & w7131) | (~w271 & w7132) | (w7131 & w7132);
assign w3223 = w271 & w7133;
assign w3224 = ~w3222 & ~w3223;
assign w3225 = w11 & w7134;
assign w3226 = ~w526 & w7135;
assign w3227 = w11 & w7136;
assign w3228 = pi0937 & w526;
assign w3229 = ~w3225 & ~w3227;
assign w3230 = ~w3228 & w3229;
assign w3231 = ~w3226 & w3230;
assign w3232 = pi0303 & pi0478;
assign w3233 = ~pi0478 & pi1043;
assign w3234 = ~w3232 & ~w3233;
assign w3235 = pi0304 & pi0478;
assign w3236 = ~pi0478 & pi1042;
assign w3237 = ~w3235 & ~w3236;
assign w3238 = pi0305 & pi0478;
assign w3239 = ~pi0478 & pi1078;
assign w3240 = ~w3238 & ~w3239;
assign w3241 = pi0306 & pi0478;
assign w3242 = ~pi0478 & pi1053;
assign w3243 = ~w3241 & ~w3242;
assign w3244 = pi0307 & pi0478;
assign w3245 = ~pi0478 & pi1047;
assign w3246 = ~w3244 & ~w3245;
assign w3247 = pi0308 & pi0478;
assign w3248 = ~pi0478 & pi1031;
assign w3249 = ~w3247 & ~w3248;
assign w3250 = pi0309 & pi0478;
assign w3251 = ~pi0478 & pi1066;
assign w3252 = ~w3250 & ~w3251;
assign w3253 = w11 & w7137;
assign w3254 = ~w526 & w7138;
assign w3255 = w11 & w7139;
assign w3256 = pi0934 & w526;
assign w3257 = ~w3253 & ~w3255;
assign w3258 = ~w3256 & w3257;
assign w3259 = ~w3254 & w3258;
assign w3260 = (pi0311 & ~w271) | (pi0311 & w7140) | (~w271 & w7140);
assign w3261 = (~pi0055 & ~w271) | (~pi0055 & w7141) | (~w271 & w7141);
assign w3262 = ~pi0311 & ~w3261;
assign w3263 = ~w3260 & ~w3262;
assign w3264 = ~pi0055 & pi0312;
assign w3265 = (w3264 & ~w271) | (w3264 & w7142) | (~w271 & w7142);
assign w3266 = ~w3218 & ~w3265;
assign w3267 = pi0313 & pi0954;
assign w3268 = w265 & ~w1757;
assign w3269 = ~w144 & ~w3268;
assign w3270 = ~pi0954 & ~w3269;
assign w3271 = ~w3267 & ~w3270;
assign w3272 = w1835 & w1884;
assign w3273 = ~w678 & w3272;
assign w3274 = w1825 & w3273;
assign w3275 = ~pi0340 & ~w1442;
assign w3276 = pi0315 & ~w3275;
assign w3277 = pi1074 & w3275;
assign w3278 = ~w3276 & ~w3277;
assign w3279 = pi0316 & ~w3275;
assign w3280 = pi1041 & w3275;
assign w3281 = ~w3279 & ~w3280;
assign w3282 = ~pi0330 & ~w1442;
assign w3283 = pi0317 & ~w3282;
assign w3284 = pi1072 & w3282;
assign w3285 = ~w3283 & ~w3284;
assign w3286 = ~pi0341 & ~w1442;
assign w3287 = pi0318 & ~w3286;
assign w3288 = pi1068 & w3286;
assign w3289 = ~w3287 & ~w3288;
assign w3290 = pi0319 & ~w3286;
assign w3291 = pi1066 & w3286;
assign w3292 = ~w3290 & ~w3291;
assign w3293 = pi0320 & ~w3275;
assign w3294 = pi1042 & w3275;
assign w3295 = ~w3293 & ~w3294;
assign w3296 = pi0321 & ~w3275;
assign w3297 = pi1052 & w3275;
assign w3298 = ~w3296 & ~w3297;
assign w3299 = pi0322 & ~w3275;
assign w3300 = pi1045 & w3275;
assign w3301 = ~w3299 & ~w3300;
assign w3302 = pi0323 & ~w3275;
assign w3303 = pi1059 & w3275;
assign w3304 = ~w3302 & ~w3303;
assign w3305 = pi0324 & ~w3286;
assign w3306 = pi1080 & w3286;
assign w3307 = ~w3305 & ~w3306;
assign w3308 = pi0325 & ~w3286;
assign w3309 = pi1057 & w3286;
assign w3310 = ~w3308 & ~w3309;
assign w3311 = pi0326 & ~w3286;
assign w3312 = pi1051 & w3286;
assign w3313 = ~w3311 & ~w3312;
assign w3314 = pi0327 & ~w3275;
assign w3315 = pi1034 & w3275;
assign w3316 = ~w3314 & ~w3315;
assign w3317 = pi0328 & ~w3286;
assign w3318 = pi1052 & w3286;
assign w3319 = ~w3317 & ~w3318;
assign w3320 = pi0329 & ~w3286;
assign w3321 = pi1037 & w3286;
assign w3322 = ~w3320 & ~w3321;
assign w3323 = pi1086 & ~w253;
assign w3324 = ~pi0330 & w1442;
assign w3325 = ~w3275 & ~w3324;
assign w3326 = w3323 & ~w3325;
assign w3327 = ~pi0331 & w1442;
assign w3328 = ~w3286 & ~w3327;
assign w3329 = w3323 & ~w3328;
assign w3330 = pi0333 & ~w3286;
assign w3331 = pi1034 & w3286;
assign w3332 = ~w3330 & ~w3331;
assign w3333 = pi0334 & ~w3286;
assign w3334 = pi1059 & w3286;
assign w3335 = ~w3333 & ~w3334;
assign w3336 = pi0335 & ~w3286;
assign w3337 = pi1063 & w3286;
assign w3338 = ~w3336 & ~w3337;
assign w3339 = pi0336 & ~w3282;
assign w3340 = pi1064 & w3282;
assign w3341 = ~w3339 & ~w3340;
assign w3342 = pi0337 & ~w3282;
assign w3343 = pi1038 & w3282;
assign w3344 = ~w3342 & ~w3343;
assign w3345 = pi0338 & ~w3282;
assign w3346 = pi1066 & w3282;
assign w3347 = ~w3345 & ~w3346;
assign w3348 = pi0339 & ~w3282;
assign w3349 = pi1080 & w3282;
assign w3350 = ~w3348 & ~w3349;
assign w3351 = ~pi0331 & ~w1442;
assign w3352 = ~pi0340 & w1442;
assign w3353 = w3323 & ~w3351;
assign w3354 = ~w3352 & w3353;
assign w3355 = ~pi0341 & w1442;
assign w3356 = ~w3282 & ~w3355;
assign w3357 = w3323 & ~w3356;
assign w3358 = pi0342 & ~w3275;
assign w3359 = pi1043 & w3275;
assign w3360 = ~w3358 & ~w3359;
assign w3361 = pi0343 & ~w3275;
assign w3362 = pi1056 & w3275;
assign w3363 = ~w3361 & ~w3362;
assign w3364 = pi0344 & ~w3275;
assign w3365 = pi1063 & w3275;
assign w3366 = ~w3364 & ~w3365;
assign w3367 = pi0345 & ~w3275;
assign w3368 = pi1033 & w3275;
assign w3369 = ~w3367 & ~w3368;
assign w3370 = pi0346 & ~w3275;
assign w3371 = pi1061 & w3275;
assign w3372 = ~w3370 & ~w3371;
assign w3373 = pi0347 & ~w3275;
assign w3374 = pi1049 & w3275;
assign w3375 = ~w3373 & ~w3374;
assign w3376 = pi0348 & ~w3275;
assign w3377 = pi1081 & w3275;
assign w3378 = ~w3376 & ~w3377;
assign w3379 = pi0349 & ~w3275;
assign w3380 = pi1037 & w3275;
assign w3381 = ~w3379 & ~w3380;
assign w3382 = pi0350 & ~w3275;
assign w3383 = pi1029 & w3275;
assign w3384 = ~w3382 & ~w3383;
assign w3385 = pi0351 & ~w3275;
assign w3386 = pi1073 & w3275;
assign w3387 = ~w3385 & ~w3386;
assign w3388 = pi0352 & ~w3275;
assign w3389 = pi1072 & w3275;
assign w3390 = ~w3388 & ~w3389;
assign w3391 = pi0353 & ~w3275;
assign w3392 = pi1057 & w3275;
assign w3393 = ~w3391 & ~w3392;
assign w3394 = pi0354 & ~w3275;
assign w3395 = pi1039 & w3275;
assign w3396 = ~w3394 & ~w3395;
assign w3397 = pi0355 & ~w3275;
assign w3398 = pi1078 & w3275;
assign w3399 = ~w3397 & ~w3398;
assign w3400 = pi0356 & ~w3275;
assign w3401 = pi1075 & w3275;
assign w3402 = ~w3400 & ~w3401;
assign w3403 = pi0357 & ~w3275;
assign w3404 = pi1070 & w3275;
assign w3405 = ~w3403 & ~w3404;
assign w3406 = pi0358 & ~w3275;
assign w3407 = pi1065 & w3275;
assign w3408 = ~w3406 & ~w3407;
assign w3409 = pi0359 & ~w3275;
assign w3410 = pi1062 & w3275;
assign w3411 = ~w3409 & ~w3410;
assign w3412 = pi0360 & ~w3275;
assign w3413 = pi1036 & w3275;
assign w3414 = ~w3412 & ~w3413;
assign w3415 = pi0361 & ~w3275;
assign w3416 = pi1053 & w3275;
assign w3417 = ~w3415 & ~w3416;
assign w3418 = pi0362 & ~w3275;
assign w3419 = pi1064 & w3275;
assign w3420 = ~w3418 & ~w3419;
assign w3421 = pi0363 & ~w3282;
assign w3422 = pi1043 & w3282;
assign w3423 = ~w3421 & ~w3422;
assign w3424 = pi0364 & ~w3282;
assign w3425 = pi1056 & w3282;
assign w3426 = ~w3424 & ~w3425;
assign w3427 = pi0365 & ~w3282;
assign w3428 = pi1059 & w3282;
assign w3429 = ~w3427 & ~w3428;
assign w3430 = pi0366 & ~w3282;
assign w3431 = pi1063 & w3282;
assign w3432 = ~w3430 & ~w3431;
assign w3433 = pi0367 & ~w3282;
assign w3434 = pi1033 & w3282;
assign w3435 = ~w3433 & ~w3434;
assign w3436 = pi0368 & ~w3282;
assign w3437 = pi1061 & w3282;
assign w3438 = ~w3436 & ~w3437;
assign w3439 = pi0369 & ~w3282;
assign w3440 = pi1074 & w3282;
assign w3441 = ~w3439 & ~w3440;
assign w3442 = pi0370 & ~w3282;
assign w3443 = pi1049 & w3282;
assign w3444 = ~w3442 & ~w3443;
assign w3445 = pi0371 & ~w3282;
assign w3446 = pi1045 & w3282;
assign w3447 = ~w3445 & ~w3446;
assign w3448 = pi0372 & ~w3282;
assign w3449 = pi1042 & w3282;
assign w3450 = ~w3448 & ~w3449;
assign w3451 = pi0373 & ~w3282;
assign w3452 = pi1081 & w3282;
assign w3453 = ~w3451 & ~w3452;
assign w3454 = pi0374 & ~w3282;
assign w3455 = pi1029 & w3282;
assign w3456 = ~w3454 & ~w3455;
assign w3457 = pi0375 & ~w3282;
assign w3458 = pi1041 & w3282;
assign w3459 = ~w3457 & ~w3458;
assign w3460 = pi0376 & ~w3282;
assign w3461 = pi1073 & w3282;
assign w3462 = ~w3460 & ~w3461;
assign w3463 = pi0377 & ~w3282;
assign w3464 = pi1068 & w3282;
assign w3465 = ~w3463 & ~w3464;
assign w3466 = pi0378 & ~w3282;
assign w3467 = pi1057 & w3282;
assign w3468 = ~w3466 & ~w3467;
assign w3469 = pi0379 & ~w3282;
assign w3470 = pi1039 & w3282;
assign w3471 = ~w3469 & ~w3470;
assign w3472 = pi0380 & ~w3282;
assign w3473 = pi1078 & w3282;
assign w3474 = ~w3472 & ~w3473;
assign w3475 = pi0381 & ~w3282;
assign w3476 = pi1075 & w3282;
assign w3477 = ~w3475 & ~w3476;
assign w3478 = pi0382 & ~w3282;
assign w3479 = pi1070 & w3282;
assign w3480 = ~w3478 & ~w3479;
assign w3481 = pi0383 & ~w3282;
assign w3482 = pi1065 & w3282;
assign w3483 = ~w3481 & ~w3482;
assign w3484 = pi0384 & ~w3282;
assign w3485 = pi1062 & w3282;
assign w3486 = ~w3484 & ~w3485;
assign w3487 = pi0385 & ~w3282;
assign w3488 = pi1036 & w3282;
assign w3489 = ~w3487 & ~w3488;
assign w3490 = pi0386 & ~w3282;
assign w3491 = pi1053 & w3282;
assign w3492 = ~w3490 & ~w3491;
assign w3493 = pi0387 & ~w3282;
assign w3494 = pi1047 & w3282;
assign w3495 = ~w3493 & ~w3494;
assign w3496 = pi0388 & ~w3282;
assign w3497 = pi1031 & w3282;
assign w3498 = ~w3496 & ~w3497;
assign w3499 = pi0389 & ~w3282;
assign w3500 = pi1030 & w3282;
assign w3501 = ~w3499 & ~w3500;
assign w3502 = pi0390 & ~w3286;
assign w3503 = pi1043 & w3286;
assign w3504 = ~w3502 & ~w3503;
assign w3505 = pi0391 & ~w3286;
assign w3506 = pi1056 & w3286;
assign w3507 = ~w3505 & ~w3506;
assign w3508 = pi0392 & ~w3286;
assign w3509 = pi1033 & w3286;
assign w3510 = ~w3508 & ~w3509;
assign w3511 = pi0393 & ~w3286;
assign w3512 = pi1061 & w3286;
assign w3513 = ~w3511 & ~w3512;
assign w3514 = pi0394 & ~w3286;
assign w3515 = pi1074 & w3286;
assign w3516 = ~w3514 & ~w3515;
assign w3517 = pi0395 & ~w3286;
assign w3518 = pi1049 & w3286;
assign w3519 = ~w3517 & ~w3518;
assign w3520 = pi0396 & ~w3286;
assign w3521 = pi1045 & w3286;
assign w3522 = ~w3520 & ~w3521;
assign w3523 = pi0397 & ~w3286;
assign w3524 = pi1042 & w3286;
assign w3525 = ~w3523 & ~w3524;
assign w3526 = pi0398 & ~w3286;
assign w3527 = pi1081 & w3286;
assign w3528 = ~w3526 & ~w3527;
assign w3529 = pi0399 & ~w3286;
assign w3530 = pi1041 & w3286;
assign w3531 = ~w3529 & ~w3530;
assign w3532 = pi0400 & ~w3286;
assign w3533 = pi1029 & w3286;
assign w3534 = ~w3532 & ~w3533;
assign w3535 = pi0401 & ~w3286;
assign w3536 = pi1073 & w3286;
assign w3537 = ~w3535 & ~w3536;
assign w3538 = pi0402 & ~w3286;
assign w3539 = pi1072 & w3286;
assign w3540 = ~w3538 & ~w3539;
assign w3541 = pi0403 & ~w3286;
assign w3542 = pi1039 & w3286;
assign w3543 = ~w3541 & ~w3542;
assign w3544 = pi0404 & ~w3286;
assign w3545 = pi1078 & w3286;
assign w3546 = ~w3544 & ~w3545;
assign w3547 = pi0405 & ~w3286;
assign w3548 = pi1075 & w3286;
assign w3549 = ~w3547 & ~w3548;
assign w3550 = pi0406 & ~w3286;
assign w3551 = pi1070 & w3286;
assign w3552 = ~w3550 & ~w3551;
assign w3553 = pi0407 & ~w3286;
assign w3554 = pi1065 & w3286;
assign w3555 = ~w3553 & ~w3554;
assign w3556 = pi0408 & ~w3286;
assign w3557 = pi1062 & w3286;
assign w3558 = ~w3556 & ~w3557;
assign w3559 = pi0409 & ~w3286;
assign w3560 = pi1036 & w3286;
assign w3561 = ~w3559 & ~w3560;
assign w3562 = pi0410 & ~w3286;
assign w3563 = pi1053 & w3286;
assign w3564 = ~w3562 & ~w3563;
assign w3565 = pi0411 & ~w3286;
assign w3566 = pi1047 & w3286;
assign w3567 = ~w3565 & ~w3566;
assign w3568 = pi0412 & ~w3286;
assign w3569 = pi1031 & w3286;
assign w3570 = ~w3568 & ~w3569;
assign w3571 = pi0413 & ~w3286;
assign w3572 = pi1030 & w3286;
assign w3573 = ~w3571 & ~w3572;
assign w3574 = pi0414 & ~w3351;
assign w3575 = pi1043 & w3351;
assign w3576 = ~w3574 & ~w3575;
assign w3577 = pi0415 & ~w3351;
assign w3578 = pi1056 & w3351;
assign w3579 = ~w3577 & ~w3578;
assign w3580 = pi0416 & ~w3351;
assign w3581 = pi1063 & w3351;
assign w3582 = ~w3580 & ~w3581;
assign w3583 = pi0417 & ~w3351;
assign w3584 = pi1033 & w3351;
assign w3585 = ~w3583 & ~w3584;
assign w3586 = pi0418 & ~w3351;
assign w3587 = pi1061 & w3351;
assign w3588 = ~w3586 & ~w3587;
assign w3589 = pi0419 & ~w3351;
assign w3590 = pi1074 & w3351;
assign w3591 = ~w3589 & ~w3590;
assign w3592 = pi0420 & ~w3351;
assign w3593 = pi1049 & w3351;
assign w3594 = ~w3592 & ~w3593;
assign w3595 = pi0421 & ~w3351;
assign w3596 = pi1045 & w3351;
assign w3597 = ~w3595 & ~w3596;
assign w3598 = pi0422 & ~w3351;
assign w3599 = pi1042 & w3351;
assign w3600 = ~w3598 & ~w3599;
assign w3601 = pi0423 & ~w3351;
assign w3602 = pi1081 & w3351;
assign w3603 = ~w3601 & ~w3602;
assign w3604 = pi0424 & ~w3351;
assign w3605 = pi1041 & w3351;
assign w3606 = ~w3604 & ~w3605;
assign w3607 = pi0425 & ~w3351;
assign w3608 = pi1029 & w3351;
assign w3609 = ~w3607 & ~w3608;
assign w3610 = pi0426 & ~w3351;
assign w3611 = pi1073 & w3351;
assign w3612 = ~w3610 & ~w3611;
assign w3613 = pi0427 & ~w3351;
assign w3614 = pi1072 & w3351;
assign w3615 = ~w3613 & ~w3614;
assign w3616 = pi0428 & ~w3351;
assign w3617 = pi1039 & w3351;
assign w3618 = ~w3616 & ~w3617;
assign w3619 = pi0429 & ~w3351;
assign w3620 = pi1078 & w3351;
assign w3621 = ~w3619 & ~w3620;
assign w3622 = pi0430 & ~w3351;
assign w3623 = pi1070 & w3351;
assign w3624 = ~w3622 & ~w3623;
assign w3625 = pi0431 & ~w3351;
assign w3626 = pi1065 & w3351;
assign w3627 = ~w3625 & ~w3626;
assign w3628 = pi0432 & ~w3351;
assign w3629 = pi1062 & w3351;
assign w3630 = ~w3628 & ~w3629;
assign w3631 = pi0433 & ~w3351;
assign w3632 = pi1036 & w3351;
assign w3633 = ~w3631 & ~w3632;
assign w3634 = pi0434 & ~w3351;
assign w3635 = pi1053 & w3351;
assign w3636 = ~w3634 & ~w3635;
assign w3637 = pi0435 & ~w3351;
assign w3638 = pi1047 & w3351;
assign w3639 = ~w3637 & ~w3638;
assign w3640 = pi0436 & ~w3351;
assign w3641 = pi1031 & w3351;
assign w3642 = ~w3640 & ~w3641;
assign w3643 = pi0437 & ~w3351;
assign w3644 = pi1064 & w3351;
assign w3645 = ~w3643 & ~w3644;
assign w3646 = pi0438 & ~w3351;
assign w3647 = pi1030 & w3351;
assign w3648 = ~w3646 & ~w3647;
assign w3649 = pi0439 & ~w3282;
assign w3650 = pi1051 & w3282;
assign w3651 = ~w3649 & ~w3650;
assign w3652 = pi0440 & ~w3282;
assign w3653 = pi1037 & w3282;
assign w3654 = ~w3652 & ~w3653;
assign w3655 = pi0441 & ~w3275;
assign w3656 = pi1038 & w3275;
assign w3657 = ~w3655 & ~w3656;
assign w3658 = pi0442 & ~w3282;
assign w3659 = pi1052 & w3282;
assign w3660 = ~w3658 & ~w3659;
assign w3661 = pi0443 & ~w3351;
assign w3662 = pi1038 & w3351;
assign w3663 = ~w3661 & ~w3662;
assign w3664 = pi0444 & ~w3351;
assign w3665 = pi1066 & w3351;
assign w3666 = ~w3664 & ~w3665;
assign w3667 = pi0445 & ~w3351;
assign w3668 = pi1075 & w3351;
assign w3669 = ~w3667 & ~w3668;
assign w3670 = pi0446 & ~w3351;
assign w3671 = pi1080 & w3351;
assign w3672 = ~w3670 & ~w3671;
assign w3673 = pi0447 & ~w3282;
assign w3674 = pi1034 & w3282;
assign w3675 = ~w3673 & ~w3674;
assign w3676 = pi0448 & ~w3351;
assign w3677 = pi1068 & w3351;
assign w3678 = ~w3676 & ~w3677;
assign w3679 = pi0449 & ~w3351;
assign w3680 = pi1051 & w3351;
assign w3681 = ~w3679 & ~w3680;
assign w3682 = pi0450 & ~w3275;
assign w3683 = pi1030 & w3275;
assign w3684 = ~w3682 & ~w3683;
assign w3685 = pi0451 & ~w3351;
assign w3686 = pi1057 & w3351;
assign w3687 = ~w3685 & ~w3686;
assign w3688 = pi0452 & ~w3275;
assign w3689 = pi1047 & w3275;
assign w3690 = ~w3688 & ~w3689;
assign w3691 = pi0453 & ~w3351;
assign w3692 = pi1034 & w3351;
assign w3693 = ~w3691 & ~w3692;
assign w3694 = pi0454 & ~w3351;
assign w3695 = pi1037 & w3351;
assign w3696 = ~w3694 & ~w3695;
assign w3697 = pi0455 & ~w3275;
assign w3698 = pi1031 & w3275;
assign w3699 = ~w3697 & ~w3698;
assign w3700 = pi0456 & ~w3286;
assign w3701 = pi1038 & w3286;
assign w3702 = ~w3700 & ~w3701;
assign w3703 = ~pi0599 & pi0810;
assign w3704 = pi0596 & ~w3703;
assign w3705 = pi0815 & ~w3704;
assign w3706 = ~pi0594 & pi0810;
assign w3707 = pi0600 & ~w3706;
assign w3708 = ~w3705 & w3707;
assign w3709 = pi0804 & ~w3708;
assign w3710 = ~pi0595 & pi0815;
assign w3711 = pi0601 & ~w3710;
assign w3712 = ~pi0804 & ~pi0810;
assign w3713 = ~w3711 & ~w3712;
assign w3714 = pi0594 & pi0597;
assign w3715 = pi0600 & pi0601;
assign w3716 = w3714 & w3715;
assign w3717 = pi0815 & ~w3716;
assign w3718 = pi0605 & pi0821;
assign w3719 = ~w3713 & w3718;
assign w3720 = ~w3717 & w3719;
assign w3721 = ~w3709 & w3720;
assign w3722 = pi0458 & ~w3275;
assign w3723 = pi1066 & w3275;
assign w3724 = ~w3722 & ~w3723;
assign w3725 = pi0459 & ~w3351;
assign w3726 = pi1052 & w3351;
assign w3727 = ~w3725 & ~w3726;
assign w3728 = pi0460 & ~w3275;
assign w3729 = pi1080 & w3275;
assign w3730 = ~w3728 & ~w3729;
assign w3731 = pi0461 & ~w3275;
assign w3732 = pi1051 & w3275;
assign w3733 = ~w3731 & ~w3732;
assign w3734 = pi0462 & ~w3275;
assign w3735 = pi1068 & w3275;
assign w3736 = ~w3734 & ~w3735;
assign w3737 = pi0463 & ~w3286;
assign w3738 = pi1064 & w3286;
assign w3739 = ~w3737 & ~w3738;
assign w3740 = pi0464 & ~w3351;
assign w3741 = pi1059 & w3351;
assign w3742 = ~w3740 & ~w3741;
assign w3743 = ~pi0243 & w522;
assign w3744 = pi1151 & w527;
assign w3745 = pi0926 & w526;
assign w3746 = ~w3743 & ~w3745;
assign w3747 = ~w3744 & w3746;
assign w3748 = pi0275 & w522;
assign w3749 = pi1145 & w527;
assign w3750 = pi0943 & w526;
assign w3751 = ~w3748 & ~w3750;
assign w3752 = ~w3749 & w3751;
assign w3753 = ~pi0979 & ~pi0984;
assign w3754 = pi0040 & ~pi0287;
assign w3755 = pi0995 & w3754;
assign w3756 = w3753 & w3755;
assign w3757 = w264 & w3756;
assign w3758 = ~w341 & ~w3757;
assign w3759 = ~pi0024 & w462;
assign w3760 = pi0468 & ~w3759;
assign w3761 = ~w1550 & ~w3760;
assign w3762 = ~pi0263 & w522;
assign w3763 = pi1150 & w527;
assign w3764 = pi0942 & w526;
assign w3765 = ~w3762 & ~w3764;
assign w3766 = ~w3763 & w3765;
assign w3767 = pi0267 & w522;
assign w3768 = pi1149 & w527;
assign w3769 = pi0925 & w526;
assign w3770 = ~w3767 & ~w3769;
assign w3771 = ~w3768 & w3770;
assign w3772 = pi0253 & w522;
assign w3773 = pi1147 & w527;
assign w3774 = pi0941 & w526;
assign w3775 = ~w3772 & ~w3774;
assign w3776 = ~w3773 & w3775;
assign w3777 = pi0254 & w522;
assign w3778 = pi1148 & w527;
assign w3779 = pi0923 & w526;
assign w3780 = ~w3777 & ~w3779;
assign w3781 = ~w3778 & w3780;
assign w3782 = pi0268 & w522;
assign w3783 = pi1146 & w527;
assign w3784 = pi0922 & w526;
assign w3785 = ~w3782 & ~w3784;
assign w3786 = ~w3783 & w3785;
assign w3787 = pi0272 & w522;
assign w3788 = pi1144 & w527;
assign w3789 = pi0931 & w526;
assign w3790 = ~w3787 & ~w3789;
assign w3791 = ~w3788 & w3790;
assign w3792 = pi0283 & w522;
assign w3793 = pi1143 & w527;
assign w3794 = pi0936 & w526;
assign w3795 = ~w3792 & ~w3794;
assign w3796 = ~w3793 & w3795;
assign w3797 = pi0071 & w1468;
assign w3798 = ~w1675 & ~w3797;
assign w3799 = pi0071 & w1477;
assign w3800 = pi0481 & ~w2533;
assign w3801 = pi0248 & w2533;
assign w3802 = ~w3800 & ~w3801;
assign w3803 = pi0482 & ~w2554;
assign w3804 = pi0249 & w2554;
assign w3805 = ~w3803 & ~w3804;
assign w3806 = pi0483 & ~w2569;
assign w3807 = pi0242 & w2569;
assign w3808 = ~w3806 & ~w3807;
assign w3809 = pi0484 & ~w2569;
assign w3810 = pi0249 & w2569;
assign w3811 = ~w3809 & ~w3810;
assign w3812 = pi0485 & ~w2639;
assign w3813 = pi0234 & w2639;
assign w3814 = ~w3812 & ~w3813;
assign w3815 = pi0486 & ~w2639;
assign w3816 = pi0244 & w2639;
assign w3817 = ~w3815 & ~w3816;
assign w3818 = pi0487 & ~w2533;
assign w3819 = pi0246 & w2533;
assign w3820 = ~w3818 & ~w3819;
assign w3821 = pi0488 & ~w2533;
assign w3822 = ~pi0239 & w2533;
assign w3823 = ~w3821 & ~w3822;
assign w3824 = pi0489 & ~w2639;
assign w3825 = pi0242 & w2639;
assign w3826 = ~w3824 & ~w3825;
assign w3827 = pi0490 & ~w2569;
assign w3828 = pi0241 & w2569;
assign w3829 = ~w3827 & ~w3828;
assign w3830 = pi0491 & ~w2569;
assign w3831 = pi0238 & w2569;
assign w3832 = ~w3830 & ~w3831;
assign w3833 = pi0492 & ~w2569;
assign w3834 = pi0240 & w2569;
assign w3835 = ~w3833 & ~w3834;
assign w3836 = pi0493 & ~w2569;
assign w3837 = pi0244 & w2569;
assign w3838 = ~w3836 & ~w3837;
assign w3839 = pi0494 & ~w2569;
assign w3840 = ~pi0239 & w2569;
assign w3841 = ~w3839 & ~w3840;
assign w3842 = pi0495 & ~w2569;
assign w3843 = pi0235 & w2569;
assign w3844 = ~w3842 & ~w3843;
assign w3845 = pi0496 & ~w2564;
assign w3846 = pi0249 & w2564;
assign w3847 = ~w3845 & ~w3846;
assign w3848 = pi0497 & ~w2564;
assign w3849 = ~pi0239 & w2564;
assign w3850 = ~w3848 & ~w3849;
assign w3851 = pi0498 & ~w2554;
assign w3852 = pi0238 & w2554;
assign w3853 = ~w3851 & ~w3852;
assign w3854 = pi0499 & ~w2564;
assign w3855 = pi0246 & w2564;
assign w3856 = ~w3854 & ~w3855;
assign w3857 = pi0500 & ~w2564;
assign w3858 = pi0241 & w2564;
assign w3859 = ~w3857 & ~w3858;
assign w3860 = pi0501 & ~w2564;
assign w3861 = pi0248 & w2564;
assign w3862 = ~w3860 & ~w3861;
assign w3863 = pi0502 & ~w2564;
assign w3864 = pi0247 & w2564;
assign w3865 = ~w3863 & ~w3864;
assign w3866 = pi0503 & ~w2564;
assign w3867 = pi0245 & w2564;
assign w3868 = ~w3866 & ~w3867;
assign w3869 = pi0504 & ~w2559;
assign w3870 = pi0242 & w2559;
assign w3871 = ~w3869 & ~w3870;
assign w3872 = pi0505 & ~w2564;
assign w3873 = pi0234 & w2564;
assign w3874 = ~w3872 & ~w3873;
assign w3875 = pi0506 & ~w2559;
assign w3876 = pi0241 & w2559;
assign w3877 = ~w3875 & ~w3876;
assign w3878 = pi0507 & ~w2559;
assign w3879 = pi0238 & w2559;
assign w3880 = ~w3878 & ~w3879;
assign w3881 = pi0508 & ~w2559;
assign w3882 = pi0247 & w2559;
assign w3883 = ~w3881 & ~w3882;
assign w3884 = pi0509 & ~w2559;
assign w3885 = pi0245 & w2559;
assign w3886 = ~w3884 & ~w3885;
assign w3887 = pi0510 & ~w2533;
assign w3888 = pi0242 & w2533;
assign w3889 = ~w3887 & ~w3888;
assign w3890 = pi0511 & ~w2533;
assign w3891 = pi0234 & w2533;
assign w3892 = ~w3890 & ~w3891;
assign w3893 = pi0512 & ~w2533;
assign w3894 = pi0235 & w2533;
assign w3895 = ~w3893 & ~w3894;
assign w3896 = pi0513 & ~w2533;
assign w3897 = pi0244 & w2533;
assign w3898 = ~w3896 & ~w3897;
assign w3899 = pi0514 & ~w2533;
assign w3900 = pi0245 & w2533;
assign w3901 = ~w3899 & ~w3900;
assign w3902 = pi0515 & ~w2533;
assign w3903 = pi0240 & w2533;
assign w3904 = ~w3902 & ~w3903;
assign w3905 = pi0516 & ~w2533;
assign w3906 = pi0247 & w2533;
assign w3907 = ~w3905 & ~w3906;
assign w3908 = pi0517 & ~w2533;
assign w3909 = pi0238 & w2533;
assign w3910 = ~w3908 & ~w3909;
assign w3911 = pi0518 & ~w2549;
assign w3912 = pi0234 & w2549;
assign w3913 = ~w3911 & ~w3912;
assign w3914 = pi0519 & ~w2549;
assign w3915 = ~pi0239 & w2549;
assign w3916 = ~w3914 & ~w3915;
assign w3917 = pi0520 & ~w2549;
assign w3918 = pi0246 & w2549;
assign w3919 = ~w3917 & ~w3918;
assign w3920 = pi0521 & ~w2549;
assign w3921 = pi0248 & w2549;
assign w3922 = ~w3920 & ~w3921;
assign w3923 = pi0522 & ~w2549;
assign w3924 = pi0238 & w2549;
assign w3925 = ~w3923 & ~w3924;
assign w3926 = pi0523 & ~w2650;
assign w3927 = pi0234 & w2650;
assign w3928 = ~w3926 & ~w3927;
assign w3929 = pi0524 & ~w2650;
assign w3930 = ~pi0239 & w2650;
assign w3931 = ~w3929 & ~w3930;
assign w3932 = pi0525 & ~w2650;
assign w3933 = pi0245 & w2650;
assign w3934 = ~w3932 & ~w3933;
assign w3935 = pi0526 & ~w2650;
assign w3936 = pi0246 & w2650;
assign w3937 = ~w3935 & ~w3936;
assign w3938 = pi0527 & ~w2650;
assign w3939 = pi0247 & w2650;
assign w3940 = ~w3938 & ~w3939;
assign w3941 = pi0528 & ~w2650;
assign w3942 = pi0249 & w2650;
assign w3943 = ~w3941 & ~w3942;
assign w3944 = pi0529 & ~w2650;
assign w3945 = pi0238 & w2650;
assign w3946 = ~w3944 & ~w3945;
assign w3947 = pi0530 & ~w2650;
assign w3948 = pi0240 & w2650;
assign w3949 = ~w3947 & ~w3948;
assign w3950 = pi0531 & ~w2554;
assign w3951 = pi0235 & w2554;
assign w3952 = ~w3950 & ~w3951;
assign w3953 = pi0532 & ~w2554;
assign w3954 = pi0247 & w2554;
assign w3955 = ~w3953 & ~w3954;
assign w3956 = pi0533 & ~w2559;
assign w3957 = pi0235 & w2559;
assign w3958 = ~w3956 & ~w3957;
assign w3959 = pi0534 & ~w2559;
assign w3960 = ~pi0239 & w2559;
assign w3961 = ~w3959 & ~w3960;
assign w3962 = pi0535 & ~w2559;
assign w3963 = pi0240 & w2559;
assign w3964 = ~w3962 & ~w3963;
assign w3965 = pi0536 & ~w2559;
assign w3966 = pi0246 & w2559;
assign w3967 = ~w3965 & ~w3966;
assign w3968 = pi0537 & ~w2559;
assign w3969 = pi0248 & w2559;
assign w3970 = ~w3968 & ~w3969;
assign w3971 = pi0538 & ~w2559;
assign w3972 = pi0249 & w2559;
assign w3973 = ~w3971 & ~w3972;
assign w3974 = pi0539 & ~w2564;
assign w3975 = pi0242 & w2564;
assign w3976 = ~w3974 & ~w3975;
assign w3977 = pi0540 & ~w2564;
assign w3978 = pi0235 & w2564;
assign w3979 = ~w3977 & ~w3978;
assign w3980 = pi0541 & ~w2564;
assign w3981 = pi0244 & w2564;
assign w3982 = ~w3980 & ~w3981;
assign w3983 = pi0542 & ~w2564;
assign w3984 = pi0240 & w2564;
assign w3985 = ~w3983 & ~w3984;
assign w3986 = pi0543 & ~w2564;
assign w3987 = pi0238 & w2564;
assign w3988 = ~w3986 & ~w3987;
assign w3989 = pi0544 & ~w2569;
assign w3990 = pi0234 & w2569;
assign w3991 = ~w3989 & ~w3990;
assign w3992 = pi0545 & ~w2569;
assign w3993 = pi0245 & w2569;
assign w3994 = ~w3992 & ~w3993;
assign w3995 = pi0546 & ~w2569;
assign w3996 = pi0246 & w2569;
assign w3997 = ~w3995 & ~w3996;
assign w3998 = pi0547 & ~w2569;
assign w3999 = pi0247 & w2569;
assign w4000 = ~w3998 & ~w3999;
assign w4001 = pi0548 & ~w2569;
assign w4002 = pi0248 & w2569;
assign w4003 = ~w4001 & ~w4002;
assign w4004 = pi0549 & ~w2639;
assign w4005 = pi0235 & w2639;
assign w4006 = ~w4004 & ~w4005;
assign w4007 = pi0550 & ~w2639;
assign w4008 = ~pi0239 & w2639;
assign w4009 = ~w4007 & ~w4008;
assign w4010 = pi0551 & ~w2639;
assign w4011 = pi0240 & w2639;
assign w4012 = ~w4010 & ~w4011;
assign w4013 = pi0552 & ~w2639;
assign w4014 = pi0247 & w2639;
assign w4015 = ~w4013 & ~w4014;
assign w4016 = pi0553 & ~w2639;
assign w4017 = pi0241 & w2639;
assign w4018 = ~w4016 & ~w4017;
assign w4019 = pi0554 & ~w2639;
assign w4020 = pi0248 & w2639;
assign w4021 = ~w4019 & ~w4020;
assign w4022 = pi0555 & ~w2639;
assign w4023 = pi0249 & w2639;
assign w4024 = ~w4022 & ~w4023;
assign w4025 = pi0556 & ~w2554;
assign w4026 = pi0242 & w2554;
assign w4027 = ~w4025 & ~w4026;
assign w4028 = pi0557 & ~w2559;
assign w4029 = pi0234 & w2559;
assign w4030 = ~w4028 & ~w4029;
assign w4031 = pi0558 & ~w2559;
assign w4032 = pi0244 & w2559;
assign w4033 = ~w4031 & ~w4032;
assign w4034 = pi0559 & ~w2533;
assign w4035 = pi0241 & w2533;
assign w4036 = ~w4034 & ~w4035;
assign w4037 = pi0560 & ~w2554;
assign w4038 = pi0240 & w2554;
assign w4039 = ~w4037 & ~w4038;
assign w4040 = pi0561 & ~w2549;
assign w4041 = pi0247 & w2549;
assign w4042 = ~w4040 & ~w4041;
assign w4043 = pi0562 & ~w2554;
assign w4044 = pi0241 & w2554;
assign w4045 = ~w4043 & ~w4044;
assign w4046 = pi0563 & ~w2639;
assign w4047 = pi0246 & w2639;
assign w4048 = ~w4046 & ~w4047;
assign w4049 = pi0564 & ~w2554;
assign w4050 = pi0246 & w2554;
assign w4051 = ~w4049 & ~w4050;
assign w4052 = pi0565 & ~w2554;
assign w4053 = pi0248 & w2554;
assign w4054 = ~w4052 & ~w4053;
assign w4055 = pi0566 & ~w2554;
assign w4056 = pi0244 & w2554;
assign w4057 = ~w4055 & ~w4056;
assign w4058 = pi0230 & w1254;
assign w4059 = ~pi0567 & pi1086;
assign w4060 = ~w4058 & w4059;
assign w4061 = pi0621 & w2063;
assign w4062 = pi0665 & w2106;
assign w4063 = ~w4061 & ~w4062;
assign w4064 = pi1085 & w1254;
assign w4065 = pi0230 & w4064;
assign w4066 = ~w4063 & w4065;
assign w4067 = ~w4060 & ~w4066;
assign w4068 = pi0568 & ~w2554;
assign w4069 = pi0245 & w2554;
assign w4070 = ~w4068 & ~w4069;
assign w4071 = pi0569 & ~w2554;
assign w4072 = ~pi0239 & w2554;
assign w4073 = ~w4071 & ~w4072;
assign w4074 = pi0570 & ~w2554;
assign w4075 = pi0234 & w2554;
assign w4076 = ~w4074 & ~w4075;
assign w4077 = pi0571 & ~w2650;
assign w4078 = pi0241 & w2650;
assign w4079 = ~w4077 & ~w4078;
assign w4080 = pi0572 & ~w2650;
assign w4081 = pi0244 & w2650;
assign w4082 = ~w4080 & ~w4081;
assign w4083 = pi0573 & ~w2650;
assign w4084 = pi0242 & w2650;
assign w4085 = ~w4083 & ~w4084;
assign w4086 = pi0574 & ~w2549;
assign w4087 = pi0241 & w2549;
assign w4088 = ~w4086 & ~w4087;
assign w4089 = pi0575 & ~w2650;
assign w4090 = pi0235 & w2650;
assign w4091 = ~w4089 & ~w4090;
assign w4092 = pi0576 & ~w2650;
assign w4093 = pi0248 & w2650;
assign w4094 = ~w4092 & ~w4093;
assign w4095 = pi0577 & ~w2639;
assign w4096 = pi0238 & w2639;
assign w4097 = ~w4095 & ~w4096;
assign w4098 = pi0578 & ~w2549;
assign w4099 = pi0249 & w2549;
assign w4100 = ~w4098 & ~w4099;
assign w4101 = pi0579 & ~w2533;
assign w4102 = pi0249 & w2533;
assign w4103 = ~w4101 & ~w4102;
assign w4104 = pi0580 & ~w2639;
assign w4105 = pi0245 & w2639;
assign w4106 = ~w4104 & ~w4105;
assign w4107 = pi0581 & ~w2549;
assign w4108 = pi0235 & w2549;
assign w4109 = ~w4107 & ~w4108;
assign w4110 = pi0582 & ~w2549;
assign w4111 = pi0240 & w2549;
assign w4112 = ~w4110 & ~w4111;
assign w4113 = pi0584 & ~w2549;
assign w4114 = pi0245 & w2549;
assign w4115 = ~w4113 & ~w4114;
assign w4116 = pi0585 & ~w2549;
assign w4117 = pi0244 & w2549;
assign w4118 = ~w4116 & ~w4117;
assign w4119 = pi0586 & ~w2549;
assign w4120 = pi0242 & w2549;
assign w4121 = ~w4119 & ~w4120;
assign w4122 = pi0230 & ~w2064;
assign w4123 = ~pi0230 & ~pi0587;
assign w4124 = ~w4122 & ~w4123;
assign w4125 = ~pi0123 & w259;
assign w4126 = w3323 & w4125;
assign w4127 = pi0591 & w4126;
assign w4128 = w3323 & ~w4125;
assign w4129 = pi0588 & w4128;
assign w4130 = ~w4127 & ~w4129;
assign w4131 = ~pi0206 & w2568;
assign w4132 = ~pi0205 & w2548;
assign w4133 = ~pi0204 & w2530;
assign w4134 = ~pi0218 & w2553;
assign w4135 = ~w4131 & ~w4132;
assign w4136 = ~w4133 & ~w4134;
assign w4137 = w4135 & w4136;
assign w4138 = ~w710 & ~w4137;
assign w4139 = ~pi0203 & w2553;
assign w4140 = ~pi0201 & w2530;
assign w4141 = ~pi0220 & w2568;
assign w4142 = ~pi0202 & w2548;
assign w4143 = ~w4139 & ~w4140;
assign w4144 = ~w4141 & ~w4142;
assign w4145 = w4143 & w4144;
assign w4146 = ~w702 & ~w4145;
assign w4147 = ~w4138 & ~w4146;
assign w4148 = ~pi0588 & w4126;
assign w4149 = ~pi0590 & w4128;
assign w4150 = ~w4148 & ~w4149;
assign w4151 = pi0592 & w4126;
assign w4152 = pi0591 & w4128;
assign w4153 = ~w4151 & ~w4152;
assign w4154 = pi0590 & w4126;
assign w4155 = pi0592 & w4128;
assign w4156 = ~w4154 & ~w4155;
assign w4157 = ~pi0241 & pi0559;
assign w4158 = ~pi0244 & ~pi0513;
assign w4159 = pi0244 & pi0513;
assign w4160 = ~w4158 & ~w4159;
assign w4161 = pi0241 & ~pi0559;
assign w4162 = pi0235 & ~pi0512;
assign w4163 = pi0239 & pi0488;
assign w4164 = ~pi0245 & pi0514;
assign w4165 = ~pi0235 & pi0512;
assign w4166 = ~pi0246 & pi0487;
assign w4167 = pi0246 & ~pi0487;
assign w4168 = pi0240 & pi0515;
assign w4169 = ~pi0240 & ~pi0515;
assign w4170 = ~w4168 & ~w4169;
assign w4171 = pi0248 & ~pi0481;
assign w4172 = pi0245 & ~pi0514;
assign w4173 = ~pi0242 & pi0510;
assign w4174 = ~pi0247 & pi0516;
assign w4175 = ~pi0239 & ~pi0488;
assign w4176 = pi0238 & ~pi0517;
assign w4177 = pi0247 & ~pi0516;
assign w4178 = pi0234 & pi0511;
assign w4179 = ~pi0234 & ~pi0511;
assign w4180 = ~w4178 & ~w4179;
assign w4181 = pi0242 & ~pi0510;
assign w4182 = ~pi0249 & pi0579;
assign w4183 = pi0249 & ~pi0579;
assign w4184 = ~pi0238 & pi0517;
assign w4185 = ~pi0248 & pi0481;
assign w4186 = w2530 & ~w4157;
assign w4187 = ~w4161 & ~w4162;
assign w4188 = ~w4163 & ~w4164;
assign w4189 = ~w4165 & ~w4166;
assign w4190 = ~w4167 & ~w4171;
assign w4191 = ~w4172 & ~w4173;
assign w4192 = ~w4174 & ~w4175;
assign w4193 = ~w4176 & ~w4177;
assign w4194 = ~w4181 & ~w4182;
assign w4195 = ~w4183 & ~w4184;
assign w4196 = ~w4185 & w4195;
assign w4197 = w4193 & w4194;
assign w4198 = w4191 & w4192;
assign w4199 = w4189 & w4190;
assign w4200 = w4187 & w4188;
assign w4201 = ~w4160 & w4186;
assign w4202 = ~w4170 & ~w4180;
assign w4203 = w4201 & w4202;
assign w4204 = w4199 & w4200;
assign w4205 = w4197 & w4198;
assign w4206 = w4196 & w4205;
assign w4207 = w4203 & w4204;
assign w4208 = w4206 & w4207;
assign w4209 = ~pi0238 & pi0529;
assign w4210 = ~pi0245 & pi0525;
assign w4211 = pi0246 & ~pi0526;
assign w4212 = ~pi0234 & pi0523;
assign w4213 = pi0234 & ~pi0523;
assign w4214 = ~pi0248 & pi0576;
assign w4215 = ~pi0241 & pi0571;
assign w4216 = pi0241 & ~pi0571;
assign w4217 = pi0245 & ~pi0525;
assign w4218 = pi0244 & ~pi0572;
assign w4219 = pi0248 & ~pi0576;
assign w4220 = ~pi0242 & pi0573;
assign w4221 = ~pi0244 & pi0572;
assign w4222 = pi0247 & ~pi0527;
assign w4223 = pi0249 & ~pi0528;
assign w4224 = ~pi0239 & ~pi0524;
assign w4225 = pi0235 & pi0575;
assign w4226 = ~pi0235 & ~pi0575;
assign w4227 = ~w4225 & ~w4226;
assign w4228 = ~pi0247 & pi0527;
assign w4229 = pi0239 & pi0524;
assign w4230 = ~pi0246 & pi0526;
assign w4231 = ~pi0249 & pi0528;
assign w4232 = pi0240 & ~pi0530;
assign w4233 = ~pi0240 & pi0530;
assign w4234 = pi0238 & ~pi0529;
assign w4235 = pi0242 & ~pi0573;
assign w4236 = w2568 & ~w4209;
assign w4237 = ~w4210 & ~w4211;
assign w4238 = ~w4212 & ~w4213;
assign w4239 = ~w4214 & ~w4215;
assign w4240 = ~w4216 & ~w4217;
assign w4241 = ~w4218 & ~w4219;
assign w4242 = ~w4220 & ~w4221;
assign w4243 = ~w4222 & ~w4223;
assign w4244 = ~w4224 & ~w4228;
assign w4245 = ~w4229 & ~w4230;
assign w4246 = ~w4231 & ~w4232;
assign w4247 = ~w4233 & ~w4234;
assign w4248 = ~w4235 & w4247;
assign w4249 = w4245 & w4246;
assign w4250 = w4243 & w4244;
assign w4251 = w4241 & w4242;
assign w4252 = w4239 & w4240;
assign w4253 = w4237 & w4238;
assign w4254 = ~w4227 & w4236;
assign w4255 = w4253 & w4254;
assign w4256 = w4251 & w4252;
assign w4257 = w4249 & w4250;
assign w4258 = w4248 & w4257;
assign w4259 = w4255 & w4256;
assign w4260 = w4258 & w4259;
assign w4261 = ~pi0244 & pi0566;
assign w4262 = pi0246 & ~pi0564;
assign w4263 = ~pi0238 & pi0498;
assign w4264 = ~pi0235 & pi0531;
assign w4265 = pi0249 & ~pi0482;
assign w4266 = ~pi0248 & pi0565;
assign w4267 = pi0245 & ~pi0568;
assign w4268 = ~pi0247 & pi0532;
assign w4269 = pi0238 & ~pi0498;
assign w4270 = pi0235 & ~pi0531;
assign w4271 = pi0240 & ~pi0560;
assign w4272 = ~pi0239 & pi0569;
assign w4273 = pi0239 & ~pi0569;
assign w4274 = ~w4272 & ~w4273;
assign w4275 = pi0234 & ~pi0570;
assign w4276 = pi0242 & ~pi0556;
assign w4277 = ~pi0245 & pi0568;
assign w4278 = pi0241 & ~pi0562;
assign w4279 = ~pi0242 & pi0556;
assign w4280 = ~pi0240 & pi0560;
assign w4281 = ~pi0234 & pi0570;
assign w4282 = ~pi0241 & pi0562;
assign w4283 = pi0247 & ~pi0532;
assign w4284 = pi0244 & ~pi0566;
assign w4285 = ~pi0249 & pi0482;
assign w4286 = ~pi0246 & pi0564;
assign w4287 = pi0248 & ~pi0565;
assign w4288 = w2553 & ~w4261;
assign w4289 = ~w4262 & ~w4263;
assign w4290 = ~w4264 & ~w4265;
assign w4291 = ~w4266 & ~w4267;
assign w4292 = ~w4268 & ~w4269;
assign w4293 = ~w4270 & ~w4271;
assign w4294 = ~w4275 & ~w4276;
assign w4295 = ~w4277 & ~w4278;
assign w4296 = ~w4279 & ~w4280;
assign w4297 = ~w4281 & ~w4282;
assign w4298 = ~w4283 & ~w4284;
assign w4299 = ~w4285 & ~w4286;
assign w4300 = ~w4287 & w4299;
assign w4301 = w4297 & w4298;
assign w4302 = w4295 & w4296;
assign w4303 = w4293 & w4294;
assign w4304 = w4291 & w4292;
assign w4305 = w4289 & w4290;
assign w4306 = ~w4274 & w4288;
assign w4307 = w4305 & w4306;
assign w4308 = w4303 & w4304;
assign w4309 = w4301 & w4302;
assign w4310 = w4300 & w4309;
assign w4311 = w4307 & w4308;
assign w4312 = w4310 & w4311;
assign w4313 = pi0248 & ~pi0521;
assign w4314 = ~pi0242 & pi0586;
assign w4315 = ~pi0248 & pi0521;
assign w4316 = pi0245 & ~pi0584;
assign w4317 = ~pi0249 & pi0578;
assign w4318 = ~pi0234 & pi0518;
assign w4319 = ~pi0247 & pi0561;
assign w4320 = ~pi0239 & ~pi0519;
assign w4321 = pi0247 & ~pi0561;
assign w4322 = pi0244 & ~pi0585;
assign w4323 = pi0238 & ~pi0522;
assign w4324 = ~pi0245 & pi0584;
assign w4325 = pi0246 & pi0520;
assign w4326 = ~pi0246 & ~pi0520;
assign w4327 = ~w4325 & ~w4326;
assign w4328 = ~pi0240 & pi0582;
assign w4329 = pi0235 & ~pi0581;
assign w4330 = ~pi0238 & pi0522;
assign w4331 = ~pi0235 & pi0581;
assign w4332 = ~pi0244 & pi0585;
assign w4333 = pi0241 & ~pi0574;
assign w4334 = pi0239 & pi0519;
assign w4335 = pi0242 & ~pi0586;
assign w4336 = ~pi0241 & pi0574;
assign w4337 = pi0249 & ~pi0578;
assign w4338 = pi0234 & ~pi0518;
assign w4339 = pi0240 & ~pi0582;
assign w4340 = w2548 & ~w4313;
assign w4341 = ~w4314 & ~w4315;
assign w4342 = ~w4316 & ~w4317;
assign w4343 = ~w4318 & ~w4319;
assign w4344 = ~w4320 & ~w4321;
assign w4345 = ~w4322 & ~w4323;
assign w4346 = ~w4324 & ~w4328;
assign w4347 = ~w4329 & ~w4330;
assign w4348 = ~w4331 & ~w4332;
assign w4349 = ~w4333 & ~w4334;
assign w4350 = ~w4335 & ~w4336;
assign w4351 = ~w4337 & ~w4338;
assign w4352 = ~w4339 & w4351;
assign w4353 = w4349 & w4350;
assign w4354 = w4347 & w4348;
assign w4355 = w4345 & w4346;
assign w4356 = w4343 & w4344;
assign w4357 = w4341 & w4342;
assign w4358 = ~w4327 & w4340;
assign w4359 = w4357 & w4358;
assign w4360 = w4355 & w4356;
assign w4361 = w4353 & w4354;
assign w4362 = w4352 & w4361;
assign w4363 = w4359 & w4360;
assign w4364 = w4362 & w4363;
assign w4365 = ~w4208 & ~w4260;
assign w4366 = ~w4312 & ~w4364;
assign w4367 = w4365 & w4366;
assign w4368 = ~w702 & ~w4367;
assign w4369 = ~pi0240 & pi0551;
assign w4370 = pi0239 & pi0550;
assign w4371 = ~pi0242 & pi0489;
assign w4372 = pi0241 & ~pi0553;
assign w4373 = pi0235 & ~pi0549;
assign w4374 = pi0248 & ~pi0554;
assign w4375 = ~pi0246 & pi0563;
assign w4376 = pi0240 & ~pi0551;
assign w4377 = pi0234 & ~pi0485;
assign w4378 = pi0245 & ~pi0580;
assign w4379 = ~pi0235 & pi0549;
assign w4380 = pi0246 & ~pi0563;
assign w4381 = pi0247 & pi0552;
assign w4382 = ~pi0247 & ~pi0552;
assign w4383 = ~w4381 & ~w4382;
assign w4384 = pi0238 & ~pi0577;
assign w4385 = ~pi0238 & pi0577;
assign w4386 = pi0249 & ~pi0555;
assign w4387 = ~pi0244 & pi0486;
assign w4388 = ~pi0245 & pi0580;
assign w4389 = ~pi0234 & pi0485;
assign w4390 = pi0242 & ~pi0489;
assign w4391 = ~pi0249 & pi0555;
assign w4392 = ~pi0239 & ~pi0550;
assign w4393 = ~pi0241 & pi0553;
assign w4394 = pi0244 & ~pi0486;
assign w4395 = ~pi0248 & pi0554;
assign w4396 = w2553 & ~w4369;
assign w4397 = ~w4370 & ~w4371;
assign w4398 = ~w4372 & ~w4373;
assign w4399 = ~w4374 & ~w4375;
assign w4400 = ~w4376 & ~w4377;
assign w4401 = ~w4378 & ~w4379;
assign w4402 = ~w4380 & ~w4384;
assign w4403 = ~w4385 & ~w4386;
assign w4404 = ~w4387 & ~w4388;
assign w4405 = ~w4389 & ~w4390;
assign w4406 = ~w4391 & ~w4392;
assign w4407 = ~w4393 & ~w4394;
assign w4408 = ~w4395 & w4407;
assign w4409 = w4405 & w4406;
assign w4410 = w4403 & w4404;
assign w4411 = w4401 & w4402;
assign w4412 = w4399 & w4400;
assign w4413 = w4397 & w4398;
assign w4414 = ~w4383 & w4396;
assign w4415 = w4413 & w4414;
assign w4416 = w4411 & w4412;
assign w4417 = w4409 & w4410;
assign w4418 = w4408 & w4417;
assign w4419 = w4415 & w4416;
assign w4420 = w4418 & w4419;
assign w4421 = ~pi0234 & ~pi0505;
assign w4422 = pi0234 & pi0505;
assign w4423 = ~w4421 & ~w4422;
assign w4424 = pi0245 & ~pi0503;
assign w4425 = pi0235 & ~pi0540;
assign w4426 = pi0242 & ~pi0539;
assign w4427 = ~pi0238 & pi0543;
assign w4428 = ~pi0239 & ~pi0497;
assign w4429 = pi0238 & ~pi0543;
assign w4430 = ~pi0242 & pi0539;
assign w4431 = pi0249 & ~pi0496;
assign w4432 = pi0239 & pi0497;
assign w4433 = ~pi0245 & pi0503;
assign w4434 = pi0241 & ~pi0500;
assign w4435 = ~pi0235 & pi0540;
assign w4436 = ~pi0248 & pi0501;
assign w4437 = ~pi0249 & pi0496;
assign w4438 = pi0248 & ~pi0501;
assign w4439 = pi0240 & pi0542;
assign w4440 = ~pi0240 & ~pi0542;
assign w4441 = ~w4439 & ~w4440;
assign w4442 = pi0244 & ~pi0541;
assign w4443 = ~pi0247 & pi0502;
assign w4444 = pi0247 & ~pi0502;
assign w4445 = ~pi0241 & pi0500;
assign w4446 = ~pi0244 & pi0541;
assign w4447 = pi0246 & ~pi0499;
assign w4448 = ~pi0246 & pi0499;
assign w4449 = w2548 & ~w4424;
assign w4450 = ~w4425 & ~w4426;
assign w4451 = ~w4427 & ~w4428;
assign w4452 = ~w4429 & ~w4430;
assign w4453 = ~w4431 & ~w4432;
assign w4454 = ~w4433 & ~w4434;
assign w4455 = ~w4435 & ~w4436;
assign w4456 = ~w4437 & ~w4438;
assign w4457 = ~w4442 & ~w4443;
assign w4458 = ~w4444 & ~w4445;
assign w4459 = ~w4446 & ~w4447;
assign w4460 = ~w4448 & w4459;
assign w4461 = w4457 & w4458;
assign w4462 = w4455 & w4456;
assign w4463 = w4453 & w4454;
assign w4464 = w4451 & w4452;
assign w4465 = w4449 & w4450;
assign w4466 = ~w4423 & ~w4441;
assign w4467 = w4465 & w4466;
assign w4468 = w4463 & w4464;
assign w4469 = w4461 & w4462;
assign w4470 = w4460 & w4469;
assign w4471 = w4467 & w4468;
assign w4472 = w4470 & w4471;
assign w4473 = pi0245 & ~pi0509;
assign w4474 = pi0242 & ~pi0504;
assign w4475 = ~pi0248 & pi0537;
assign w4476 = pi0239 & pi0534;
assign w4477 = ~pi0239 & ~pi0534;
assign w4478 = pi0235 & ~pi0533;
assign w4479 = pi0234 & ~pi0557;
assign w4480 = ~pi0249 & pi0538;
assign w4481 = pi0246 & ~pi0536;
assign w4482 = ~pi0238 & pi0507;
assign w4483 = ~pi0245 & pi0509;
assign w4484 = pi0244 & ~pi0558;
assign w4485 = pi0247 & pi0508;
assign w4486 = ~pi0247 & ~pi0508;
assign w4487 = ~w4485 & ~w4486;
assign w4488 = pi0241 & ~pi0506;
assign w4489 = pi0240 & ~pi0535;
assign w4490 = pi0248 & ~pi0537;
assign w4491 = ~pi0235 & pi0533;
assign w4492 = ~pi0240 & pi0535;
assign w4493 = pi0238 & ~pi0507;
assign w4494 = ~pi0246 & pi0536;
assign w4495 = ~pi0244 & pi0558;
assign w4496 = ~pi0242 & pi0504;
assign w4497 = pi0249 & ~pi0538;
assign w4498 = ~pi0234 & pi0557;
assign w4499 = ~pi0241 & pi0506;
assign w4500 = w2530 & ~w4473;
assign w4501 = ~w4474 & ~w4475;
assign w4502 = ~w4476 & ~w4477;
assign w4503 = ~w4478 & ~w4479;
assign w4504 = ~w4480 & ~w4481;
assign w4505 = ~w4482 & ~w4483;
assign w4506 = ~w4484 & ~w4488;
assign w4507 = ~w4489 & ~w4490;
assign w4508 = ~w4491 & ~w4492;
assign w4509 = ~w4493 & ~w4494;
assign w4510 = ~w4495 & ~w4496;
assign w4511 = ~w4497 & ~w4498;
assign w4512 = ~w4499 & w4511;
assign w4513 = w4509 & w4510;
assign w4514 = w4507 & w4508;
assign w4515 = w4505 & w4506;
assign w4516 = w4503 & w4504;
assign w4517 = w4501 & w4502;
assign w4518 = ~w4487 & w4500;
assign w4519 = w4517 & w4518;
assign w4520 = w4515 & w4516;
assign w4521 = w4513 & w4514;
assign w4522 = w4512 & w4521;
assign w4523 = w4519 & w4520;
assign w4524 = w4522 & w4523;
assign w4525 = ~pi0234 & pi0544;
assign w4526 = ~pi0245 & pi0545;
assign w4527 = ~pi0246 & pi0546;
assign w4528 = pi0247 & ~pi0547;
assign w4529 = pi0246 & ~pi0546;
assign w4530 = pi0242 & pi0483;
assign w4531 = ~pi0242 & ~pi0483;
assign w4532 = ~w4530 & ~w4531;
assign w4533 = ~pi0235 & pi0495;
assign w4534 = ~pi0238 & pi0491;
assign w4535 = pi0241 & ~pi0490;
assign w4536 = ~pi0247 & pi0547;
assign w4537 = pi0235 & ~pi0495;
assign w4538 = pi0238 & ~pi0491;
assign w4539 = ~pi0240 & pi0492;
assign w4540 = pi0234 & ~pi0544;
assign w4541 = ~pi0239 & ~pi0494;
assign w4542 = pi0239 & pi0494;
assign w4543 = pi0245 & ~pi0545;
assign w4544 = ~pi0241 & pi0490;
assign w4545 = pi0244 & ~pi0493;
assign w4546 = ~pi0244 & pi0493;
assign w4547 = pi0240 & ~pi0492;
assign w4548 = ~pi0249 & pi0484;
assign w4549 = pi0249 & ~pi0484;
assign w4550 = pi0248 & ~pi0548;
assign w4551 = ~pi0248 & pi0548;
assign w4552 = w2568 & ~w4525;
assign w4553 = ~w4526 & ~w4527;
assign w4554 = ~w4528 & ~w4529;
assign w4555 = ~w4533 & ~w4534;
assign w4556 = ~w4535 & ~w4536;
assign w4557 = ~w4537 & ~w4538;
assign w4558 = ~w4539 & ~w4540;
assign w4559 = ~w4541 & ~w4542;
assign w4560 = ~w4543 & ~w4544;
assign w4561 = ~w4545 & ~w4546;
assign w4562 = ~w4547 & ~w4548;
assign w4563 = ~w4549 & ~w4550;
assign w4564 = ~w4551 & w4563;
assign w4565 = w4561 & w4562;
assign w4566 = w4559 & w4560;
assign w4567 = w4557 & w4558;
assign w4568 = w4555 & w4556;
assign w4569 = w4553 & w4554;
assign w4570 = ~w4532 & w4552;
assign w4571 = w4569 & w4570;
assign w4572 = w4567 & w4568;
assign w4573 = w4565 & w4566;
assign w4574 = w4564 & w4573;
assign w4575 = w4571 & w4572;
assign w4576 = w4574 & w4575;
assign w4577 = ~w4420 & ~w4472;
assign w4578 = ~w4524 & ~w4576;
assign w4579 = w4577 & w4578;
assign w4580 = ~w710 & ~w4579;
assign w4581 = ~w4368 & ~w4580;
assign w4582 = pi0605 & ~pi0806;
assign w4583 = pi0601 & w4582;
assign w4584 = pi0600 & w4583;
assign w4585 = ~pi0594 & ~w4584;
assign w4586 = pi0594 & w4584;
assign w4587 = ~pi0332 & ~w4585;
assign w4588 = ~w4586 & w4587;
assign w4589 = w3716 & w4582;
assign w4590 = ~pi0595 & ~w4589;
assign w4591 = pi0595 & w4589;
assign w4592 = ~pi0332 & ~w4590;
assign w4593 = ~w4591 & w4592;
assign w4594 = ~pi0596 & ~w4591;
assign w4595 = pi0596 & w4591;
assign w4596 = ~pi0332 & ~w4594;
assign w4597 = ~w4595 & w4596;
assign w4598 = ~pi0597 & ~w4586;
assign w4599 = ~pi0332 & ~w4589;
assign w4600 = ~w4598 & w4599;
assign w4601 = ~pi0059 & w2;
assign w4602 = ~pi0882 & w4601;
assign w4603 = pi0947 & w4602;
assign w4604 = pi0598 & ~w4603;
assign w4605 = pi0740 & pi0780;
assign w4606 = w700 & w4605;
assign w4607 = ~w4604 & ~w4606;
assign w4608 = ~pi0599 & ~w4595;
assign w4609 = pi0599 & w4595;
assign w4610 = ~pi0332 & ~w4608;
assign w4611 = ~w4609 & w4610;
assign w4612 = ~pi0600 & ~w4583;
assign w4613 = ~pi0332 & ~w4584;
assign w4614 = ~w4612 & w4613;
assign w4615 = ~pi0601 & ~w4582;
assign w4616 = ~pi0332 & ~w4583;
assign w4617 = ~w4615 & w4616;
assign w4618 = pi0230 & ~w2107;
assign w4619 = ~pi0230 & ~pi0602;
assign w4620 = ~w4618 & ~w4619;
assign w4621 = pi0832 & ~pi0980;
assign w4622 = pi1032 & pi1054;
assign w4623 = ~pi1055 & w4622;
assign w4624 = w4621 & w4623;
assign w4625 = pi0952 & w4624;
assign w4626 = ~pi0966 & ~w4625;
assign w4627 = pi0603 & w4626;
assign w4628 = pi0872 & pi0966;
assign w4629 = ~pi0966 & w4625;
assign w4630 = pi1094 & w4629;
assign w4631 = pi0871 & pi0966;
assign w4632 = ~w4628 & ~w4631;
assign w4633 = ~w4627 & w4632;
assign w4634 = ~w4630 & w4633;
assign w4635 = pi0823 & w707;
assign w4636 = ~pi0779 & w4635;
assign w4637 = ~pi0299 & pi0983;
assign w4638 = pi0907 & w4637;
assign w4639 = pi0604 & ~w4638;
assign w4640 = ~w4635 & w4639;
assign w4641 = ~w4636 & ~w4640;
assign w4642 = ~pi0605 & pi0806;
assign w4643 = ~pi0332 & ~w4582;
assign w4644 = ~w4642 & w4643;
assign w4645 = pi1098 & w4629;
assign w4646 = pi0606 & w4626;
assign w4647 = pi0837 & pi0966;
assign w4648 = ~w4645 & ~w4647;
assign w4649 = ~w4646 & w4648;
assign w4650 = pi0607 & w4626;
assign w4651 = pi1101 & w4629;
assign w4652 = ~w4650 & ~w4651;
assign w4653 = pi0608 & w4626;
assign w4654 = pi1110 & w4629;
assign w4655 = ~w4653 & ~w4654;
assign w4656 = pi0609 & w4626;
assign w4657 = pi1112 & w4629;
assign w4658 = ~w4656 & ~w4657;
assign w4659 = pi0610 & w4626;
assign w4660 = pi1107 & w4629;
assign w4661 = ~w4659 & ~w4660;
assign w4662 = pi0611 & w4626;
assign w4663 = pi1108 & w4629;
assign w4664 = ~w4662 & ~w4663;
assign w4665 = pi0612 & w4626;
assign w4666 = pi1105 & w4629;
assign w4667 = ~w4665 & ~w4666;
assign w4668 = pi0613 & w4626;
assign w4669 = pi1109 & w4629;
assign w4670 = ~w4668 & ~w4669;
assign w4671 = pi1096 & w4629;
assign w4672 = pi0614 & w4626;
assign w4673 = ~w4631 & ~w4671;
assign w4674 = ~w4672 & w4673;
assign w4675 = pi0907 & w4602;
assign w4676 = ~pi0615 & ~w4675;
assign w4677 = pi0779 & pi0797;
assign w4678 = w708 & w4677;
assign w4679 = ~w4676 & ~w4678;
assign w4680 = pi1095 & w4629;
assign w4681 = pi0616 & w4626;
assign w4682 = ~w4628 & ~w4680;
assign w4683 = ~w4681 & w4682;
assign w4684 = pi1099 & w4629;
assign w4685 = pi0617 & w4626;
assign w4686 = pi0850 & pi0966;
assign w4687 = ~w4684 & ~w4686;
assign w4688 = ~w4685 & w4687;
assign w4689 = pi0618 & w4626;
assign w4690 = pi1111 & w4629;
assign w4691 = ~w4689 & ~w4690;
assign w4692 = pi0619 & w4626;
assign w4693 = pi1116 & w4629;
assign w4694 = ~w4692 & ~w4693;
assign w4695 = pi0620 & w4626;
assign w4696 = pi1106 & w4629;
assign w4697 = ~w4695 & ~w4696;
assign w4698 = pi0621 & w4626;
assign w4699 = pi1102 & w4629;
assign w4700 = ~w4698 & ~w4699;
assign w4701 = pi0622 & w4626;
assign w4702 = pi1103 & w4629;
assign w4703 = ~w4701 & ~w4702;
assign w4704 = pi0623 & w4626;
assign w4705 = pi1100 & w4629;
assign w4706 = ~w4704 & ~w4705;
assign w4707 = pi0831 & w699;
assign w4708 = ~pi0780 & w4707;
assign w4709 = pi0947 & w4637;
assign w4710 = pi0624 & ~w4709;
assign w4711 = ~w4707 & w4710;
assign w4712 = ~w4708 & ~w4711;
assign w4713 = pi0832 & ~pi0973;
assign w4714 = ~pi1048 & pi1060;
assign w4715 = pi1082 & w4714;
assign w4716 = w4713 & w4715;
assign w4717 = ~pi0953 & w4716;
assign w4718 = ~pi0962 & w4717;
assign w4719 = pi1110 & w4718;
assign w4720 = ~pi0962 & ~w4717;
assign w4721 = pi0625 & w4720;
assign w4722 = ~w4719 & ~w4721;
assign w4723 = pi0626 & w4626;
assign w4724 = pi1115 & w4629;
assign w4725 = ~w4723 & ~w4724;
assign w4726 = pi1111 & w4718;
assign w4727 = pi0627 & w4720;
assign w4728 = ~w4726 & ~w4727;
assign w4729 = pi1113 & w4718;
assign w4730 = pi0628 & w4720;
assign w4731 = ~w4729 & ~w4730;
assign w4732 = pi0629 & w4626;
assign w4733 = pi1113 & w4629;
assign w4734 = ~w4732 & ~w4733;
assign w4735 = pi0630 & w4626;
assign w4736 = pi1114 & w4629;
assign w4737 = ~w4735 & ~w4736;
assign w4738 = pi1107 & w4718;
assign w4739 = ~pi0631 & w4720;
assign w4740 = ~w4738 & ~w4739;
assign w4741 = pi1109 & w4718;
assign w4742 = ~pi0632 & w4720;
assign w4743 = ~w4741 & ~w4742;
assign w4744 = pi0633 & w4626;
assign w4745 = pi1104 & w4629;
assign w4746 = ~w4744 & ~w4745;
assign w4747 = pi1104 & w4718;
assign w4748 = pi0634 & w4720;
assign w4749 = ~w4747 & ~w4748;
assign w4750 = pi1106 & w4718;
assign w4751 = ~pi0635 & w4720;
assign w4752 = ~w4750 & ~w4751;
assign w4753 = pi0636 & w4626;
assign w4754 = pi1121 & w4629;
assign w4755 = ~w4753 & ~w4754;
assign w4756 = pi1099 & w4718;
assign w4757 = pi0637 & w4720;
assign w4758 = ~w4756 & ~w4757;
assign w4759 = pi1101 & w4718;
assign w4760 = pi0638 & w4720;
assign w4761 = ~w4759 & ~w4760;
assign w4762 = pi1103 & w4718;
assign w4763 = pi0639 & w4720;
assign w4764 = ~w4762 & ~w4763;
assign w4765 = pi0640 & w4626;
assign w4766 = pi1122 & w4629;
assign w4767 = ~w4765 & ~w4766;
assign w4768 = pi1115 & w4718;
assign w4769 = pi0641 & w4720;
assign w4770 = ~w4768 & ~w4769;
assign w4771 = pi0642 & w4626;
assign w4772 = pi1097 & w4629;
assign w4773 = ~w4771 & ~w4772;
assign w4774 = pi1098 & w4718;
assign w4775 = pi0643 & w4720;
assign w4776 = ~w4774 & ~w4775;
assign w4777 = pi0644 & w4626;
assign w4778 = pi1117 & w4629;
assign w4779 = ~w4777 & ~w4778;
assign w4780 = pi0645 & w4626;
assign w4781 = pi1119 & w4629;
assign w4782 = ~w4780 & ~w4781;
assign w4783 = pi1108 & w4718;
assign w4784 = ~pi0646 & w4720;
assign w4785 = ~w4783 & ~w4784;
assign w4786 = pi1114 & w4718;
assign w4787 = pi0647 & w4720;
assign w4788 = ~w4786 & ~w4787;
assign w4789 = pi1116 & w4718;
assign w4790 = pi0648 & w4720;
assign w4791 = ~w4789 & ~w4790;
assign w4792 = pi1120 & w4718;
assign w4793 = ~pi0649 & w4720;
assign w4794 = ~w4792 & ~w4793;
assign w4795 = pi1121 & w4718;
assign w4796 = ~pi0650 & w4720;
assign w4797 = ~w4795 & ~w4796;
assign w4798 = pi0651 & w4626;
assign w4799 = pi1124 & w4629;
assign w4800 = ~w4798 & ~w4799;
assign w4801 = pi0652 & w4626;
assign w4802 = pi1125 & w4629;
assign w4803 = ~w4801 & ~w4802;
assign w4804 = pi0653 & w4626;
assign w4805 = pi1123 & w4629;
assign w4806 = ~w4804 & ~w4805;
assign w4807 = pi1124 & w4718;
assign w4808 = ~pi0654 & w4720;
assign w4809 = ~w4807 & ~w4808;
assign w4810 = pi1118 & w4718;
assign w4811 = ~pi0655 & w4720;
assign w4812 = ~w4810 & ~w4811;
assign w4813 = pi0656 & w4626;
assign w4814 = pi1120 & w4629;
assign w4815 = ~w4813 & ~w4814;
assign w4816 = pi1125 & w4718;
assign w4817 = ~pi0657 & w4720;
assign w4818 = ~w4816 & ~w4817;
assign w4819 = pi0658 & w4626;
assign w4820 = pi1118 & w4629;
assign w4821 = ~w4819 & ~w4820;
assign w4822 = pi0278 & pi0279;
assign w4823 = pi0266 & w4822;
assign w4824 = ~pi0280 & w4823;
assign w4825 = ~pi0269 & w4824;
assign w4826 = ~pi0281 & w4825;
assign w4827 = ~pi0282 & w4826;
assign w4828 = ~pi0270 & w4827;
assign w4829 = ~pi0277 & w4828;
assign w4830 = ~pi0264 & w4829;
assign w4831 = ~pi0265 & w4830;
assign w4832 = pi0274 & ~w4831;
assign w4833 = ~pi0274 & w4831;
assign w4834 = ~w4832 & ~w4833;
assign w4835 = pi1112 & w4718;
assign w4836 = pi0660 & w4720;
assign w4837 = ~w4835 & ~w4836;
assign w4838 = pi1095 & w4718;
assign w4839 = pi0661 & w4720;
assign w4840 = ~w4838 & ~w4839;
assign w4841 = pi1096 & w4718;
assign w4842 = pi0662 & w4720;
assign w4843 = ~w4841 & ~w4842;
assign w4844 = ~pi1128 & ~pi1130;
assign w4845 = ~pi1131 & ~pi1132;
assign w4846 = ~w886 & w4845;
assign w4847 = pi1129 & w4846;
assign w4848 = w4844 & w4847;
assign w4849 = pi0784 & w4848;
assign w4850 = ~pi1129 & w4846;
assign w4851 = pi1128 & ~pi1130;
assign w4852 = w4850 & w4851;
assign w4853 = pi0855 & w4852;
assign w4854 = ~pi1128 & pi1130;
assign w4855 = w4850 & w4854;
assign w4856 = pi0633 & w4855;
assign w4857 = ~pi0223 & ~pi0224;
assign w4858 = w886 & ~w4857;
assign w4859 = ~pi0199 & w4858;
assign w4860 = pi0257 & w4859;
assign w4861 = pi1128 & pi1130;
assign w4862 = w4850 & w4861;
assign w4863 = pi0766 & w4862;
assign w4864 = w4844 & w4850;
assign w4865 = pi0815 & w4864;
assign w4866 = w4847 & w4861;
assign w4867 = pi0700 & w4866;
assign w4868 = w886 & w4857;
assign w4869 = ~w965 & w4868;
assign w4870 = w4847 & w4854;
assign w4871 = pi0634 & w4870;
assign w4872 = pi0199 & w4858;
assign w4873 = pi1059 & w4872;
assign w4874 = ~w4860 & ~w4873;
assign w4875 = ~w4849 & w4874;
assign w4876 = ~w4853 & ~w4856;
assign w4877 = ~w4863 & ~w4865;
assign w4878 = ~w4867 & ~w4869;
assign w4879 = ~w4871 & w4878;
assign w4880 = w4876 & w4877;
assign w4881 = w4875 & w4880;
assign w4882 = w4879 & w4881;
assign w4883 = ~w1085 & w4868;
assign w4884 = pi0872 & w4852;
assign w4885 = pi0785 & w4848;
assign w4886 = pi1078 & w4872;
assign w4887 = pi0772 & w4862;
assign w4888 = pi0614 & w4855;
assign w4889 = pi0662 & w4870;
assign w4890 = pi0811 & w4864;
assign w4891 = pi0727 & w4866;
assign w4892 = pi0292 & w4859;
assign w4893 = ~w4886 & ~w4892;
assign w4894 = ~w4883 & w4893;
assign w4895 = ~w4884 & ~w4885;
assign w4896 = ~w4887 & ~w4888;
assign w4897 = ~w4889 & ~w4890;
assign w4898 = ~w4891 & w4897;
assign w4899 = w4895 & w4896;
assign w4900 = w4894 & w4899;
assign w4901 = w4898 & w4900;
assign w4902 = pi1102 & w4718;
assign w4903 = pi0665 & w4720;
assign w4904 = ~w4902 & ~w4903;
assign w4905 = ~pi0799 & w4864;
assign w4906 = pi0873 & w4852;
assign w4907 = ~w1078 & w4868;
assign w4908 = pi0297 & w4859;
assign w4909 = pi0764 & w4862;
assign w4910 = pi0638 & w4870;
assign w4911 = pi0691 & w4866;
assign w4912 = pi0790 & w4848;
assign w4913 = pi0607 & w4855;
assign w4914 = pi1038 & w4872;
assign w4915 = ~w4908 & ~w4914;
assign w4916 = ~w4905 & w4915;
assign w4917 = ~w4906 & ~w4907;
assign w4918 = ~w4909 & ~w4910;
assign w4919 = ~w4911 & ~w4912;
assign w4920 = ~w4913 & w4919;
assign w4921 = w4917 & w4918;
assign w4922 = w4916 & w4921;
assign w4923 = w4920 & w4922;
assign w4924 = pi0699 & w4866;
assign w4925 = pi0763 & w4862;
assign w4926 = pi0792 & w4848;
assign w4927 = pi1066 & w4872;
assign w4928 = pi0871 & w4852;
assign w4929 = pi0681 & w4870;
assign w4930 = ~pi0809 & w4864;
assign w4931 = ~w1102 & w4868;
assign w4932 = pi0642 & w4855;
assign w4933 = pi0294 & w4859;
assign w4934 = ~w4927 & ~w4933;
assign w4935 = ~w4924 & w4934;
assign w4936 = ~w4925 & ~w4926;
assign w4937 = ~w4928 & ~w4929;
assign w4938 = ~w4930 & ~w4931;
assign w4939 = ~w4932 & w4938;
assign w4940 = w4936 & w4937;
assign w4941 = w4935 & w4940;
assign w4942 = w4939 & w4941;
assign w4943 = pi1043 & w4872;
assign w4944 = pi0837 & w4852;
assign w4945 = pi0778 & w4848;
assign w4946 = pi0291 & w4859;
assign w4947 = pi0759 & w4862;
assign w4948 = pi0696 & w4866;
assign w4949 = pi0603 & w4855;
assign w4950 = ~w1112 & w4868;
assign w4951 = pi0680 & w4870;
assign w4952 = pi0981 & w4864;
assign w4953 = ~w4943 & ~w4946;
assign w4954 = ~w4944 & w4953;
assign w4955 = ~w4945 & ~w4947;
assign w4956 = ~w4948 & ~w4949;
assign w4957 = ~w4950 & ~w4951;
assign w4958 = ~w4952 & w4957;
assign w4959 = w4955 & w4956;
assign w4960 = w4954 & w4959;
assign w4961 = w4958 & w4960;
assign w4962 = pi1119 & w4718;
assign w4963 = ~pi0669 & w4720;
assign w4964 = ~w4962 & ~w4963;
assign w4965 = pi0852 & w4852;
assign w4966 = ~pi0723 & w4866;
assign w4967 = ~pi0695 & w4870;
assign w4968 = pi0612 & w4855;
assign w4969 = ~w948 & w4868;
assign w4970 = pi0258 & w4859;
assign w4971 = pi1056 & w4872;
assign w4972 = ~pi0745 & w4862;
assign w4973 = ~w4970 & ~w4971;
assign w4974 = ~w4965 & w4973;
assign w4975 = ~w4966 & ~w4967;
assign w4976 = ~w4968 & ~w4969;
assign w4977 = ~w4972 & w4976;
assign w4978 = w4974 & w4975;
assign w4979 = w4977 & w4978;
assign w4980 = pi0865 & w4852;
assign w4981 = ~pi0646 & w4870;
assign w4982 = pi0611 & w4855;
assign w4983 = ~pi0724 & w4866;
assign w4984 = ~w975 & w4868;
assign w4985 = pi1034 & w4872;
assign w4986 = pi0261 & w4859;
assign w4987 = ~pi0741 & w4862;
assign w4988 = ~w4985 & ~w4986;
assign w4989 = ~w4980 & w4988;
assign w4990 = ~w4981 & ~w4982;
assign w4991 = ~w4983 & ~w4984;
assign w4992 = ~w4987 & w4991;
assign w4993 = w4989 & w4990;
assign w4994 = w4992 & w4993;
assign w4995 = pi0808 & w4864;
assign w4996 = pi0758 & w4862;
assign w4997 = pi0661 & w4870;
assign w4998 = pi1042 & w4872;
assign w4999 = pi0850 & w4852;
assign w5000 = ~w1132 & w4868;
assign w5001 = pi0781 & w4848;
assign w5002 = pi0736 & w4866;
assign w5003 = pi0616 & w4855;
assign w5004 = pi0290 & w4859;
assign w5005 = ~w4998 & ~w5004;
assign w5006 = ~w4995 & w5005;
assign w5007 = ~w4996 & ~w4997;
assign w5008 = ~w4999 & ~w5000;
assign w5009 = ~w5001 & ~w5002;
assign w5010 = ~w5003 & w5009;
assign w5011 = w5007 & w5008;
assign w5012 = w5006 & w5011;
assign w5013 = w5010 & w5012;
assign w5014 = pi0637 & w4870;
assign w5015 = pi0749 & w4862;
assign w5016 = ~pi0814 & w4864;
assign w5017 = pi1047 & w4872;
assign w5018 = pi0866 & w4852;
assign w5019 = pi0617 & w4855;
assign w5020 = ~w1142 & w4868;
assign w5021 = pi0706 & w4866;
assign w5022 = pi0788 & w4848;
assign w5023 = pi0295 & w4859;
assign w5024 = ~w5017 & ~w5023;
assign w5025 = ~w5014 & w5024;
assign w5026 = ~w5015 & ~w5016;
assign w5027 = ~w5018 & ~w5019;
assign w5028 = ~w5020 & ~w5021;
assign w5029 = ~w5022 & w5028;
assign w5030 = w5026 & w5027;
assign w5031 = w5025 & w5030;
assign w5032 = w5029 & w5031;
assign w5033 = pi0783 & w4848;
assign w5034 = pi0743 & w4862;
assign w5035 = pi0735 & w4866;
assign w5036 = pi0256 & w4859;
assign w5037 = pi0859 & w4852;
assign w5038 = pi0622 & w4855;
assign w5039 = pi0639 & w4870;
assign w5040 = ~w941 & w4868;
assign w5041 = pi0804 & w4864;
assign w5042 = pi1064 & w4872;
assign w5043 = ~w5036 & ~w5042;
assign w5044 = ~w5033 & w5043;
assign w5045 = ~w5034 & ~w5035;
assign w5046 = ~w5037 & ~w5038;
assign w5047 = ~w5039 & ~w5040;
assign w5048 = ~w5041 & w5047;
assign w5049 = w5045 & w5046;
assign w5050 = w5044 & w5049;
assign w5051 = w5048 & w5050;
assign w5052 = pi0789 & w4848;
assign w5053 = pi0748 & w4862;
assign w5054 = ~pi0803 & w4864;
assign w5055 = pi1031 & w4872;
assign w5056 = pi0876 & w4852;
assign w5057 = pi0623 & w4855;
assign w5058 = pi0710 & w4870;
assign w5059 = pi0730 & w4866;
assign w5060 = ~w1125 & w4868;
assign w5061 = pi0296 & w4859;
assign w5062 = ~w5055 & ~w5061;
assign w5063 = ~w5052 & w5062;
assign w5064 = ~w5053 & ~w5054;
assign w5065 = ~w5056 & ~w5057;
assign w5066 = ~w5058 & ~w5059;
assign w5067 = ~w5060 & w5066;
assign w5068 = w5064 & w5065;
assign w5069 = w5063 & w5068;
assign w5070 = w5067 & w5069;
assign w5071 = pi0729 & w4866;
assign w5072 = pi0746 & w4862;
assign w5073 = pi0787 & w4848;
assign w5074 = pi0293 & w4859;
assign w5075 = pi0881 & w4852;
assign w5076 = pi0606 & w4855;
assign w5077 = pi0643 & w4870;
assign w5078 = ~w1149 & w4868;
assign w5079 = ~pi0812 & w4864;
assign w5080 = pi1053 & w4872;
assign w5081 = ~w5074 & ~w5080;
assign w5082 = ~w5071 & w5081;
assign w5083 = ~w5072 & ~w5073;
assign w5084 = ~w5075 & ~w5076;
assign w5085 = ~w5077 & ~w5078;
assign w5086 = ~w5079 & w5085;
assign w5087 = w5083 & w5084;
assign w5088 = w5082 & w5087;
assign w5089 = w5086 & w5088;
assign w5090 = pi0870 & w4852;
assign w5091 = pi0620 & w4855;
assign w5092 = ~w911 & w4868;
assign w5093 = ~pi0704 & w4866;
assign w5094 = ~pi0635 & w4870;
assign w5095 = pi1063 & w4872;
assign w5096 = pi0259 & w4859;
assign w5097 = ~pi0742 & w4862;
assign w5098 = ~w5095 & ~w5096;
assign w5099 = ~w5090 & w5098;
assign w5100 = ~w5091 & ~w5092;
assign w5101 = ~w5093 & ~w5094;
assign w5102 = ~w5097 & w5101;
assign w5103 = w5099 & w5100;
assign w5104 = w5102 & w5103;
assign w5105 = pi0856 & w4852;
assign w5106 = ~pi0632 & w4870;
assign w5107 = ~pi0688 & w4866;
assign w5108 = ~w928 & w4868;
assign w5109 = pi0613 & w4855;
assign w5110 = pi1061 & w4872;
assign w5111 = pi0260 & w4859;
assign w5112 = ~pi0760 & w4862;
assign w5113 = ~w5110 & ~w5111;
assign w5114 = ~w5105 & w5113;
assign w5115 = ~w5106 & ~w5107;
assign w5116 = ~w5108 & ~w5109;
assign w5117 = ~w5112 & w5116;
assign w5118 = w5114 & w5115;
assign w5119 = w5117 & w5118;
assign w5120 = ~w921 & w4868;
assign w5121 = pi0874 & w4852;
assign w5122 = pi0665 & w4870;
assign w5123 = pi1030 & w4872;
assign w5124 = pi0739 & w4862;
assign w5125 = pi0690 & w4866;
assign w5126 = pi0791 & w4848;
assign w5127 = pi0621 & w4855;
assign w5128 = pi0810 & w4864;
assign w5129 = pi0255 & w4859;
assign w5130 = ~w5123 & ~w5129;
assign w5131 = ~w5120 & w5130;
assign w5132 = ~w5121 & ~w5122;
assign w5133 = ~w5124 & ~w5125;
assign w5134 = ~w5126 & ~w5127;
assign w5135 = ~w5128 & w5134;
assign w5136 = w5132 & w5133;
assign w5137 = w5131 & w5136;
assign w5138 = w5135 & w5137;
assign w5139 = pi1094 & w4718;
assign w5140 = pi0680 & w4720;
assign w5141 = ~w5139 & ~w5140;
assign w5142 = pi1097 & w4718;
assign w5143 = pi0681 & w4720;
assign w5144 = ~w5142 & ~w5143;
assign w5145 = pi0848 & w4852;
assign w5146 = pi0610 & w4855;
assign w5147 = ~pi0686 & w4866;
assign w5148 = ~pi0631 & w4870;
assign w5149 = ~w904 & w4868;
assign w5150 = pi0251 & w4859;
assign w5151 = pi1033 & w4872;
assign w5152 = ~pi0757 & w4862;
assign w5153 = ~w5150 & ~w5151;
assign w5154 = ~w5145 & w5153;
assign w5155 = ~w5146 & ~w5147;
assign w5156 = ~w5148 & ~w5149;
assign w5157 = ~w5152 & w5156;
assign w5158 = w5154 & w5155;
assign w5159 = w5157 & w5158;
assign w5160 = pi0953 & w4716;
assign w5161 = ~pi0962 & w5160;
assign w5162 = pi1124 & w5161;
assign w5163 = ~pi0962 & ~w5160;
assign w5164 = ~pi0684 & w5163;
assign w5165 = ~w5162 & ~w5164;
assign w5166 = ~w1236 & w4868;
assign w5167 = ~pi0744 & w4862;
assign w5168 = pi0813 & w4864;
assign w5169 = ~pi0200 & w4859;
assign w5170 = pi1038 & w5169;
assign w5171 = pi0860 & w4852;
assign w5172 = pi0200 & w4859;
assign w5173 = pi1061 & w5172;
assign w5174 = ~pi0728 & w4866;
assign w5175 = ~pi0657 & w4870;
assign w5176 = pi0652 & w4855;
assign w5177 = pi1070 & w4872;
assign w5178 = ~w5166 & ~w5177;
assign w5179 = ~w5167 & ~w5168;
assign w5180 = ~w5170 & ~w5171;
assign w5181 = ~w5173 & ~w5174;
assign w5182 = ~w5175 & ~w5176;
assign w5183 = w5181 & w5182;
assign w5184 = w5179 & w5180;
assign w5185 = w5178 & w5184;
assign w5186 = w5183 & w5185;
assign w5187 = pi1107 & w5161;
assign w5188 = ~pi0686 & w5163;
assign w5189 = ~w5187 & ~w5188;
assign w5190 = pi1121 & w5161;
assign w5191 = pi0687 & w5163;
assign w5192 = ~w5190 & ~w5191;
assign w5193 = pi1109 & w5161;
assign w5194 = ~pi0688 & w5163;
assign w5195 = ~w5193 & ~w5194;
assign w5196 = pi0703 & w4866;
assign w5197 = pi0843 & w4852;
assign w5198 = pi0798 & w4864;
assign w5199 = pi1030 & w5172;
assign w5200 = ~pi0752 & w4862;
assign w5201 = pi1043 & w5169;
assign w5202 = ~w1209 & w4868;
assign w5203 = pi0658 & w4855;
assign w5204 = ~pi0655 & w4870;
assign w5205 = pi1073 & w4872;
assign w5206 = ~w5196 & ~w5205;
assign w5207 = ~w5197 & ~w5198;
assign w5208 = ~w5199 & ~w5200;
assign w5209 = ~w5201 & ~w5202;
assign w5210 = ~w5203 & ~w5204;
assign w5211 = w5209 & w5210;
assign w5212 = w5207 & w5208;
assign w5213 = w5206 & w5212;
assign w5214 = w5211 & w5213;
assign w5215 = pi1102 & w5161;
assign w5216 = pi0690 & w5163;
assign w5217 = ~w5215 & ~w5216;
assign w5218 = pi1101 & w5161;
assign w5219 = pi0691 & w5163;
assign w5220 = ~w5218 & ~w5219;
assign w5221 = ~w1202 & w4868;
assign w5222 = ~pi0770 & w4862;
assign w5223 = pi0801 & w4864;
assign w5224 = pi1059 & w5172;
assign w5225 = pi0844 & w4852;
assign w5226 = pi1078 & w5169;
assign w5227 = ~pi0649 & w4870;
assign w5228 = pi0656 & w4855;
assign w5229 = pi0726 & w4866;
assign w5230 = pi1072 & w4872;
assign w5231 = ~w5221 & ~w5230;
assign w5232 = ~w5222 & ~w5223;
assign w5233 = ~w5224 & ~w5225;
assign w5234 = ~w5226 & ~w5227;
assign w5235 = ~w5228 & ~w5229;
assign w5236 = w5234 & w5235;
assign w5237 = w5232 & w5233;
assign w5238 = w5231 & w5237;
assign w5239 = w5236 & w5238;
assign w5240 = pi1123 & w4718;
assign w5241 = ~pi0693 & w4720;
assign w5242 = ~w5240 & ~w5241;
assign w5243 = pi1122 & w5161;
assign w5244 = ~pi0694 & w5163;
assign w5245 = ~w5243 & ~w5244;
assign w5246 = pi1105 & w4718;
assign w5247 = ~pi0695 & w4720;
assign w5248 = ~w5246 & ~w5247;
assign w5249 = pi1094 & w5161;
assign w5250 = pi0696 & w5163;
assign w5251 = ~w5249 & ~w5250;
assign w5252 = pi1123 & w5161;
assign w5253 = ~pi0697 & w5163;
assign w5254 = ~w5252 & ~w5253;
assign w5255 = pi1110 & w5161;
assign w5256 = ~pi0698 & w5163;
assign w5257 = ~w5255 & ~w5256;
assign w5258 = pi1097 & w5161;
assign w5259 = pi0699 & w5163;
assign w5260 = ~w5258 & ~w5259;
assign w5261 = pi1104 & w5161;
assign w5262 = pi0700 & w5163;
assign w5263 = ~w5261 & ~w5262;
assign w5264 = pi1117 & w5161;
assign w5265 = ~pi0701 & w5163;
assign w5266 = ~w5264 & ~w5265;
assign w5267 = pi1111 & w5161;
assign w5268 = ~pi0702 & w5163;
assign w5269 = ~w5267 & ~w5268;
assign w5270 = pi1118 & w5161;
assign w5271 = pi0703 & w5163;
assign w5272 = ~w5270 & ~w5271;
assign w5273 = pi1106 & w5161;
assign w5274 = ~pi0704 & w5163;
assign w5275 = ~w5273 & ~w5274;
assign w5276 = pi1119 & w5161;
assign w5277 = pi0705 & w5163;
assign w5278 = ~w5276 & ~w5277;
assign w5279 = pi1099 & w5161;
assign w5280 = pi0706 & w5163;
assign w5281 = ~w5279 & ~w5280;
assign w5282 = ~pi0753 & w4862;
assign w5283 = pi1042 & w5172;
assign w5284 = pi0304 & w5169;
assign w5285 = pi1049 & w4872;
assign w5286 = pi0618 & w4855;
assign w5287 = ~pi0702 & w4866;
assign w5288 = pi0627 & w4870;
assign w5289 = ~w1028 & w4868;
assign w5290 = pi0847 & w4852;
assign w5291 = ~w5282 & ~w5285;
assign w5292 = ~w5283 & ~w5284;
assign w5293 = ~w5286 & ~w5287;
assign w5294 = ~w5288 & ~w5289;
assign w5295 = ~w5290 & w5294;
assign w5296 = w5292 & w5293;
assign w5297 = w5291 & w5296;
assign w5298 = w5295 & w5297;
assign w5299 = ~pi0754 & w4862;
assign w5300 = pi0305 & w5169;
assign w5301 = pi1078 & w5172;
assign w5302 = pi1052 & w4872;
assign w5303 = pi0660 & w4870;
assign w5304 = ~w1062 & w4868;
assign w5305 = pi0609 & w4855;
assign w5306 = ~pi0709 & w4866;
assign w5307 = pi0857 & w4852;
assign w5308 = ~w5299 & ~w5302;
assign w5309 = ~w5300 & ~w5301;
assign w5310 = ~w5303 & ~w5304;
assign w5311 = ~w5305 & ~w5306;
assign w5312 = ~w5307 & w5311;
assign w5313 = w5309 & w5310;
assign w5314 = w5308 & w5313;
assign w5315 = w5312 & w5314;
assign w5316 = pi1112 & w5161;
assign w5317 = ~pi0709 & w5163;
assign w5318 = ~w5316 & ~w5317;
assign w5319 = pi1100 & w4718;
assign w5320 = pi0710 & w4720;
assign w5321 = ~w5319 & ~w5320;
assign w5322 = ~pi0755 & w4862;
assign w5323 = pi1053 & w5172;
assign w5324 = pi0306 & w5169;
assign w5325 = pi1081 & w4872;
assign w5326 = ~w1052 & w4868;
assign w5327 = pi0647 & w4870;
assign w5328 = pi0630 & w4855;
assign w5329 = ~pi0725 & w4866;
assign w5330 = pi0858 & w4852;
assign w5331 = ~w5322 & ~w5325;
assign w5332 = ~w5323 & ~w5324;
assign w5333 = ~w5326 & ~w5327;
assign w5334 = ~w5328 & ~w5329;
assign w5335 = ~w5330 & w5334;
assign w5336 = w5332 & w5333;
assign w5337 = w5331 & w5336;
assign w5338 = w5335 & w5337;
assign w5339 = ~pi0751 & w4862;
assign w5340 = pi0298 & w5169;
assign w5341 = pi1038 & w5172;
assign w5342 = pi1029 & w4872;
assign w5343 = ~w1035 & w4868;
assign w5344 = ~pi0701 & w4866;
assign w5345 = pi0644 & w4855;
assign w5346 = pi0715 & w4870;
assign w5347 = pi0842 & w4852;
assign w5348 = ~w5339 & ~w5342;
assign w5349 = ~w5340 & ~w5341;
assign w5350 = ~w5343 & ~w5344;
assign w5351 = ~w5345 & ~w5346;
assign w5352 = ~w5347 & w5351;
assign w5353 = w5349 & w5350;
assign w5354 = w5348 & w5353;
assign w5355 = w5352 & w5354;
assign w5356 = ~pi0756 & w4862;
assign w5357 = pi0309 & w5169;
assign w5358 = pi1066 & w5172;
assign w5359 = pi1045 & w4872;
assign w5360 = pi0628 & w4870;
assign w5361 = ~pi0734 & w4866;
assign w5362 = pi0629 & w4855;
assign w5363 = ~w1015 & w4868;
assign w5364 = pi0854 & w4852;
assign w5365 = ~w5356 & ~w5359;
assign w5366 = ~w5357 & ~w5358;
assign w5367 = ~w5360 & ~w5361;
assign w5368 = ~w5362 & ~w5363;
assign w5369 = ~w5364 & w5368;
assign w5370 = w5366 & w5367;
assign w5371 = w5365 & w5370;
assign w5372 = w5369 & w5371;
assign w5373 = ~w1226 & w4868;
assign w5374 = ~pi0762 & w4862;
assign w5375 = pi0653 & w4855;
assign w5376 = pi1047 & w5169;
assign w5377 = pi0867 & w4852;
assign w5378 = pi1033 & w5172;
assign w5379 = ~pi0693 & w4870;
assign w5380 = pi0816 & w4864;
assign w5381 = ~pi0697 & w4866;
assign w5382 = pi1051 & w4872;
assign w5383 = ~w5373 & ~w5382;
assign w5384 = ~w5374 & ~w5375;
assign w5385 = ~w5376 & ~w5377;
assign w5386 = ~w5378 & ~w5379;
assign w5387 = ~w5380 & ~w5381;
assign w5388 = w5386 & w5387;
assign w5389 = w5384 & w5385;
assign w5390 = w5383 & w5389;
assign w5391 = w5388 & w5390;
assign w5392 = pi1117 & w4718;
assign w5393 = pi0715 & w4720;
assign w5394 = ~w5392 & ~w5393;
assign w5395 = ~pi0761 & w4862;
assign w5396 = pi0307 & w5169;
assign w5397 = pi1047 & w5172;
assign w5398 = pi1037 & w4872;
assign w5399 = pi0641 & w4870;
assign w5400 = ~pi0738 & w4866;
assign w5401 = pi0626 & w4855;
assign w5402 = ~w998 & w4868;
assign w5403 = pi0845 & w4852;
assign w5404 = ~w5395 & ~w5398;
assign w5405 = ~w5396 & ~w5397;
assign w5406 = ~w5399 & ~w5400;
assign w5407 = ~w5401 & ~w5402;
assign w5408 = ~w5403 & w5407;
assign w5409 = w5405 & w5406;
assign w5410 = w5404 & w5409;
assign w5411 = w5408 & w5410;
assign w5412 = ~pi0669 & w4870;
assign w5413 = ~pi0768 & w4862;
assign w5414 = pi0800 & w4864;
assign w5415 = pi1064 & w5172;
assign w5416 = pi0839 & w4852;
assign w5417 = pi1042 & w5169;
assign w5418 = pi0645 & w4855;
assign w5419 = ~w1182 & w4868;
assign w5420 = pi0705 & w4866;
assign w5421 = pi1068 & w4872;
assign w5422 = ~w5412 & ~w5421;
assign w5423 = ~w5413 & ~w5414;
assign w5424 = ~w5415 & ~w5416;
assign w5425 = ~w5417 & ~w5418;
assign w5426 = ~w5419 & ~w5420;
assign w5427 = w5425 & w5426;
assign w5428 = w5423 & w5424;
assign w5429 = w5422 & w5428;
assign w5430 = w5427 & w5429;
assign w5431 = ~pi0767 & w4862;
assign w5432 = pi1043 & w5172;
assign w5433 = pi0303 & w5169;
assign w5434 = pi1074 & w4872;
assign w5435 = pi0608 & w4855;
assign w5436 = ~pi0698 & w4866;
assign w5437 = pi0625 & w4870;
assign w5438 = ~w991 & w4868;
assign w5439 = pi0853 & w4852;
assign w5440 = ~w5431 & ~w5434;
assign w5441 = ~w5432 & ~w5433;
assign w5442 = ~w5435 & ~w5436;
assign w5443 = ~w5437 & ~w5438;
assign w5444 = ~w5439 & w5443;
assign w5445 = w5441 & w5442;
assign w5446 = w5440 & w5445;
assign w5447 = w5444 & w5446;
assign w5448 = pi0636 & w4855;
assign w5449 = ~pi0774 & w4862;
assign w5450 = pi0687 & w4866;
assign w5451 = pi1056 & w5172;
assign w5452 = pi0868 & w4852;
assign w5453 = pi1066 & w5169;
assign w5454 = ~w1189 & w4868;
assign w5455 = pi0807 & w4864;
assign w5456 = ~pi0650 & w4870;
assign w5457 = pi1057 & w4872;
assign w5458 = ~w5448 & ~w5457;
assign w5459 = ~w5449 & ~w5450;
assign w5460 = ~w5451 & ~w5452;
assign w5461 = ~w5453 & ~w5454;
assign w5462 = ~w5455 & ~w5456;
assign w5463 = w5461 & w5462;
assign w5464 = w5459 & w5460;
assign w5465 = w5458 & w5464;
assign w5466 = w5463 & w5465;
assign w5467 = pi0651 & w4855;
assign w5468 = pi0880 & w4852;
assign w5469 = ~w1165 & w4868;
assign w5470 = pi1034 & w5172;
assign w5471 = ~pi0750 & w4862;
assign w5472 = pi1031 & w5169;
assign w5473 = ~pi0654 & w4870;
assign w5474 = ~pi0684 & w4866;
assign w5475 = pi0794 & w4864;
assign w5476 = pi1075 & w4872;
assign w5477 = ~w5467 & ~w5476;
assign w5478 = ~w5468 & ~w5469;
assign w5479 = ~w5470 & ~w5471;
assign w5480 = ~w5472 & ~w5473;
assign w5481 = ~w5474 & ~w5475;
assign w5482 = w5480 & w5481;
assign w5483 = w5478 & w5479;
assign w5484 = w5477 & w5483;
assign w5485 = w5482 & w5484;
assign w5486 = pi0775 & ~pi0816;
assign w5487 = ~pi0721 & pi0813;
assign w5488 = pi0773 & ~pi0801;
assign w5489 = pi0771 & ~pi0800;
assign w5490 = ~pi0773 & pi0801;
assign w5491 = ~pi0771 & pi0800;
assign w5492 = pi0769 & pi0794;
assign w5493 = ~pi0769 & ~pi0794;
assign w5494 = ~w5492 & ~w5493;
assign w5495 = pi0747 & pi0807;
assign w5496 = ~pi0747 & ~pi0807;
assign w5497 = ~w5495 & ~w5496;
assign w5498 = pi0731 & ~pi0795;
assign w5499 = ~pi0775 & pi0816;
assign w5500 = pi0765 & ~pi0798;
assign w5501 = pi0721 & ~pi0813;
assign w5502 = ~pi0765 & pi0798;
assign w5503 = ~pi0731 & pi0795;
assign w5504 = ~w5486 & ~w5487;
assign w5505 = ~w5488 & ~w5489;
assign w5506 = ~w5490 & ~w5491;
assign w5507 = ~w5498 & ~w5499;
assign w5508 = ~w5500 & ~w5501;
assign w5509 = ~w5502 & ~w5503;
assign w5510 = w5508 & w5509;
assign w5511 = w5506 & w5507;
assign w5512 = w5504 & w5505;
assign w5513 = ~w5494 & ~w5497;
assign w5514 = w5512 & w5513;
assign w5515 = w5510 & w5511;
assign w5516 = w5514 & w5515;
assign w5517 = ~pi0794 & ~pi0795;
assign w5518 = ~pi0798 & ~pi0800;
assign w5519 = ~pi0801 & ~pi0807;
assign w5520 = ~pi0813 & ~pi0816;
assign w5521 = w5519 & w5520;
assign w5522 = w5517 & w5518;
assign w5523 = w5521 & w5522;
assign w5524 = w5516 & ~w5523;
assign w5525 = pi0765 & ~pi0945;
assign w5526 = pi0771 & w5525;
assign w5527 = pi0773 & w5526;
assign w5528 = pi0747 & w5527;
assign w5529 = pi0731 & w5528;
assign w5530 = pi0775 & w5529;
assign w5531 = pi0769 & w5530;
assign w5532 = ~pi0721 & ~w5531;
assign w5533 = pi0721 & w5531;
assign w5534 = ~w5524 & ~w5532;
assign w5535 = ~w5533 & w5534;
assign w5536 = pi0640 & w4855;
assign w5537 = pi0851 & w4852;
assign w5538 = ~w1172 & w4868;
assign w5539 = pi1063 & w5172;
assign w5540 = ~pi0776 & w4862;
assign w5541 = pi1053 & w5169;
assign w5542 = ~pi0732 & w4870;
assign w5543 = pi0795 & w4864;
assign w5544 = ~pi0694 & w4866;
assign w5545 = pi1039 & w4872;
assign w5546 = ~w5536 & ~w5545;
assign w5547 = ~w5537 & ~w5538;
assign w5548 = ~w5539 & ~w5540;
assign w5549 = ~w5541 & ~w5542;
assign w5550 = ~w5543 & ~w5544;
assign w5551 = w5549 & w5550;
assign w5552 = w5547 & w5548;
assign w5553 = w5546 & w5552;
assign w5554 = w5551 & w5553;
assign w5555 = pi1105 & w5161;
assign w5556 = ~pi0723 & w5163;
assign w5557 = ~w5555 & ~w5556;
assign w5558 = pi1108 & w5161;
assign w5559 = ~pi0724 & w5163;
assign w5560 = ~w5558 & ~w5559;
assign w5561 = pi1114 & w5161;
assign w5562 = ~pi0725 & w5163;
assign w5563 = ~w5561 & ~w5562;
assign w5564 = pi1120 & w5161;
assign w5565 = pi0726 & w5163;
assign w5566 = ~w5564 & ~w5565;
assign w5567 = pi1096 & w5161;
assign w5568 = pi0727 & w5163;
assign w5569 = ~w5567 & ~w5568;
assign w5570 = pi1125 & w5161;
assign w5571 = ~pi0728 & w5163;
assign w5572 = ~w5570 & ~w5571;
assign w5573 = pi1098 & w5161;
assign w5574 = pi0729 & w5163;
assign w5575 = ~w5573 & ~w5574;
assign w5576 = pi1100 & w5161;
assign w5577 = pi0730 & w5163;
assign w5578 = ~w5576 & ~w5577;
assign w5579 = ~pi0731 & ~w5528;
assign w5580 = ~w5529 & ~w5579;
assign w5581 = ~w5524 & w5580;
assign w5582 = pi1122 & w4718;
assign w5583 = ~pi0732 & w4720;
assign w5584 = ~w5582 & ~w5583;
assign w5585 = pi0838 & w4852;
assign w5586 = pi1031 & w5172;
assign w5587 = pi0308 & w5169;
assign w5588 = pi1041 & w4872;
assign w5589 = ~w1008 & w4868;
assign w5590 = ~pi0737 & w4866;
assign w5591 = pi0648 & w4870;
assign w5592 = pi0619 & w4855;
assign w5593 = ~pi0777 & w4862;
assign w5594 = ~w5585 & ~w5588;
assign w5595 = ~w5586 & ~w5587;
assign w5596 = ~w5589 & ~w5590;
assign w5597 = ~w5591 & ~w5592;
assign w5598 = ~w5593 & w5597;
assign w5599 = w5595 & w5596;
assign w5600 = w5594 & w5599;
assign w5601 = w5598 & w5600;
assign w5602 = pi1113 & w5161;
assign w5603 = ~pi0734 & w5163;
assign w5604 = ~w5602 & ~w5603;
assign w5605 = pi1103 & w5161;
assign w5606 = pi0735 & w5163;
assign w5607 = ~w5605 & ~w5606;
assign w5608 = pi1095 & w5161;
assign w5609 = pi0736 & w5163;
assign w5610 = ~w5608 & ~w5609;
assign w5611 = pi1116 & w5161;
assign w5612 = ~pi0737 & w5163;
assign w5613 = ~w5611 & ~w5612;
assign w5614 = pi1115 & w5161;
assign w5615 = ~pi0738 & w5163;
assign w5616 = ~w5614 & ~w5615;
assign w5617 = ~pi0952 & w4624;
assign w5618 = pi1102 & w5617;
assign w5619 = pi0739 & ~w5617;
assign w5620 = ~pi0966 & ~w5618;
assign w5621 = ~w5619 & w5620;
assign w5622 = ~pi0741 & ~w5617;
assign w5623 = pi1108 & w5617;
assign w5624 = ~pi0966 & ~w5622;
assign w5625 = ~w5623 & w5624;
assign w5626 = ~pi0742 & ~w5617;
assign w5627 = pi1106 & w5617;
assign w5628 = ~pi0966 & ~w5626;
assign w5629 = ~w5627 & w5628;
assign w5630 = pi1103 & w5617;
assign w5631 = pi0743 & ~w5617;
assign w5632 = ~pi0966 & ~w5630;
assign w5633 = ~w5631 & w5632;
assign w5634 = ~pi0744 & ~w5617;
assign w5635 = pi1125 & w5617;
assign w5636 = ~pi0966 & ~w5634;
assign w5637 = ~w5635 & w5636;
assign w5638 = ~pi0745 & ~w5617;
assign w5639 = pi1105 & w5617;
assign w5640 = ~pi0966 & ~w5638;
assign w5641 = ~w5639 & w5640;
assign w5642 = pi1098 & w5617;
assign w5643 = pi0746 & ~w5617;
assign w5644 = ~pi0966 & ~w5642;
assign w5645 = ~w5643 & w5644;
assign w5646 = ~pi0747 & ~w5527;
assign w5647 = ~w5528 & ~w5646;
assign w5648 = ~w5524 & w5647;
assign w5649 = pi1100 & w5617;
assign w5650 = pi0748 & ~w5617;
assign w5651 = ~pi0966 & ~w5649;
assign w5652 = ~w5650 & w5651;
assign w5653 = pi1099 & w5617;
assign w5654 = pi0749 & ~w5617;
assign w5655 = ~pi0966 & ~w5653;
assign w5656 = ~w5654 & w5655;
assign w5657 = ~pi0750 & ~w5617;
assign w5658 = pi1124 & w5617;
assign w5659 = ~pi0966 & ~w5657;
assign w5660 = ~w5658 & w5659;
assign w5661 = ~pi0751 & ~w5617;
assign w5662 = pi1117 & w5617;
assign w5663 = ~pi0966 & ~w5661;
assign w5664 = ~w5662 & w5663;
assign w5665 = ~pi0752 & ~w5617;
assign w5666 = pi1118 & w5617;
assign w5667 = ~pi0966 & ~w5665;
assign w5668 = ~w5666 & w5667;
assign w5669 = ~pi0753 & ~w5617;
assign w5670 = pi1111 & w5617;
assign w5671 = ~pi0966 & ~w5669;
assign w5672 = ~w5670 & w5671;
assign w5673 = ~pi0754 & ~w5617;
assign w5674 = pi1112 & w5617;
assign w5675 = ~pi0966 & ~w5673;
assign w5676 = ~w5674 & w5675;
assign w5677 = ~pi0755 & ~w5617;
assign w5678 = pi1114 & w5617;
assign w5679 = ~pi0966 & ~w5677;
assign w5680 = ~w5678 & w5679;
assign w5681 = ~pi0756 & ~w5617;
assign w5682 = pi1113 & w5617;
assign w5683 = ~pi0966 & ~w5681;
assign w5684 = ~w5682 & w5683;
assign w5685 = ~pi0757 & ~w5617;
assign w5686 = pi1107 & w5617;
assign w5687 = ~pi0966 & ~w5685;
assign w5688 = ~w5686 & w5687;
assign w5689 = pi1095 & w5617;
assign w5690 = pi0758 & ~w5617;
assign w5691 = ~pi0966 & ~w5689;
assign w5692 = ~w5690 & w5691;
assign w5693 = pi1094 & w5617;
assign w5694 = pi0759 & ~w5617;
assign w5695 = ~pi0966 & ~w5693;
assign w5696 = ~w5694 & w5695;
assign w5697 = ~pi0760 & ~w5617;
assign w5698 = pi1109 & w5617;
assign w5699 = ~pi0966 & ~w5697;
assign w5700 = ~w5698 & w5699;
assign w5701 = ~pi0761 & ~w5617;
assign w5702 = pi1115 & w5617;
assign w5703 = ~pi0966 & ~w5701;
assign w5704 = ~w5702 & w5703;
assign w5705 = ~pi0762 & ~w5617;
assign w5706 = pi1123 & w5617;
assign w5707 = ~pi0966 & ~w5705;
assign w5708 = ~w5706 & w5707;
assign w5709 = pi1097 & w5617;
assign w5710 = pi0763 & ~w5617;
assign w5711 = ~pi0966 & ~w5709;
assign w5712 = ~w5710 & w5711;
assign w5713 = pi1101 & w5617;
assign w5714 = pi0764 & ~w5617;
assign w5715 = ~pi0966 & ~w5713;
assign w5716 = ~w5714 & w5715;
assign w5717 = ~pi0765 & pi0945;
assign w5718 = ~w5525 & ~w5717;
assign w5719 = ~w5524 & w5718;
assign w5720 = pi1104 & w5617;
assign w5721 = pi0766 & ~w5617;
assign w5722 = ~pi0966 & ~w5720;
assign w5723 = ~w5721 & w5722;
assign w5724 = ~pi0767 & ~w5617;
assign w5725 = pi1110 & w5617;
assign w5726 = ~pi0966 & ~w5724;
assign w5727 = ~w5725 & w5726;
assign w5728 = ~pi0768 & ~w5617;
assign w5729 = pi1119 & w5617;
assign w5730 = ~pi0966 & ~w5728;
assign w5731 = ~w5729 & w5730;
assign w5732 = ~pi0769 & ~w5530;
assign w5733 = ~w5524 & ~w5531;
assign w5734 = ~w5732 & w5733;
assign w5735 = ~pi0770 & ~w5617;
assign w5736 = pi1120 & w5617;
assign w5737 = ~pi0966 & ~w5735;
assign w5738 = ~w5736 & w5737;
assign w5739 = ~pi0771 & ~w5525;
assign w5740 = ~w5526 & ~w5739;
assign w5741 = ~w5524 & w5740;
assign w5742 = pi1096 & w5617;
assign w5743 = pi0772 & ~w5617;
assign w5744 = ~pi0966 & ~w5742;
assign w5745 = ~w5743 & w5744;
assign w5746 = ~pi0773 & ~w5526;
assign w5747 = ~w5527 & ~w5746;
assign w5748 = ~w5524 & w5747;
assign w5749 = ~pi0774 & ~w5617;
assign w5750 = pi1121 & w5617;
assign w5751 = ~pi0966 & ~w5749;
assign w5752 = ~w5750 & w5751;
assign w5753 = ~pi0775 & ~w5529;
assign w5754 = ~w5524 & ~w5530;
assign w5755 = ~w5753 & w5754;
assign w5756 = ~pi0776 & ~w5617;
assign w5757 = pi1122 & w5617;
assign w5758 = ~pi0966 & ~w5756;
assign w5759 = ~w5757 & w5758;
assign w5760 = ~pi0777 & ~w5617;
assign w5761 = pi1116 & w5617;
assign w5762 = ~pi0966 & ~w5760;
assign w5763 = ~w5761 & w5762;
assign w5764 = pi0832 & pi0956;
assign w5765 = ~pi1040 & ~pi1077;
assign w5766 = pi1079 & w5765;
assign w5767 = w5764 & w5766;
assign w5768 = ~pi0968 & w5767;
assign w5769 = pi0778 & ~w5768;
assign w5770 = pi1094 & w5768;
assign w5771 = ~w5769 & ~w5770;
assign w5772 = pi0779 & ~w4675;
assign w5773 = pi0780 & ~w4603;
assign w5774 = pi0781 & ~w5768;
assign w5775 = pi1095 & w5768;
assign w5776 = ~w5774 & ~w5775;
assign w5777 = ~w3753 & ~w4637;
assign w5778 = ~w4602 & w5777;
assign w5779 = pi0783 & ~w5768;
assign w5780 = pi1103 & w5768;
assign w5781 = ~w5779 & ~w5780;
assign w5782 = pi0784 & ~w5768;
assign w5783 = pi1104 & w5768;
assign w5784 = ~w5782 & ~w5783;
assign w5785 = pi0785 & ~w5768;
assign w5786 = pi1096 & w5768;
assign w5787 = ~w5785 & ~w5786;
assign w5788 = pi0786 & pi0954;
assign w5789 = pi0024 & ~pi0954;
assign w5790 = ~w5788 & ~w5789;
assign w5791 = pi0787 & ~w5768;
assign w5792 = pi1098 & w5768;
assign w5793 = ~w5791 & ~w5792;
assign w5794 = pi0788 & ~w5768;
assign w5795 = pi1099 & w5768;
assign w5796 = ~w5794 & ~w5795;
assign w5797 = pi0789 & ~w5768;
assign w5798 = pi1100 & w5768;
assign w5799 = ~w5797 & ~w5798;
assign w5800 = pi0790 & ~w5768;
assign w5801 = pi1101 & w5768;
assign w5802 = ~w5800 & ~w5801;
assign w5803 = pi0791 & ~w5768;
assign w5804 = pi1102 & w5768;
assign w5805 = ~w5803 & ~w5804;
assign w5806 = pi0792 & ~w5768;
assign w5807 = pi1097 & w5768;
assign w5808 = ~w5806 & ~w5807;
assign w5809 = pi0968 & w5767;
assign w5810 = pi0794 & ~w5809;
assign w5811 = pi1124 & w5809;
assign w5812 = ~w5810 & ~w5811;
assign w5813 = pi0795 & ~w5809;
assign w5814 = pi1122 & w5809;
assign w5815 = ~w5813 & ~w5814;
assign w5816 = pi0264 & ~w4829;
assign w5817 = ~w4830 & ~w5816;
assign w5818 = pi0798 & ~w5809;
assign w5819 = pi1118 & w5809;
assign w5820 = ~w5818 & ~w5819;
assign w5821 = pi0799 & ~w5809;
assign w5822 = ~pi1101 & w5809;
assign w5823 = ~w5821 & ~w5822;
assign w5824 = pi0800 & ~w5809;
assign w5825 = pi1119 & w5809;
assign w5826 = ~w5824 & ~w5825;
assign w5827 = pi0801 & ~w5809;
assign w5828 = pi1120 & w5809;
assign w5829 = ~w5827 & ~w5828;
assign w5830 = pi0803 & ~w5809;
assign w5831 = ~pi1100 & w5809;
assign w5832 = ~w5830 & ~w5831;
assign w5833 = pi0804 & ~w5809;
assign w5834 = pi1103 & w5809;
assign w5835 = ~w5833 & ~w5834;
assign w5836 = pi0270 & ~w4827;
assign w5837 = ~w4828 & ~w5836;
assign w5838 = pi0807 & ~w5809;
assign w5839 = pi1121 & w5809;
assign w5840 = ~w5838 & ~w5839;
assign w5841 = pi0808 & ~w5809;
assign w5842 = pi1095 & w5809;
assign w5843 = ~w5841 & ~w5842;
assign w5844 = pi0809 & ~w5809;
assign w5845 = ~pi1097 & w5809;
assign w5846 = ~w5844 & ~w5845;
assign w5847 = pi0810 & ~w5809;
assign w5848 = pi1102 & w5809;
assign w5849 = ~w5847 & ~w5848;
assign w5850 = pi0811 & ~w5809;
assign w5851 = pi1096 & w5809;
assign w5852 = ~w5850 & ~w5851;
assign w5853 = pi0812 & ~w5809;
assign w5854 = ~pi1098 & w5809;
assign w5855 = ~w5853 & ~w5854;
assign w5856 = pi0813 & ~w5809;
assign w5857 = pi1125 & w5809;
assign w5858 = ~w5856 & ~w5857;
assign w5859 = pi0814 & ~w5809;
assign w5860 = ~pi1099 & w5809;
assign w5861 = ~w5859 & ~w5860;
assign w5862 = pi0815 & ~w5809;
assign w5863 = pi1104 & w5809;
assign w5864 = ~w5862 & ~w5863;
assign w5865 = pi0816 & ~w5809;
assign w5866 = pi1123 & w5809;
assign w5867 = ~w5865 & ~w5866;
assign w5868 = pi0269 & ~w4824;
assign w5869 = ~w4825 & ~w5868;
assign w5870 = pi0265 & ~w4830;
assign w5871 = ~w4831 & ~w5870;
assign w5872 = pi0277 & ~w4828;
assign w5873 = ~w4829 & ~w5872;
assign w5874 = ~pi0811 & ~pi0893;
assign w5875 = ~pi0982 & pi1086;
assign w5876 = ~pi1085 & w1666;
assign w5877 = ~w5875 & ~w5876;
assign w5878 = w257 & ~w5877;
assign w5879 = pi0123 & ~pi0222;
assign w5880 = w4857 & w5879;
assign w5881 = ~pi0825 & w5880;
assign w5882 = pi1120 & ~pi1121;
assign w5883 = ~pi1120 & pi1121;
assign w5884 = ~w5882 & ~w5883;
assign w5885 = pi1122 & ~pi1125;
assign w5886 = ~pi1122 & pi1125;
assign w5887 = ~w5885 & ~w5886;
assign w5888 = ~pi1123 & ~pi1124;
assign w5889 = pi1123 & pi1124;
assign w5890 = ~w5888 & ~w5889;
assign w5891 = ~pi1118 & ~pi1119;
assign w5892 = pi1118 & pi1119;
assign w5893 = ~w5891 & ~w5892;
assign w5894 = w5890 & ~w5893;
assign w5895 = ~w5890 & w5893;
assign w5896 = ~w5894 & ~w5895;
assign w5897 = w5887 & w5896;
assign w5898 = ~w5887 & ~w5896;
assign w5899 = ~w5897 & ~w5898;
assign w5900 = ~w5884 & w5899;
assign w5901 = w5884 & ~w5899;
assign w5902 = ~w5880 & ~w5900;
assign w5903 = ~w5901 & w5902;
assign w5904 = ~w5881 & ~w5903;
assign w5905 = ~pi0826 & w5880;
assign w5906 = pi1115 & ~pi1117;
assign w5907 = ~pi1115 & pi1117;
assign w5908 = ~w5906 & ~w5907;
assign w5909 = pi1112 & ~pi1113;
assign w5910 = ~pi1112 & pi1113;
assign w5911 = ~w5909 & ~w5910;
assign w5912 = ~pi1110 & ~pi1111;
assign w5913 = pi1110 & pi1111;
assign w5914 = ~w5912 & ~w5913;
assign w5915 = ~pi1114 & ~pi1116;
assign w5916 = pi1114 & pi1116;
assign w5917 = ~w5915 & ~w5916;
assign w5918 = w5914 & ~w5917;
assign w5919 = ~w5914 & w5917;
assign w5920 = ~w5918 & ~w5919;
assign w5921 = w5911 & w5920;
assign w5922 = ~w5911 & ~w5920;
assign w5923 = ~w5921 & ~w5922;
assign w5924 = ~w5908 & w5923;
assign w5925 = w5908 & ~w5923;
assign w5926 = ~w5880 & ~w5924;
assign w5927 = ~w5925 & w5926;
assign w5928 = ~w5905 & ~w5927;
assign w5929 = ~pi0827 & w5880;
assign w5930 = pi1094 & ~pi1095;
assign w5931 = ~pi1094 & pi1095;
assign w5932 = ~w5930 & ~w5931;
assign w5933 = pi1100 & ~pi1101;
assign w5934 = ~pi1100 & pi1101;
assign w5935 = ~w5933 & ~w5934;
assign w5936 = ~pi1096 & ~pi1097;
assign w5937 = pi1096 & pi1097;
assign w5938 = ~w5936 & ~w5937;
assign w5939 = ~pi1098 & ~pi1099;
assign w5940 = pi1098 & pi1099;
assign w5941 = ~w5939 & ~w5940;
assign w5942 = w5938 & ~w5941;
assign w5943 = ~w5938 & w5941;
assign w5944 = ~w5942 & ~w5943;
assign w5945 = w5935 & w5944;
assign w5946 = ~w5935 & ~w5944;
assign w5947 = ~w5945 & ~w5946;
assign w5948 = ~w5932 & w5947;
assign w5949 = w5932 & ~w5947;
assign w5950 = ~w5880 & ~w5948;
assign w5951 = ~w5949 & w5950;
assign w5952 = ~w5929 & ~w5951;
assign w5953 = ~pi0828 & w5880;
assign w5954 = pi1107 & ~pi1108;
assign w5955 = ~pi1107 & pi1108;
assign w5956 = ~w5954 & ~w5955;
assign w5957 = pi1102 & ~pi1103;
assign w5958 = ~pi1102 & pi1103;
assign w5959 = ~w5957 & ~w5958;
assign w5960 = ~pi1104 & ~pi1105;
assign w5961 = pi1104 & pi1105;
assign w5962 = ~w5960 & ~w5961;
assign w5963 = ~pi1106 & ~pi1109;
assign w5964 = pi1106 & pi1109;
assign w5965 = ~w5963 & ~w5964;
assign w5966 = w5962 & ~w5965;
assign w5967 = ~w5962 & w5965;
assign w5968 = ~w5966 & ~w5967;
assign w5969 = w5959 & w5968;
assign w5970 = ~w5959 & ~w5968;
assign w5971 = ~w5969 & ~w5970;
assign w5972 = ~w5956 & w5971;
assign w5973 = w5956 & ~w5971;
assign w5974 = ~w5880 & ~w5972;
assign w5975 = ~w5973 & w5974;
assign w5976 = ~w5953 & ~w5975;
assign w5977 = ~pi0951 & pi1086;
assign w5978 = w886 & w4064;
assign w5979 = ~w5977 & ~w5978;
assign w5980 = pi0281 & ~w4825;
assign w5981 = ~w4826 & ~w5980;
assign w5982 = ~pi0832 & w1256;
assign w5983 = w4064 & w5982;
assign w5984 = pi0833 & ~w1254;
assign w5985 = ~w4064 & ~w5984;
assign w5986 = pi0946 & w1254;
assign w5987 = pi0282 & ~w4826;
assign w5988 = ~w4827 & ~w5987;
assign w5989 = pi0837 & pi0955;
assign w5990 = ~pi0955 & pi1043;
assign w5991 = ~w5989 & ~w5990;
assign w5992 = pi0838 & pi0955;
assign w5993 = ~pi0955 & pi1041;
assign w5994 = ~w5992 & ~w5993;
assign w5995 = pi0839 & pi0955;
assign w5996 = ~pi0955 & pi1068;
assign w5997 = ~w5995 & ~w5996;
assign w5998 = pi0840 & ~w1254;
assign w5999 = pi1190 & w1254;
assign w6000 = ~w5998 & ~w5999;
assign w6001 = pi0842 & pi0955;
assign w6002 = ~pi0955 & pi1029;
assign w6003 = ~w6001 & ~w6002;
assign w6004 = pi0843 & pi0955;
assign w6005 = ~pi0955 & pi1073;
assign w6006 = ~w6004 & ~w6005;
assign w6007 = pi0844 & pi0955;
assign w6008 = ~pi0955 & pi1072;
assign w6009 = ~w6007 & ~w6008;
assign w6010 = pi0845 & pi0955;
assign w6011 = ~pi0955 & pi1037;
assign w6012 = ~w6010 & ~w6011;
assign w6013 = pi1128 & ~w2979;
assign w6014 = pi0846 & w2979;
assign w6015 = ~w6013 & ~w6014;
assign w6016 = pi0847 & pi0955;
assign w6017 = ~pi0955 & pi1049;
assign w6018 = ~w6016 & ~w6017;
assign w6019 = pi0848 & pi0955;
assign w6020 = ~pi0955 & pi1033;
assign w6021 = ~w6019 & ~w6020;
assign w6022 = pi0849 & ~w1254;
assign w6023 = pi1192 & w1254;
assign w6024 = ~w6022 & ~w6023;
assign w6025 = pi0850 & pi0955;
assign w6026 = ~pi0955 & pi1042;
assign w6027 = ~w6025 & ~w6026;
assign w6028 = pi0851 & pi0955;
assign w6029 = ~pi0955 & pi1039;
assign w6030 = ~w6028 & ~w6029;
assign w6031 = pi0852 & pi0955;
assign w6032 = ~pi0955 & pi1056;
assign w6033 = ~w6031 & ~w6032;
assign w6034 = pi0853 & pi0955;
assign w6035 = ~pi0955 & pi1074;
assign w6036 = ~w6034 & ~w6035;
assign w6037 = pi0854 & pi0955;
assign w6038 = ~pi0955 & pi1045;
assign w6039 = ~w6037 & ~w6038;
assign w6040 = pi0855 & pi0955;
assign w6041 = ~pi0955 & pi1059;
assign w6042 = ~w6040 & ~w6041;
assign w6043 = pi0856 & pi0955;
assign w6044 = ~pi0955 & pi1061;
assign w6045 = ~w6043 & ~w6044;
assign w6046 = pi0857 & pi0955;
assign w6047 = ~pi0955 & pi1052;
assign w6048 = ~w6046 & ~w6047;
assign w6049 = pi0858 & pi0955;
assign w6050 = ~pi0955 & pi1081;
assign w6051 = ~w6049 & ~w6050;
assign w6052 = pi0859 & pi0955;
assign w6053 = ~pi0955 & pi1064;
assign w6054 = ~w6052 & ~w6053;
assign w6055 = pi0860 & pi0955;
assign w6056 = ~pi0955 & pi1070;
assign w6057 = ~w6055 & ~w6056;
assign w6058 = pi1135 & ~w2979;
assign w6059 = pi0861 & w2979;
assign w6060 = ~w6058 & ~w6059;
assign w6061 = pi1133 & ~w2979;
assign w6062 = pi0862 & w2979;
assign w6063 = ~w6061 & ~w6062;
assign w6064 = pi0863 & ~w1254;
assign w6065 = pi1193 & w1254;
assign w6066 = ~w6064 & ~w6065;
assign w6067 = pi0864 & ~w1254;
assign w6068 = pi1191 & w1254;
assign w6069 = ~w6067 & ~w6068;
assign w6070 = pi0865 & pi0955;
assign w6071 = ~pi0955 & pi1034;
assign w6072 = ~w6070 & ~w6071;
assign w6073 = pi0866 & pi0955;
assign w6074 = ~pi0955 & pi1047;
assign w6075 = ~w6073 & ~w6074;
assign w6076 = pi0867 & pi0955;
assign w6077 = ~pi0955 & pi1051;
assign w6078 = ~w6076 & ~w6077;
assign w6079 = pi0868 & pi0955;
assign w6080 = ~pi0955 & pi1057;
assign w6081 = ~w6079 & ~w6080;
assign w6082 = pi1134 & ~w2979;
assign w6083 = pi0869 & w2979;
assign w6084 = ~w6082 & ~w6083;
assign w6085 = pi0870 & pi0955;
assign w6086 = ~pi0955 & pi1063;
assign w6087 = ~w6085 & ~w6086;
assign w6088 = pi0871 & pi0955;
assign w6089 = ~pi0955 & pi1066;
assign w6090 = ~w6088 & ~w6089;
assign w6091 = pi0872 & pi0955;
assign w6092 = ~pi0955 & pi1078;
assign w6093 = ~w6091 & ~w6092;
assign w6094 = pi0873 & pi0955;
assign w6095 = ~pi0955 & pi1038;
assign w6096 = ~w6094 & ~w6095;
assign w6097 = pi0874 & pi0955;
assign w6098 = ~pi0955 & pi1030;
assign w6099 = ~w6097 & ~w6098;
assign w6100 = pi1130 & ~w2979;
assign w6101 = pi0875 & w2979;
assign w6102 = ~w6100 & ~w6101;
assign w6103 = pi0876 & pi0955;
assign w6104 = ~pi0955 & pi1031;
assign w6105 = ~w6103 & ~w6104;
assign w6106 = pi1132 & ~w2979;
assign w6107 = pi0877 & w2979;
assign w6108 = ~w6106 & ~w6107;
assign w6109 = pi1131 & ~w2979;
assign w6110 = pi0878 & w2979;
assign w6111 = ~w6109 & ~w6110;
assign w6112 = pi1129 & ~w2979;
assign w6113 = pi0879 & w2979;
assign w6114 = ~w6112 & ~w6113;
assign w6115 = pi0880 & pi0955;
assign w6116 = ~pi0955 & pi1075;
assign w6117 = ~w6115 & ~w6116;
assign w6118 = pi0881 & pi0955;
assign w6119 = ~pi0955 & pi1053;
assign w6120 = ~w6118 & ~w6119;
assign w6121 = pi1101 & ~w5880;
assign w6122 = ~pi0883 & w5880;
assign w6123 = ~w6121 & ~w6122;
assign w6124 = pi1118 & ~w5880;
assign w6125 = ~pi0884 & w5880;
assign w6126 = ~w6124 & ~w6125;
assign w6127 = pi1119 & ~w5880;
assign w6128 = ~pi0885 & w5880;
assign w6129 = ~w6127 & ~w6128;
assign w6130 = pi1103 & ~w5880;
assign w6131 = ~pi0886 & w5880;
assign w6132 = ~w6130 & ~w6131;
assign w6133 = pi1094 & ~w5880;
assign w6134 = ~pi0887 & w5880;
assign w6135 = ~w6133 & ~w6134;
assign w6136 = pi1114 & ~w5880;
assign w6137 = ~pi0888 & w5880;
assign w6138 = ~w6136 & ~w6137;
assign w6139 = pi1097 & ~w5880;
assign w6140 = ~pi0889 & w5880;
assign w6141 = ~w6139 & ~w6140;
assign w6142 = pi1120 & ~w5880;
assign w6143 = ~pi0890 & w5880;
assign w6144 = ~w6142 & ~w6143;
assign w6145 = pi1110 & ~w5880;
assign w6146 = ~pi0891 & w5880;
assign w6147 = ~w6145 & ~w6146;
assign w6148 = pi1095 & ~w5880;
assign w6149 = ~pi0892 & w5880;
assign w6150 = ~w6148 & ~w6149;
assign w6151 = pi1113 & ~w5880;
assign w6152 = ~pi0894 & w5880;
assign w6153 = ~w6151 & ~w6152;
assign w6154 = pi1107 & ~w5880;
assign w6155 = ~pi0895 & w5880;
assign w6156 = ~w6154 & ~w6155;
assign w6157 = pi1112 & ~w5880;
assign w6158 = ~pi0896 & w5880;
assign w6159 = ~w6157 & ~w6158;
assign w6160 = pi1123 & ~w5880;
assign w6161 = ~pi0898 & w5880;
assign w6162 = ~w6160 & ~w6161;
assign w6163 = pi1109 & ~w5880;
assign w6164 = ~pi0899 & w5880;
assign w6165 = ~w6163 & ~w6164;
assign w6166 = pi1104 & ~w5880;
assign w6167 = ~pi0900 & w5880;
assign w6168 = ~w6166 & ~w6167;
assign w6169 = pi1105 & ~w5880;
assign w6170 = ~pi0902 & w5880;
assign w6171 = ~w6169 & ~w6170;
assign w6172 = pi1115 & ~w5880;
assign w6173 = ~pi0903 & w5880;
assign w6174 = ~w6172 & ~w6173;
assign w6175 = pi1121 & ~w5880;
assign w6176 = ~pi0904 & w5880;
assign w6177 = ~w6175 & ~w6176;
assign w6178 = pi1125 & ~w5880;
assign w6179 = ~pi0905 & w5880;
assign w6180 = ~w6178 & ~w6179;
assign w6181 = pi1122 & ~w5880;
assign w6182 = ~pi0906 & w5880;
assign w6183 = ~w6181 & ~w6182;
assign w6184 = ~pi0782 & pi0907;
assign w6185 = pi0624 & ~pi0979;
assign w6186 = pi0598 & pi0979;
assign w6187 = pi0782 & ~w6185;
assign w6188 = ~w6186 & w6187;
assign w6189 = ~pi0604 & ~pi0979;
assign w6190 = pi0615 & pi0979;
assign w6191 = ~w6189 & ~w6190;
assign w6192 = w6188 & w6191;
assign w6193 = ~w6184 & ~w6192;
assign w6194 = pi1116 & ~w5880;
assign w6195 = ~pi0908 & w5880;
assign w6196 = ~w6194 & ~w6195;
assign w6197 = pi1099 & ~w5880;
assign w6198 = ~pi0909 & w5880;
assign w6199 = ~w6197 & ~w6198;
assign w6200 = pi1111 & ~w5880;
assign w6201 = ~pi0910 & w5880;
assign w6202 = ~w6200 & ~w6201;
assign w6203 = pi1124 & ~w5880;
assign w6204 = ~pi0911 & w5880;
assign w6205 = ~w6203 & ~w6204;
assign w6206 = pi1108 & ~w5880;
assign w6207 = ~pi0912 & w5880;
assign w6208 = ~w6206 & ~w6207;
assign w6209 = pi1100 & ~w5880;
assign w6210 = ~pi0913 & w5880;
assign w6211 = ~w6209 & ~w6210;
assign w6212 = pi0280 & ~w4823;
assign w6213 = ~w4824 & ~w6212;
assign w6214 = pi1102 & ~w5880;
assign w6215 = ~pi0915 & w5880;
assign w6216 = ~w6214 & ~w6215;
assign w6217 = pi1117 & ~w5880;
assign w6218 = ~pi0916 & w5880;
assign w6219 = ~w6217 & ~w6218;
assign w6220 = pi1106 & ~w5880;
assign w6221 = ~pi0917 & w5880;
assign w6222 = ~w6220 & ~w6221;
assign w6223 = pi1098 & ~w5880;
assign w6224 = ~pi0918 & w5880;
assign w6225 = ~w6223 & ~w6224;
assign w6226 = pi1096 & ~w5880;
assign w6227 = ~pi0919 & w5880;
assign w6228 = ~w6226 & ~w6227;
assign w6229 = pi1087 & pi1133;
assign w6230 = pi0920 & ~pi1087;
assign w6231 = ~w6229 & ~w6230;
assign w6232 = pi1087 & pi1134;
assign w6233 = pi0921 & ~pi1087;
assign w6234 = ~w6232 & ~w6233;
assign w6235 = pi1087 & pi1146;
assign w6236 = pi0922 & ~pi1087;
assign w6237 = ~w6235 & ~w6236;
assign w6238 = pi1087 & pi1148;
assign w6239 = pi0923 & ~pi1087;
assign w6240 = ~w6238 & ~w6239;
assign w6241 = ~pi0300 & pi0301;
assign w6242 = pi0311 & ~pi0312;
assign w6243 = w6241 & w6242;
assign w6244 = pi1087 & pi1149;
assign w6245 = pi0925 & ~pi1087;
assign w6246 = ~w6244 & ~w6245;
assign w6247 = pi1087 & pi1151;
assign w6248 = pi0926 & ~pi1087;
assign w6249 = ~w6247 & ~w6248;
assign w6250 = pi1087 & pi1139;
assign w6251 = pi0927 & ~pi1087;
assign w6252 = ~w6250 & ~w6251;
assign w6253 = pi1087 & pi1130;
assign w6254 = pi0928 & ~pi1087;
assign w6255 = ~w6253 & ~w6254;
assign w6256 = pi1087 & pi1138;
assign w6257 = pi0929 & ~pi1087;
assign w6258 = ~w6256 & ~w6257;
assign w6259 = pi1087 & pi1128;
assign w6260 = pi0930 & ~pi1087;
assign w6261 = ~w6259 & ~w6260;
assign w6262 = pi1087 & pi1144;
assign w6263 = pi0931 & ~pi1087;
assign w6264 = ~w6262 & ~w6263;
assign w6265 = pi1087 & pi1136;
assign w6266 = pi0932 & ~pi1087;
assign w6267 = ~w6265 & ~w6266;
assign w6268 = pi1087 & pi1131;
assign w6269 = pi0933 & ~pi1087;
assign w6270 = ~w6268 & ~w6269;
assign w6271 = pi1087 & pi1141;
assign w6272 = pi0934 & ~pi1087;
assign w6273 = ~w6271 & ~w6272;
assign w6274 = pi1087 & pi1135;
assign w6275 = pi0935 & ~pi1087;
assign w6276 = ~w6274 & ~w6275;
assign w6277 = pi1087 & pi1143;
assign w6278 = pi0936 & ~pi1087;
assign w6279 = ~w6277 & ~w6278;
assign w6280 = pi1087 & pi1142;
assign w6281 = pi0937 & ~pi1087;
assign w6282 = ~w6280 & ~w6281;
assign w6283 = pi1087 & pi1129;
assign w6284 = pi0938 & ~pi1087;
assign w6285 = ~w6283 & ~w6284;
assign w6286 = pi1087 & pi1140;
assign w6287 = pi0939 & ~pi1087;
assign w6288 = ~w6286 & ~w6287;
assign w6289 = pi1087 & pi1132;
assign w6290 = pi0940 & ~pi1087;
assign w6291 = ~w6289 & ~w6290;
assign w6292 = pi1087 & pi1147;
assign w6293 = pi0941 & ~pi1087;
assign w6294 = ~w6292 & ~w6293;
assign w6295 = pi1087 & pi1150;
assign w6296 = pi0942 & ~pi1087;
assign w6297 = ~w6295 & ~w6296;
assign w6298 = pi1087 & pi1145;
assign w6299 = pi0943 & ~pi1087;
assign w6300 = ~w6298 & ~w6299;
assign w6301 = pi1087 & pi1137;
assign w6302 = pi0944 & ~pi1087;
assign w6303 = ~w6301 & ~w6302;
assign w6304 = ~w700 & ~w708;
assign w6305 = ~pi0782 & ~pi0947;
assign w6306 = ~w6188 & ~w6305;
assign w6307 = ~pi0266 & ~w4822;
assign w6308 = ~w4823 & ~w6307;
assign w6309 = pi0313 & ~pi0954;
assign w6310 = ~pi0949 & pi0954;
assign w6311 = ~w6309 & ~w6310;
assign w6312 = ~pi0031 & ~w254;
assign w6313 = ~pi0278 & ~pi0279;
assign w6314 = ~w4822 & ~w6313;
assign w6315 = ~pi0782 & pi0960;
assign w6316 = ~pi0230 & pi0961;
assign w6317 = ~pi0782 & pi0963;
assign w6318 = ~pi0230 & pi0967;
assign w6319 = ~pi0230 & pi0969;
assign w6320 = ~pi0782 & pi0970;
assign w6321 = ~pi0230 & pi0971;
assign w6322 = ~pi0782 & pi0972;
assign w6323 = ~pi0230 & pi0974;
assign w6324 = ~pi0782 & pi0975;
assign w6325 = ~pi0230 & pi0977;
assign w6326 = ~pi0782 & pi0978;
assign w6327 = ~pi0598 & pi0615;
assign w6328 = ~pi0604 & ~pi0624;
assign w6329 = w21 & w23;
assign w6330 = w56 & w61;
assign w6331 = w41 & w103;
assign w6332 = w71 & w115;
assign w6333 = w31 & w120;
assign w6334 = w2 & w131;
assign w6335 = w113 & w137;
assign w6336 = w89 & w142;
assign w6337 = w89 & w139;
assign w6338 = ~pi0083 & w82;
assign w6339 = w60 & w165;
assign w6340 = w64 & ~pi0109;
assign w6341 = w71 & w171;
assign w6342 = ~pi0083 & ~w186;
assign w6343 = w35 & w197;
assign w6344 = w26 & w199;
assign w6345 = w26 & w204;
assign w6346 = w89 & w211;
assign w6347 = ~w3 & pi0166;
assign w6348 = w3 & pi0189;
assign w6349 = ~w3 & pi0161;
assign w6350 = w3 & pi0144;
assign w6351 = ~w3 & pi0152;
assign w6352 = w3 & pi0174;
assign w6353 = w35 & w277;
assign w6354 = w89 & w300;
assign w6355 = w28 & w306;
assign w6356 = w38 & w311;
assign w6357 = w119 & w316;
assign w6358 = w71 & w321;
assign w6359 = w71 & w331;
assign w6360 = w32 & w356;
assign w6361 = w55 & w361;
assign w6362 = w67 & w70;
assign w6363 = w368 & w372;
assign w6364 = w89 & w376;
assign w6365 = w47 & w385;
assign w6366 = w38 & w401;
assign w6367 = w47 & w407;
assign w6368 = w41 & w412;
assign w6369 = w60 & w423;
assign w6370 = ~w18 & w442;
assign w6371 = w368 & w86;
assign w6372 = ~w480 & pi0054;
assign w6373 = w512 & w6422;
assign w6374 = ~w18 & w516;
assign w6375 = w18 & ~pi0153;
assign w6376 = ~w18 & ~w442;
assign w6377 = w18 & ~pi0146;
assign w6378 = w18 & pi0172;
assign w6379 = w18 & pi0171;
assign w6380 = w18 & pi0170;
assign w6381 = w18 & pi0148;
assign w6382 = w18 & pi0169;
assign w6383 = w18 & pi0168;
assign w6384 = w18 & ~pi0166;
assign w6385 = w18 & ~pi0161;
assign w6386 = w18 & ~pi0152;
assign w6387 = w3 & ~pi0967;
assign w6388 = ~w3 & pi0947;
assign w6389 = w3 & pi0587;
assign w6390 = ~w462 & w6423;
assign w6391 = ~w462 & w6424;
assign w6392 = ~w462 & w6425;
assign w6393 = ~w462 & w6426;
assign w6394 = ~w462 & w6427;
assign w6395 = ~w462 & w6428;
assign w6396 = w244 & w6429;
assign w6397 = w244 & w6430;
assign w6398 = ~w868 & ~w859;
assign w6399 = ~w869 & ~w264;
assign w6400 = ~w934 & pi1191;
assign w6401 = ~w1021 & pi1192;
assign w6402 = w1155 & pi1190;
assign w6403 = w1195 & pi1193;
assign w6404 = (~w725 & w462) | (~w725 & w6431) | (w462 & w6431);
assign w6405 = ~w462 & w6432;
assign w6406 = ~w462 & w6433;
assign w6407 = ~w462 & w740;
assign w6408 = ~w869 & ~w1443;
assign w6409 = ~w3 & pi0219;
assign w6410 = w3 & pi0199;
assign w6411 = ~w462 & w6434;
assign w6412 = ~w462 & w6435;
assign w6413 = ~w462 & w6436;
assign w6414 = ~w462 & w6437;
assign w6415 = ~w462 & w6438;
assign w6416 = ~w462 & w6439;
assign w6417 = w378 & w1811;
assign w6418 = pi1087 & ~w1807;
assign w6419 = w435 & ~pi0841;
assign w6420 = w2011 & ~w265;
assign w6421 = ~pi0081 & w2842;
assign w6422 = ~w509 & ~pi0137;
assign w6423 = w747 & pi0160;
assign w6424 = w750 & pi0182;
assign w6425 = w747 & pi0158;
assign w6426 = w750 & pi0180;
assign w6427 = w747 & pi0159;
assign w6428 = w750 & pi0181;
assign w6429 = w452 & w863;
assign w6430 = w245 & pi0228;
assign w6431 = ~w860 & ~w725;
assign w6432 = w747 & pi0169;
assign w6433 = w750 & pi0191;
assign w6434 = w747 & pi0163;
assign w6435 = w750 & pi0184;
assign w6436 = w747 & pi0150;
assign w6437 = w750 & pi0185;
assign w6438 = w747 & pi0151;
assign w6439 = w750 & pi0173;
assign w6440 = w6376 & pi0239;
assign w6441 = w18 & ~pi0154;
assign w6442 = w6376 & pi0235;
assign w6443 = w18 & ~pi0151;
assign w6444 = w6376 & ~pi0238;
assign w6445 = w15 & pi0146;
assign w6446 = w15 & ~w6377;
assign w6447 = w6376 & ~pi0249;
assign w6448 = w15 & ~pi0172;
assign w6449 = w15 & ~w6378;
assign w6450 = w6370 & ~pi0861;
assign w6451 = w15 & ~pi0171;
assign w6452 = w15 & ~w6379;
assign w6453 = w6376 & ~pi0248;
assign w6454 = w15 & ~pi0170;
assign w6455 = w15 & ~w6380;
assign w6456 = w6376 & ~pi0247;
assign w6457 = w15 & ~pi0148;
assign w6458 = w15 & ~w6381;
assign w6459 = w6376 & ~pi0246;
assign w6460 = w15 & ~pi0169;
assign w6461 = w15 & ~w6382;
assign w6462 = w6376 & ~pi0240;
assign w6463 = w15 & ~pi0168;
assign w6464 = w15 & ~w6383;
assign w6465 = w6370 & ~pi0875;
assign w6466 = w15 & pi0166;
assign w6467 = w15 & ~w6384;
assign w6468 = w6376 & ~pi0244;
assign w6469 = w15 & pi0161;
assign w6470 = w15 & ~w6385;
assign w6471 = w6376 & ~pi0242;
assign w6472 = w15 & pi0152;
assign w6473 = w15 & ~w6386;
assign w6474 = ~w3 & ~pi0970;
assign w6475 = ~w3 & pi0907;
assign w6476 = w3 & pi0602;
assign w6477 = ~w112 & w378;
assign w6478 = w712 & pi1087;
assign w6479 = ~w711 & w525;
assign w6480 = ~w870 & ~w882;
assign w6481 = w1249 & ~w264;
assign w6482 = w1249 & ~w883;
assign w6483 = ~w1250 & w1251;
assign w6484 = w748 & pi0164;
assign w6485 = w751 & pi0186;
assign w6486 = ~w678 & ~w377;
assign w6487 = w748 & pi0167;
assign w6488 = w751 & pi0188;
assign w6489 = w6407 & ~w1356;
assign w6490 = w748 & pi0148;
assign w6491 = w751 & pi0141;
assign w6492 = w259 & ~w725;
assign w6493 = w259 & w6404;
assign w6494 = ~w870 & pi0228;
assign w6495 = ~pi0044 & ~w1443;
assign w6496 = ~pi0044 & ~w1435;
assign w6497 = w717 & ~w1443;
assign w6498 = w717 & ~w1435;
assign w6499 = w723 & ~w1443;
assign w6500 = w723 & ~w1435;
assign w6501 = w722 & ~w1443;
assign w6502 = w722 & ~w1435;
assign w6503 = w748 & pi0153;
assign w6504 = w751 & pi0175;
assign w6505 = w6407 & w1645;
assign w6506 = w1646 & ~w25;
assign w6507 = w748 & pi0147;
assign w6508 = w718 & ~w1443;
assign w6509 = w718 & ~w1435;
assign w6510 = w720 & ~w1443;
assign w6511 = w720 & ~w1435;
assign w6512 = w751 & pi0143;
assign w6513 = w6407 & ~w1331;
assign w6514 = ~w1791 & ~w1795;
assign w6515 = ~w3 & pi0221;
assign w6516 = w3 & pi0222;
assign w6517 = ~w3 & pi0215;
assign w6518 = w3 & pi0223;
assign w6519 = ~w3 & pi0216;
assign w6520 = w3 & pi0224;
assign w6521 = ~w3 & ~w16;
assign w6522 = ~pi0072 & pi0111;
assign w6523 = w71 & w136;
assign w6524 = w2 & w196;
assign w6525 = ~w3 & pi0146;
assign w6526 = w3 & pi0142;
assign w6527 = w28 & ~pi0094;
assign w6528 = w119 & w246;
assign w6529 = ~w250 & pi0129;
assign w6530 = ~w254 & pi0950;
assign w6531 = ~pi0111 & pi0072;
assign w6532 = w71 & w295;
assign w6533 = w55 & w299;
assign w6534 = w31 & w315;
assign w6535 = w71 & ~w371;
assign w6536 = w32 & ~pi0050;
assign w6537 = w6536 & w390;
assign w6538 = w119 & w391;
assign w6539 = w26 & w447;
assign w6540 = w119 & w453;
assign w6541 = w6536 & w460;
assign w6542 = ~w3 & pi0210;
assign w6543 = w3 & pi0198;
assign w6544 = ~pi0095 & pi0332;
assign w6545 = ~w235 & w240;
assign w6546 = w262 & pi1087;
assign w6547 = w262 & ~pi0841;
assign w6548 = ~w455 & w508;
assign w6549 = w441 & pi0234;
assign w6550 = ~w14 & ~pi0265;
assign w6551 = w14 & pi0833;
assign w6552 = ~w11 & pi1138;
assign w6553 = ~w14 & pi0276;
assign w6554 = ~w11 & pi1140;
assign w6555 = ~w14 & ~pi0274;
assign w6556 = ~w11 & pi1139;
assign w6557 = w6370 & pi0284;
assign w6558 = ~w14 & ~pi0264;
assign w6559 = ~w11 & pi1137;
assign w6560 = w6370 & pi0262;
assign w6561 = ~w14 & ~pi0277;
assign w6562 = ~w11 & pi1136;
assign w6563 = w6376 & ~pi0241;
assign w6564 = ~w14 & ~pi0270;
assign w6565 = ~w11 & pi1135;
assign w6566 = w6370 & ~pi0869;
assign w6567 = ~w14 & ~pi0282;
assign w6568 = ~w11 & pi1134;
assign w6569 = w6370 & ~pi0862;
assign w6570 = ~w14 & ~pi0281;
assign w6571 = ~w11 & pi1133;
assign w6572 = w6370 & ~pi0877;
assign w6573 = ~w14 & ~pi0269;
assign w6574 = ~w11 & pi1132;
assign w6575 = w6370 & ~pi0878;
assign w6576 = ~w14 & ~pi0280;
assign w6577 = ~w11 & pi1131;
assign w6578 = w6376 & ~pi0245;
assign w6579 = ~w14 & pi0266;
assign w6580 = ~w11 & pi1130;
assign w6581 = w6370 & ~pi0879;
assign w6582 = ~w14 & pi0279;
assign w6583 = ~w11 & pi1129;
assign w6584 = w6370 & ~pi0846;
assign w6585 = ~w14 & pi0278;
assign w6586 = ~w11 & pi1128;
assign w6587 = w524 & ~w14;
assign w6588 = w6587 & ~w503;
assign w6589 = ~pi0642 & pi0603;
assign w6590 = ~w680 & ~w701;
assign w6591 = ~pi0681 & pi0680;
assign w6592 = ~w680 & ~w709;
assign w6593 = w702 & w710;
assign w6594 = ~w714 & w350;
assign w6595 = ~pi0101 & ~pi0099;
assign w6596 = w719 & w721;
assign w6597 = ~pi0042 & w724;
assign w6598 = ~w725 & pi0683;
assign w6599 = ~w461 & w747;
assign w6600 = ~w461 & w750;
assign w6601 = ~w3 & pi0197;
assign w6602 = w3 & pi0145;
assign w6603 = ~w359 & ~w482;
assign w6604 = w668 & w778;
assign w6605 = w252 & w247;
assign w6606 = ~w783 & w727;
assign w6607 = w775 & w802;
assign w6608 = w803 & ~pi0228;
assign w6609 = ~w3 & ~pi0972;
assign w6610 = w3 & ~pi0961;
assign w6611 = ~w3 & ~pi0960;
assign w6612 = w3 & ~pi0977;
assign w6613 = ~w3 & ~pi0963;
assign w6614 = w3 & ~pi0969;
assign w6615 = ~w3 & ~pi0975;
assign w6616 = w3 & ~pi0971;
assign w6617 = ~w3 & ~pi0978;
assign w6618 = w3 & ~pi0974;
assign w6619 = ~w803 & ~pi0954;
assign w6620 = pi0119 & ~pi0468;
assign w6621 = ~pi0024 & w858;
assign w6622 = w235 & w740;
assign w6623 = ~w461 & w860;
assign w6624 = w119 & w6396;
assign w6625 = w119 & w6397;
assign w6626 = pi1087 & ~pi0122;
assign w6627 = w258 & ~w879;
assign w6628 = w886 & ~w264;
assign w6629 = w886 & ~w883;
assign w6630 = w1254 & ~w1258;
assign w6631 = pi0252 & w725;
assign w6632 = pi0252 & ~w6404;
assign w6633 = ~pi0024 & ~w263;
assign w6634 = ~w262 & ~w879;
assign w6635 = ~w1271 & w1270;
assign w6636 = ~pi0024 & ~pi0841;
assign w6637 = w771 & ~w14;
assign w6638 = ~w168 & w1279;
assign w6639 = ~w359 & ~w788;
assign w6640 = ~pi0040 & w40;
assign w6641 = w1291 & ~w1305;
assign w6642 = w1289 & w1306;
assign w6643 = ~w3 & pi0149;
assign w6644 = w3 & pi0183;
assign w6645 = w6407 & ~w1316;
assign w6646 = ~w1318 & ~w1307;
assign w6647 = w6407 & w235;
assign w6648 = w748 & pi0172;
assign w6649 = w751 & pi0193;
assign w6650 = ~w3 & pi0157;
assign w6651 = w3 & pi0178;
assign w6652 = w6407 & w1335;
assign w6653 = w1337 & ~w1324;
assign w6654 = w748 & pi0154;
assign w6655 = w751 & pi0176;
assign w6656 = w1294 & ~pi0034;
assign w6657 = w1291 & ~w1348;
assign w6658 = w1289 & w1352;
assign w6659 = w3 & pi0140;
assign w6660 = ~w1363 & ~w1353;
assign w6661 = w748 & pi0155;
assign w6662 = w751 & pi0177;
assign w6663 = w6407 & w231;
assign w6664 = w6407 & ~w1379;
assign w6665 = w6407 & w240;
assign w6666 = ~w1372 & ~w1322;
assign w6667 = ~w726 & pi0137;
assign w6668 = ~w6667 & ~w864;
assign w6669 = pi0683 & w1390;
assign w6670 = ~w1271 & ~w1270;
assign w6671 = w435 & pi0841;
assign w6672 = ~w1398 & ~w1399;
assign w6673 = ~w1397 & ~w1389;
assign w6674 = w278 & ~pi0841;
assign w6675 = pi1087 & ~pi0986;
assign w6676 = pi0252 & pi0986;
assign w6677 = pi0252 & ~w6675;
assign w6678 = ~w712 & w1419;
assign w6679 = w712 & ~w10;
assign w6680 = w1426 & ~pi0841;
assign w6681 = pi0101 & pi0041;
assign w6682 = w6407 & w228;
assign w6683 = ~w231 & w235;
assign w6684 = ~w6683 & w1451;
assign w6685 = ~w3 & pi0214;
assign w6686 = w3 & pi0207;
assign w6687 = ~w3 & pi0212;
assign w6688 = w3 & pi0208;
assign w6689 = ~w3 & pi0211;
assign w6690 = w3 & pi0200;
assign w6691 = w1451 & ~w1470;
assign w6692 = w1472 & w1447;
assign w6693 = w1457 & ~w1479;
assign w6694 = w1478 & ~w1481;
assign w6695 = w1451 & ~w1482;
assign w6696 = w861 & w1451;
assign w6697 = pi0044 & w1443;
assign w6698 = pi0044 & w1435;
assign w6699 = w484 & pi0024;
assign w6700 = pi1087 & ~w263;
assign w6701 = w6670 & ~w876;
assign w6702 = ~w278 & ~w291;
assign w6703 = ~pi0841 & ~w1504;
assign w6704 = w448 & ~pi0024;
assign w6705 = w262 & pi0252;
assign w6706 = ~pi0252 & ~w725;
assign w6707 = ~pi0252 & w6404;
assign w6708 = w1513 & w309;
assign w6709 = w1451 & w1478;
assign w6710 = w1521 & ~w1443;
assign w6711 = w1521 & ~w1435;
assign w6712 = pi0043 & w1523;
assign w6713 = pi0056 & w1504;
assign w6714 = pi0056 & ~w6703;
assign w6715 = w454 & pi0024;
assign w6716 = w472 & pi0024;
assign w6717 = ~w668 & w667;
assign w6718 = pi0841 & pi0061;
assign w6719 = w465 & ~pi0024;
assign w6720 = w484 & ~pi0024;
assign w6721 = pi0064 & w1504;
assign w6722 = pi0064 & ~w6703;
assign w6723 = pi0081 & pi0314;
assign w6724 = w668 & w522;
assign w6725 = w113 & w1576;
assign w6726 = ~w665 & ~pi0593;
assign w6727 = pi0589 & w1585;
assign w6728 = w15 & w1586;
assign w6729 = ~w6728 & ~pi0287;
assign w6730 = pi0081 & w1468;
assign w6731 = w258 & pi1087;
assign w6732 = w149 & w1594;
assign w6733 = w771 & w14;
assign w6734 = w448 & pi0024;
assign w6735 = ~w262 & ~pi0841;
assign w6736 = w1604 & ~pi0479;
assign w6737 = ~w1606 & w1499;
assign w6738 = ~w783 & ~w727;
assign w6739 = pi0252 & ~w725;
assign w6740 = pi0252 & w6404;
assign w6741 = ~w1612 & ~w1539;
assign w6742 = w1614 & w725;
assign w6743 = w1614 & ~w6404;
assign w6744 = w138 & ~pi0314;
assign w6745 = w1496 & pi0077;
assign w6746 = w748 & pi0156;
assign w6747 = w751 & pi0179;
assign w6748 = w1279 & w1322;
assign w6749 = ~w1635 & ~w1282;
assign w6750 = ~w1333 & ~w1374;
assign w6751 = w1291 & w25;
assign w6752 = ~w6656 & pi0079;
assign w6753 = pi0079 & w40;
assign w6754 = w1652 & w1292;
assign w6755 = w751 & pi0187;
assign w6756 = ~w6507 & ~w1289;
assign w6757 = w1654 & w1651;
assign w6758 = ~w1658 & w1640;
assign w6759 = w1254 & ~pi0080;
assign w6760 = pi0081 & ~pi0314;
assign w6761 = w157 & ~pi0314;
assign w6762 = w149 & ~pi1087;
assign w6763 = w147 & w879;
assign w6764 = pi0841 & pi0089;
assign w6765 = pi0090 & w1504;
assign w6766 = pi0090 & ~w6703;
assign w6767 = w364 & ~w1695;
assign w6768 = ~w678 & ~w1600;
assign w6769 = w777 & ~w1581;
assign w6770 = w345 & w1706;
assign w6771 = w1604 & pi0479;
assign w6772 = w1711 & pi0096;
assign w6773 = pi0589 & pi0593;
assign w6774 = w777 & w1717;
assign w6775 = w1724 & w1447;
assign w6776 = ~w231 & w1726;
assign w6777 = pi0314 & ~w6676;
assign w6778 = pi0314 & ~w6677;
assign w6779 = ~w252 & w247;
assign w6780 = ~w1612 & w1732;
assign w6781 = ~pi0024 & w263;
assign w6782 = w147 & w880;
assign w6783 = w370 & pi0314;
assign w6784 = pi0115 & pi0114;
assign w6785 = pi0113 & pi0116;
assign w6786 = pi0079 & pi0118;
assign w6787 = w1282 & ~w1778;
assign w6788 = ~w1290 & w1784;
assign w6789 = w748 & pi0165;
assign w6790 = ~w6512 & ~w1289;
assign w6791 = w748 & pi0168;
assign w6792 = w751 & pi0190;
assign w6793 = w6514 & ~w1785;
assign w6794 = ~w711 & ~w1807;
assign w6795 = w1694 & ~w1808;
assign w6796 = ~w6417 & ~pi0228;
assign w6797 = w1254 & w1817;
assign w6798 = w1816 & pi1087;
assign w6799 = ~w369 & ~pi0024;
assign w6800 = ~pi0121 & ~pi0126;
assign w6801 = ~pi0132 & ~pi0130;
assign w6802 = w6801 & ~pi0136;
assign w6803 = ~pi0135 & ~pi0134;
assign w6804 = w1837 & w1829;
assign w6805 = w1829 & w1839;
assign w6806 = ~pi0087 & w1825;
assign w6807 = ~w1824 & w1847;
assign w6808 = ~w263 & w1854;
assign w6809 = ~w6808 & pi0039;
assign w6810 = w169 & ~w1857;
assign w6811 = w87 & ~w1859;
assign w6812 = w1858 & w71;
assign w6813 = ~w162 & w155;
assign w6814 = w1866 & ~w155;
assign w6815 = w1866 & ~w6813;
assign w6816 = w1856 & w1870;
assign w6817 = w6407 & ~w757;
assign w6818 = w1847 & w1884;
assign w6819 = ~w1835 & ~w1887;
assign w6820 = ~w6803 & w1832;
assign w6821 = pi0121 & pi0126;
assign w6822 = w1847 & ~w1903;
assign w6823 = ~w1845 & ~w678;
assign w6824 = w450 & w437;
assign w6825 = ~w350 & ~w392;
assign w6826 = ~pi0250 & pi0127;
assign w6827 = pi0250 & ~w265;
assign w6828 = w485 & pi0129;
assign w6829 = w247 & ~pi0250;
assign w6830 = ~w265 & ~pi0250;
assign w6831 = ~w265 & w6829;
assign w6832 = ~pi0129 & ~w455;
assign w6833 = pi0132 & pi0130;
assign w6834 = ~w1835 & ~w1934;
assign w6835 = ~w6803 & ~pi0133;
assign w6836 = w1847 & ~w1957;
assign w6837 = w751 & pi0192;
assign w6838 = w748 & pi0171;
assign w6839 = pi0135 & pi0134;
assign w6840 = ~pi0135 & pi0134;
assign w6841 = ~pi0135 & w1829;
assign w6842 = w748 & pi0170;
assign w6843 = w1976 & ~w1829;
assign w6844 = w1847 & w1980;
assign w6845 = ~w6801 & pi0136;
assign w6846 = ~w1835 & ~w1986;
assign w6847 = w861 & w1992;
assign w6848 = w1296 & ~pi0139;
assign w6849 = ~w6848 & pi0138;
assign w6850 = w6848 & ~pi0138;
assign w6851 = w1282 & ~w1998;
assign w6852 = ~w1296 & pi0139;
assign w6853 = w1282 & ~w2003;
assign w6854 = pi0287 & pi0120;
assign w6855 = ~w1584 & ~pi0287;
assign w6856 = w2007 & w350;
assign w6857 = w1416 & pi0252;
assign w6858 = ~w495 & w2015;
assign w6859 = w2017 & ~w1595;
assign w6860 = ~pi0832 & ~w2010;
assign w6861 = ~w1254 & ~pi0140;
assign w6862 = w2026 & pi0603;
assign w6863 = w2060 & ~w2024;
assign w6864 = w2069 & pi0680;
assign w6865 = w2103 & ~w2067;
assign w6866 = ~w1254 & ~pi0141;
assign w6867 = ~w1254 & pi0142;
assign w6868 = ~w1254 & ~pi0143;
assign w6869 = ~w1254 & pi0144;
assign w6870 = ~w1254 & ~pi0145;
assign w6871 = ~w1254 & pi0146;
assign w6872 = pi0743 & pi0947;
assign w6873 = ~w1254 & ~pi0147;
assign w6874 = ~pi0770 & pi0947;
assign w6875 = ~w1254 & ~pi0148;
assign w6876 = pi0749 & pi0947;
assign w6877 = ~w1254 & ~pi0149;
assign w6878 = ~pi0755 & pi0947;
assign w6879 = ~w1254 & ~pi0150;
assign w6880 = ~pi0751 & pi0947;
assign w6881 = ~w1254 & ~pi0151;
assign w6882 = ~pi0745 & pi0947;
assign w6883 = ~w1254 & pi0152;
assign w6884 = pi0759 & pi0947;
assign w6885 = ~w1254 & ~pi0153;
assign w6886 = pi0766 & pi0947;
assign w6887 = ~w1254 & ~pi0154;
assign w6888 = ~pi0742 & pi0947;
assign w6889 = ~w1254 & ~pi0155;
assign w6890 = ~pi0757 & pi0947;
assign w6891 = ~w1254 & ~pi0156;
assign w6892 = ~pi0741 & pi0947;
assign w6893 = ~w1254 & ~pi0157;
assign w6894 = ~pi0760 & pi0947;
assign w6895 = ~w1254 & ~pi0158;
assign w6896 = ~pi0753 & pi0947;
assign w6897 = ~w1254 & ~pi0159;
assign w6898 = ~pi0754 & pi0947;
assign w6899 = ~w1254 & ~pi0160;
assign w6900 = ~pi0756 & pi0947;
assign w6901 = ~w1254 & pi0161;
assign w6902 = pi0758 & pi0947;
assign w6903 = ~w1254 & ~pi0162;
assign w6904 = ~pi0761 & pi0947;
assign w6905 = ~w1254 & ~pi0163;
assign w6906 = ~pi0777 & pi0947;
assign w6907 = ~w1254 & ~pi0164;
assign w6908 = ~pi0752 & pi0947;
assign w6909 = ~w1254 & ~pi0165;
assign w6910 = ~pi0774 & pi0947;
assign w6911 = ~w1254 & pi0166;
assign w6912 = pi0772 & pi0947;
assign w6913 = ~w1254 & ~pi0167;
assign w6914 = ~pi0768 & pi0947;
assign w6915 = ~w1254 & ~pi0168;
assign w6916 = pi0763 & pi0947;
assign w6917 = ~w1254 & ~pi0169;
assign w6918 = pi0746 & pi0947;
assign w6919 = ~w1254 & ~pi0170;
assign w6920 = pi0748 & pi0947;
assign w6921 = ~w1254 & ~pi0171;
assign w6922 = pi0764 & pi0947;
assign w6923 = ~w1254 & ~pi0172;
assign w6924 = pi0739 & pi0947;
assign w6925 = ~w1254 & ~pi0173;
assign w6926 = ~w1254 & pi0174;
assign w6927 = ~w1254 & ~pi0175;
assign w6928 = ~w1254 & ~pi0176;
assign w6929 = ~w1254 & ~pi0177;
assign w6930 = ~w1254 & ~pi0178;
assign w6931 = ~w1254 & ~pi0179;
assign w6932 = ~w1254 & ~pi0180;
assign w6933 = ~w1254 & ~pi0181;
assign w6934 = ~w1254 & ~pi0182;
assign w6935 = ~w1254 & ~pi0183;
assign w6936 = ~w1254 & ~pi0184;
assign w6937 = ~w1254 & ~pi0185;
assign w6938 = ~w1254 & ~pi0186;
assign w6939 = ~w1254 & ~pi0187;
assign w6940 = ~w1254 & ~pi0188;
assign w6941 = ~w1254 & pi0189;
assign w6942 = ~w1254 & ~pi0190;
assign w6943 = ~w1254 & ~pi0191;
assign w6944 = ~w1254 & ~pi0192;
assign w6945 = ~w1254 & ~pi0193;
assign w6946 = ~w1254 & ~pi0194;
assign w6947 = w6850 & ~pi0196;
assign w6948 = w1282 & w2496;
assign w6949 = ~w6850 & pi0196;
assign w6950 = w1282 & ~w2500;
assign w6951 = ~w1254 & ~pi0197;
assign w6952 = w2010 & w1254;
assign w6953 = w702 & ~pi0332;
assign w6954 = ~pi0841 & w2542;
assign w6955 = ~w6954 & ~w2541;
assign w6956 = ~pi0201 & ~pi0332;
assign w6957 = ~pi0201 & w6953;
assign w6958 = ~w2545 & w6956;
assign w6959 = ~w2545 & w6957;
assign w6960 = ~pi0202 & ~pi0332;
assign w6961 = ~pi0202 & w6953;
assign w6962 = ~w2550 & w6960;
assign w6963 = ~w2550 & w6961;
assign w6964 = ~pi0203 & ~pi0332;
assign w6965 = ~pi0203 & w6953;
assign w6966 = ~w2555 & w6964;
assign w6967 = ~w2555 & w6965;
assign w6968 = w710 & ~pi0332;
assign w6969 = ~pi0204 & ~pi0332;
assign w6970 = ~pi0204 & w6968;
assign w6971 = ~w2561 & w6969;
assign w6972 = ~w2561 & w6970;
assign w6973 = ~pi0205 & ~pi0332;
assign w6974 = ~pi0205 & w6968;
assign w6975 = ~w2565 & w6973;
assign w6976 = ~w2565 & w6974;
assign w6977 = ~pi0206 & ~pi0332;
assign w6978 = ~pi0206 & w6968;
assign w6979 = ~w2570 & w6977;
assign w6980 = ~w2570 & w6978;
assign w6981 = ~pi0218 & ~pi0332;
assign w6982 = ~pi0218 & w6968;
assign w6983 = ~pi0220 & ~pi0332;
assign w6984 = ~pi0220 & w6953;
assign w6985 = w6824 & w458;
assign w6986 = ~w459 & ~w497;
assign w6987 = ~w2685 & ~pi0228;
assign w6988 = ~w262 & ~w253;
assign w6989 = ~w777 & w208;
assign w6990 = w775 & ~w1421;
assign w6991 = ~w3 & pi0213;
assign w6992 = w3 & pi0209;
assign w6993 = ~w1478 & pi1137;
assign w6994 = ~w2719 & w2709;
assign w6995 = w2734 & w2712;
assign w6996 = ~w2711 & w2737;
assign w6997 = w2741 & ~w2736;
assign w6998 = ~w1463 & ~w2731;
assign w6999 = ~w1478 & pi1147;
assign w7000 = w2752 & w2737;
assign w7001 = ~w2709 & ~w2745;
assign w7002 = ~w1478 & pi1148;
assign w7003 = ~w2762 & w2737;
assign w7004 = w2734 & w2711;
assign w7005 = ~w1478 & pi1138;
assign w7006 = ~w2776 & w2709;
assign w7007 = w2782 & w2712;
assign w7008 = ~w1464 & w2737;
assign w7009 = ~w2762 & ~w2739;
assign w7010 = ~w1478 & pi1146;
assign w7011 = w2796 & w2737;
assign w7012 = ~w2709 & ~w2801;
assign w7013 = ~w1478 & pi1140;
assign w7014 = w2809 & w2737;
assign w7015 = ~w1478 & pi1142;
assign w7016 = w2815 & w2709;
assign w7017 = w2796 & w2709;
assign w7018 = ~w1478 & pi1144;
assign w7019 = w2825 & w2737;
assign w7020 = ~w1478 & pi1139;
assign w7021 = w2835 & w2709;
assign w7022 = w2719 & w2737;
assign w7023 = pi0314 & ~w2842;
assign w7024 = pi0314 & ~w6421;
assign w7025 = pi0802 & pi0276;
assign w7026 = w7025 & pi0271;
assign w7027 = w7026 & pi0273;
assign w7028 = w7027 & pi0283;
assign w7029 = w7028 & pi0272;
assign w7030 = pi0275 & pi0268;
assign w7031 = pi0267 & ~pi0263;
assign w7032 = w7030 & w2852;
assign w7033 = ~w7032 & w2853;
assign w7034 = pi0243 & w2853;
assign w7035 = pi0243 & w7033;
assign w7036 = w7032 & w2856;
assign w7037 = ~pi1149 & ~w2853;
assign w7038 = w2809 & w2709;
assign w7039 = w2835 & w2737;
assign w7040 = ~w1478 & pi1141;
assign w7041 = w2873 & w2709;
assign w7042 = ~w1478 & pi1143;
assign w7043 = w2882 & w2709;
assign w7044 = w2873 & w2737;
assign w7045 = w2815 & w2737;
assign w7046 = w2882 & w2737;
assign w7047 = ~w1478 & pi1145;
assign w7048 = w2898 & w2709;
assign w7049 = w2898 & w2737;
assign w7050 = ~pi0476 & pi1033;
assign w7051 = pi0897 & pi1047;
assign w7052 = pi1157 & pi1087;
assign w7053 = w7030 & pi0253;
assign w7054 = ~w7030 & ~pi0253;
assign w7055 = ~pi1147 & ~w2853;
assign w7056 = ~w7053 & ~pi0254;
assign w7057 = w7030 & w2850;
assign w7058 = ~w7057 & w2853;
assign w7059 = w2938 & ~w2853;
assign w7060 = pi0897 & pi1043;
assign w7061 = ~pi0476 & pi1030;
assign w7062 = pi0897 & pi1042;
assign w7063 = ~pi0476 & pi1064;
assign w7064 = ~pi0476 & pi1059;
assign w7065 = pi0897 & pi1078;
assign w7066 = ~pi0476 & pi1056;
assign w7067 = pi0897 & pi1066;
assign w7068 = ~pi0476 & pi1063;
assign w7069 = pi0897 & pi1053;
assign w7070 = pi0897 & pi1038;
assign w7071 = ~pi0476 & pi1061;
assign w7072 = ~pi0476 & pi1034;
assign w7073 = pi0897 & pi1031;
assign w7074 = w7030 & w2851;
assign w7075 = ~w7074 & pi0263;
assign w7076 = w2781 & ~w2853;
assign w7077 = w2853 & ~w7023;
assign w7078 = w2853 & ~w7024;
assign w7079 = w2853 & w7023;
assign w7080 = w2853 & w7024;
assign w7081 = ~pi1137 & ~w2853;
assign w7082 = ~w2996 & ~w2991;
assign w7083 = ~pi1138 & ~w2853;
assign w7084 = ~w3004 & ~w3000;
assign w7085 = ~pi1130 & ~w2853;
assign w7086 = ~w3012 & ~w3008;
assign w7087 = ~w7057 & ~pi0267;
assign w7088 = w2793 & ~w2853;
assign w7089 = ~pi0275 & ~pi0268;
assign w7090 = ~pi1144 & ~w2853;
assign w7091 = ~pi1132 & ~w2853;
assign w7092 = ~w3035 & ~w3031;
assign w7093 = ~pi1135 & ~w2853;
assign w7094 = ~w3043 & ~w3039;
assign w7095 = ~w7025 & ~pi0271;
assign w7096 = ~pi1139 & ~w2853;
assign w7097 = ~w7028 & ~pi0272;
assign w7098 = ~pi1142 & ~w2853;
assign w7099 = w3066 & ~w2853;
assign w7100 = ~w7027 & w2853;
assign w7101 = ~w3078 & ~w3073;
assign w7102 = ~pi1143 & ~w2853;
assign w7103 = ~pi0802 & ~pi0276;
assign w7104 = ~pi1136 & ~w2853;
assign w7105 = ~w3104 & ~w3100;
assign w7106 = ~pi1127 & ~w2853;
assign w7107 = ~w3112 & ~w3108;
assign w7108 = ~pi1129 & ~w2853;
assign w7109 = ~w3120 & ~w3116;
assign w7110 = ~pi1131 & ~w2853;
assign w7111 = ~w3128 & ~w3124;
assign w7112 = ~pi1133 & ~w2853;
assign w7113 = ~w3136 & ~w3132;
assign w7114 = ~pi1134 & ~w2853;
assign w7115 = ~w3144 & ~w3140;
assign w7116 = ~w7027 & ~pi0283;
assign w7117 = ~pi1141 & ~w2853;
assign w7118 = w882 & w877;
assign w7119 = w7118 & ~pi0289;
assign w7120 = ~w882 & w3164;
assign w7121 = w7120 & pi0289;
assign w7122 = ~w882 & ~w3173;
assign w7123 = w882 & w3173;
assign w7124 = ~w7122 & ~pi0793;
assign w7125 = ~pi0288 & ~pi0793;
assign w7126 = pi0289 & ~pi0793;
assign w7127 = w6719 & ~pi0312;
assign w7128 = w7127 & ~pi0300;
assign w7129 = ~w7128 & ~pi0055;
assign w7130 = ~w7127 & pi0300;
assign w7131 = ~pi0301 & ~pi0055;
assign w7132 = ~pi0301 & w7129;
assign w7133 = w7128 & pi0301;
assign w7134 = ~w14 & pi0273;
assign w7135 = ~w11 & pi1142;
assign w7136 = w14 & ~pi0237;
assign w7137 = ~w14 & pi0271;
assign w7138 = ~w11 & pi1141;
assign w7139 = w14 & ~pi0233;
assign w7140 = ~w7133 & pi0311;
assign w7141 = ~w7133 & ~pi0055;
assign w7142 = ~w6719 & w3264;
assign one = 1;
assign po0000 = pi0668;// level 0
assign po0001 = pi0672;// level 0
assign po0002 = pi0664;// level 0
assign po0003 = pi0667;// level 0
assign po0004 = pi0676;// level 0
assign po0005 = pi0673;// level 0
assign po0006 = pi0675;// level 0
assign po0007 = pi0666;// level 0
assign po0008 = pi0679;// level 0
assign po0009 = pi0674;// level 0
assign po0010 = pi0663;// level 0
assign po0011 = pi0670;// level 0
assign po0012 = pi0677;// level 0
assign po0013 = pi0682;// level 0
assign po0014 = pi0671;// level 0
assign po0015 = pi0678;// level 0
assign po0016 = pi0718;// level 0
assign po0017 = pi0707;// level 0
assign po0018 = pi0708;// level 0
assign po0019 = pi0713;// level 0
assign po0020 = pi0711;// level 0
assign po0021 = pi0716;// level 0
assign po0022 = pi0733;// level 0
assign po0023 = pi0712;// level 0
assign po0024 = pi0689;// level 0
assign po0025 = pi0717;// level 0
assign po0026 = pi0692;// level 0
assign po0027 = pi0719;// level 0
assign po0028 = pi0722;// level 0
assign po0029 = pi0714;// level 0
assign po0030 = pi0720;// level 0
assign po0031 = pi0685;// level 0
assign po0032 = pi0837;// level 0
assign po0033 = pi0850;// level 0
assign po0034 = pi0872;// level 0
assign po0035 = pi0871;// level 0
assign po0036 = pi0881;// level 0
assign po0037 = pi0866;// level 0
assign po0038 = pi0876;// level 0
assign po0039 = pi0873;// level 0
assign po0040 = pi0874;// level 0
assign po0041 = pi0859;// level 0
assign po0042 = pi0855;// level 0
assign po0043 = pi0852;// level 0
assign po0044 = pi0870;// level 0
assign po0045 = pi0848;// level 0
assign po0046 = pi0865;// level 0
assign po0047 = pi0856;// level 0
assign po0048 = pi0853;// level 0
assign po0049 = pi0847;// level 0
assign po0050 = pi0857;// level 0
assign po0051 = pi0854;// level 0
assign po0052 = pi0858;// level 0
assign po0053 = pi0845;// level 0
assign po0054 = pi0838;// level 0
assign po0055 = pi0842;// level 0
assign po0056 = pi0843;// level 0
assign po0057 = pi0839;// level 0
assign po0058 = pi0844;// level 0
assign po0059 = pi0868;// level 0
assign po0060 = pi0851;// level 0
assign po0061 = pi0867;// level 0
assign po0062 = pi0880;// level 0
assign po0063 = pi0860;// level 0
assign po0064 = pi1024;// level 0
assign po0065 = pi1028;// level 0
assign po0066 = pi1009;// level 0
assign po0067 = pi1014;// level 0
assign po0068 = pi1019;// level 0
assign po0069 = pi0999;// level 0
assign po0070 = pi0990;// level 0
assign po0071 = pi1006;// level 0
assign po0072 = pi0987;// level 0
assign po0073 = pi1010;// level 0
assign po0074 = pi1015;// level 0
assign po0075 = pi1004;// level 0
assign po0076 = pi1021;// level 0
assign po0077 = pi1012;// level 0
assign po0078 = pi1011;// level 0
assign po0079 = pi1018;// level 0
assign po0080 = pi1003;// level 0
assign po0081 = pi1026;// level 0
assign po0082 = pi0997;// level 0
assign po0083 = pi0991;// level 0
assign po0084 = pi1007;// level 0
assign po0085 = pi1005;// level 0
assign po0086 = pi1002;// level 0
assign po0087 = pi1013;// level 0
assign po0088 = pi1025;// level 0
assign po0089 = pi1016;// level 0
assign po0090 = pi0994;// level 0
assign po0091 = pi1017;// level 0
assign po0092 = pi0996;// level 0
assign po0093 = pi1020;// level 0
assign po0094 = pi1000;// level 0
assign po0095 = pi0992;// level 0
assign po0096 = pi0031;// level 0
assign po0097 = pi0080;// level 0
assign po0098 = pi0893;// level 0
assign po0099 = pi0467;// level 0
assign po0100 = pi0078;// level 0
assign po0101 = pi0112;// level 0
assign po0102 = pi0013;// level 0
assign po0103 = pi0025;// level 0
assign po0104 = pi0226;// level 0
assign po0105 = pi0127;// level 0
assign po0106 = pi0822;// level 0
assign po0107 = pi0808;// level 0
assign po0108 = pi0227;// level 0
assign po0109 = pi0477;// level 0
assign po0110 = pi0834;// level 0
assign po0111 = pi0229;// level 0
assign po0112 = pi0012;// level 0
assign po0113 = pi0011;// level 0
assign po0114 = pi0010;// level 0
assign po0115 = pi0009;// level 0
assign po0116 = pi0008;// level 0
assign po0117 = pi0007;// level 0
assign po0118 = pi0006;// level 0
assign po0119 = pi0005;// level 0
assign po0120 = pi0004;// level 0
assign po0121 = pi0003;// level 0
assign po0122 = pi0000;// level 0
assign po0123 = pi0002;// level 0
assign po0124 = pi0001;// level 0
assign po0125 = pi0310;// level 0
assign po0126 = pi0302;// level 0
assign po0127 = pi0475;// level 0
assign po0128 = pi0474;// level 0
assign po0129 = pi0466;// level 0
assign po0130 = pi0473;// level 0
assign po0131 = pi0471;// level 0
assign po0132 = pi0472;// level 0
assign po0133 = pi0470;// level 0
assign po0134 = pi0469;// level 0
assign po0135 = pi0465;// level 0
assign po0136 = pi1022;// level 0
assign po0137 = pi1027;// level 0
assign po0138 = pi0989;// level 0
assign po0139 = pi0988;// level 0
assign po0140 = pi0028;// level 0
assign po0141 = pi0027;// level 0
assign po0142 = pi0026;// level 0
assign po0143 = pi0029;// level 0
assign po0144 = pi0015;// level 0
assign po0145 = pi0014;// level 0
assign po0146 = pi0021;// level 0
assign po0147 = pi0020;// level 0
assign po0148 = pi0019;// level 0
assign po0149 = pi0018;// level 0
assign po0150 = pi0017;// level 0
assign po0151 = pi0016;// level 0
assign po0152 = pi1090;// level 0
assign po0153 = ~w533;// level 19
assign po0154 = ~w543;// level 18
assign po0155 = ~w553;// level 18
assign po0156 = ~w564;// level 18
assign po0157 = ~w575;// level 18
assign po0158 = ~w586;// level 18
assign po0159 = ~w597;// level 18
assign po0160 = ~w608;// level 18
assign po0161 = ~w619;// level 18
assign po0162 = ~w630;// level 18
assign po0163 = ~w641;// level 18
assign po0164 = ~w652;// level 18
assign po0165 = ~w663;// level 18
assign po0166 = one;// level 0
assign po0167 = ~w739;// level 15
assign po0168 = pi0228;// level 0
assign po0169 = pi0022;// level 0
assign po0170 = ~pi1084;// level 0
assign po0171 = ~w808;// level 17
assign po0172 = ~w810;// level 17
assign po0173 = ~w814;// level 17
assign po0174 = ~w819;// level 17
assign po0175 = ~w824;// level 17
assign po0176 = ~w829;// level 17
assign po0177 = ~w834;// level 17
assign po0178 = ~w839;// level 17
assign po0179 = pi1083;// level 0
assign po0180 = pi0023;// level 0
assign po0181 = ~w739;// level 15
assign po0182 = ~w842;// level 17
assign po0183 = ~w846;// level 16
assign po0184 = ~w850;// level 3
assign po0185 = ~w852;// level 3
assign po0186 = ~w854;// level 3
assign po0187 = ~w856;// level 3
assign po0188 = pi0037;// level 0
assign po0189 = ~w1260;// level 18
assign po0190 = ~w1277;// level 15
assign po0191 = w1344;// level 18
assign po0192 = w1388;// level 18
assign po0193 = ~w1410;// level 15
assign po0194 = w1412;// level 10
assign po0195 = ~w804;// level 16
assign po0196 = ~w1415;// level 10
assign po0197 = ~w1431;// level 12
assign po0198 = ~w1434;// level 9
assign po0199 = w1454;// level 17
assign po0200 = ~w1476;// level 17
assign po0201 = ~w1488;// level 18
assign po0202 = ~w1493;// level 17
assign po0203 = w1495;// level 8
assign po0204 = ~w1498;// level 9
assign po0205 = ~w1503;// level 10
assign po0206 = w1508;// level 12
assign po0207 = ~w1511;// level 9
assign po0208 = ~w1519;// level 13
assign po0209 = w382;// level 7
assign po0210 = ~w1526;// level 16
assign po0211 = ~w1530;// level 9
assign po0212 = ~w1533;// level 10
assign po0213 = ~w1535;// level 9
assign po0214 = ~w1538;// level 12
assign po0215 = ~w1544;// level 11
assign po0216 = w1278;// level 8
assign po0217 = ~w1548;// level 9
assign po0218 = ~w1551;// level 9
assign po0219 = ~w1557;// level 11
assign po0220 = ~w1560;// level 9
assign po0221 = ~w1563;// level 9
assign po0222 = ~w1565;// level 12
assign po0223 = w1566;// level 9
assign po0224 = w1568;// level 9
assign po0225 = w1572;// level 8
assign po0226 = w1574;// level 10
assign po0227 = ~w1579;// level 9
assign po0228 = ~w1589;// level 11
assign po0229 = w1593;// level 10
assign po0230 = ~w1599;// level 11
assign po0231 = w1602;// level 12
assign po0232 = ~w1609;// level 10
assign po0233 = ~w1621;// level 17
assign po0234 = ~w1625;// level 12
assign po0235 = ~w1628;// level 11
assign po0236 = w1630;// level 2
assign po0237 = w1665;// level 17
assign po0238 = w1668;// level 17
assign po0239 = ~w1670;// level 9
assign po0240 = ~w1674;// level 9
assign po0241 = ~w1677;// level 9
assign po0242 = w1678;// level 9
assign po0243 = ~w1680;// level 9
assign po0244 = w1681;// level 10
assign po0245 = w1682;// level 8
assign po0246 = w1686;// level 10
assign po0247 = ~w1689;// level 11
assign po0248 = ~w1692;// level 12
assign po0249 = ~w1697;// level 10
assign po0250 = w1699;// level 11
assign po0251 = ~w1701;// level 9
assign po0252 = ~w1703;// level 13
assign po0253 = ~w1709;// level 11
assign po0254 = ~w1713;// level 12
assign po0255 = ~w1719;// level 11
assign po0256 = w1722;// level 9
assign po0257 = ~w1728;// level 17
assign po0258 = ~w1737;// level 17
assign po0259 = ~w1743;// level 18
assign po0260 = w1744;// level 8
assign po0261 = ~w1745;// level 9
assign po0262 = ~w1748;// level 13
assign po0263 = pi0117;// level 0
assign po0264 = ~w1751;// level 9
assign po0265 = w1752;// level 8
assign po0266 = ~w1753;// level 10
assign po0267 = w1754;// level 8
assign po0268 = ~w1756;// level 13
assign po0269 = ~w1759;// level 11
assign po0270 = ~w1760;// level 1
assign po0271 = w1764;// level 17
assign po0272 = w1769;// level 17
assign po0273 = w1772;// level 17
assign po0274 = w1775;// level 17
assign po0275 = ~w844;// level 14
assign po0276 = ~w1805;// level 17
assign po0277 = ~w1814;// level 17
assign po0278 = w1822;// level 15
assign po0279 = w1852;// level 17
assign po0280 = w884;// level 14
assign po0281 = ~w1873;// level 14
assign po0282 = ~w1894;// level 17
assign po0283 = w1911;// level 16
assign po0284 = w1923;// level 16
assign po0285 = pi0131;// level 0
assign po0286 = w1930;// level 16
assign po0287 = ~w1939;// level 16
assign po0288 = ~w1812;// level 16
assign po0289 = ~w1953;// level 16
assign po0290 = ~w1962;// level 15
assign po0291 = ~w1971;// level 15
assign po0292 = ~w1983;// level 15
assign po0293 = ~w1990;// level 15
assign po0294 = ~w1994;// level 12
assign po0295 = ~w2001;// level 14
assign po0296 = ~w2006;// level 14
assign po0297 = ~w2113;// level 15
assign po0298 = ~w2121;// level 15
assign po0299 = ~w2129;// level 15
assign po0300 = ~w2137;// level 15
assign po0301 = ~w2145;// level 15
assign po0302 = ~w2153;// level 15
assign po0303 = ~w2161;// level 15
assign po0304 = ~w2168;// level 15
assign po0305 = ~w2174;// level 15
assign po0306 = ~w2181;// level 15
assign po0307 = ~w2188;// level 15
assign po0308 = ~w2195;// level 15
assign po0309 = ~w2202;// level 15
assign po0310 = ~w2209;// level 15
assign po0311 = ~w2216;// level 15
assign po0312 = ~w2223;// level 15
assign po0313 = ~w2230;// level 15
assign po0314 = ~w2237;// level 15
assign po0315 = ~w2244;// level 15
assign po0316 = ~w2251;// level 15
assign po0317 = ~w2258;// level 15
assign po0318 = ~w2264;// level 15
assign po0319 = ~w2270;// level 15
assign po0320 = ~w2277;// level 15
assign po0321 = ~w2284;// level 15
assign po0322 = ~w2290;// level 15
assign po0323 = ~w2297;// level 15
assign po0324 = ~w2304;// level 15
assign po0325 = ~w2311;// level 15
assign po0326 = ~w2318;// level 15
assign po0327 = ~w2325;// level 15
assign po0328 = ~w2332;// level 15
assign po0329 = ~w2339;// level 15
assign po0330 = ~w2346;// level 15
assign po0331 = ~w2353;// level 15
assign po0332 = ~w2360;// level 15
assign po0333 = ~w2367;// level 15
assign po0334 = ~w2374;// level 15
assign po0335 = ~w2381;// level 15
assign po0336 = ~w2388;// level 15
assign po0337 = ~w2395;// level 15
assign po0338 = ~w2402;// level 15
assign po0339 = ~w2409;// level 15
assign po0340 = ~w2416;// level 15
assign po0341 = ~w2423;// level 15
assign po0342 = ~w2430;// level 15
assign po0343 = ~w2437;// level 15
assign po0344 = ~w2444;// level 15
assign po0345 = ~w2451;// level 15
assign po0346 = ~w2458;// level 15
assign po0347 = ~w2465;// level 15
assign po0348 = ~w2472;// level 15
assign po0349 = ~w2479;// level 15
assign po0350 = ~w2486;// level 15
assign po0351 = ~w2493;// level 15
assign po0352 = ~w2498;// level 14
assign po0353 = ~w2503;// level 15
assign po0354 = ~w2509;// level 15
assign po0355 = ~w2517;// level 15
assign po0356 = ~w2523;// level 15
assign po0357 = ~w2529;// level 15
assign po0358 = ~w2547;// level 10
assign po0359 = ~w2552;// level 10
assign po0360 = ~w2557;// level 10
assign po0361 = ~w2563;// level 10
assign po0362 = ~w2567;// level 10
assign po0363 = ~w2572;// level 10
assign po0364 = ~w2578;// level 15
assign po0365 = ~w2584;// level 15
assign po0366 = ~w2590;// level 15
assign po0367 = ~w2596;// level 15
assign po0368 = ~w2602;// level 15
assign po0369 = w2608;// level 15
assign po0370 = w2614;// level 15
assign po0371 = w2620;// level 15
assign po0372 = ~w2626;// level 15
assign po0373 = ~w2632;// level 15
assign po0374 = ~w2638;// level 15
assign po0375 = ~w2643;// level 11
assign po0376 = ~w2649;// level 15
assign po0377 = ~w2654;// level 11
assign po0378 = ~w2660;// level 15
assign po0379 = ~w2666;// level 15
assign po0380 = ~w2672;// level 15
assign po0381 = ~w2678;// level 15
assign po0382 = ~w514;// level 15
assign po0383 = ~w2688;// level 15
assign po0384 = w2693;// level 11
assign po0385 = ~w2698;// level 12
assign po0386 = pi0232;// level 0
assign po0387 = ~w2510;// level 13
assign po0388 = pi0236;// level 0
assign po0389 = ~w2704;// level 14
assign po0390 = w2744;// level 12
assign po0391 = ~w2757;// level 12
assign po0392 = w2771;// level 12
assign po0393 = ~w2686;// level 14
assign po0394 = w2789;// level 12
assign po0395 = ~w2800;// level 12
assign po0396 = ~w2805;// level 10
assign po0397 = ~w2820;// level 12
assign po0398 = ~w2831;// level 12
assign po0399 = ~w2841;// level 12
assign po0400 = w2863;// level 10
assign po0401 = ~w2868;// level 12
assign po0402 = ~w2878;// level 12
assign po0403 = ~w2888;// level 12
assign po0404 = ~w2893;// level 12
assign po0405 = ~w2903;// level 12
assign po0406 = ~w2908;// level 12
assign po0407 = w2910;// level 10
assign po0408 = ~w2920;// level 5
assign po0409 = ~w2925;// level 10
assign po0410 = w2934;// level 10
assign po0411 = ~w2941;// level 9
assign po0412 = ~w2946;// level 5
assign po0413 = ~w2951;// level 5
assign po0414 = ~w2956;// level 5
assign po0415 = ~w2961;// level 5
assign po0416 = ~w2966;// level 5
assign po0417 = ~w2971;// level 5
assign po0418 = ~w2976;// level 5
assign po0419 = ~w2983;// level 9
assign po0420 = ~w2989;// level 9
assign po0421 = w2999;// level 9
assign po0422 = w3007;// level 9
assign po0423 = w3015;// level 9
assign po0424 = ~w3021;// level 10
assign po0425 = w3030;// level 10
assign po0426 = w3038;// level 9
assign po0427 = w3046;// level 9
assign po0428 = w3055;// level 9
assign po0429 = w3064;// level 9
assign po0430 = ~w3072;// level 9
assign po0431 = w3081;// level 9
assign po0432 = w3090;// level 10
assign po0433 = w3099;// level 9
assign po0434 = w3107;// level 9
assign po0435 = w3115;// level 9
assign po0436 = w3123;// level 9
assign po0437 = w3131;// level 9
assign po0438 = w3139;// level 9
assign po0439 = w3147;// level 9
assign po0440 = w3156;// level 9
assign po0441 = ~w3160;// level 9
assign po0442 = w3172;// level 13
assign po0443 = w3179;// level 13
assign po0444 = w3181;// level 2
assign po0445 = w3184;// level 13
assign po0446 = w3188;// level 13
assign po0447 = ~w3191;// level 2
assign po0448 = ~w3194;// level 2
assign po0449 = ~w3197;// level 2
assign po0450 = ~w3200;// level 2
assign po0451 = ~w3203;// level 2
assign po0452 = ~w3206;// level 2
assign po0453 = ~w3209;// level 2
assign po0454 = ~w3212;// level 2
assign po0455 = ~w3215;// level 2
assign po0456 = ~w3217;// level 9
assign po0457 = ~w3221;// level 9
assign po0458 = ~w3224;// level 9
assign po0459 = ~w3231;// level 9
assign po0460 = ~w3234;// level 2
assign po0461 = ~w3237;// level 2
assign po0462 = ~w3240;// level 2
assign po0463 = ~w3243;// level 2
assign po0464 = ~w3246;// level 2
assign po0465 = ~w3249;// level 2
assign po0466 = ~w3252;// level 2
assign po0467 = ~w3259;// level 9
assign po0468 = w3263;// level 10
assign po0469 = ~w3266;// level 9
assign po0470 = w3271;// level 14
assign po0471 = w3274;// level 11
assign po0472 = ~w3278;// level 12
assign po0473 = ~w3281;// level 12
assign po0474 = ~w3285;// level 12
assign po0475 = ~w3289;// level 12
assign po0476 = ~w3292;// level 12
assign po0477 = ~w3295;// level 12
assign po0478 = ~w3298;// level 12
assign po0479 = ~w3301;// level 12
assign po0480 = ~w3304;// level 12
assign po0481 = ~w3307;// level 12
assign po0482 = ~w3310;// level 12
assign po0483 = ~w3313;// level 12
assign po0484 = ~w3316;// level 12
assign po0485 = ~w3319;// level 12
assign po0486 = ~w3322;// level 12
assign po0487 = w3326;// level 12
assign po0488 = w3329;// level 12
assign po0489 = ~w1313;// level 11
assign po0490 = ~w3332;// level 12
assign po0491 = ~w3335;// level 12
assign po0492 = ~w3338;// level 12
assign po0493 = ~w3341;// level 12
assign po0494 = ~w3344;// level 12
assign po0495 = ~w3347;// level 12
assign po0496 = ~w3350;// level 12
assign po0497 = ~w3354;// level 12
assign po0498 = w3357;// level 12
assign po0499 = ~w3360;// level 12
assign po0500 = ~w3363;// level 12
assign po0501 = ~w3366;// level 12
assign po0502 = ~w3369;// level 12
assign po0503 = ~w3372;// level 12
assign po0504 = ~w3375;// level 12
assign po0505 = ~w3378;// level 12
assign po0506 = ~w3381;// level 12
assign po0507 = ~w3384;// level 12
assign po0508 = ~w3387;// level 12
assign po0509 = ~w3390;// level 12
assign po0510 = ~w3393;// level 12
assign po0511 = ~w3396;// level 12
assign po0512 = ~w3399;// level 12
assign po0513 = ~w3402;// level 12
assign po0514 = ~w3405;// level 12
assign po0515 = ~w3408;// level 12
assign po0516 = ~w3411;// level 12
assign po0517 = ~w3414;// level 12
assign po0518 = ~w3417;// level 12
assign po0519 = ~w3420;// level 12
assign po0520 = ~w3423;// level 12
assign po0521 = ~w3426;// level 12
assign po0522 = ~w3429;// level 12
assign po0523 = ~w3432;// level 12
assign po0524 = ~w3435;// level 12
assign po0525 = ~w3438;// level 12
assign po0526 = ~w3441;// level 12
assign po0527 = ~w3444;// level 12
assign po0528 = ~w3447;// level 12
assign po0529 = ~w3450;// level 12
assign po0530 = ~w3453;// level 12
assign po0531 = ~w3456;// level 12
assign po0532 = ~w3459;// level 12
assign po0533 = ~w3462;// level 12
assign po0534 = ~w3465;// level 12
assign po0535 = ~w3468;// level 12
assign po0536 = ~w3471;// level 12
assign po0537 = ~w3474;// level 12
assign po0538 = ~w3477;// level 12
assign po0539 = ~w3480;// level 12
assign po0540 = ~w3483;// level 12
assign po0541 = ~w3486;// level 12
assign po0542 = ~w3489;// level 12
assign po0543 = ~w3492;// level 12
assign po0544 = ~w3495;// level 12
assign po0545 = ~w3498;// level 12
assign po0546 = ~w3501;// level 12
assign po0547 = ~w3504;// level 12
assign po0548 = ~w3507;// level 12
assign po0549 = ~w3510;// level 12
assign po0550 = ~w3513;// level 12
assign po0551 = ~w3516;// level 12
assign po0552 = ~w3519;// level 12
assign po0553 = ~w3522;// level 12
assign po0554 = ~w3525;// level 12
assign po0555 = ~w3528;// level 12
assign po0556 = ~w3531;// level 12
assign po0557 = ~w3534;// level 12
assign po0558 = ~w3537;// level 12
assign po0559 = ~w3540;// level 12
assign po0560 = ~w3543;// level 12
assign po0561 = ~w3546;// level 12
assign po0562 = ~w3549;// level 12
assign po0563 = ~w3552;// level 12
assign po0564 = ~w3555;// level 12
assign po0565 = ~w3558;// level 12
assign po0566 = ~w3561;// level 12
assign po0567 = ~w3564;// level 12
assign po0568 = ~w3567;// level 12
assign po0569 = ~w3570;// level 12
assign po0570 = ~w3573;// level 12
assign po0571 = ~w3576;// level 12
assign po0572 = ~w3579;// level 12
assign po0573 = ~w3582;// level 12
assign po0574 = ~w3585;// level 12
assign po0575 = ~w3588;// level 12
assign po0576 = ~w3591;// level 12
assign po0577 = ~w3594;// level 12
assign po0578 = ~w3597;// level 12
assign po0579 = ~w3600;// level 12
assign po0580 = ~w3603;// level 12
assign po0581 = ~w3606;// level 12
assign po0582 = ~w3609;// level 12
assign po0583 = ~w3612;// level 12
assign po0584 = ~w3615;// level 12
assign po0585 = ~w3618;// level 12
assign po0586 = ~w3621;// level 12
assign po0587 = ~w3624;// level 12
assign po0588 = ~w3627;// level 12
assign po0589 = ~w3630;// level 12
assign po0590 = ~w3633;// level 12
assign po0591 = ~w3636;// level 12
assign po0592 = ~w3639;// level 12
assign po0593 = ~w3642;// level 12
assign po0594 = ~w3645;// level 12
assign po0595 = ~w3648;// level 12
assign po0596 = ~w3651;// level 12
assign po0597 = ~w3654;// level 12
assign po0598 = ~w3657;// level 12
assign po0599 = ~w3660;// level 12
assign po0600 = ~w3663;// level 12
assign po0601 = ~w3666;// level 12
assign po0602 = ~w3669;// level 12
assign po0603 = ~w3672;// level 12
assign po0604 = ~w3675;// level 12
assign po0605 = ~w3678;// level 12
assign po0606 = ~w3681;// level 12
assign po0607 = ~w3684;// level 12
assign po0608 = ~w3687;// level 12
assign po0609 = ~w3690;// level 12
assign po0610 = ~w3693;// level 12
assign po0611 = ~w3696;// level 12
assign po0612 = ~w3699;// level 12
assign po0613 = ~w3702;// level 12
assign po0614 = w3721;// level 6
assign po0615 = ~w3724;// level 12
assign po0616 = ~w3727;// level 12
assign po0617 = ~w3730;// level 12
assign po0618 = ~w3733;// level 12
assign po0619 = ~w3736;// level 12
assign po0620 = ~w3739;// level 12
assign po0621 = ~w3742;// level 12
assign po0622 = ~w3747;// level 9
assign po0623 = ~w3752;// level 9
assign po0624 = ~w3758;// level 8
assign po0625 = ~w3761;// level 11
assign po0626 = ~w3766;// level 9
assign po0627 = ~w3771;// level 9
assign po0628 = ~w3776;// level 9
assign po0629 = ~w3781;// level 9
assign po0630 = ~w3786;// level 9
assign po0631 = ~w3791;// level 9
assign po0632 = ~w3796;// level 9
assign po0633 = ~w3798;// level 9
assign po0634 = ~w3269;// level 12
assign po0635 = w3799;// level 6
assign po0636 = pi0583;// level 0
assign po0637 = ~w1442;// level 9
assign po0638 = ~w3802;// level 9
assign po0639 = ~w3805;// level 9
assign po0640 = ~w3808;// level 9
assign po0641 = ~w3811;// level 9
assign po0642 = ~w3814;// level 9
assign po0643 = ~w3817;// level 9
assign po0644 = ~w3820;// level 9
assign po0645 = w3823;// level 9
assign po0646 = ~w3826;// level 9
assign po0647 = ~w3829;// level 9
assign po0648 = ~w3832;// level 9
assign po0649 = ~w3835;// level 9
assign po0650 = ~w3838;// level 9
assign po0651 = w3841;// level 9
assign po0652 = ~w3844;// level 9
assign po0653 = ~w3847;// level 9
assign po0654 = w3850;// level 9
assign po0655 = ~w3853;// level 9
assign po0656 = ~w3856;// level 9
assign po0657 = ~w3859;// level 9
assign po0658 = ~w3862;// level 9
assign po0659 = ~w3865;// level 9
assign po0660 = ~w3868;// level 9
assign po0661 = ~w3871;// level 9
assign po0662 = ~w3874;// level 9
assign po0663 = ~w3877;// level 9
assign po0664 = ~w3880;// level 9
assign po0665 = ~w3883;// level 9
assign po0666 = ~w3886;// level 9
assign po0667 = ~w3889;// level 9
assign po0668 = ~w3892;// level 9
assign po0669 = ~w3895;// level 9
assign po0670 = ~w3898;// level 9
assign po0671 = ~w3901;// level 9
assign po0672 = ~w3904;// level 9
assign po0673 = ~w3907;// level 9
assign po0674 = ~w3910;// level 9
assign po0675 = ~w3913;// level 9
assign po0676 = w3916;// level 9
assign po0677 = ~w3919;// level 9
assign po0678 = ~w3922;// level 9
assign po0679 = ~w3925;// level 9
assign po0680 = ~w3928;// level 9
assign po0681 = w3931;// level 9
assign po0682 = ~w3934;// level 9
assign po0683 = ~w3937;// level 9
assign po0684 = ~w3940;// level 9
assign po0685 = ~w3943;// level 9
assign po0686 = ~w3946;// level 9
assign po0687 = ~w3949;// level 9
assign po0688 = ~w3952;// level 9
assign po0689 = ~w3955;// level 9
assign po0690 = ~w3958;// level 9
assign po0691 = w3961;// level 9
assign po0692 = ~w3964;// level 9
assign po0693 = ~w3967;// level 9
assign po0694 = ~w3970;// level 9
assign po0695 = ~w3973;// level 9
assign po0696 = ~w3976;// level 9
assign po0697 = ~w3979;// level 9
assign po0698 = ~w3982;// level 9
assign po0699 = ~w3985;// level 9
assign po0700 = ~w3988;// level 9
assign po0701 = ~w3991;// level 9
assign po0702 = ~w3994;// level 9
assign po0703 = ~w3997;// level 9
assign po0704 = ~w4000;// level 9
assign po0705 = ~w4003;// level 9
assign po0706 = ~w4006;// level 9
assign po0707 = w4009;// level 9
assign po0708 = ~w4012;// level 9
assign po0709 = ~w4015;// level 9
assign po0710 = ~w4018;// level 9
assign po0711 = ~w4021;// level 9
assign po0712 = ~w4024;// level 9
assign po0713 = ~w4027;// level 9
assign po0714 = ~w4030;// level 9
assign po0715 = ~w4033;// level 9
assign po0716 = ~w4036;// level 9
assign po0717 = ~w4039;// level 9
assign po0718 = ~w4042;// level 9
assign po0719 = ~w4045;// level 9
assign po0720 = ~w4048;// level 9
assign po0721 = ~w4051;// level 9
assign po0722 = ~w4054;// level 9
assign po0723 = ~w4057;// level 9
assign po0724 = ~w4067;// level 11
assign po0725 = ~w4070;// level 9
assign po0726 = w4073;// level 9
assign po0727 = ~w4076;// level 9
assign po0728 = ~w4079;// level 9
assign po0729 = ~w4082;// level 9
assign po0730 = ~w4085;// level 9
assign po0731 = ~w4088;// level 9
assign po0732 = ~w4091;// level 9
assign po0733 = ~w4094;// level 9
assign po0734 = ~w4097;// level 9
assign po0735 = ~w4100;// level 9
assign po0736 = ~w4103;// level 9
assign po0737 = ~w4106;// level 9
assign po0738 = ~w4109;// level 9
assign po0739 = ~w4112;// level 9
assign po0740 = w265;// level 6
assign po0741 = ~w4115;// level 9
assign po0742 = ~w4118;// level 9
assign po0743 = ~w4121;// level 9
assign po0744 = w4124;// level 9
assign po0745 = ~w4130;// level 8
assign po0746 = ~w4147;// level 7
assign po0747 = w4150;// level 8
assign po0748 = ~w4153;// level 8
assign po0749 = ~w4156;// level 8
assign po0750 = ~w4581;// level 10
assign po0751 = w4588;// level 6
assign po0752 = w4593;// level 6
assign po0753 = w4597;// level 7
assign po0754 = w4600;// level 6
assign po0755 = ~w4607;// level 7
assign po0756 = w4611;// level 8
assign po0757 = w4614;// level 5
assign po0758 = w4617;// level 4
assign po0759 = w4620;// level 9
assign po0760 = ~w4634;// level 8
assign po0761 = ~w4641;// level 5
assign po0762 = w4644;// level 3
assign po0763 = ~w4649;// level 8
assign po0764 = ~w4652;// level 7
assign po0765 = ~w4655;// level 7
assign po0766 = ~w4658;// level 7
assign po0767 = ~w4661;// level 7
assign po0768 = ~w4664;// level 7
assign po0769 = ~w4667;// level 7
assign po0770 = ~w4670;// level 7
assign po0771 = ~w4674;// level 8
assign po0772 = ~w4679;// level 7
assign po0773 = ~w4683;// level 8
assign po0774 = ~w4688;// level 8
assign po0775 = ~w4691;// level 7
assign po0776 = ~w4694;// level 7
assign po0777 = ~w4697;// level 7
assign po0778 = ~w4700;// level 7
assign po0779 = ~w4703;// level 7
assign po0780 = ~w4706;// level 7
assign po0781 = ~w4712;// level 5
assign po0782 = ~w4722;// level 7
assign po0783 = ~w4725;// level 7
assign po0784 = ~w4728;// level 7
assign po0785 = ~w4731;// level 7
assign po0786 = ~w4734;// level 7
assign po0787 = ~w4737;// level 7
assign po0788 = ~w4740;// level 7
assign po0789 = ~w4743;// level 7
assign po0790 = ~w4746;// level 7
assign po0791 = ~w4749;// level 7
assign po0792 = ~w4752;// level 7
assign po0793 = ~w4755;// level 7
assign po0794 = ~w4758;// level 7
assign po0795 = ~w4761;// level 7
assign po0796 = ~w4764;// level 7
assign po0797 = ~w4767;// level 7
assign po0798 = ~w4770;// level 7
assign po0799 = ~w4773;// level 7
assign po0800 = ~w4776;// level 7
assign po0801 = ~w4779;// level 7
assign po0802 = ~w4782;// level 7
assign po0803 = ~w4785;// level 7
assign po0804 = ~w4788;// level 7
assign po0805 = ~w4791;// level 7
assign po0806 = ~w4794;// level 7
assign po0807 = ~w4797;// level 7
assign po0808 = ~w4800;// level 7
assign po0809 = ~w4803;// level 7
assign po0810 = ~w4806;// level 7
assign po0811 = ~w4809;// level 7
assign po0812 = ~w4812;// level 7
assign po0813 = ~w4815;// level 7
assign po0814 = ~w4818;// level 7
assign po0815 = ~w4821;// level 7
assign po0816 = w4834;// level 12
assign po0817 = ~w4837;// level 7
assign po0818 = ~w4840;// level 7
assign po0819 = ~w4843;// level 7
assign po0820 = ~w4882;// level 10
assign po0821 = ~w4901;// level 10
assign po0822 = ~w4904;// level 7
assign po0823 = ~w4923;// level 10
assign po0824 = ~w4942;// level 10
assign po0825 = ~w4961;// level 10
assign po0826 = ~w4964;// level 7
assign po0827 = ~w4979;// level 9
assign po0828 = ~w4994;// level 9
assign po0829 = ~w5013;// level 10
assign po0830 = ~w5032;// level 10
assign po0831 = ~w5051;// level 10
assign po0832 = ~w5070;// level 10
assign po0833 = ~w5089;// level 10
assign po0834 = ~w5104;// level 9
assign po0835 = ~w5119;// level 9
assign po0836 = ~w5138;// level 10
assign po0837 = ~w5141;// level 7
assign po0838 = ~w5144;// level 7
assign po0839 = ~w5159;// level 9
assign po0840 = w263;// level 4
assign po0841 = ~w5165;// level 7
assign po0842 = ~w5186;// level 10
assign po0843 = ~w5189;// level 7
assign po0844 = ~w5192;// level 7
assign po0845 = ~w5195;// level 7
assign po0846 = ~w5214;// level 10
assign po0847 = ~w5217;// level 7
assign po0848 = ~w5220;// level 7
assign po0849 = ~w5239;// level 10
assign po0850 = ~w5242;// level 7
assign po0851 = ~w5245;// level 7
assign po0852 = ~w5248;// level 7
assign po0853 = ~w5251;// level 7
assign po0854 = ~w5254;// level 7
assign po0855 = ~w5257;// level 7
assign po0856 = ~w5260;// level 7
assign po0857 = ~w5263;// level 7
assign po0858 = ~w5266;// level 7
assign po0859 = ~w5269;// level 7
assign po0860 = ~w5272;// level 7
assign po0861 = ~w5275;// level 7
assign po0862 = ~w5278;// level 7
assign po0863 = ~w5281;// level 7
assign po0864 = ~w5298;// level 10
assign po0865 = ~w5315;// level 10
assign po0866 = ~w5318;// level 7
assign po0867 = ~w5321;// level 7
assign po0868 = ~w5338;// level 10
assign po0869 = ~w5355;// level 10
assign po0870 = ~w5372;// level 10
assign po0871 = ~w5391;// level 10
assign po0872 = ~w5394;// level 7
assign po0873 = ~w5411;// level 10
assign po0874 = ~w5430;// level 10
assign po0875 = ~w5447;// level 10
assign po0876 = ~w5466;// level 10
assign po0877 = ~w5485;// level 10
assign po0878 = w5535;// level 10
assign po0879 = ~w5554;// level 10
assign po0880 = ~w5557;// level 7
assign po0881 = ~w5560;// level 7
assign po0882 = ~w5563;// level 7
assign po0883 = ~w5566;// level 7
assign po0884 = ~w5569;// level 7
assign po0885 = ~w5572;// level 7
assign po0886 = ~w5575;// level 7
assign po0887 = ~w5578;// level 7
assign po0888 = w5581;// level 7
assign po0889 = ~w5584;// level 7
assign po0890 = ~w5601;// level 10
assign po0891 = ~w5604;// level 7
assign po0892 = ~w5607;// level 7
assign po0893 = ~w5610;// level 7
assign po0894 = ~w5613;// level 7
assign po0895 = ~w5616;// level 7
assign po0896 = ~w5621;// level 7
assign po0897 = w4625;// level 4
assign po0898 = ~w5625;// level 7
assign po0899 = ~w5629;// level 7
assign po0900 = ~w5633;// level 7
assign po0901 = ~w5637;// level 7
assign po0902 = ~w5641;// level 7
assign po0903 = ~w5645;// level 7
assign po0904 = w5648;// level 7
assign po0905 = ~w5652;// level 7
assign po0906 = ~w5656;// level 7
assign po0907 = ~w5660;// level 7
assign po0908 = ~w5664;// level 7
assign po0909 = ~w5668;// level 7
assign po0910 = ~w5672;// level 7
assign po0911 = ~w5676;// level 7
assign po0912 = ~w5680;// level 7
assign po0913 = ~w5684;// level 7
assign po0914 = ~w5688;// level 7
assign po0915 = ~w5692;// level 7
assign po0916 = ~w5696;// level 7
assign po0917 = ~w5700;// level 7
assign po0918 = ~w5704;// level 7
assign po0919 = ~w5708;// level 7
assign po0920 = ~w5712;// level 7
assign po0921 = ~w5716;// level 7
assign po0922 = w5719;// level 7
assign po0923 = ~w5723;// level 7
assign po0924 = ~w5727;// level 7
assign po0925 = ~w5731;// level 7
assign po0926 = w5734;// level 9
assign po0927 = ~w5738;// level 7
assign po0928 = w5741;// level 7
assign po0929 = ~w5745;// level 7
assign po0930 = w5748;// level 7
assign po0931 = ~w5752;// level 7
assign po0932 = w5755;// level 8
assign po0933 = ~w5759;// level 7
assign po0934 = ~w5763;// level 7
assign po0935 = ~w5771;// level 6
assign po0936 = ~w5772;// level 6
assign po0937 = ~w5773;// level 6
assign po0938 = ~w5776;// level 6
assign po0939 = ~w5778;// level 5
assign po0940 = ~w5781;// level 6
assign po0941 = ~w5784;// level 6
assign po0942 = ~w5787;// level 6
assign po0943 = w5790;// level 2
assign po0944 = ~w5793;// level 6
assign po0945 = ~w5796;// level 6
assign po0946 = ~w5799;// level 6
assign po0947 = ~w5802;// level 6
assign po0948 = ~w5805;// level 6
assign po0949 = ~w5808;// level 6
assign po0950 = w264;// level 5
assign po0951 = ~w5812;// level 6
assign po0952 = ~w5815;// level 6
assign po0953 = w5817;// level 10
assign po0954 = w4717;// level 4
assign po0955 = ~w5820;// level 6
assign po0956 = w5823;// level 6
assign po0957 = ~w5826;// level 6
assign po0958 = ~w5829;// level 6
assign po0959 = w4833;// level 11
assign po0960 = w5832;// level 6
assign po0961 = ~w5835;// level 6
assign po0962 = w5837;// level 8
assign po0963 = w5524;// level 6
assign po0964 = ~w5840;// level 6
assign po0965 = ~w5843;// level 6
assign po0966 = w5846;// level 6
assign po0967 = ~w5849;// level 6
assign po0968 = ~w5852;// level 6
assign po0969 = w5855;// level 6
assign po0970 = ~w5858;// level 6
assign po0971 = w5861;// level 6
assign po0972 = ~w5864;// level 6
assign po0973 = ~w5867;// level 6
assign po0974 = w5869;// level 5
assign po0975 = ~w1819;// level 4
assign po0976 = w5871;// level 11
assign po0977 = w5873;// level 9
assign po0978 = w5516;// level 5
assign po0979 = w5874;// level 1
assign po0980 = w5160;// level 4
assign po0981 = w5878;// level 6
assign po0982 = ~w5904;// level 10
assign po0983 = ~w5928;// level 10
assign po0984 = ~w5952;// level 10
assign po0985 = ~w5976;// level 10
assign po0986 = ~w5979;// level 4
assign po0987 = w5981;// level 6
assign po0988 = w5617;// level 4
assign po0989 = w5983;// level 4
assign po0990 = ~w5985;// level 3
assign po0991 = w5986;// level 2
assign po0992 = w5988;// level 7
assign po0993 = ~w5991;// level 2
assign po0994 = ~w5994;// level 2
assign po0995 = ~w5997;// level 2
assign po0996 = ~w6000;// level 3
assign po0997 = w1301;// level 3
assign po0998 = ~w6003;// level 2
assign po0999 = ~w6006;// level 2
assign po1000 = ~w6009;// level 2
assign po1001 = ~w6012;// level 2
assign po1002 = ~w6015;// level 4
assign po1003 = ~w6018;// level 2
assign po1004 = ~w6021;// level 2
assign po1005 = ~w6024;// level 3
assign po1006 = ~w6027;// level 2
assign po1007 = ~w6030;// level 2
assign po1008 = ~w6033;// level 2
assign po1009 = ~w6036;// level 2
assign po1010 = ~w6039;// level 2
assign po1011 = ~w6042;// level 2
assign po1012 = ~w6045;// level 2
assign po1013 = ~w6048;// level 2
assign po1014 = ~w6051;// level 2
assign po1015 = ~w6054;// level 2
assign po1016 = ~w6057;// level 2
assign po1017 = ~w6060;// level 4
assign po1018 = ~w6063;// level 4
assign po1019 = ~w6066;// level 3
assign po1020 = ~w6069;// level 3
assign po1021 = ~w6072;// level 2
assign po1022 = ~w6075;// level 2
assign po1023 = ~w6078;// level 2
assign po1024 = ~w6081;// level 2
assign po1025 = ~w6084;// level 4
assign po1026 = ~w6087;// level 2
assign po1027 = ~w6090;// level 2
assign po1028 = ~w6093;// level 2
assign po1029 = ~w6096;// level 2
assign po1030 = ~w6099;// level 2
assign po1031 = ~w6102;// level 4
assign po1032 = ~w6105;// level 2
assign po1033 = ~w6108;// level 4
assign po1034 = ~w6111;// level 4
assign po1035 = ~w6114;// level 4
assign po1036 = ~w6117;// level 2
assign po1037 = ~w6120;// level 2
assign po1038 = ~w4601;// level 3
assign po1039 = ~w6123;// level 4
assign po1040 = ~w6126;// level 4
assign po1041 = ~w6129;// level 4
assign po1042 = ~w6132;// level 4
assign po1043 = ~w6135;// level 4
assign po1044 = ~w6138;// level 4
assign po1045 = ~w6141;// level 4
assign po1046 = ~w6144;// level 4
assign po1047 = ~w6147;// level 4
assign po1048 = ~w6150;// level 4
assign po1049 = ~w41;// level 2
assign po1050 = ~w6153;// level 4
assign po1051 = ~w6156;// level 4
assign po1052 = ~w6159;// level 4
assign po1053 = pi0067;// level 0
assign po1054 = ~w6162;// level 4
assign po1055 = ~w6165;// level 4
assign po1056 = ~w6168;// level 4
assign po1057 = ~w725;// level 4
assign po1058 = ~w6171;// level 4
assign po1059 = ~w6174;// level 4
assign po1060 = ~w6177;// level 4
assign po1061 = ~w6180;// level 4
assign po1062 = ~w6183;// level 4
assign po1063 = ~w6193;// level 5
assign po1064 = ~w6196;// level 4
assign po1065 = ~w6199;// level 4
assign po1066 = ~w6202;// level 4
assign po1067 = ~w6205;// level 4
assign po1068 = ~w6208;// level 4
assign po1069 = ~w6211;// level 4
assign po1070 = w6213;// level 4
assign po1071 = ~w6216;// level 4
assign po1072 = ~w6219;// level 4
assign po1073 = ~w6222;// level 4
assign po1074 = ~w6225;// level 4
assign po1075 = ~w6228;// level 4
assign po1076 = ~w6231;// level 2
assign po1077 = ~w6234;// level 2
assign po1078 = ~w6237;// level 2
assign po1079 = ~w6240;// level 2
assign po1080 = w6243;// level 2
assign po1081 = ~w6246;// level 2
assign po1082 = ~w6249;// level 2
assign po1083 = ~w6252;// level 2
assign po1084 = ~w6255;// level 2
assign po1085 = ~w6258;// level 2
assign po1086 = ~w6261;// level 2
assign po1087 = ~w6264;// level 2
assign po1088 = ~w6267;// level 2
assign po1089 = ~w6270;// level 2
assign po1090 = ~w6273;// level 2
assign po1091 = ~w6276;// level 2
assign po1092 = ~w6279;// level 2
assign po1093 = ~w6282;// level 2
assign po1094 = ~w6285;// level 2
assign po1095 = ~w6288;// level 2
assign po1096 = ~w6291;// level 2
assign po1097 = ~w6294;// level 2
assign po1098 = ~w6297;// level 2
assign po1099 = ~w6300;// level 2
assign po1100 = ~w6303;// level 2
assign po1101 = ~w6304;// level 3
assign po1102 = w4058;// level 2
assign po1103 = w6306;// level 4
assign po1104 = w6308;// level 3
assign po1105 = w6311;// level 2
assign po1106 = w256;// level 3
assign po1107 = w262;// level 2
assign po1108 = pi1128;// level 0
assign po1109 = pi0964;// level 0
assign po1110 = ~pi0954;// level 0
assign po1111 = pi0965;// level 0
assign po1112 = ~w6312;// level 2
assign po1113 = w6314;// level 2
assign po1114 = pi0985;// level 0
assign po1115 = w6315;// level 1
assign po1116 = w6316;// level 1
assign po1117 = pi1008;// level 0
assign po1118 = w6317;// level 1
assign po1119 = pi1023;// level 0
assign po1120 = pi0998;// level 0
assign po1121 = pi1001;// level 0
assign po1122 = w6318;// level 1
assign po1123 = pi1129;// level 0
assign po1124 = w6319;// level 1
assign po1125 = w6320;// level 1
assign po1126 = w6321;// level 1
assign po1127 = w6322;// level 1
assign po1128 = w6323;// level 1
assign po1129 = w6324;// level 1
assign po1130 = ~pi0278;// level 0
assign po1131 = w6325;// level 1
assign po1132 = w6326;// level 1
assign po1133 = ~w6327;// level 1
assign po1134 = pi1058;// level 0
assign po1135 = w258;// level 1
assign po1136 = pi0299;// level 0
assign po1137 = ~w6328;// level 1
assign po1138 = pi1069;// level 0
assign po1139 = pi1046;// level 0
assign po1140 = ~pi0915;// level 0
assign po1141 = ~pi0825;// level 0
assign po1142 = ~pi0826;// level 0
assign po1143 = ~pi0913;// level 0
assign po1144 = ~pi0894;// level 0
assign po1145 = ~pi0905;// level 0
assign po1146 = pi1089;// level 0
assign po1147 = ~pi0890;// level 0
assign po1148 = pi1088;// level 0
assign po1149 = ~pi0906;// level 0
assign po1150 = ~pi0896;// level 0
assign po1151 = ~pi0909;// level 0
assign po1152 = ~pi0911;// level 0
assign po1153 = ~pi0908;// level 0
assign po1154 = ~pi0891;// level 0
assign po1155 = ~pi0902;// level 0
assign po1156 = ~pi0903;// level 0
assign po1157 = ~pi0883;// level 0
assign po1158 = ~pi0888;// level 0
assign po1159 = ~pi0919;// level 0
assign po1160 = ~pi0886;// level 0
assign po1161 = ~pi0912;// level 0
assign po1162 = ~pi0895;// level 0
assign po1163 = ~pi0916;// level 0
assign po1164 = ~pi0889;// level 0
assign po1165 = ~pi0900;// level 0
assign po1166 = ~pi0885;// level 0
assign po1167 = ~pi0904;// level 0
assign po1168 = ~pi0899;// level 0
assign po1169 = ~pi0918;// level 0
assign po1170 = ~pi0898;// level 0
assign po1171 = ~pi0917;// level 0
assign po1172 = ~pi0827;// level 0
assign po1173 = ~pi0887;// level 0
assign po1174 = ~pi0884;// level 0
assign po1175 = ~pi0910;// level 0
assign po1176 = ~pi0828;// level 0
assign po1177 = ~pi0892;// level 0
assign po1178 = pi1181;// level 0
assign po1179 = pi1166;// level 0
assign po1180 = pi1164;// level 0
assign po1181 = pi1132;// level 0
assign po1182 = pi1171;// level 0
assign po1183 = pi1172;// level 0
assign po1184 = pi0863;// level 0
assign po1185 = pi1197;// level 0
assign po1186 = pi1179;// level 0
assign po1187 = pi1165;// level 0
assign po1188 = pi1186;// level 0
assign po1189 = pi1131;// level 0
assign po1190 = pi1180;// level 0
assign po1191 = pi1159;// level 0
assign po1192 = pi1158;// level 0
assign po1193 = pi1092;// level 0
assign po1194 = pi1177;// level 0
assign po1195 = pi0230;// level 0
assign po1196 = pi1163;// level 0
assign po1197 = pi1130;// level 0
assign po1198 = pi1175;// level 0
assign po1199 = pi0849;// level 0
assign po1200 = pi1187;// level 0
assign po1201 = pi1176;// level 0
assign po1202 = pi1162;// level 0
assign po1203 = pi1169;// level 0
assign po1204 = pi1185;// level 0
assign po1205 = pi1093;// level 0
assign po1206 = pi1168;// level 0
assign po1207 = pi1173;// level 0
assign po1208 = pi1196;// level 0
assign po1209 = pi1170;// level 0
assign po1210 = pi1167;// level 0
assign po1211 = pi1195;// level 0
assign po1212 = pi1161;// level 0
assign po1213 = pi0840;// level 0
assign po1214 = pi1183;// level 0
assign po1215 = pi1189;// level 0
assign po1216 = pi0864;// level 0
assign po1217 = pi1184;// level 0
assign po1218 = pi1182;// level 0
assign po1219 = pi1174;// level 0
assign po1220 = pi1188;// level 0
assign po1221 = pi1091;// level 0
assign po1222 = pi1160;// level 0
assign po1223 = pi1194;// level 0
assign po1224 = pi1178;// level 0
endmodule
