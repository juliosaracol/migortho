module mem_ctrl ( 
    pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007, pi0008,
    pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016, pi0017,
    pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025, pi0026,
    pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034, pi0035,
    pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043, pi0044,
    pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052, pi0053,
    pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061, pi0062,
    pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070, pi0071,
    pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079, pi0080,
    pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088, pi0089,
    pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097, pi0098,
    pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106, pi0107,
    pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115, pi0116,
    pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124, pi0125,
    pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133, pi0134,
    pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142, pi0143,
    pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151, pi0152,
    pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160, pi0161,
    pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169, pi0170,
    pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178, pi0179,
    pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187, pi0188,
    pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196, pi0197,
    pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205, pi0206,
    pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214, pi0215,
    pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223, pi0224,
    pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232, pi0233,
    pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241, pi0242,
    pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250, pi0251,
    pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259, pi0260,
    pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268, pi0269,
    pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277, pi0278,
    pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286, pi0287,
    pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295, pi0296,
    pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304, pi0305,
    pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313, pi0314,
    pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322, pi0323,
    pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331, pi0332,
    pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340, pi0341,
    pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349, pi0350,
    pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358, pi0359,
    pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367, pi0368,
    pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376, pi0377,
    pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385, pi0386,
    pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394, pi0395,
    pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403, pi0404,
    pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412, pi0413,
    pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421, pi0422,
    pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430, pi0431,
    pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439, pi0440,
    pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448, pi0449,
    pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457, pi0458,
    pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466, pi0467,
    pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475, pi0476,
    pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484, pi0485,
    pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493, pi0494,
    pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502, pi0503,
    pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511, pi0512,
    pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520, pi0521,
    pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529, pi0530,
    pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538, pi0539,
    pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547, pi0548,
    pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556, pi0557,
    pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565, pi0566,
    pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574, pi0575,
    pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583, pi0584,
    pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592, pi0593,
    pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601, pi0602,
    pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610, pi0611,
    pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619, pi0620,
    pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628, pi0629,
    pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637, pi0638,
    pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646, pi0647,
    pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655, pi0656,
    pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664, pi0665,
    pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673, pi0674,
    pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682, pi0683,
    pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691, pi0692,
    pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700, pi0701,
    pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709, pi0710,
    pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718, pi0719,
    pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727, pi0728,
    pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736, pi0737,
    pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745, pi0746,
    pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754, pi0755,
    pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763, pi0764,
    pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772, pi0773,
    pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781, pi0782,
    pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790, pi0791,
    pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799, pi0800,
    pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808, pi0809,
    pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817, pi0818,
    pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826, pi0827,
    pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835, pi0836,
    pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844, pi0845,
    pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853, pi0854,
    pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862, pi0863,
    pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871, pi0872,
    pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880, pi0881,
    pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889, pi0890,
    pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898, pi0899,
    pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907, pi0908,
    pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916, pi0917,
    pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925, pi0926,
    pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934, pi0935,
    pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943, pi0944,
    pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952, pi0953,
    pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961, pi0962,
    pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970, pi0971,
    pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979, pi0980,
    pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988, pi0989,
    pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997, pi0998,
    pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197,
    po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007, po0008,
    po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016, po0017,
    po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025, po0026,
    po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034, po0035,
    po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043, po0044,
    po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052, po0053,
    po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061, po0062,
    po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070, po0071,
    po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079, po0080,
    po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088, po0089,
    po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097, po0098,
    po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106, po0107,
    po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115, po0116,
    po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124, po0125,
    po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133, po0134,
    po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142, po0143,
    po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151, po0152,
    po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160, po0161,
    po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169, po0170,
    po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178, po0179,
    po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187, po0188,
    po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196, po0197,
    po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205, po0206,
    po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214, po0215,
    po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223, po0224,
    po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232, po0233,
    po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241, po0242,
    po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250, po0251,
    po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259, po0260,
    po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268, po0269,
    po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277, po0278,
    po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286, po0287,
    po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295, po0296,
    po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304, po0305,
    po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313, po0314,
    po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322, po0323,
    po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331, po0332,
    po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340, po0341,
    po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349, po0350,
    po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358, po0359,
    po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367, po0368,
    po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376, po0377,
    po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385, po0386,
    po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394, po0395,
    po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403, po0404,
    po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412, po0413,
    po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421, po0422,
    po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430, po0431,
    po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439, po0440,
    po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448, po0449,
    po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457, po0458,
    po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466, po0467,
    po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475, po0476,
    po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484, po0485,
    po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493, po0494,
    po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502, po0503,
    po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511, po0512,
    po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520, po0521,
    po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529, po0530,
    po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538, po0539,
    po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547, po0548,
    po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556, po0557,
    po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565, po0566,
    po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574, po0575,
    po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583, po0584,
    po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592, po0593,
    po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601, po0602,
    po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610, po0611,
    po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619, po0620,
    po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628, po0629,
    po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637, po0638,
    po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646, po0647,
    po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655, po0656,
    po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664, po0665,
    po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673, po0674,
    po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682, po0683,
    po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691, po0692,
    po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700, po0701,
    po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709, po0710,
    po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718, po0719,
    po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727, po0728,
    po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736, po0737,
    po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745, po0746,
    po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754, po0755,
    po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763, po0764,
    po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772, po0773,
    po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781, po0782,
    po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790, po0791,
    po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799, po0800,
    po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808, po0809,
    po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817, po0818,
    po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826, po0827,
    po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835, po0836,
    po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844, po0845,
    po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853, po0854,
    po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862, po0863,
    po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871, po0872,
    po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880, po0881,
    po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889, po0890,
    po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898, po0899,
    po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907, po0908,
    po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916, po0917,
    po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925, po0926,
    po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934, po0935,
    po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943, po0944,
    po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952, po0953,
    po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961, po0962,
    po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970, po0971,
    po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979, po0980,
    po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988, po0989,
    po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997, po0998,
    po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224  );
  input  pi0000, pi0001, pi0002, pi0003, pi0004, pi0005, pi0006, pi0007,
    pi0008, pi0009, pi0010, pi0011, pi0012, pi0013, pi0014, pi0015, pi0016,
    pi0017, pi0018, pi0019, pi0020, pi0021, pi0022, pi0023, pi0024, pi0025,
    pi0026, pi0027, pi0028, pi0029, pi0030, pi0031, pi0032, pi0033, pi0034,
    pi0035, pi0036, pi0037, pi0038, pi0039, pi0040, pi0041, pi0042, pi0043,
    pi0044, pi0045, pi0046, pi0047, pi0048, pi0049, pi0050, pi0051, pi0052,
    pi0053, pi0054, pi0055, pi0056, pi0057, pi0058, pi0059, pi0060, pi0061,
    pi0062, pi0063, pi0064, pi0065, pi0066, pi0067, pi0068, pi0069, pi0070,
    pi0071, pi0072, pi0073, pi0074, pi0075, pi0076, pi0077, pi0078, pi0079,
    pi0080, pi0081, pi0082, pi0083, pi0084, pi0085, pi0086, pi0087, pi0088,
    pi0089, pi0090, pi0091, pi0092, pi0093, pi0094, pi0095, pi0096, pi0097,
    pi0098, pi0099, pi0100, pi0101, pi0102, pi0103, pi0104, pi0105, pi0106,
    pi0107, pi0108, pi0109, pi0110, pi0111, pi0112, pi0113, pi0114, pi0115,
    pi0116, pi0117, pi0118, pi0119, pi0120, pi0121, pi0122, pi0123, pi0124,
    pi0125, pi0126, pi0127, pi0128, pi0129, pi0130, pi0131, pi0132, pi0133,
    pi0134, pi0135, pi0136, pi0137, pi0138, pi0139, pi0140, pi0141, pi0142,
    pi0143, pi0144, pi0145, pi0146, pi0147, pi0148, pi0149, pi0150, pi0151,
    pi0152, pi0153, pi0154, pi0155, pi0156, pi0157, pi0158, pi0159, pi0160,
    pi0161, pi0162, pi0163, pi0164, pi0165, pi0166, pi0167, pi0168, pi0169,
    pi0170, pi0171, pi0172, pi0173, pi0174, pi0175, pi0176, pi0177, pi0178,
    pi0179, pi0180, pi0181, pi0182, pi0183, pi0184, pi0185, pi0186, pi0187,
    pi0188, pi0189, pi0190, pi0191, pi0192, pi0193, pi0194, pi0195, pi0196,
    pi0197, pi0198, pi0199, pi0200, pi0201, pi0202, pi0203, pi0204, pi0205,
    pi0206, pi0207, pi0208, pi0209, pi0210, pi0211, pi0212, pi0213, pi0214,
    pi0215, pi0216, pi0217, pi0218, pi0219, pi0220, pi0221, pi0222, pi0223,
    pi0224, pi0225, pi0226, pi0227, pi0228, pi0229, pi0230, pi0231, pi0232,
    pi0233, pi0234, pi0235, pi0236, pi0237, pi0238, pi0239, pi0240, pi0241,
    pi0242, pi0243, pi0244, pi0245, pi0246, pi0247, pi0248, pi0249, pi0250,
    pi0251, pi0252, pi0253, pi0254, pi0255, pi0256, pi0257, pi0258, pi0259,
    pi0260, pi0261, pi0262, pi0263, pi0264, pi0265, pi0266, pi0267, pi0268,
    pi0269, pi0270, pi0271, pi0272, pi0273, pi0274, pi0275, pi0276, pi0277,
    pi0278, pi0279, pi0280, pi0281, pi0282, pi0283, pi0284, pi0285, pi0286,
    pi0287, pi0288, pi0289, pi0290, pi0291, pi0292, pi0293, pi0294, pi0295,
    pi0296, pi0297, pi0298, pi0299, pi0300, pi0301, pi0302, pi0303, pi0304,
    pi0305, pi0306, pi0307, pi0308, pi0309, pi0310, pi0311, pi0312, pi0313,
    pi0314, pi0315, pi0316, pi0317, pi0318, pi0319, pi0320, pi0321, pi0322,
    pi0323, pi0324, pi0325, pi0326, pi0327, pi0328, pi0329, pi0330, pi0331,
    pi0332, pi0333, pi0334, pi0335, pi0336, pi0337, pi0338, pi0339, pi0340,
    pi0341, pi0342, pi0343, pi0344, pi0345, pi0346, pi0347, pi0348, pi0349,
    pi0350, pi0351, pi0352, pi0353, pi0354, pi0355, pi0356, pi0357, pi0358,
    pi0359, pi0360, pi0361, pi0362, pi0363, pi0364, pi0365, pi0366, pi0367,
    pi0368, pi0369, pi0370, pi0371, pi0372, pi0373, pi0374, pi0375, pi0376,
    pi0377, pi0378, pi0379, pi0380, pi0381, pi0382, pi0383, pi0384, pi0385,
    pi0386, pi0387, pi0388, pi0389, pi0390, pi0391, pi0392, pi0393, pi0394,
    pi0395, pi0396, pi0397, pi0398, pi0399, pi0400, pi0401, pi0402, pi0403,
    pi0404, pi0405, pi0406, pi0407, pi0408, pi0409, pi0410, pi0411, pi0412,
    pi0413, pi0414, pi0415, pi0416, pi0417, pi0418, pi0419, pi0420, pi0421,
    pi0422, pi0423, pi0424, pi0425, pi0426, pi0427, pi0428, pi0429, pi0430,
    pi0431, pi0432, pi0433, pi0434, pi0435, pi0436, pi0437, pi0438, pi0439,
    pi0440, pi0441, pi0442, pi0443, pi0444, pi0445, pi0446, pi0447, pi0448,
    pi0449, pi0450, pi0451, pi0452, pi0453, pi0454, pi0455, pi0456, pi0457,
    pi0458, pi0459, pi0460, pi0461, pi0462, pi0463, pi0464, pi0465, pi0466,
    pi0467, pi0468, pi0469, pi0470, pi0471, pi0472, pi0473, pi0474, pi0475,
    pi0476, pi0477, pi0478, pi0479, pi0480, pi0481, pi0482, pi0483, pi0484,
    pi0485, pi0486, pi0487, pi0488, pi0489, pi0490, pi0491, pi0492, pi0493,
    pi0494, pi0495, pi0496, pi0497, pi0498, pi0499, pi0500, pi0501, pi0502,
    pi0503, pi0504, pi0505, pi0506, pi0507, pi0508, pi0509, pi0510, pi0511,
    pi0512, pi0513, pi0514, pi0515, pi0516, pi0517, pi0518, pi0519, pi0520,
    pi0521, pi0522, pi0523, pi0524, pi0525, pi0526, pi0527, pi0528, pi0529,
    pi0530, pi0531, pi0532, pi0533, pi0534, pi0535, pi0536, pi0537, pi0538,
    pi0539, pi0540, pi0541, pi0542, pi0543, pi0544, pi0545, pi0546, pi0547,
    pi0548, pi0549, pi0550, pi0551, pi0552, pi0553, pi0554, pi0555, pi0556,
    pi0557, pi0558, pi0559, pi0560, pi0561, pi0562, pi0563, pi0564, pi0565,
    pi0566, pi0567, pi0568, pi0569, pi0570, pi0571, pi0572, pi0573, pi0574,
    pi0575, pi0576, pi0577, pi0578, pi0579, pi0580, pi0581, pi0582, pi0583,
    pi0584, pi0585, pi0586, pi0587, pi0588, pi0589, pi0590, pi0591, pi0592,
    pi0593, pi0594, pi0595, pi0596, pi0597, pi0598, pi0599, pi0600, pi0601,
    pi0602, pi0603, pi0604, pi0605, pi0606, pi0607, pi0608, pi0609, pi0610,
    pi0611, pi0612, pi0613, pi0614, pi0615, pi0616, pi0617, pi0618, pi0619,
    pi0620, pi0621, pi0622, pi0623, pi0624, pi0625, pi0626, pi0627, pi0628,
    pi0629, pi0630, pi0631, pi0632, pi0633, pi0634, pi0635, pi0636, pi0637,
    pi0638, pi0639, pi0640, pi0641, pi0642, pi0643, pi0644, pi0645, pi0646,
    pi0647, pi0648, pi0649, pi0650, pi0651, pi0652, pi0653, pi0654, pi0655,
    pi0656, pi0657, pi0658, pi0659, pi0660, pi0661, pi0662, pi0663, pi0664,
    pi0665, pi0666, pi0667, pi0668, pi0669, pi0670, pi0671, pi0672, pi0673,
    pi0674, pi0675, pi0676, pi0677, pi0678, pi0679, pi0680, pi0681, pi0682,
    pi0683, pi0684, pi0685, pi0686, pi0687, pi0688, pi0689, pi0690, pi0691,
    pi0692, pi0693, pi0694, pi0695, pi0696, pi0697, pi0698, pi0699, pi0700,
    pi0701, pi0702, pi0703, pi0704, pi0705, pi0706, pi0707, pi0708, pi0709,
    pi0710, pi0711, pi0712, pi0713, pi0714, pi0715, pi0716, pi0717, pi0718,
    pi0719, pi0720, pi0721, pi0722, pi0723, pi0724, pi0725, pi0726, pi0727,
    pi0728, pi0729, pi0730, pi0731, pi0732, pi0733, pi0734, pi0735, pi0736,
    pi0737, pi0738, pi0739, pi0740, pi0741, pi0742, pi0743, pi0744, pi0745,
    pi0746, pi0747, pi0748, pi0749, pi0750, pi0751, pi0752, pi0753, pi0754,
    pi0755, pi0756, pi0757, pi0758, pi0759, pi0760, pi0761, pi0762, pi0763,
    pi0764, pi0765, pi0766, pi0767, pi0768, pi0769, pi0770, pi0771, pi0772,
    pi0773, pi0774, pi0775, pi0776, pi0777, pi0778, pi0779, pi0780, pi0781,
    pi0782, pi0783, pi0784, pi0785, pi0786, pi0787, pi0788, pi0789, pi0790,
    pi0791, pi0792, pi0793, pi0794, pi0795, pi0796, pi0797, pi0798, pi0799,
    pi0800, pi0801, pi0802, pi0803, pi0804, pi0805, pi0806, pi0807, pi0808,
    pi0809, pi0810, pi0811, pi0812, pi0813, pi0814, pi0815, pi0816, pi0817,
    pi0818, pi0819, pi0820, pi0821, pi0822, pi0823, pi0824, pi0825, pi0826,
    pi0827, pi0828, pi0829, pi0830, pi0831, pi0832, pi0833, pi0834, pi0835,
    pi0836, pi0837, pi0838, pi0839, pi0840, pi0841, pi0842, pi0843, pi0844,
    pi0845, pi0846, pi0847, pi0848, pi0849, pi0850, pi0851, pi0852, pi0853,
    pi0854, pi0855, pi0856, pi0857, pi0858, pi0859, pi0860, pi0861, pi0862,
    pi0863, pi0864, pi0865, pi0866, pi0867, pi0868, pi0869, pi0870, pi0871,
    pi0872, pi0873, pi0874, pi0875, pi0876, pi0877, pi0878, pi0879, pi0880,
    pi0881, pi0882, pi0883, pi0884, pi0885, pi0886, pi0887, pi0888, pi0889,
    pi0890, pi0891, pi0892, pi0893, pi0894, pi0895, pi0896, pi0897, pi0898,
    pi0899, pi0900, pi0901, pi0902, pi0903, pi0904, pi0905, pi0906, pi0907,
    pi0908, pi0909, pi0910, pi0911, pi0912, pi0913, pi0914, pi0915, pi0916,
    pi0917, pi0918, pi0919, pi0920, pi0921, pi0922, pi0923, pi0924, pi0925,
    pi0926, pi0927, pi0928, pi0929, pi0930, pi0931, pi0932, pi0933, pi0934,
    pi0935, pi0936, pi0937, pi0938, pi0939, pi0940, pi0941, pi0942, pi0943,
    pi0944, pi0945, pi0946, pi0947, pi0948, pi0949, pi0950, pi0951, pi0952,
    pi0953, pi0954, pi0955, pi0956, pi0957, pi0958, pi0959, pi0960, pi0961,
    pi0962, pi0963, pi0964, pi0965, pi0966, pi0967, pi0968, pi0969, pi0970,
    pi0971, pi0972, pi0973, pi0974, pi0975, pi0976, pi0977, pi0978, pi0979,
    pi0980, pi0981, pi0982, pi0983, pi0984, pi0985, pi0986, pi0987, pi0988,
    pi0989, pi0990, pi0991, pi0992, pi0993, pi0994, pi0995, pi0996, pi0997,
    pi0998, pi0999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197;
  output po0000, po0001, po0002, po0003, po0004, po0005, po0006, po0007,
    po0008, po0009, po0010, po0011, po0012, po0013, po0014, po0015, po0016,
    po0017, po0018, po0019, po0020, po0021, po0022, po0023, po0024, po0025,
    po0026, po0027, po0028, po0029, po0030, po0031, po0032, po0033, po0034,
    po0035, po0036, po0037, po0038, po0039, po0040, po0041, po0042, po0043,
    po0044, po0045, po0046, po0047, po0048, po0049, po0050, po0051, po0052,
    po0053, po0054, po0055, po0056, po0057, po0058, po0059, po0060, po0061,
    po0062, po0063, po0064, po0065, po0066, po0067, po0068, po0069, po0070,
    po0071, po0072, po0073, po0074, po0075, po0076, po0077, po0078, po0079,
    po0080, po0081, po0082, po0083, po0084, po0085, po0086, po0087, po0088,
    po0089, po0090, po0091, po0092, po0093, po0094, po0095, po0096, po0097,
    po0098, po0099, po0100, po0101, po0102, po0103, po0104, po0105, po0106,
    po0107, po0108, po0109, po0110, po0111, po0112, po0113, po0114, po0115,
    po0116, po0117, po0118, po0119, po0120, po0121, po0122, po0123, po0124,
    po0125, po0126, po0127, po0128, po0129, po0130, po0131, po0132, po0133,
    po0134, po0135, po0136, po0137, po0138, po0139, po0140, po0141, po0142,
    po0143, po0144, po0145, po0146, po0147, po0148, po0149, po0150, po0151,
    po0152, po0153, po0154, po0155, po0156, po0157, po0158, po0159, po0160,
    po0161, po0162, po0163, po0164, po0165, po0166, po0167, po0168, po0169,
    po0170, po0171, po0172, po0173, po0174, po0175, po0176, po0177, po0178,
    po0179, po0180, po0181, po0182, po0183, po0184, po0185, po0186, po0187,
    po0188, po0189, po0190, po0191, po0192, po0193, po0194, po0195, po0196,
    po0197, po0198, po0199, po0200, po0201, po0202, po0203, po0204, po0205,
    po0206, po0207, po0208, po0209, po0210, po0211, po0212, po0213, po0214,
    po0215, po0216, po0217, po0218, po0219, po0220, po0221, po0222, po0223,
    po0224, po0225, po0226, po0227, po0228, po0229, po0230, po0231, po0232,
    po0233, po0234, po0235, po0236, po0237, po0238, po0239, po0240, po0241,
    po0242, po0243, po0244, po0245, po0246, po0247, po0248, po0249, po0250,
    po0251, po0252, po0253, po0254, po0255, po0256, po0257, po0258, po0259,
    po0260, po0261, po0262, po0263, po0264, po0265, po0266, po0267, po0268,
    po0269, po0270, po0271, po0272, po0273, po0274, po0275, po0276, po0277,
    po0278, po0279, po0280, po0281, po0282, po0283, po0284, po0285, po0286,
    po0287, po0288, po0289, po0290, po0291, po0292, po0293, po0294, po0295,
    po0296, po0297, po0298, po0299, po0300, po0301, po0302, po0303, po0304,
    po0305, po0306, po0307, po0308, po0309, po0310, po0311, po0312, po0313,
    po0314, po0315, po0316, po0317, po0318, po0319, po0320, po0321, po0322,
    po0323, po0324, po0325, po0326, po0327, po0328, po0329, po0330, po0331,
    po0332, po0333, po0334, po0335, po0336, po0337, po0338, po0339, po0340,
    po0341, po0342, po0343, po0344, po0345, po0346, po0347, po0348, po0349,
    po0350, po0351, po0352, po0353, po0354, po0355, po0356, po0357, po0358,
    po0359, po0360, po0361, po0362, po0363, po0364, po0365, po0366, po0367,
    po0368, po0369, po0370, po0371, po0372, po0373, po0374, po0375, po0376,
    po0377, po0378, po0379, po0380, po0381, po0382, po0383, po0384, po0385,
    po0386, po0387, po0388, po0389, po0390, po0391, po0392, po0393, po0394,
    po0395, po0396, po0397, po0398, po0399, po0400, po0401, po0402, po0403,
    po0404, po0405, po0406, po0407, po0408, po0409, po0410, po0411, po0412,
    po0413, po0414, po0415, po0416, po0417, po0418, po0419, po0420, po0421,
    po0422, po0423, po0424, po0425, po0426, po0427, po0428, po0429, po0430,
    po0431, po0432, po0433, po0434, po0435, po0436, po0437, po0438, po0439,
    po0440, po0441, po0442, po0443, po0444, po0445, po0446, po0447, po0448,
    po0449, po0450, po0451, po0452, po0453, po0454, po0455, po0456, po0457,
    po0458, po0459, po0460, po0461, po0462, po0463, po0464, po0465, po0466,
    po0467, po0468, po0469, po0470, po0471, po0472, po0473, po0474, po0475,
    po0476, po0477, po0478, po0479, po0480, po0481, po0482, po0483, po0484,
    po0485, po0486, po0487, po0488, po0489, po0490, po0491, po0492, po0493,
    po0494, po0495, po0496, po0497, po0498, po0499, po0500, po0501, po0502,
    po0503, po0504, po0505, po0506, po0507, po0508, po0509, po0510, po0511,
    po0512, po0513, po0514, po0515, po0516, po0517, po0518, po0519, po0520,
    po0521, po0522, po0523, po0524, po0525, po0526, po0527, po0528, po0529,
    po0530, po0531, po0532, po0533, po0534, po0535, po0536, po0537, po0538,
    po0539, po0540, po0541, po0542, po0543, po0544, po0545, po0546, po0547,
    po0548, po0549, po0550, po0551, po0552, po0553, po0554, po0555, po0556,
    po0557, po0558, po0559, po0560, po0561, po0562, po0563, po0564, po0565,
    po0566, po0567, po0568, po0569, po0570, po0571, po0572, po0573, po0574,
    po0575, po0576, po0577, po0578, po0579, po0580, po0581, po0582, po0583,
    po0584, po0585, po0586, po0587, po0588, po0589, po0590, po0591, po0592,
    po0593, po0594, po0595, po0596, po0597, po0598, po0599, po0600, po0601,
    po0602, po0603, po0604, po0605, po0606, po0607, po0608, po0609, po0610,
    po0611, po0612, po0613, po0614, po0615, po0616, po0617, po0618, po0619,
    po0620, po0621, po0622, po0623, po0624, po0625, po0626, po0627, po0628,
    po0629, po0630, po0631, po0632, po0633, po0634, po0635, po0636, po0637,
    po0638, po0639, po0640, po0641, po0642, po0643, po0644, po0645, po0646,
    po0647, po0648, po0649, po0650, po0651, po0652, po0653, po0654, po0655,
    po0656, po0657, po0658, po0659, po0660, po0661, po0662, po0663, po0664,
    po0665, po0666, po0667, po0668, po0669, po0670, po0671, po0672, po0673,
    po0674, po0675, po0676, po0677, po0678, po0679, po0680, po0681, po0682,
    po0683, po0684, po0685, po0686, po0687, po0688, po0689, po0690, po0691,
    po0692, po0693, po0694, po0695, po0696, po0697, po0698, po0699, po0700,
    po0701, po0702, po0703, po0704, po0705, po0706, po0707, po0708, po0709,
    po0710, po0711, po0712, po0713, po0714, po0715, po0716, po0717, po0718,
    po0719, po0720, po0721, po0722, po0723, po0724, po0725, po0726, po0727,
    po0728, po0729, po0730, po0731, po0732, po0733, po0734, po0735, po0736,
    po0737, po0738, po0739, po0740, po0741, po0742, po0743, po0744, po0745,
    po0746, po0747, po0748, po0749, po0750, po0751, po0752, po0753, po0754,
    po0755, po0756, po0757, po0758, po0759, po0760, po0761, po0762, po0763,
    po0764, po0765, po0766, po0767, po0768, po0769, po0770, po0771, po0772,
    po0773, po0774, po0775, po0776, po0777, po0778, po0779, po0780, po0781,
    po0782, po0783, po0784, po0785, po0786, po0787, po0788, po0789, po0790,
    po0791, po0792, po0793, po0794, po0795, po0796, po0797, po0798, po0799,
    po0800, po0801, po0802, po0803, po0804, po0805, po0806, po0807, po0808,
    po0809, po0810, po0811, po0812, po0813, po0814, po0815, po0816, po0817,
    po0818, po0819, po0820, po0821, po0822, po0823, po0824, po0825, po0826,
    po0827, po0828, po0829, po0830, po0831, po0832, po0833, po0834, po0835,
    po0836, po0837, po0838, po0839, po0840, po0841, po0842, po0843, po0844,
    po0845, po0846, po0847, po0848, po0849, po0850, po0851, po0852, po0853,
    po0854, po0855, po0856, po0857, po0858, po0859, po0860, po0861, po0862,
    po0863, po0864, po0865, po0866, po0867, po0868, po0869, po0870, po0871,
    po0872, po0873, po0874, po0875, po0876, po0877, po0878, po0879, po0880,
    po0881, po0882, po0883, po0884, po0885, po0886, po0887, po0888, po0889,
    po0890, po0891, po0892, po0893, po0894, po0895, po0896, po0897, po0898,
    po0899, po0900, po0901, po0902, po0903, po0904, po0905, po0906, po0907,
    po0908, po0909, po0910, po0911, po0912, po0913, po0914, po0915, po0916,
    po0917, po0918, po0919, po0920, po0921, po0922, po0923, po0924, po0925,
    po0926, po0927, po0928, po0929, po0930, po0931, po0932, po0933, po0934,
    po0935, po0936, po0937, po0938, po0939, po0940, po0941, po0942, po0943,
    po0944, po0945, po0946, po0947, po0948, po0949, po0950, po0951, po0952,
    po0953, po0954, po0955, po0956, po0957, po0958, po0959, po0960, po0961,
    po0962, po0963, po0964, po0965, po0966, po0967, po0968, po0969, po0970,
    po0971, po0972, po0973, po0974, po0975, po0976, po0977, po0978, po0979,
    po0980, po0981, po0982, po0983, po0984, po0985, po0986, po0987, po0988,
    po0989, po0990, po0991, po0992, po0993, po0994, po0995, po0996, po0997,
    po0998, po0999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224;
  wire n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
    n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635,
    n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665,
    n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
    n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2721, n2722, n2723, n2725, n2726, n2727,
    n2728, n2730, n2733, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
    n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
    n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
    n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
    n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
    n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2951, n2952, n2953,
    n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
    n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
    n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
    n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
    n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
    n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
    n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
    n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
    n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3140, n3141, n3142, n3143, n3144, n3145,
    n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
    n3167, n3168, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3218, n3219, n3220,
    n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
    n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
    n3263, n3264, n3265, n3266, n3267, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3314, n3315, n3316,
    n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
    n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
    n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
    n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
    n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
    n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
    n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3504, n3505, n3506, n3509, n3511, n3513,
    n3515, n3517, n3519, n3521, n3522, n3524, n3525, n3526, n3527, n3529,
    n3530, n3532, n3533, n3535, n3536, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
    n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
    n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
    n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
    n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
    n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
    n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
    n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
    n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
    n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
    n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
    n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
    n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
    n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
    n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
    n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
    n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
    n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
    n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
    n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
    n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
    n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
    n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
    n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
    n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
    n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
    n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
    n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
    n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
    n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
    n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
    n4802, n4803, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
    n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
    n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4950, n4951, n4952, n4953, n4954, n4955,
    n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996,
    n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
    n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
    n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
    n5129, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
    n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
    n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
    n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
    n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
    n5240, n5241, n5242, n5243, n5244, n5245, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
    n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
    n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
    n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
    n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
    n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
    n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
    n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
    n5472, n5473, n5474, n5475, n5477, n5478, n5479, n5480, n5481, n5482,
    n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
    n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
    n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5592, n5593,
    n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
    n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
    n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
    n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
    n5714, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
    n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
    n5846, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
    n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
    n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
    n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
    n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
    n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
    n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
    n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
    n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
    n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
    n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
    n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
    n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
    n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
    n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305, n6307, n6308, n6309, n6310,
    n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
    n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
    n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
    n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6430, n6431,
    n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
    n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
    n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
    n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
    n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
    n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
    n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
    n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
    n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
    n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
    n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
    n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
    n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
    n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
    n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
    n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
    n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
    n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
    n6774, n6775, n6776, n6777, n6779, n6780, n6781, n6782, n6783, n6784,
    n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
    n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
    n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
    n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
    n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7006,
    n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096,
    n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127,
    n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157,
    n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187,
    n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
    n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7348, n7349,
    n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
    n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
    n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
    n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
    n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
    n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
    n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
    n7460, n7461, n7462, n7463, n7464, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591,
    n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601,
    n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621,
    n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631,
    n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651,
    n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661,
    n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681,
    n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691,
    n7692, n7693, n7694, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
    n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
    n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808, n7810, n7811, n7812, n7813,
    n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
    n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
    n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
    n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
    n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
    n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
    n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
    n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
    n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
    n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
    n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
    n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
    n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
    n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
    n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
    n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8164, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297,
    n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307,
    n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
    n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337,
    n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357,
    n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367,
    n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387,
    n8388, n8389, n8390, n8391, n8392, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
    n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
    n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
    n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
    n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
    n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
    n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
    n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
    n8620, n8621, n8622, n8623, n8624, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736, n8738, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788, n8790, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
    n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
    n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
    n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
    n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
    n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
    n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
    n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
    n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
    n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
    n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9137,
    n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147,
    n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167,
    n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177,
    n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197,
    n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207,
    n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
    n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237,
    n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9367, n9368, n9369,
    n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
    n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
    n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
    n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
    n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
    n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
    n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
    n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
    n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9596, n9597, n9598, n9599, n9600, n9601,
    n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621,
    n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631,
    n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651,
    n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661,
    n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681,
    n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691,
    n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9703, n9704, n9705, n9707, n9708, n9709, n9710, n9711, n9712,
    n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
    n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
    n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
    n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9822, n9823,
    n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
    n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
    n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
    n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
    n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
    n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
    n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
    n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
    n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
    n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
    n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
    n9934, n9935, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
    n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
    n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
    n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
    n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
    n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030,
    n10031, n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
    n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
    n10049, n10050, n10051, n10052, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
    n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
    n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
    n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
    n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
    n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
    n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293, n10294,
    n10295, n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
    n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
    n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
    n10394, n10395, n10396, n10398, n10399, n10400, n10401, n10402, n10403,
    n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
    n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
    n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
    n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
    n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
    n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10521,
    n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
    n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
    n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
    n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
    n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
    n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
    n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
    n10630, n10631, n10632, n10633, n10634, n10636, n10637, n10638, n10639,
    n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
    n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
    n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
    n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
    n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10752, n10753, n10754, n10755, n10756, n10757,
    n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
    n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
    n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
    n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
    n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
    n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
    n10866, n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
    n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893, n10894,
    n10895, n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
    n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
    n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
    n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
    n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
    n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
    n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
    n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965, n10966,
    n10967, n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
    n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
    n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
    n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11003, n11004,
    n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
    n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021, n11022,
    n11023, n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
    n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
    n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
    n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
    n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
    n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
    n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
    n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
    n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11117, n11118, n11119, n11120, n11121, n11122,
    n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
    n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157, n11158,
    n11159, n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
    n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229, n11231,
    n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
    n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
    n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11345, n11346, n11347, n11348, n11349,
    n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357, n11358,
    n11359, n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
    n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
    n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
    n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
    n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
    n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
    n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
    n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
    n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
    n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
    n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
    n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
    n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565, n11566,
    n11567, n11568, n11569, n11570, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
    n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
    n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
    n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11688, n11689, n11690, n11691, n11692, n11693, n11694,
    n11695, n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
    n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
    n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
    n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
    n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
    n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765, n11766,
    n11767, n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
    n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
    n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
    n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
    n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
    n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
    n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829, n11830,
    n11831, n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
    n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
    n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
    n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901, n11902,
    n11903, n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12033, n12034, n12035, n12036, n12037, n12038, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12048, n12049, n12050, n12051,
    n12052, n12053, n12055, n12056, n12057, n12058, n12059, n12060, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068, n12070, n12071, n12072,
    n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
    n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
    n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
    n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
    n12109, n12110, n12112, n12113, n12114, n12115, n12116, n12117, n12118,
    n12119, n12120, n12121, n12122, n12123, n12124, n12125, n12127, n12129,
    n12130, n12131, n12132, n12133, n12135, n12136, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182, n12184, n12185, n12186,
    n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
    n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
    n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
    n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221, n12222,
    n12223, n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
    n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
    n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
    n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
    n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
    n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275, n12276,
    n12277, n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
    n12286, n12287, n12288, n12289, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
    n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
    n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
    n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12342,
    n12343, n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
    n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
    n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
    n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
    n12379, n12381, n12382, n12383, n12384, n12385, n12386, n12387, n12388,
    n12389, n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
    n12398, n12399, n12400, n12401, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
    n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
    n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443, n12444,
    n12445, n12447, n12448, n12449, n12450, n12451, n12452, n12453, n12454,
    n12455, n12456, n12457, n12458, n12459, n12460, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
    n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12482, n12483,
    n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491, n12492,
    n12493, n12494, n12495, n12496, n12497, n12498, n12500, n12501, n12502,
    n12503, n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12517, n12518, n12520, n12521, n12522,
    n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
    n12532, n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
    n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
    n12570, n12571, n12572, n12573, n12575, n12576, n12577, n12578, n12579,
    n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587, n12588,
    n12589, n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
    n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605, n12606,
    n12607, n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
    n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
    n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
    n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
    n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
    n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659, n12660,
    n12661, n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
    n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677, n12678,
    n12679, n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
    n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
    n12697, n12698, n12699, n12701, n12702, n12703, n12704, n12705, n12706,
    n12708, n12709, n12710, n12711, n12712, n12713, n12715, n12716, n12717,
    n12718, n12719, n12720, n12722, n12723, n12724, n12725, n12726, n12727,
    n12729, n12730, n12731, n12732, n12733, n12734, n12736, n12737, n12738,
    n12739, n12740, n12741, n12743, n12744, n12745, n12746, n12747, n12748,
    n12750, n12751, n12752, n12753, n12754, n12756, n12757, n12758, n12759,
    n12760, n12761, n12763, n12764, n12765, n12766, n12767, n12768, n12770,
    n12771, n12772, n12773, n12774, n12775, n12777, n12778, n12779, n12780,
    n12781, n12782, n12784, n12785, n12786, n12787, n12788, n12789, n12791,
    n12792, n12793, n12794, n12795, n12796, n12798, n12799, n12800, n12801,
    n12802, n12803, n12805, n12806, n12807, n12808, n12809, n12810, n12812,
    n12813, n12814, n12815, n12816, n12817, n12819, n12820, n12821, n12822,
    n12823, n12824, n12826, n12827, n12828, n12829, n12830, n12831, n12833,
    n12834, n12835, n12836, n12837, n12838, n12840, n12841, n12842, n12843,
    n12844, n12846, n12847, n12848, n12849, n12850, n12852, n12853, n12854,
    n12855, n12856, n12857, n12859, n12860, n12861, n12862, n12863, n12864,
    n12866, n12867, n12868, n12869, n12870, n12872, n12873, n12874, n12875,
    n12876, n12877, n12879, n12880, n12881, n12882, n12883, n12884, n12886,
    n12887, n12888, n12889, n12890, n12891, n12893, n12894, n12895, n12896,
    n12897, n12898, n12900, n12901, n12902, n12903, n12904, n12905, n12907,
    n12908, n12909, n12910, n12911, n12912, n12914, n12915, n12916, n12917,
    n12918, n12919, n12921, n12922, n12923, n12924, n12925, n12927, n12928,
    n12929, n12930, n12931, n12933, n12934, n12935, n12936, n12937, n12939,
    n12940, n12941, n12942, n12943, n12945, n12946, n12947, n12948, n12949,
    n12951, n12952, n12953, n12954, n12955, n12957, n12958, n12959, n12960,
    n12961, n12963, n12964, n12965, n12966, n12967, n12969, n12970, n12971,
    n12972, n12973, n12975, n12976, n12977, n12978, n12979, n12981, n12982,
    n12983, n12984, n12985, n12987, n12988, n12989, n12990, n12991, n12993,
    n12994, n12995, n12996, n12997, n12999, n13000, n13001, n13002, n13003,
    n13005, n13006, n13007, n13008, n13009, n13011, n13012, n13013, n13014,
    n13015, n13017, n13018, n13019, n13020, n13021, n13023, n13024, n13025,
    n13026, n13027, n13029, n13030, n13031, n13032, n13033, n13035, n13036,
    n13037, n13038, n13039, n13041, n13042, n13043, n13044, n13045, n13047,
    n13048, n13049, n13050, n13051, n13053, n13054, n13055, n13056, n13057,
    n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
    n13067, n13068, n13069, n13070, n13071, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
    n13086, n13087, n13089, n13090, n13091, n13092, n13093, n13095, n13096,
    n13097, n13098, n13099, n13100, n13102, n13103, n13104, n13105, n13106,
    n13108, n13109, n13110, n13111, n13112, n13114, n13115, n13116, n13117,
    n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125, n13126,
    n13127, n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
    n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
    n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
    n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
    n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
    n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179, n13180,
    n13181, n13182, n13183, n13185, n13186, n13187, n13188, n13189, n13190,
    n13192, n13193, n13194, n13195, n13196, n13198, n13199, n13200, n13201,
    n13202, n13203, n13204, n13205, n13207, n13208, n13209, n13210, n13211,
    n13213, n13214, n13215, n13216, n13217, n13219, n13220, n13221, n13222,
    n13223, n13224, n13226, n13227, n13228, n13229, n13230, n13231, n13233,
    n13234, n13235, n13236, n13237, n13238, n13240, n13241, n13242, n13243,
    n13244, n13246, n13247, n13248, n13249, n13250, n13252, n13253, n13254,
    n13255, n13256, n13258, n13259, n13260, n13261, n13262, n13264, n13265,
    n13266, n13267, n13268, n13270, n13271, n13272, n13273, n13274, n13275,
    n13276, n13278, n13279, n13280, n13281, n13282, n13284, n13285, n13286,
    n13287, n13288, n13290, n13291, n13292, n13293, n13295, n13296, n13297,
    n13298, n13299, n13301, n13302, n13303, n13304, n13306, n13307, n13308,
    n13309, n13310, n13312, n13313, n13314, n13315, n13316, n13318, n13319,
    n13320, n13321, n13322, n13324, n13325, n13326, n13327, n13328, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336, n13338, n13340, n13341,
    n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349, n13350,
    n13351, n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
    n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
    n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
    n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
    n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403, n13404,
    n13405, n13406, n13407, n13408, n13409, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
    n13424, n13425, n13426, n13427, n13428, n13430, n13431, n13432, n13433,
    n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
    n13453, n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
    n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469, n13470,
    n13471, n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
    n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
    n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
    n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
    n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515, n13516,
    n13517, n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
    n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13534, n13535,
    n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
    n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13563,
    n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571, n13572,
    n13573, n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
    n13582, n13583, n13584, n13585, n13586, n13587, n13589, n13590, n13591,
    n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13607, n13608, n13609, n13610,
    n13611, n13613, n13614, n13615, n13616, n13617, n13618, n13619, n13620,
    n13621, n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
    n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637, n13638,
    n13639, n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
    n13668, n13669, n13670, n13671, n13672, n13673, n13675, n13676, n13677,
    n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685, n13686,
    n13687, n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
    n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
    n13705, n13706, n13708, n13709, n13710, n13711, n13712, n13714, n13715,
    n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13731, n13732, n13733, n13734,
    n13735, n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13748, n13749, n13750, n13751, n13752, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
    n13764, n13765, n13766, n13767, n13768, n13769, n13771, n13772, n13773,
    n13774, n13775, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
    n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
    n13795, n13796, n13797, n13798, n13800, n13801, n13802, n13803, n13804,
    n13805, n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13832, n13833,
    n13834, n13835, n13836, n13838, n13839, n13840, n13841, n13842, n13844,
    n13845, n13846, n13847, n13848, n13850, n13851, n13852, n13853, n13854,
    n13856, n13857, n13858, n13859, n13860, n13862, n13863, n13864, n13865,
    n13866, n13868, n13869, n13870, n13871, n13872, n13874, n13875, n13876,
    n13877, n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13904, n13905,
    n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13915,
    n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923, n13924,
    n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
    n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
    n13954, n13955, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
    n13964, n13965, n13966, n13967, n13968, n13969, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13982, n13983,
    n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13993,
    n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
    n14003, n14004, n14005, n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018, n14019, n14021, n14022,
    n14023, n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
    n14032, n14033, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
    n14042, n14043, n14044, n14046, n14047, n14048, n14049, n14050, n14051,
    n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14060, n14061,
    n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069, n14070,
    n14071, n14072, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
    n14081, n14082, n14083, n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14107, n14108, n14109, n14110,
    n14111, n14112, n14113, n14114, n14115, n14116, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14129, n14130,
    n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14140,
    n14141, n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
    n14150, n14151, n14152, n14154, n14155, n14156, n14157, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
    n14170, n14171, n14172, n14173, n14175, n14176, n14177, n14178, n14179,
    n14180, n14181, n14182, n14183, n14184, n14186, n14188, n14189, n14190,
    n14191, n14192, n14193, n14195, n14196, n14197, n14198, n14199, n14200,
    n14201, n14202, n14203, n14204, n14206, n14207, n14209, n14210, n14212,
    n14213, n14215, n14216, n14218, n14219, n14221, n14222, n14224, n14225,
    n14227, n14228, n14230, n14231, n14233, n14234, n14235, n14236, n14237,
    n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
    n14256, n14257, n14258, n14260, n14261, n14262, n14263, n14264, n14265,
    n14267, n14268, n14269, n14270, n14271, n14272, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14282, n14283, n14285, n14286, n14288,
    n14289, n14291, n14292, n14294, n14295, n14297, n14298, n14300, n14301,
    n14303, n14304, n14305, n14306, n14307, n14308, n14309, n14311, n14312,
    n14313, n14314, n14315, n14316, n14318, n14319, n14320, n14322, n14323,
    n14324, n14325, n14326, n14328, n14329, n14331, n14332, n14333, n14334,
    n14336, n14337, n14338, n14340, n14341, n14343, n14344, n14345, n14347,
    n14348, n14349, n14351, n14352, n14354, n14355, n14357, n14358, n14360,
    n14361, n14363, n14364, n14366, n14367, n14369, n14370, n14372, n14373,
    n14375, n14376, n14378, n14379, n14381, n14382, n14384, n14385, n14386,
    n14388, n14389, n14391, n14393, n14394, n14396, n14397, n14399, n14400,
    n14402, n14403, n14405, n14406, n14408, n14409, n14411, n14412, n14414,
    n14415, n14416, n14418, n14419, n14421, n14422, n14424, n14425, n14427,
    n14428, n14430, n14431, n14433, n14434, n14436, n14437, n14439, n14440,
    n14442, n14443, n14445, n14446, n14448, n14449, n14451, n14452, n14454,
    n14455, n14457, n14458, n14460, n14461, n14463, n14464, n14466, n14467,
    n14469, n14470, n14472, n14473, n14475, n14476, n14478, n14479, n14481,
    n14482, n14484, n14485, n14487, n14488, n14490, n14491, n14493, n14494,
    n14496, n14497, n14499, n14500, n14502, n14503, n14505, n14506, n14508,
    n14509, n14511, n14512, n14514, n14515, n14517, n14518, n14520, n14521,
    n14523, n14524, n14526, n14527, n14529, n14530, n14532, n14533, n14535,
    n14536, n14538, n14539, n14541, n14542, n14544, n14545, n14547, n14548,
    n14550, n14551, n14553, n14554, n14556, n14557, n14559, n14560, n14562,
    n14563, n14565, n14566, n14568, n14569, n14571, n14572, n14574, n14575,
    n14577, n14578, n14580, n14581, n14583, n14584, n14586, n14587, n14589,
    n14590, n14592, n14593, n14595, n14596, n14598, n14599, n14601, n14602,
    n14604, n14605, n14607, n14608, n14610, n14611, n14613, n14614, n14616,
    n14617, n14619, n14620, n14622, n14623, n14625, n14626, n14628, n14629,
    n14631, n14632, n14634, n14635, n14637, n14638, n14640, n14641, n14643,
    n14644, n14646, n14647, n14649, n14650, n14652, n14653, n14655, n14656,
    n14658, n14659, n14661, n14662, n14664, n14665, n14667, n14668, n14670,
    n14671, n14673, n14674, n14676, n14677, n14679, n14680, n14682, n14683,
    n14685, n14686, n14688, n14689, n14691, n14692, n14694, n14695, n14697,
    n14698, n14700, n14701, n14703, n14704, n14706, n14707, n14709, n14710,
    n14712, n14713, n14715, n14716, n14718, n14719, n14721, n14722, n14724,
    n14725, n14727, n14728, n14730, n14731, n14733, n14734, n14736, n14737,
    n14739, n14740, n14742, n14743, n14745, n14746, n14748, n14749, n14751,
    n14752, n14754, n14755, n14757, n14758, n14760, n14761, n14763, n14764,
    n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
    n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
    n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14819, n14820,
    n14822, n14823, n14825, n14826, n14828, n14829, n14831, n14832, n14834,
    n14835, n14837, n14838, n14840, n14841, n14842, n14843, n14844, n14846,
    n14847, n14848, n14849, n14850, n14852, n14853, n14854, n14855, n14856,
    n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
    n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
    n14875, n14876, n14877, n14878, n14880, n14881, n14882, n14884, n14885,
    n14886, n14887, n14888, n14890, n14891, n14892, n14893, n14894, n14896,
    n14897, n14898, n14899, n14900, n14902, n14903, n14904, n14905, n14906,
    n14908, n14909, n14910, n14911, n14912, n14914, n14915, n14916, n14917,
    n14918, n14920, n14921, n14922, n14923, n14924, n14926, n14927, n14928,
    n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
    n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
    n14947, n14948, n14949, n14952, n14953, n14955, n14956, n14958, n14959,
    n14961, n14962, n14964, n14965, n14967, n14968, n14970, n14971, n14973,
    n14974, n14976, n14977, n14979, n14980, n14982, n14983, n14985, n14986,
    n14988, n14989, n14991, n14992, n14994, n14995, n14997, n14998, n15000,
    n15001, n15003, n15004, n15006, n15007, n15009, n15010, n15012, n15013,
    n15015, n15016, n15018, n15019, n15021, n15022, n15024, n15025, n15027,
    n15028, n15030, n15031, n15033, n15034, n15036, n15037, n15039, n15040,
    n15042, n15043, n15045, n15046, n15048, n15049, n15051, n15052, n15054,
    n15055, n15057, n15058, n15060, n15061, n15063, n15064, n15066, n15067,
    n15069, n15070, n15072, n15073, n15075, n15076, n15078, n15079, n15081,
    n15082, n15084, n15085, n15087, n15088, n15090, n15091, n15093, n15094,
    n15096, n15097, n15099, n15100, n15102, n15103, n15105, n15106, n15108,
    n15109, n15111, n15112, n15114, n15115, n15117, n15118, n15120, n15121,
    n15123, n15124, n15126, n15127, n15129, n15130, n15132, n15133, n15135,
    n15136, n15138, n15139, n15141, n15142, n15144, n15145, n15147, n15148,
    n15150, n15151, n15153, n15154, n15156, n15157, n15159, n15160, n15162,
    n15163, n15165, n15166, n15168, n15169, n15171, n15172, n15174, n15175,
    n15177, n15178, n15180, n15181, n15183, n15184, n15186, n15187, n15189,
    n15190, n15192, n15193, n15195, n15196, n15198, n15199, n15201, n15202,
    n15204, n15205, n15207, n15208, n15211, n15212, n15213, n15214, n15215,
    n15216, n15217, n15219, n15220, n15222, n15223, n15225, n15226, n15228,
    n15229, n15231, n15232, n15234, n15235, n15237, n15238, n15240, n15241,
    n15243, n15244, n15246, n15247, n15249, n15250, n15252, n15253, n15255,
    n15256, n15258, n15259, n15261, n15262, n15264, n15265, n15267, n15268,
    n15270, n15271, n15273, n15274, n15276, n15277, n15278, n15279, n15281,
    n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296, n15298, n15299, n15300,
    n15302, n15303, n15304, n15306, n15307, n15308, n15310, n15311, n15312,
    n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
    n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347, n15348,
    n15349, n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365, n15366,
    n15367, n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
    n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
    n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419, n15420,
    n15421, n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437, n15438,
    n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
    n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
    n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
    n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492,
    n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
    n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509, n15510,
    n15511, n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
    n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
    n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
    n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
    n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
    n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563, n15564,
    n15565, n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
    n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581, n15582,
    n15583, n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
    n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
    n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
    n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
    n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635, n15636,
    n15637, n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
    n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653, n15654,
    n15655, n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
    n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
    n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
    n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
    n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
    n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707, n15708,
    n15709, n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
    n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725, n15726,
    n15727, n15728, n15729, n15730, n15731, n15732, n15733, n15735, n15736,
    n15737, n15738, n15739, n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15750, n15751, n15752, n15753, n15754, n15755, n15756,
    n15757, n15759, n15760, n15761, n15762, n15763, n15764, n15767, n15768,
    n15769, n15770, n15771, n15772, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15783, n15784, n15785, n15786, n15787, n15789,
    n15790, n15791, n15792, n15793, n15794, n15796, n15797, n15799, n15800,
    n15801, n15802, n15803, n15804, n15806, n15807, n15808, n15809, n15810,
    n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15820, n15821,
    n15822, n15824, n15825, n15826, n15827, n15828, n15830, n15831, n15832,
    n15834, n15835, n15836, n15838, n15839, n15840, n15842, n15843, n15844,
    n15846, n15847, n15848, n15850, n15851, n15852, n15854, n15855, n15856,
    n15858, n15859, n15860, n15861, n15863, n15864, n15865, n15866, n15867,
    n15869, n15870, n15871, n15872, n15874, n15875, n15876, n15877, n15878,
    n15880, n15881, n15882, n15884, n15885, n15886, n15888, n15889, n15890,
    n15892, n15893, n15894, n15896, n15897, n15898, n15900, n15901, n15902,
    n15904, n15905, n15906, n15907, n15908, n15910, n15911, n15912, n15913,
    n15915, n15916, n15917, n15919, n15920, n15921, n15923, n15924, n15925,
    n15927, n15928, n15929, n15931, n15932, n15933, n15935, n15936, n15937,
    n15939, n15940, n15941, n15943, n15944, n15945, n15947, n15948, n15949,
    n15951, n15952, n15953, n15955, n15956, n15957, n15959, n15960, n15961,
    n15963, n15964, n15965, n15967, n15968, n15969, n15971, n15972, n15973,
    n15975, n15976, n15977, n15979, n15980, n15981, n15983, n15984, n15985,
    n15987, n15988, n15989, n15991, n15992, n15993, n15995, n15996, n15997,
    n15999, n16000, n16001, n16003, n16004, n16005, n16007, n16008, n16009,
    n16011, n16012, n16013, n16015, n16016, n16017, n16019, n16020, n16021,
    n16023, n16024, n16025, n16027, n16028, n16029, n16031, n16032, n16033,
    n16035, n16036, n16037, n16039, n16040, n16041, n16043, n16044, n16045,
    n16047, n16048, n16049, n16051, n16052, n16053, n16054, n16055, n16056,
    n16057, n16058, n16059, n16060, n16061, n16062, n16064, n16065, n16066,
    n16068, n16069, n16070, n16072, n16073, n16074, n16076, n16077, n16078,
    n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
    n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
    n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
    n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
    n16115, n16116, n16117, n16118, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
    n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16142, n16143,
    n16144, n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
    n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
    n16163, n16164, n16165, n16166, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16190, n16191,
    n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
    n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
    n16210, n16212, n16213, n16214, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
    n16249, n16250, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
    n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
    n16268, n16269, n16270, n16271, n16272, n16274, n16275, n16276, n16277,
    n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16296,
    n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
    n16315, n16316, n16318, n16319, n16320, n16321, n16322, n16323, n16324,
    n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
    n16334, n16335, n16336, n16337, n16338, n16340, n16341, n16342, n16343,
    n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16362,
    n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
    n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16380, n16381,
    n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389, n16390,
    n16391, n16392, n16393, n16394, n16395, n16396, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
    n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
    n16420, n16421, n16422, n16424, n16425, n16426, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
    n16440, n16441, n16442, n16443, n16444, n16447, n16448, n16449, n16451,
    n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
    n16470, n16471, n16473, n16474, n16475, n16477, n16478, n16479, n16481,
    n16482, n16483, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
    n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16507, n16508, n16509, n16511,
    n16512, n16513, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
    n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
    n16531, n16532, n16533, n16534, n16535, n16537, n16538, n16539, n16541,
    n16542, n16543, n16545, n16546, n16547, n16549, n16550, n16551, n16553,
    n16554, n16555, n16557, n16558, n16559, n16561, n16562, n16563, n16565,
    n16566, n16567, n16569, n16570, n16571, n16573, n16574, n16575, n16577,
    n16578, n16579, n16581, n16582, n16583, n16585, n16586, n16587, n16589,
    n16590, n16591, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
    n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
    n16609, n16610, n16611, n16613, n16614, n16615, n16616, n16617, n16618,
    n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
    n16628, n16629, n16630, n16631, n16633, n16634, n16635, n16637, n16638,
    n16639, n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
    n16658, n16659, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
    n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16681, n16682, n16683, n16684, n16685, n16686,
    n16687, n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
    n16696, n16697, n16698, n16699, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16723, n16724,
    n16725, n16727, n16728, n16729, n16730, n16731, n16732, n16733, n16734,
    n16735, n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
    n16744, n16745, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
    n16782, n16783, n16784, n16785, n16786, n16787, n16789, n16790, n16791,
    n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
    n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
    n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
    n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
    n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
    n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
    n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16907, n16908, n16909, n16911, n16912, n16913, n16915, n16916,
    n16917, n16919, n16920, n16921, n16923, n16924, n16925, n16927, n16928,
    n16929, n16931, n16932, n16933, n16935, n16936, n16937, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16947, n16948, n16949, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
    n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
    n16971, n16972, n16973, n16975, n16976, n16977, n16979, n16980, n16981,
    n16983, n16984, n16985, n16987, n16988, n16989, n16992, n16993, n16994,
    n16996, n16997, n16998, n17000, n17001, n17002, n17004, n17005, n17006,
    n17008, n17009, n17010, n17012, n17013, n17014, n17016, n17017, n17018,
    n17020, n17021, n17022, n17023, n17024, n17026, n17027, n17028, n17030,
    n17031, n17032, n17034, n17035, n17036, n17038, n17039, n17040, n17042,
    n17043, n17044, n17046, n17047, n17048, n17050, n17051, n17052, n17054,
    n17055, n17056, n17058, n17059, n17060, n17062, n17063, n17064, n17066,
    n17067, n17068, n17070, n17071, n17072, n17074, n17075, n17076, n17078,
    n17079, n17080, n17082, n17083, n17084, n17086, n17087, n17088, n17090,
    n17091, n17092, n17094, n17095, n17096, n17098, n17099, n17100, n17102,
    n17103, n17104, n17106, n17107, n17108, n17110, n17111, n17112, n17113,
    n17114, n17115, n17116, n17117, n17118, n17120, n17121, n17122, n17124,
    n17125, n17126, n17127, n17128, n17129, n17131, n17132, n17133, n17135,
    n17136, n17137, n17138, n17139, n17141, n17142, n17143, n17145, n17146,
    n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17155, n17156,
    n17157, n17159, n17160, n17161, n17163, n17164, n17165, n17166, n17167,
    n17168, n17169, n17173, n17174, n17176, n17177, n17179, n17180, n17182,
    n17183, n17185, n17186, n17188, n17189, n17191, n17192, n17194, n17195,
    n17197, n17198, n17200, n17201, n17203, n17204, n17206, n17207, n17209,
    n17210, n17211, n17212, n17214, n17215, n17217, n17218, n17219, n17220,
    n17221, n17222, n17223, n17224, n17225, n17226, n17228, n17229, n17231,
    n17232, n17234, n17235, n17237, n17238, n17240, n17241, n17242, n17243,
    n17244, n17245, n17247, n17248, n17250, n17251, n17253, n17254, n17256,
    n17257, n17259, n17260, n17262, n17263, n17265, n17266, n17268, n17269,
    n17271, n17272, n17274, n17275, n17277, n17278, n17280, n17281, n17283,
    n17284, n17286, n17287, n17289, n17290, n17291, n17292, n17293, n17294,
    n17296, n17297, n17298, n17301, n17302, n17303, n17305, n17306, n17307,
    n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315, n17316,
    n17317, n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
    n17326, n17327, n17328, n17330, n17331, n17332, n17333, n17334, n17335,
    n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
    n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
    n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17378, n17379, n17380, n17381, n17382,
    n17383, n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
    n17402, n17403, n17405, n17406, n17407, n17409, n17410, n17412, n17415,
    n17416, n17418, n17419, n17421, n17422, n17424, n17425, n17427, n17428,
    n17430, n17431, n17433, n17434, n17436, n17437, n17439, n17440, n17442,
    n17443, n17445, n17446, n17448, n17449, n17451, n17452, n17454, n17455,
    n17457, n17458, n17460, n17461, n17463, n17464, n17466, n17467, n17469,
    n17470, n17472, n17473, n17475, n17476, n17478, n17479, n17481, n17482,
    n17484, n17485, n17487, n17488, n17490, n17491, n17493, n17494, n17496,
    n17497, n17499, n17500, n17502, n17503, n17505, n17506, n17508, n17509,
    n17511, n17512, n17514, n17515, n17517, n17518, n17520, n17521, n17523,
    n17524, n17526, n17527, n17529, n17530, n17532, n17533, n17535, n17536,
    n17538, n17539, n17541, n17542, n17544, n17545, n17547, n17548, n17550,
    n17551, n17553, n17554, n17556, n17557, n17559, n17560, n17562, n17563,
    n17565, n17566, n17568, n17569, n17571, n17572, n17574, n17575, n17577,
    n17578, n17580, n17581, n17583, n17584, n17586, n17587, n17589, n17590,
    n17592, n17593, n17595, n17596, n17598, n17599, n17601, n17602, n17604,
    n17605, n17607, n17608, n17610, n17611, n17613, n17614, n17615, n17616,
    n17617, n17618, n17619, n17620, n17621, n17623, n17624, n17626, n17627,
    n17629, n17630, n17632, n17633, n17635, n17636, n17638, n17639, n17641,
    n17642, n17644, n17645, n17647, n17648, n17650, n17651, n17653, n17654,
    n17656, n17657, n17659, n17660, n17662, n17663, n17665, n17666, n17668,
    n17669, n17671, n17673, n17674, n17676, n17677, n17679, n17680, n17682,
    n17683, n17685, n17686, n17688, n17689, n17691, n17692, n17694, n17695,
    n17697, n17698, n17700, n17701, n17703, n17704, n17706, n17707, n17709,
    n17710, n17712, n17713, n17715, n17716, n17718, n17719, n17721, n17722,
    n17724, n17725, n17727, n17728, n17730, n17731, n17734, n17735, n17737,
    n17738, n17740, n17741, n17743, n17745, n17746;
  assign n2425 = ~pi0056 & ~pi0062;
  assign n2426 = ~pi0057 & ~pi0059;
  assign n2427 = ~pi0055 & ~pi0299;
  assign n2428 = n2426 & n2427;
  assign n2429 = n2425 & n2428;
  assign n2430 = pi0224 & n2429;
  assign n2431 = pi0216 & ~n2429;
  assign n2432 = ~n2430 & ~n2431;
  assign n2433 = pi0222 & n2429;
  assign n2434 = pi0221 & ~n2429;
  assign n2435 = ~n2433 & ~n2434;
  assign n2436 = pi0215 & ~n2429;
  assign n2437 = pi0223 & n2429;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = n2435 & n2438;
  assign n2440 = ~n2432 & n2439;
  assign n2441 = ~pi0265 & n2440;
  assign n2442 = ~pi0153 & ~n2429;
  assign n2443 = ~pi0175 & n2429;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = ~pi0045 & ~pi0053;
  assign n2446 = ~pi0054 & ~pi0106;
  assign n2447 = n2445 & n2446;
  assign n2448 = ~pi0055 & ~pi0057;
  assign n2449 = n2425 & n2448;
  assign n2450 = n2447 & n2449;
  assign n2451 = ~pi0064 & ~pi0065;
  assign n2452 = ~pi0063 & ~pi0107;
  assign n2453 = n2451 & n2452;
  assign n2454 = ~pi0046 & ~pi0061;
  assign n2455 = ~pi0059 & ~pi0060;
  assign n2456 = n2454 & n2455;
  assign n2457 = n2453 & n2456;
  assign n2458 = n2450 & n2457;
  assign n2459 = ~pi0095 & ~pi0097;
  assign n2460 = ~pi0074 & ~pi0096;
  assign n2461 = n2459 & n2460;
  assign n2462 = ~pi0035 & ~pi0070;
  assign n2463 = ~pi0089 & ~pi0108;
  assign n2464 = n2462 & n2463;
  assign n2465 = n2461 & n2464;
  assign n2466 = ~pi0032 & ~pi0038;
  assign n2467 = ~pi0050 & ~pi0100;
  assign n2468 = ~pi0049 & ~pi0076;
  assign n2469 = ~pi0075 & ~pi0094;
  assign n2470 = n2468 & n2469;
  assign n2471 = n2467 & n2470;
  assign n2472 = n2466 & n2471;
  assign n2473 = n2465 & n2472;
  assign n2474 = n2458 & n2473;
  assign n2475 = ~pi0039 & ~pi0048;
  assign n2476 = ~pi0067 & ~pi0071;
  assign n2477 = ~pi0083 & ~pi0085;
  assign n2478 = n2476 & n2477;
  assign n2479 = ~pi0066 & ~pi0082;
  assign n2480 = ~pi0051 & ~pi0084;
  assign n2481 = n2479 & n2480;
  assign n2482 = ~pi0040 & ~pi0081;
  assign n2483 = ~pi0068 & ~pi0102;
  assign n2484 = n2482 & n2483;
  assign n2485 = n2481 & n2484;
  assign n2486 = ~pi0077 & ~pi0086;
  assign n2487 = ~pi0069 & ~pi0109;
  assign n2488 = n2486 & n2487;
  assign n2489 = n2485 & n2488;
  assign n2490 = n2478 & n2489;
  assign n2491 = n2475 & n2490;
  assign n2492 = n2474 & n2491;
  assign n2493 = ~pi0092 & ~pi0093;
  assign n2494 = ~pi0087 & ~pi0111;
  assign n2495 = ~pi0072 & ~pi0103;
  assign n2496 = n2494 & n2495;
  assign n2497 = ~pi0088 & ~pi0104;
  assign n2498 = ~pi0047 & ~pi0110;
  assign n2499 = n2497 & n2498;
  assign n2500 = n2496 & n2499;
  assign n2501 = ~pi0073 & ~pi0090;
  assign n2502 = ~pi0036 & ~pi0091;
  assign n2503 = n2501 & n2502;
  assign n2504 = pi0058 & n2503;
  assign n2505 = n2500 & n2504;
  assign n2506 = ~pi0098 & n2505;
  assign n2507 = n2493 & n2506;
  assign n2508 = n2492 & n2507;
  assign n2509 = n2496 & n2503;
  assign n2510 = ~pi0058 & ~pi0098;
  assign n2511 = n2493 & n2510;
  assign n2512 = n2498 & n2511;
  assign n2513 = n2509 & n2512;
  assign n2514 = ~pi0088 & n2513;
  assign n2515 = pi0104 & n2514;
  assign n2516 = n2492 & n2515;
  assign n2517 = ~n2508 & ~n2516;
  assign n2518 = n2503 & n2511;
  assign n2519 = n2475 & n2500;
  assign n2520 = n2518 & n2519;
  assign n2521 = n2458 & n2520;
  assign n2522 = n2473 & n2521;
  assign n2523 = n2488 & n2522;
  assign n2524 = n2485 & n2523;
  assign n2525 = ~pi0071 & n2524;
  assign n2526 = n2477 & n2525;
  assign n2527 = pi0067 & n2526;
  assign n2528 = n2476 & n2485;
  assign n2529 = ~pi0085 & n2528;
  assign n2530 = n2474 & n2520;
  assign n2531 = pi0083 & n2488;
  assign n2532 = n2530 & n2531;
  assign n2533 = n2529 & n2532;
  assign n2534 = ~n2527 & ~n2533;
  assign n2535 = ~pi0067 & pi0071;
  assign n2536 = n2477 & n2535;
  assign n2537 = n2524 & n2536;
  assign n2538 = ~pi0083 & n2488;
  assign n2539 = n2473 & n2520;
  assign n2540 = n2458 & n2539;
  assign n2541 = pi0085 & n2476;
  assign n2542 = n2485 & n2541;
  assign n2543 = n2540 & n2542;
  assign n2544 = n2538 & n2543;
  assign n2545 = ~n2537 & ~n2544;
  assign n2546 = n2534 & n2545;
  assign n2547 = n2517 & n2546;
  assign n2548 = n2450 & n2456;
  assign n2549 = n2473 & n2548;
  assign n2550 = n2500 & n2518;
  assign n2551 = n2490 & n2550;
  assign n2552 = n2475 & n2551;
  assign po1049 = pi0064 | ~n2452;
  assign n2554 = n2552 & ~po1049;
  assign n2555 = pi0065 & n2554;
  assign n2556 = n2549 & n2555;
  assign n2557 = ~pi0228 & ~n2556;
  assign n2558 = n2547 & n2557;
  assign n2559 = ~pi0036 & n2501;
  assign n2560 = pi0091 & n2511;
  assign n2561 = n2492 & n2560;
  assign n2562 = n2500 & n2561;
  assign n2563 = n2559 & n2562;
  assign n2564 = n2499 & n2503;
  assign n2565 = pi0072 & ~pi0103;
  assign n2566 = n2564 & n2565;
  assign n2567 = n2494 & n2511;
  assign n2568 = n2492 & n2567;
  assign n2569 = n2566 & n2568;
  assign n2570 = ~n2563 & ~n2569;
  assign n2571 = pi0063 & ~pi0107;
  assign n2572 = n2450 & n2552;
  assign n2573 = n2473 & n2572;
  assign n2574 = n2451 & n2456;
  assign n2575 = n2573 & n2574;
  assign n2576 = n2571 & n2575;
  assign n2577 = pi0056 & ~pi0062;
  assign n2578 = n2448 & n2453;
  assign n2579 = n2447 & n2552;
  assign n2580 = n2456 & n2579;
  assign n2581 = n2473 & n2580;
  assign n2582 = n2578 & n2581;
  assign n2583 = n2577 & n2582;
  assign n2584 = ~n2576 & ~n2583;
  assign n2585 = n2570 & n2584;
  assign n2586 = n2558 & n2585;
  assign n2587 = ~pi0057 & n2425;
  assign n2588 = n2473 & n2587;
  assign n2589 = n2453 & n2588;
  assign n2590 = pi0055 & n2589;
  assign n2591 = n2580 & n2590;
  assign n2592 = n2449 & n2456;
  assign n2593 = n2552 & n2592;
  assign n2594 = ~pi0045 & n2446;
  assign n2595 = n2453 & n2594;
  assign n2596 = pi0053 & n2595;
  assign n2597 = n2473 & n2596;
  assign n2598 = n2593 & n2597;
  assign n2599 = ~n2591 & ~n2598;
  assign n2600 = ~pi0047 & n2511;
  assign n2601 = n2509 & n2600;
  assign n2602 = pi0110 & n2601;
  assign n2603 = n2497 & n2602;
  assign n2604 = n2492 & n2603;
  assign n2605 = n2462 & n2468;
  assign n2606 = n2469 & n2605;
  assign n2607 = n2466 & n2467;
  assign n2608 = n2490 & n2520;
  assign n2609 = n2458 & n2608;
  assign n2610 = n2607 & n2609;
  assign n2611 = n2461 & n2610;
  assign n2612 = pi0108 & n2611;
  assign n2613 = ~pi0089 & n2612;
  assign n2614 = n2606 & n2613;
  assign n2615 = n2503 & n2510;
  assign n2616 = n2500 & n2615;
  assign n2617 = ~pi0093 & n2616;
  assign n2618 = pi0092 & n2617;
  assign n2619 = n2492 & n2618;
  assign n2620 = ~n2614 & ~n2619;
  assign n2621 = ~n2604 & n2620;
  assign n2622 = ~pi0110 & n2497;
  assign n2623 = n2509 & n2622;
  assign n2624 = n2511 & n2623;
  assign n2625 = pi0047 & n2624;
  assign n2626 = n2492 & n2625;
  assign n2627 = n2484 & n2488;
  assign n2628 = n2478 & n2479;
  assign n2629 = n2627 & n2628;
  assign n2630 = ~pi0084 & n2629;
  assign n2631 = pi0051 & n2630;
  assign n2632 = n2530 & n2631;
  assign n2633 = n2478 & n2486;
  assign n2634 = n2485 & n2633;
  assign n2635 = pi0109 & n2634;
  assign n2636 = ~pi0069 & n2635;
  assign n2637 = n2530 & n2636;
  assign n2638 = ~n2632 & ~n2637;
  assign n2639 = ~pi0054 & pi0106;
  assign n2640 = n2473 & n2639;
  assign n2641 = n2592 & n2640;
  assign n2642 = n2445 & n2552;
  assign n2643 = n2453 & n2642;
  assign n2644 = n2641 & n2643;
  assign n2645 = n2638 & ~n2644;
  assign n2646 = ~pi0095 & pi0097;
  assign n2647 = n2464 & n2607;
  assign n2648 = n2609 & n2647;
  assign n2649 = n2470 & n2648;
  assign n2650 = n2460 & n2649;
  assign n2651 = n2646 & n2650;
  assign n2652 = ~pi0086 & n2478;
  assign n2653 = n2485 & n2487;
  assign n2654 = n2530 & n2653;
  assign n2655 = n2652 & n2654;
  assign n2656 = pi0077 & n2655;
  assign n2657 = ~n2651 & ~n2656;
  assign n2658 = pi0111 & n2511;
  assign n2659 = n2564 & n2658;
  assign n2660 = ~pi0087 & n2659;
  assign n2661 = n2495 & n2660;
  assign n2662 = n2492 & n2661;
  assign n2663 = pi0098 & n2493;
  assign n2664 = n2492 & n2500;
  assign n2665 = ~pi0058 & n2503;
  assign n2666 = n2664 & n2665;
  assign n2667 = n2663 & n2666;
  assign n2668 = ~n2662 & ~n2667;
  assign n2669 = n2657 & n2668;
  assign n2670 = n2645 & n2669;
  assign n2671 = ~n2626 & n2670;
  assign n2672 = n2621 & n2671;
  assign n2673 = n2599 & n2672;
  assign n2674 = n2481 & n2488;
  assign n2675 = ~pi0068 & n2478;
  assign n2676 = n2674 & n2675;
  assign n2677 = n2482 & n2676;
  assign n2678 = pi0102 & n2677;
  assign n2679 = n2540 & n2678;
  assign n2680 = pi0095 & n2650;
  assign n2681 = ~pi0097 & n2680;
  assign n2682 = pi0032 & ~pi0038;
  assign n2683 = n2465 & n2609;
  assign n2684 = n2471 & n2683;
  assign n2685 = n2682 & n2684;
  assign n2686 = ~n2681 & ~n2685;
  assign n2687 = ~n2679 & n2686;
  assign n2688 = n2673 & n2687;
  assign n2689 = n2586 & n2688;
  assign n2690 = ~pi0066 & n2478;
  assign n2691 = n2627 & n2690;
  assign n2692 = n2480 & n2691;
  assign n2693 = pi0082 & n2692;
  assign n2694 = n2530 & n2693;
  assign n2695 = n2458 & n2551;
  assign n2696 = n2473 & n2695;
  assign n2697 = ~pi0039 & pi0048;
  assign n2698 = n2696 & n2697;
  assign n2699 = ~n2694 & ~n2698;
  assign n2700 = pi0142 & n2429;
  assign n2701 = pi0146 & ~n2429;
  assign n2702 = ~n2700 & ~n2701;
  assign n2703 = pi0152 & ~n2429;
  assign n2704 = pi0174 & n2429;
  assign n2705 = ~n2703 & ~n2704;
  assign n2706 = n2427 & n2587;
  assign n2707 = ~pi0059 & n2706;
  assign n2708 = pi0144 & n2707;
  assign n2709 = pi0161 & ~n2429;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2705 & n2710;
  assign n2712 = pi0189 & n2707;
  assign n2713 = pi0166 & ~n2707;
  assign n2714 = ~n2712 & ~n2713;
  assign n2715 = n2711 & n2714;
  assign n2716 = n2702 & ~n2715;
  assign n2717 = pi0252 & ~n2716;
  assign n2718 = ~pi0250 & n2716;
  assign n2719 = pi0129 & ~n2718;
  assign po1135 = pi0824 & pi1086;
  assign n2721 = pi1086 & pi1087;
  assign n2722 = pi0957 & pi1085;
  assign n2723 = ~pi0833 & n2722;
  assign po1106 = n2721 & n2723;
  assign n2725 = pi0950 & ~po1106;
  assign n2726 = po1135 & n2725;
  assign n2727 = ~pi1085 & pi1087;
  assign n2728 = pi0829 & pi1086;
  assign po1107 = ~n2727 & n2728;
  assign n2730 = pi0950 & po1107;
  assign po0840 = ~po1106 & n2730;
  assign po0950 = ~n2726 & ~po0840;
  assign n2733 = pi1086 & ~pi1087;
  assign po0740 = ~po0950 & n2733;
  assign n2735 = n2718 & ~po0740;
  assign n2736 = ~n2719 & ~n2735;
  assign n2737 = pi0100 & n2470;
  assign n2738 = ~pi0050 & n2737;
  assign n2739 = n2466 & n2683;
  assign n2740 = n2738 & n2739;
  assign n2741 = n2736 & n2740;
  assign n2742 = ~n2717 & n2741;
  assign n2743 = pi0064 & ~pi0065;
  assign n2744 = n2548 & n2552;
  assign n2745 = n2473 & n2744;
  assign n2746 = n2452 & n2745;
  assign n2747 = n2743 & n2746;
  assign n2748 = ~n2742 & ~n2747;
  assign n2749 = ~pi0252 & ~n2716;
  assign n2750 = ~n2736 & ~n2749;
  assign n2751 = ~pi0115 & ~pi0116;
  assign n2752 = ~pi0099 & ~pi0113;
  assign n2753 = n2751 & n2752;
  assign n2754 = ~pi0044 & n2753;
  assign n2755 = ~pi0042 & ~pi0043;
  assign n2756 = ~pi0041 & n2755;
  assign n2757 = ~pi0052 & n2756;
  assign n2758 = ~pi0114 & n2757;
  assign n2759 = ~pi0101 & n2758;
  assign po1057 = ~n2754 | ~n2759;
  assign n2761 = pi0683 & po1057;
  assign n2762 = ~pi0332 & ~pi0468;
  assign n2763 = pi0232 & n2762;
  assign n2764 = n2714 & n2763;
  assign n2765 = n2711 & n2764;
  assign n2766 = pi0089 & n2606;
  assign n2767 = n2461 & n2607;
  assign n2768 = ~pi0108 & n2767;
  assign n2769 = n2609 & n2768;
  assign n2770 = n2766 & n2769;
  assign n2771 = pi0070 & n2470;
  assign n2772 = n2463 & n2771;
  assign n2773 = ~pi0035 & n2772;
  assign n2774 = n2611 & n2773;
  assign n2775 = ~n2770 & ~n2774;
  assign n2776 = pi0039 & ~pi0048;
  assign n2777 = n2696 & n2776;
  assign n2778 = ~n2770 & ~n2777;
  assign n2779 = pi0332 & n2778;
  assign n2780 = ~n2775 & n2779;
  assign n2781 = pi0287 & n2775;
  assign n2782 = pi0332 & ~n2775;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = ~n2778 & ~n2783;
  assign n2785 = ~pi0032 & n2471;
  assign n2786 = pi0038 & n2465;
  assign n2787 = n2785 & n2786;
  assign n2788 = n2609 & n2787;
  assign n2789 = pi0046 & n2455;
  assign n2790 = ~pi0061 & n2453;
  assign n2791 = n2473 & n2790;
  assign n2792 = n2789 & n2791;
  assign n2793 = n2450 & n2475;
  assign n2794 = n2792 & n2793;
  assign n2795 = n2551 & n2794;
  assign n2796 = ~n2788 & ~n2795;
  assign n2797 = n2778 & ~n2796;
  assign n2798 = n2775 & n2797;
  assign n2799 = ~n2784 & ~n2798;
  assign n2800 = ~n2780 & n2799;
  assign n2801 = n2765 & n2800;
  assign n2802 = n2716 & ~n2801;
  assign n2803 = n2761 & n2802;
  assign n2804 = n2717 & ~n2803;
  assign n2805 = n2750 & ~n2804;
  assign n2806 = ~n2717 & ~n2736;
  assign n2807 = n2749 & n2806;
  assign n2808 = ~n2805 & ~n2807;
  assign n2809 = n2740 & ~n2808;
  assign n2810 = pi0094 & n2468;
  assign n2811 = ~pi0075 & n2810;
  assign n2812 = n2607 & n2683;
  assign n2813 = n2811 & n2812;
  assign n2814 = ~n2809 & ~n2813;
  assign n2815 = n2748 & n2814;
  assign n2816 = n2699 & n2815;
  assign n2817 = n2502 & n2511;
  assign n2818 = n2500 & n2817;
  assign n2819 = n2458 & n2818;
  assign n2820 = ~pi0073 & pi0090;
  assign n2821 = n2473 & n2820;
  assign n2822 = n2491 & n2821;
  assign n2823 = n2819 & n2822;
  assign n2824 = pi0093 & n2616;
  assign n2825 = ~pi0092 & n2824;
  assign n2826 = n2492 & n2825;
  assign n2827 = ~n2823 & ~n2826;
  assign n2828 = ~pi0070 & n2470;
  assign n2829 = n2463 & n2828;
  assign n2830 = pi0035 & n2829;
  assign n2831 = n2611 & n2830;
  assign n2832 = pi0073 & ~pi0090;
  assign n2833 = n2664 & n2817;
  assign n2834 = n2832 & n2833;
  assign n2835 = ~n2831 & ~n2834;
  assign n2836 = n2827 & n2835;
  assign n2837 = pi0045 & n2446;
  assign n2838 = ~pi0053 & n2453;
  assign n2839 = n2473 & n2593;
  assign n2840 = n2838 & n2839;
  assign n2841 = n2837 & n2840;
  assign n2842 = n2836 & ~n2841;
  assign n2843 = pi0049 & n2461;
  assign n2844 = n2609 & n2843;
  assign n2845 = n2469 & n2844;
  assign n2846 = ~pi0076 & n2845;
  assign n2847 = n2647 & n2846;
  assign n2848 = ~pi0072 & pi0103;
  assign n2849 = n2564 & n2848;
  assign n2850 = n2492 & n2849;
  assign n2851 = n2567 & n2850;
  assign n2852 = ~pi0035 & n2771;
  assign n2853 = n2611 & n2852;
  assign n2854 = n2463 & n2853;
  assign n2855 = ~pi0074 & n2470;
  assign n2856 = pi0096 & n2855;
  assign n2857 = n2459 & n2648;
  assign n2858 = n2856 & n2857;
  assign n2859 = ~n2854 & ~n2858;
  assign n2860 = ~n2851 & n2859;
  assign n2861 = ~n2847 & n2860;
  assign n2862 = ~pi0051 & pi0084;
  assign n2863 = n2479 & n2862;
  assign n2864 = n2473 & n2478;
  assign n2865 = n2521 & n2864;
  assign n2866 = n2627 & n2865;
  assign n2867 = n2863 & n2866;
  assign n2868 = ~pi0082 & n2480;
  assign n2869 = n2627 & n2868;
  assign n2870 = pi0066 & n2869;
  assign n2871 = n2478 & n2870;
  assign n2872 = n2530 & n2871;
  assign n2873 = ~n2867 & ~n2872;
  assign n2874 = ~pi0102 & n2482;
  assign n2875 = pi0068 & n2478;
  assign n2876 = n2530 & n2875;
  assign n2877 = n2674 & n2876;
  assign n2878 = n2874 & n2877;
  assign n2879 = ~pi0104 & n2513;
  assign n2880 = pi0088 & n2492;
  assign n2881 = n2879 & n2880;
  assign n2882 = ~n2878 & ~n2881;
  assign n2883 = n2873 & n2882;
  assign n2884 = n2861 & n2883;
  assign n2885 = ~pi0091 & n2511;
  assign n2886 = pi0036 & n2501;
  assign n2887 = n2664 & n2886;
  assign n2888 = n2885 & n2887;
  assign n2889 = ~pi0046 & n2455;
  assign n2890 = pi0061 & n2453;
  assign n2891 = n2573 & n2890;
  assign n2892 = n2889 & n2891;
  assign n2893 = ~pi0063 & pi0107;
  assign n2894 = n2573 & n2893;
  assign n2895 = n2574 & n2894;
  assign n2896 = ~n2892 & ~n2895;
  assign n2897 = n2478 & n2483;
  assign n2898 = n2674 & n2897;
  assign n2899 = ~pi0040 & n2898;
  assign n2900 = pi0081 & n2899;
  assign n2901 = n2530 & n2900;
  assign n2902 = n2896 & ~n2901;
  assign n2903 = ~n2888 & n2902;
  assign n2904 = n2778 & n2903;
  assign n2905 = n2453 & n2454;
  assign n2906 = ~pi0059 & pi0060;
  assign n2907 = n2552 & n2906;
  assign n2908 = n2473 & n2907;
  assign n2909 = n2905 & n2908;
  assign n2910 = n2450 & n2909;
  assign n2911 = pi0050 & ~pi0100;
  assign n2912 = n2470 & n2911;
  assign n2913 = n2739 & n2912;
  assign n2914 = ~pi0056 & pi0062;
  assign n2915 = n2578 & n2580;
  assign n2916 = n2473 & n2915;
  assign n2917 = n2914 & n2916;
  assign n2918 = pi0087 & n2495;
  assign n2919 = ~pi0111 & n2511;
  assign n2920 = n2564 & n2919;
  assign n2921 = n2918 & n2920;
  assign n2922 = n2492 & n2921;
  assign n2923 = ~n2917 & ~n2922;
  assign n2924 = ~pi0081 & n2898;
  assign n2925 = pi0040 & n2530;
  assign n2926 = n2924 & n2925;
  assign n2927 = n2923 & ~n2926;
  assign n2928 = pi0076 & n2469;
  assign n2929 = ~pi0049 & n2928;
  assign n2930 = n2812 & n2929;
  assign n2931 = n2927 & ~n2930;
  assign n2932 = ~n2913 & n2931;
  assign n2933 = ~n2910 & n2932;
  assign n2934 = ~pi0109 & n2634;
  assign n2935 = pi0069 & n2934;
  assign n2936 = n2530 & n2935;
  assign n2937 = pi0086 & n2478;
  assign n2938 = n2485 & n2937;
  assign n2939 = n2487 & n2938;
  assign n2940 = ~pi0077 & n2939;
  assign n2941 = n2530 & n2940;
  assign n2942 = ~n2936 & ~n2941;
  assign n2943 = n2933 & n2942;
  assign n2944 = n2904 & n2943;
  assign n2945 = n2884 & n2944;
  assign n2946 = n2842 & n2945;
  assign n2947 = n2816 & n2946;
  assign n2948 = n2689 & n2947;
  assign n2949 = ~pi0105 & pi0228;
  assign po0183 = ~n2948 & ~n2949;
  assign n2951 = ~n2444 & ~po0183;
  assign n2952 = ~n2429 & n2951;
  assign n2953 = pi0095 & ~pi0479;
  assign n2954 = ~pi0049 & ~pi0094;
  assign n2955 = ~pi0074 & ~pi0097;
  assign n2956 = ~pi0075 & ~pi0076;
  assign n2957 = ~pi0058 & ~pi0092;
  assign n2958 = ~pi0093 & ~pi0098;
  assign n2959 = n2957 & n2958;
  assign n2960 = n2956 & n2959;
  assign n2961 = n2955 & n2960;
  assign n2962 = ~pi0089 & ~pi0095;
  assign n2963 = ~pi0048 & n2962;
  assign n2964 = pi0096 & n2963;
  assign n2965 = n2961 & n2964;
  assign n2966 = ~pi0039 & ~pi0108;
  assign n2967 = n2462 & n2966;
  assign n2968 = n2965 & n2967;
  assign n2969 = ~pi0095 & n2968;
  assign n2970 = n2954 & n2969;
  assign n2971 = ~pi0071 & ~pi0085;
  assign n2972 = ~pi0067 & ~pi0083;
  assign n2973 = n2971 & n2972;
  assign n2974 = ~pi0068 & ~pi0081;
  assign n2975 = n2973 & n2974;
  assign n2976 = ~pi0065 & n2975;
  assign n2977 = ~po1049 & n2976;
  assign n2978 = ~pi0040 & ~pi0102;
  assign n2979 = n2481 & n2978;
  assign n2980 = ~pi0056 & ~pi0057;
  assign n2981 = ~pi0055 & ~pi0059;
  assign n2982 = ~pi0062 & n2981;
  assign n2983 = ~pi0060 & n2454;
  assign n2984 = n2982 & n2983;
  assign n2985 = n2447 & n2984;
  assign n2986 = n2980 & n2985;
  assign n2987 = ~pi0032 & ~pi0050;
  assign n2988 = n2986 & n2987;
  assign n2989 = n2979 & n2988;
  assign n2990 = ~pi0100 & n2989;
  assign n2991 = ~pi0038 & n2990;
  assign n2992 = ~pi0072 & ~pi0111;
  assign n2993 = ~pi0069 & ~pi0086;
  assign n2994 = ~pi0077 & ~pi0109;
  assign n2995 = n2993 & n2994;
  assign n2996 = ~pi0087 & ~pi0103;
  assign n2997 = n2995 & n2996;
  assign n2998 = ~pi0104 & ~pi0110;
  assign n2999 = ~pi0088 & n2998;
  assign n3000 = ~pi0047 & n2999;
  assign n3001 = n2997 & n3000;
  assign n3002 = n2503 & n3001;
  assign n3003 = n2992 & n3002;
  assign n3004 = n2991 & n3003;
  assign n3005 = n2977 & n3004;
  assign n3006 = n2970 & n3005;
  assign n3007 = ~n2953 & ~n3006;
  assign n3008 = pi0234 & ~n3007;
  assign n3009 = ~n2556 & ~n2679;
  assign n3010 = ~n2576 & ~n2795;
  assign n3011 = n3009 & n3010;
  assign n3012 = ~n2583 & ~n2813;
  assign n3013 = n3011 & n3012;
  assign n3014 = pi0137 & ~n3013;
  assign n3015 = pi0137 & n2747;
  assign n3016 = pi0198 & n2707;
  assign n3017 = pi0210 & ~n2707;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~n2716 & n3018;
  assign n3020 = ~pi0137 & ~n3019;
  assign n3021 = n2740 & ~n3020;
  assign n3022 = ~n3015 & ~n3021;
  assign n3023 = ~n2563 & ~n2694;
  assign n3024 = ~n2698 & n3023;
  assign n3025 = ~n2569 & n3024;
  assign n3026 = pi0137 & ~n3025;
  assign n3027 = n3022 & ~n3026;
  assign n3028 = ~n2930 & ~n2936;
  assign n3029 = ~n2922 & n3028;
  assign n3030 = pi0057 & n2425;
  assign n3031 = ~pi0055 & n2453;
  assign n3032 = n2581 & n3031;
  assign n3033 = n3030 & n3032;
  assign n3034 = n3029 & ~n3033;
  assign n3035 = ~n2917 & ~n2926;
  assign n3036 = n3034 & n3035;
  assign n3037 = n2547 & n3036;
  assign n3038 = ~n2913 & n3037;
  assign n3039 = pi0137 & ~n3038;
  assign n3040 = ~pi0094 & n2468;
  assign n3041 = pi0075 & n3040;
  assign n3042 = n2812 & n3041;
  assign n3043 = ~n3020 & n3042;
  assign n3044 = pi0137 & n2941;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = ~n3039 & n3045;
  assign n3047 = ~n2910 & n3046;
  assign n3048 = ~n2681 & n2896;
  assign n3049 = ~n2901 & n3048;
  assign n3050 = pi0137 & ~n3049;
  assign n3051 = n3047 & ~n3050;
  assign n3052 = pi0225 & n2831;
  assign n3053 = ~pi0841 & ~n3018;
  assign n3054 = pi0225 & n3053;
  assign n3055 = n2685 & n3054;
  assign n3056 = ~n3052 & ~n3055;
  assign n3057 = ~pi0841 & n3018;
  assign n3058 = ~n3053 & ~n3057;
  assign n3059 = n2685 & n3058;
  assign n3060 = pi0225 & n3059;
  assign n3061 = pi0137 & ~n2873;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n3056 & n3062;
  assign n3064 = pi0059 & ~pi0060;
  assign n3065 = n2573 & n3064;
  assign n3066 = n2905 & n3065;
  assign n3067 = ~n2851 & ~n3066;
  assign n3068 = pi0137 & ~n3067;
  assign n3069 = n2470 & n2857;
  assign n3070 = ~pi0096 & n3069;
  assign n3071 = pi0074 & n3070;
  assign n3072 = ~n2788 & ~n3071;
  assign n3073 = ~n2841 & ~n2847;
  assign n3074 = n3072 & n3073;
  assign n3075 = ~n2826 & ~n2878;
  assign n3076 = ~n2881 & n3075;
  assign n3077 = ~n2834 & n3076;
  assign n3078 = n3074 & n3077;
  assign n3079 = pi0137 & ~n3078;
  assign n3080 = pi0332 & n2854;
  assign n3081 = pi0137 & n2823;
  assign n3082 = ~n3080 & ~n3081;
  assign n3083 = ~pi0137 & pi0841;
  assign n3084 = po0840 & ~n3020;
  assign n3085 = pi0137 & ~po0840;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = ~pi0841 & n3086;
  assign n3088 = ~n3083 & ~n3087;
  assign n3089 = n2858 & n3088;
  assign n3090 = n3082 & ~n3089;
  assign n3091 = ~n3079 & n3090;
  assign n3092 = ~n3068 & n3091;
  assign n3093 = n3063 & n3092;
  assign n3094 = n2778 & ~n2888;
  assign n3095 = pi0137 & ~n3094;
  assign n3096 = n3093 & ~n3095;
  assign n3097 = n3051 & n3096;
  assign n3098 = n3027 & n3097;
  assign n3099 = ~n3014 & n3098;
  assign n3100 = ~n2637 & ~n2644;
  assign n3101 = pi0137 & ~n3100;
  assign n3102 = po0840 & ~po0740;
  assign n3103 = ~n3020 & n3102;
  assign n3104 = pi0137 & ~n3102;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = n2651 & ~n3105;
  assign n3107 = pi0054 & ~pi0106;
  assign n3108 = n2473 & n3107;
  assign n3109 = n2592 & n3108;
  assign n3110 = n2643 & n3109;
  assign n3111 = n2620 & ~n3110;
  assign n3112 = pi0137 & ~n3111;
  assign n3113 = ~n3106 & ~n3112;
  assign n3114 = ~n2604 & ~n2626;
  assign n3115 = ~n2632 & ~n2656;
  assign n3116 = n3114 & n3115;
  assign n3117 = n2668 & n3116;
  assign n3118 = pi0137 & ~n3117;
  assign n3119 = n2599 & ~n3118;
  assign n3120 = n3113 & n3119;
  assign n3121 = ~n3101 & n3120;
  assign po0382 = ~n3099 | ~n3121;
  assign n3123 = n3007 & po0382;
  assign n3124 = ~n3008 & ~n3123;
  assign n3125 = ~n2429 & ~po0183;
  assign n3126 = ~n3124 & ~n3125;
  assign n3127 = ~n2952 & ~n3126;
  assign n3128 = n2432 & n2439;
  assign n3129 = ~n3127 & n3128;
  assign n3130 = ~n2435 & n2438;
  assign n3131 = pi0833 & n3130;
  assign n3132 = n2432 & n3131;
  assign n3133 = pi0929 & n3132;
  assign n3134 = pi1138 & ~n3132;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = ~n2439 & ~n3135;
  assign n3137 = ~n3129 & ~n3136;
  assign n3138 = ~pi0332 & n3137;
  assign po0153 = n2441 | ~n3138;
  assign n3140 = pi0939 & n3132;
  assign n3141 = pi1140 & ~n3132;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = ~n2439 & ~n3142;
  assign n3144 = pi0239 & ~n3007;
  assign n3145 = ~n3125 & ~n3144;
  assign n3146 = ~pi0176 & n2429;
  assign n3147 = ~pi0154 & ~n2429;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = n3125 & n3148;
  assign n3150 = n3128 & ~n3149;
  assign n3151 = ~n3145 & n3150;
  assign n3152 = pi0276 & n2440;
  assign n3153 = ~n3151 & ~n3152;
  assign po0154 = n3143 | ~n3153;
  assign n3155 = pi0927 & n3132;
  assign n3156 = pi1139 & ~n3132;
  assign n3157 = ~n3155 & ~n3156;
  assign n3158 = ~n2439 & ~n3157;
  assign n3159 = pi0235 & ~n3007;
  assign n3160 = ~n3125 & ~n3159;
  assign n3161 = pi0173 & n2429;
  assign n3162 = pi0151 & ~n2429;
  assign n3163 = ~n3161 & ~n3162;
  assign n3164 = n3125 & ~n3163;
  assign n3165 = n3128 & ~n3164;
  assign n3166 = ~n3160 & n3165;
  assign n3167 = ~pi0274 & n2440;
  assign n3168 = ~n3166 & ~n3167;
  assign po0155 = n3158 | ~n3168;
  assign n3170 = ~n2702 & n3125;
  assign n3171 = pi0238 & ~n3007;
  assign n3172 = ~pi0284 & n3007;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3125 & ~n3173;
  assign n3175 = ~n3170 & ~n3174;
  assign n3176 = n3128 & ~n3175;
  assign n3177 = ~pi0264 & n2440;
  assign n3178 = ~n3176 & ~n3177;
  assign n3179 = pi0944 & n3132;
  assign n3180 = pi1137 & ~n3132;
  assign n3181 = ~n3179 & ~n3180;
  assign n3182 = ~n2439 & ~n3181;
  assign po0156 = ~n3178 | n3182;
  assign n3184 = ~pi0172 & ~n2429;
  assign n3185 = ~pi0193 & n2429;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = n3125 & ~n3186;
  assign n3188 = pi0249 & ~n3007;
  assign n3189 = ~pi0262 & n3007;
  assign n3190 = ~n3188 & ~n3189;
  assign n3191 = ~n3125 & ~n3190;
  assign n3192 = ~n3187 & ~n3191;
  assign n3193 = n3128 & ~n3192;
  assign n3194 = ~pi0277 & n2440;
  assign n3195 = ~n3193 & ~n3194;
  assign n3196 = pi0932 & n3132;
  assign n3197 = pi1136 & ~n3132;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = ~n2439 & ~n3198;
  assign po0157 = ~n3195 | n3199;
  assign n3201 = ~pi0171 & ~n2429;
  assign n3202 = ~pi0192 & n2429;
  assign n3203 = ~n3201 & ~n3202;
  assign n3204 = n3125 & ~n3203;
  assign n3205 = pi0241 & ~n3007;
  assign n3206 = pi0861 & n3007;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n3125 & ~n3207;
  assign n3209 = ~n3204 & ~n3208;
  assign n3210 = n3128 & ~n3209;
  assign n3211 = ~pi0270 & n2440;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = pi0935 & n3132;
  assign n3214 = pi1135 & ~n3132;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = ~n2439 & ~n3215;
  assign po0158 = ~n3212 | n3216;
  assign n3218 = ~pi0170 & ~n2429;
  assign n3219 = ~pi0194 & n2429;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = n3125 & ~n3220;
  assign n3222 = pi0248 & ~n3007;
  assign n3223 = pi0869 & n3007;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = ~n3125 & ~n3224;
  assign n3226 = ~n3221 & ~n3225;
  assign n3227 = n3128 & ~n3226;
  assign n3228 = ~pi0282 & n2440;
  assign n3229 = ~n3227 & ~n3228;
  assign n3230 = pi0921 & n3132;
  assign n3231 = pi1134 & ~n3132;
  assign n3232 = ~n3230 & ~n3231;
  assign n3233 = ~n2439 & ~n3232;
  assign po0159 = ~n3229 | n3233;
  assign n3235 = ~pi0141 & n2429;
  assign n3236 = ~pi0148 & ~n2429;
  assign n3237 = ~n3235 & ~n3236;
  assign n3238 = n3125 & ~n3237;
  assign n3239 = pi0247 & ~n3007;
  assign n3240 = pi0862 & n3007;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~n3125 & ~n3241;
  assign n3243 = ~n3238 & ~n3242;
  assign n3244 = n3128 & ~n3243;
  assign n3245 = ~pi0281 & n2440;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = pi0920 & n3132;
  assign n3248 = pi1133 & ~n3132;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n2439 & ~n3249;
  assign po0160 = ~n3246 | n3250;
  assign n3252 = ~pi0191 & n2429;
  assign n3253 = ~pi0169 & ~n2429;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = n3125 & ~n3254;
  assign n3256 = pi0246 & ~n3007;
  assign n3257 = pi0877 & n3007;
  assign n3258 = ~n3256 & ~n3257;
  assign n3259 = ~n3125 & ~n3258;
  assign n3260 = ~n3255 & ~n3259;
  assign n3261 = n3128 & ~n3260;
  assign n3262 = ~pi0269 & n2440;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = pi0940 & n3132;
  assign n3265 = pi1132 & ~n3132;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = ~n2439 & ~n3266;
  assign po0161 = ~n3263 | n3267;
  assign n3269 = ~pi0168 & ~n2429;
  assign n3270 = ~pi0190 & n2429;
  assign n3271 = ~n3269 & ~n3270;
  assign n3272 = n3125 & ~n3271;
  assign n3273 = pi0240 & ~n3007;
  assign n3274 = pi0878 & n3007;
  assign n3275 = ~n3273 & ~n3274;
  assign n3276 = ~n3125 & ~n3275;
  assign n3277 = ~n3272 & ~n3276;
  assign n3278 = n3128 & ~n3277;
  assign n3279 = ~pi0280 & n2440;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = pi0933 & n3132;
  assign n3282 = pi1131 & ~n3132;
  assign n3283 = ~n3281 & ~n3282;
  assign n3284 = ~n2439 & ~n3283;
  assign po0162 = ~n3280 | n3284;
  assign n3286 = ~n2714 & n3125;
  assign n3287 = pi0245 & ~n3007;
  assign n3288 = pi0875 & n3007;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = ~n3125 & ~n3289;
  assign n3291 = ~n3286 & ~n3290;
  assign n3292 = n3128 & ~n3291;
  assign n3293 = pi0266 & n2440;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = pi0928 & n3132;
  assign n3296 = pi1130 & ~n3132;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = ~n2439 & ~n3297;
  assign po0163 = ~n3294 | n3298;
  assign n3300 = ~n2710 & n3125;
  assign n3301 = pi0244 & ~n3007;
  assign n3302 = pi0879 & n3007;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = ~n3125 & ~n3303;
  assign n3305 = ~n3300 & ~n3304;
  assign n3306 = n3128 & ~n3305;
  assign n3307 = pi0279 & n2440;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = pi0938 & n3132;
  assign n3310 = pi1129 & ~n3132;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = ~n2439 & ~n3311;
  assign po0164 = ~n3308 | n3312;
  assign n3314 = ~n2705 & n3125;
  assign n3315 = pi0242 & ~n3007;
  assign n3316 = pi0846 & n3007;
  assign n3317 = ~n3315 & ~n3316;
  assign n3318 = ~n3125 & ~n3317;
  assign n3319 = ~n3314 & ~n3318;
  assign n3320 = n3128 & ~n3319;
  assign n3321 = pi0278 & n2440;
  assign n3322 = ~n3320 & ~n3321;
  assign n3323 = pi0930 & n3132;
  assign n3324 = pi1128 & ~n3132;
  assign n3325 = ~n3323 & ~n3324;
  assign n3326 = ~n2439 & ~n3325;
  assign po0165 = ~n3322 | n3326;
  assign n3328 = ~n2644 & n3037;
  assign n3329 = n2750 & ~n2803;
  assign n3330 = ~n2717 & n3329;
  assign n3331 = ~n2807 & ~n3330;
  assign n3332 = n2740 & ~n3331;
  assign n3333 = ~n2569 & n3012;
  assign n3334 = ~n2694 & n3333;
  assign n3335 = n2748 & n3334;
  assign n3336 = ~n3332 & n3335;
  assign n3337 = ~n2637 & ~n2651;
  assign n3338 = n3011 & n3337;
  assign n3339 = ~n2698 & n3338;
  assign n3340 = n3336 & n3339;
  assign n3341 = n3328 & n3340;
  assign n3342 = ~n2604 & ~n2614;
  assign n3343 = n2668 & n3342;
  assign n3344 = n3341 & n3343;
  assign n3345 = ~n2626 & n3344;
  assign n3346 = ~n2632 & n3345;
  assign n3347 = n2685 & n3053;
  assign n3348 = n2685 & ~n3057;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = pi0287 & n2777;
  assign n3351 = pi0961 & n2429;
  assign n3352 = pi0972 & ~n2707;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = pi0977 & n2429;
  assign n3355 = pi0960 & ~n2429;
  assign n3356 = ~n3354 & ~n3355;
  assign n3357 = pi0969 & n2707;
  assign n3358 = pi0963 & ~n2429;
  assign n3359 = ~n3357 & ~n3358;
  assign n3360 = pi0967 & n2707;
  assign n3361 = pi0970 & ~n2429;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = n3359 & n3362;
  assign n3364 = n3356 & n3363;
  assign n3365 = n3353 & n3364;
  assign n3366 = n2762 & ~n3365;
  assign n3367 = ~pi0614 & ~pi0642;
  assign n3368 = ~pi0616 & n3367;
  assign n3369 = pi0603 & n3368;
  assign n3370 = ~n2762 & ~n3369;
  assign n3371 = pi0587 & n2429;
  assign n3372 = pi0947 & ~n2707;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = n2762 & n3373;
  assign n3375 = ~n3370 & ~n3374;
  assign n3376 = ~pi0661 & pi0680;
  assign n3377 = ~pi0662 & ~pi0681;
  assign n3378 = n3376 & n3377;
  assign n3379 = ~n2762 & n3378;
  assign n3380 = pi0602 & n2429;
  assign n3381 = pi0907 & ~n2429;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = n2762 & ~n3382;
  assign n3384 = ~n3379 & ~n3383;
  assign n3385 = ~n3375 & n3384;
  assign n3386 = pi0974 & n2707;
  assign n3387 = pi0978 & ~n2707;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = pi0971 & n2707;
  assign n3390 = pi0975 & ~n2707;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = n3388 & n3391;
  assign n3393 = n2762 & ~n3392;
  assign n3394 = n3385 & ~n3393;
  assign n3395 = ~n3366 & n3394;
  assign n3396 = pi0835 & ~po0950;
  assign n3397 = ~n3395 & n3396;
  assign n3398 = ~n2432 & n3130;
  assign n3399 = ~n3102 & n3398;
  assign n3400 = n3397 & ~n3399;
  assign n3401 = n2432 & n2438;
  assign n3402 = ~n2435 & n3401;
  assign n3403 = pi0835 & pi0984;
  assign n3404 = ~pi0979 & ~n3403;
  assign n3405 = ~pi0252 & ~pi0995;
  assign n3406 = n3404 & ~n3405;
  assign n3407 = ~n2440 & ~n3128;
  assign n3408 = n3406 & n3407;
  assign n3409 = ~n3402 & n3408;
  assign n3410 = n3400 & n3409;
  assign n3411 = n2777 & ~n3410;
  assign n3412 = ~n2770 & ~n3411;
  assign n3413 = ~n3350 & n3412;
  assign n3414 = ~pi0841 & n2826;
  assign n3415 = ~n2823 & ~n2881;
  assign n3416 = ~n3414 & n3415;
  assign n3417 = ~n2841 & n3416;
  assign n3418 = ~n2847 & ~n2858;
  assign n3419 = n3072 & n3418;
  assign n3420 = n3417 & n3419;
  assign n3421 = n2873 & ~n2878;
  assign n3422 = ~n2851 & n3421;
  assign n3423 = n2835 & n3422;
  assign n3424 = ~n2681 & n2903;
  assign n3425 = n3423 & n3424;
  assign n3426 = n3420 & n3425;
  assign n3427 = n3413 & n3426;
  assign n3428 = n3349 & n3427;
  assign po0167 = ~n3346 | ~n3428;
  assign n3430 = ~n2656 & ~n3110;
  assign n3431 = n2599 & n3430;
  assign n3432 = ~n2749 & n2803;
  assign n3433 = ~n2736 & n3432;
  assign n3434 = ~n2717 & ~n3433;
  assign n3435 = n2740 & ~n3434;
  assign n3436 = ~n2569 & ~n3435;
  assign n3437 = ~n2563 & n3436;
  assign n3438 = ~n2795 & n3437;
  assign n3439 = ~n2533 & ~n2910;
  assign n3440 = ~n3033 & n3439;
  assign n3441 = ~n3071 & n3421;
  assign n3442 = ~n2913 & ~n3042;
  assign n3443 = ~n2941 & n3442;
  assign n3444 = ~n2694 & n3443;
  assign n3445 = ~n2823 & ~n2854;
  assign n3446 = ~pi0314 & n2851;
  assign n3447 = ~n2788 & ~n2834;
  assign n3448 = pi0841 & n2826;
  assign n3449 = ~n3066 & ~n3448;
  assign n3450 = n3447 & n3449;
  assign n3451 = ~n3446 & n3450;
  assign n3452 = n3445 & n3451;
  assign n3453 = n3444 & n3452;
  assign n3454 = n3441 & n3453;
  assign n3455 = ~n2544 & ~n2936;
  assign n3456 = ~n2527 & n3455;
  assign n3457 = ~n2537 & n3456;
  assign n3458 = n3454 & n3457;
  assign n3459 = n3440 & n3458;
  assign n3460 = n3438 & n3459;
  assign n3461 = ~n3053 & n3057;
  assign n3462 = n2685 & n3461;
  assign n3463 = ~pi0479 & n2681;
  assign n3464 = ~pi0287 & ~pi0979;
  assign n3465 = n2777 & n3464;
  assign n3466 = ~n3403 & ~n3405;
  assign n3467 = n3465 & n3466;
  assign n3468 = ~po0840 & ~po0740;
  assign n3469 = n3402 & n3468;
  assign n3470 = ~po0740 & n3398;
  assign n3471 = ~n3469 & ~n3470;
  assign n3472 = n3397 & ~n3471;
  assign n3473 = n3467 & n3472;
  assign n3474 = ~n3463 & ~n3473;
  assign n3475 = ~n3462 & n3474;
  assign n3476 = ~pi0145 & n2429;
  assign n3477 = ~pi0197 & ~n2429;
  assign n3478 = ~n3476 & ~n3477;
  assign n3479 = n2763 & ~n2780;
  assign n3480 = ~n2784 & n3479;
  assign n3481 = ~n2798 & n3480;
  assign n3482 = n3478 & n3481;
  assign n3483 = ~pi0181 & n2429;
  assign n3484 = ~pi0159 & ~n2429;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = n3481 & n3485;
  assign n3487 = n3482 & n3486;
  assign n3488 = ~pi0182 & n2429;
  assign n3489 = ~pi0160 & ~n2429;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = n3481 & n3490;
  assign n3492 = ~pi0180 & n2429;
  assign n3493 = ~pi0158 & ~n2429;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = n3481 & n3494;
  assign n3496 = n3491 & n3495;
  assign n3497 = n3487 & n3496;
  assign n3498 = n2637 & ~n3497;
  assign n3499 = n3475 & ~n3498;
  assign n3500 = n3460 & n3499;
  assign n3501 = ~n2619 & ~n2901;
  assign n3502 = n3500 & n3501;
  assign po0195 = ~n3431 | ~n3502;
  assign n3504 = ~pi0228 & po0195;
  assign n3505 = pi0030 & pi0228;
  assign n3506 = ~n3504 & ~n3505;
  assign po0171 = n3384 | n3506;
  assign po0172 = ~n3375 | n3506;
  assign n3509 = n2762 & ~n3362;
  assign po0173 = n3506 | ~n3509;
  assign n3511 = n2762 & ~n3353;
  assign po0174 = n3506 | ~n3511;
  assign n3513 = n2762 & ~n3356;
  assign po0175 = n3506 | ~n3513;
  assign n3515 = n2762 & ~n3359;
  assign po0176 = n3506 | ~n3515;
  assign n3517 = n2762 & ~n3391;
  assign po0177 = n3506 | ~n3517;
  assign n3519 = n2762 & ~n3388;
  assign po0178 = n3506 | ~n3519;
  assign n3521 = ~pi0024 & pi0954;
  assign n3522 = ~pi0954 & po0195;
  assign po0182 = n3521 | n3522;
  assign n3524 = ~pi0228 & pi0252;
  assign n3525 = ~pi0119 & ~n3524;
  assign n3526 = pi0119 & pi1050;
  assign n3527 = ~n3525 & ~n3526;
  assign po0184 = pi0468 | ~n3527;
  assign n3529 = pi0119 & pi1071;
  assign n3530 = ~n3525 & ~n3529;
  assign po0185 = pi0468 | ~n3530;
  assign n3532 = pi0119 & pi1067;
  assign n3533 = ~n3525 & ~n3532;
  assign po0186 = pi0468 | ~n3533;
  assign n3535 = pi0119 & pi1035;
  assign n3536 = ~n3525 & ~n3535;
  assign po0187 = pi0468 | ~n3536;
  assign n3538 = ~pi1155 & ~pi1156;
  assign n3539 = ~pi1157 & n3538;
  assign n3540 = po1057 & ~n2801;
  assign n3541 = ~pi0122 & po0840;
  assign n3542 = ~pi0024 & n3541;
  assign n3543 = pi0252 & n3542;
  assign n3544 = n3042 & n3543;
  assign n3545 = ~po0740 & n3544;
  assign n3546 = n3540 & n3545;
  assign n3547 = ~pi0287 & n2777;
  assign n3548 = n3397 & n3547;
  assign n3549 = n3102 & n3402;
  assign n3550 = n3548 & n3549;
  assign n3551 = n3406 & n3550;
  assign n3552 = ~pi0024 & n2563;
  assign n3553 = ~pi0122 & ~po0740;
  assign n3554 = n3552 & n3553;
  assign n3555 = po0840 & n3554;
  assign n3556 = ~pi0122 & n3102;
  assign n3557 = n2651 & n3556;
  assign n3558 = ~pi0841 & n2823;
  assign n3559 = ~n2922 & ~n3558;
  assign n3560 = ~n2667 & n3559;
  assign n3561 = ~n2632 & n3560;
  assign n3562 = ~n3414 & n3561;
  assign n3563 = ~n3557 & n3562;
  assign n3564 = ~n3555 & n3563;
  assign n3565 = ~po0740 & n3541;
  assign n3566 = pi0228 & n3565;
  assign n3567 = n2740 & n3566;
  assign n3568 = n3540 & n3567;
  assign n3569 = n2858 & n3541;
  assign n3570 = ~pi0841 & n3569;
  assign n3571 = ~n3568 & ~n3570;
  assign n3572 = n3564 & n3571;
  assign n3573 = ~n3551 & n3572;
  assign n3574 = ~n3546 & n3573;
  assign n3575 = ~pi0286 & ~pi0288;
  assign n3576 = ~pi0289 & n3575;
  assign n3577 = ~pi0285 & n3576;
  assign n3578 = pi1085 & pi1087;
  assign n3579 = n3553 & ~n3578;
  assign n3580 = n2726 & n3579;
  assign n3581 = ~n3577 & n3580;
  assign n3582 = n3574 & ~n3581;
  assign po0280 = ~po0950 & ~n3582;
  assign n3584 = ~pi0217 & ~pi1085;
  assign n3585 = n2721 & n3584;
  assign n3586 = ~po0950 & n3585;
  assign n3587 = ~n3582 & n3586;
  assign n3588 = ~pi0588 & ~pi0590;
  assign n3589 = ~pi0591 & n3588;
  assign n3590 = pi0592 & n3589;
  assign n3591 = pi0383 & n3590;
  assign n3592 = ~pi0588 & ~pi0591;
  assign n3593 = ~pi0592 & n3592;
  assign n3594 = pi0590 & n3593;
  assign n3595 = pi0358 & n3594;
  assign n3596 = ~n3591 & ~n3595;
  assign n3597 = ~pi0590 & ~pi0592;
  assign n3598 = ~pi0588 & n3597;
  assign n3599 = pi0591 & n3598;
  assign n3600 = pi0407 & n3599;
  assign n3601 = pi0588 & ~pi0590;
  assign n3602 = ~pi0591 & ~pi0592;
  assign n3603 = n3601 & n3602;
  assign n3604 = pi0431 & n3603;
  assign n3605 = ~n3600 & ~n3604;
  assign n3606 = n3596 & n3605;
  assign n3607 = pi0364 & n3590;
  assign n3608 = pi0343 & n3594;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = pi0391 & n3599;
  assign n3611 = pi0415 & n3603;
  assign n3612 = ~n3610 & ~n3611;
  assign n3613 = n3609 & n3612;
  assign n3614 = pi0367 & n3590;
  assign n3615 = pi0345 & n3594;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617 = pi0392 & n3599;
  assign n3618 = pi0417 & n3603;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = n3616 & n3619;
  assign n3621 = ~n3613 & n3620;
  assign n3622 = n3613 & ~n3620;
  assign n3623 = ~n3621 & ~n3622;
  assign n3624 = pi0336 & n3590;
  assign n3625 = pi0362 & n3594;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = pi0463 & n3599;
  assign n3628 = pi0437 & n3603;
  assign n3629 = ~n3627 & ~n3628;
  assign n3630 = n3626 & n3629;
  assign n3631 = pi0447 & n3590;
  assign n3632 = pi0327 & n3594;
  assign n3633 = ~n3631 & ~n3632;
  assign n3634 = pi0333 & n3599;
  assign n3635 = pi0453 & n3603;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = n3633 & n3636;
  assign n3638 = ~n3630 & n3637;
  assign n3639 = n3630 & ~n3637;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = ~n3623 & n3640;
  assign n3642 = n3623 & ~n3640;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = pi0368 & n3590;
  assign n3645 = pi0346 & n3594;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = pi0393 & n3599;
  assign n3648 = pi0418 & n3603;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = n3646 & n3649;
  assign n3651 = pi0389 & n3590;
  assign n3652 = pi0450 & n3594;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = pi0413 & n3599;
  assign n3655 = pi0438 & n3603;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = n3653 & n3656;
  assign n3658 = ~n3650 & n3657;
  assign n3659 = n3650 & ~n3657;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = pi0365 & n3590;
  assign n3662 = pi0323 & n3594;
  assign n3663 = ~n3661 & ~n3662;
  assign n3664 = pi0334 & n3599;
  assign n3665 = pi0464 & n3603;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = n3663 & n3666;
  assign n3668 = pi0366 & n3590;
  assign n3669 = pi0344 & n3594;
  assign n3670 = ~n3668 & ~n3669;
  assign n3671 = pi0335 & n3599;
  assign n3672 = pi0416 & n3603;
  assign n3673 = ~n3671 & ~n3672;
  assign n3674 = n3670 & n3673;
  assign n3675 = ~n3667 & n3674;
  assign n3676 = n3667 & ~n3674;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = ~n3660 & n3677;
  assign n3679 = n3660 & ~n3677;
  assign n3680 = ~n3678 & ~n3679;
  assign n3681 = ~n3643 & n3680;
  assign n3682 = n3643 & ~n3680;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = ~n3606 & n3683;
  assign n3685 = n3606 & ~n3683;
  assign n3686 = ~n3684 & ~n3685;
  assign n3687 = pi1191 & ~n3686;
  assign n3688 = pi0433 & n3603;
  assign n3689 = pi0385 & n3590;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = pi0409 & n3599;
  assign n3692 = pi0360 & n3594;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = n3690 & n3693;
  assign n3695 = pi0377 & n3590;
  assign n3696 = pi0462 & n3594;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = pi0318 & n3599;
  assign n3699 = pi0448 & n3603;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = n3697 & n3700;
  assign n3702 = pi0381 & n3590;
  assign n3703 = pi0356 & n3594;
  assign n3704 = ~n3702 & ~n3703;
  assign n3705 = pi0405 & n3599;
  assign n3706 = pi0445 & n3603;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = n3704 & n3707;
  assign n3709 = ~n3701 & n3708;
  assign n3710 = n3701 & ~n3708;
  assign n3711 = ~n3709 & ~n3710;
  assign n3712 = pi0326 & n3599;
  assign n3713 = pi0449 & n3603;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = pi0461 & n3594;
  assign n3716 = pi0439 & n3590;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n3714 & n3717;
  assign n3719 = pi0451 & n3603;
  assign n3720 = pi0353 & n3594;
  assign n3721 = ~n3719 & ~n3720;
  assign n3722 = pi0325 & n3599;
  assign n3723 = pi0378 & n3590;
  assign n3724 = ~n3722 & ~n3723;
  assign n3725 = n3721 & n3724;
  assign n3726 = ~n3718 & n3725;
  assign n3727 = n3718 & ~n3725;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = ~n3711 & n3728;
  assign n3730 = n3711 & ~n3728;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = pi0382 & n3590;
  assign n3733 = pi0357 & n3594;
  assign n3734 = ~n3732 & ~n3733;
  assign n3735 = pi0406 & n3599;
  assign n3736 = pi0430 & n3603;
  assign n3737 = ~n3735 & ~n3736;
  assign n3738 = n3734 & n3737;
  assign n3739 = pi0401 & n3599;
  assign n3740 = pi0351 & n3594;
  assign n3741 = ~n3739 & ~n3740;
  assign n3742 = pi0426 & n3603;
  assign n3743 = pi0376 & n3590;
  assign n3744 = ~n3742 & ~n3743;
  assign n3745 = n3741 & n3744;
  assign n3746 = ~n3738 & n3745;
  assign n3747 = n3738 & ~n3745;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = pi0317 & n3590;
  assign n3750 = pi0352 & n3594;
  assign n3751 = ~n3749 & ~n3750;
  assign n3752 = pi0402 & n3599;
  assign n3753 = pi0427 & n3603;
  assign n3754 = ~n3752 & ~n3753;
  assign n3755 = n3751 & n3754;
  assign n3756 = pi0379 & n3590;
  assign n3757 = pi0354 & n3594;
  assign n3758 = ~n3756 & ~n3757;
  assign n3759 = pi0403 & n3599;
  assign n3760 = pi0428 & n3603;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = n3758 & n3761;
  assign n3763 = ~n3755 & n3762;
  assign n3764 = n3755 & ~n3762;
  assign n3765 = ~n3763 & ~n3764;
  assign n3766 = ~n3748 & n3765;
  assign n3767 = n3748 & ~n3765;
  assign n3768 = ~n3766 & ~n3767;
  assign n3769 = ~n3731 & n3768;
  assign n3770 = n3731 & ~n3768;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n3694 & n3771;
  assign n3773 = n3694 & ~n3771;
  assign n3774 = ~n3772 & ~n3773;
  assign n3775 = pi1193 & ~n3774;
  assign n3776 = pi0324 & n3599;
  assign n3777 = pi0446 & n3603;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = pi0339 & n3590;
  assign n3780 = pi0460 & n3594;
  assign n3781 = ~n3779 & ~n3780;
  assign n3782 = n3778 & n3781;
  assign n3783 = pi0456 & n3599;
  assign n3784 = pi0443 & n3603;
  assign n3785 = ~n3783 & ~n3784;
  assign n3786 = pi0337 & n3590;
  assign n3787 = pi0441 & n3594;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = n3785 & n3788;
  assign n3790 = pi0390 & n3599;
  assign n3791 = pi0342 & n3594;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = pi0414 & n3603;
  assign n3794 = pi0363 & n3590;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = n3792 & n3795;
  assign n3797 = ~n3789 & n3796;
  assign n3798 = n3789 & ~n3796;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = pi0380 & n3590;
  assign n3801 = pi0355 & n3594;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = pi0404 & n3599;
  assign n3804 = pi0429 & n3603;
  assign n3805 = ~n3803 & ~n3804;
  assign n3806 = n3802 & n3805;
  assign n3807 = pi0386 & n3590;
  assign n3808 = pi0361 & n3594;
  assign n3809 = ~n3807 & ~n3808;
  assign n3810 = pi0410 & n3599;
  assign n3811 = pi0434 & n3603;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = n3809 & n3812;
  assign n3814 = ~n3806 & n3813;
  assign n3815 = n3806 & ~n3813;
  assign n3816 = ~n3814 & ~n3815;
  assign n3817 = ~n3799 & n3816;
  assign n3818 = n3799 & ~n3816;
  assign n3819 = ~n3817 & ~n3818;
  assign n3820 = pi0319 & n3599;
  assign n3821 = pi0458 & n3594;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = pi0444 & n3603;
  assign n3824 = pi0338 & n3590;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = n3822 & n3825;
  assign n3827 = pi0411 & n3599;
  assign n3828 = pi0435 & n3603;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = pi0387 & n3590;
  assign n3831 = pi0452 & n3594;
  assign n3832 = ~n3830 & ~n3831;
  assign n3833 = n3829 & n3832;
  assign n3834 = ~n3826 & n3833;
  assign n3835 = n3826 & ~n3833;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = pi0372 & n3590;
  assign n3838 = pi0320 & n3594;
  assign n3839 = ~n3837 & ~n3838;
  assign n3840 = pi0397 & n3599;
  assign n3841 = pi0422 & n3603;
  assign n3842 = ~n3840 & ~n3841;
  assign n3843 = n3839 & n3842;
  assign n3844 = pi0412 & n3599;
  assign n3845 = pi0388 & n3590;
  assign n3846 = ~n3844 & ~n3845;
  assign n3847 = pi0436 & n3603;
  assign n3848 = pi0455 & n3594;
  assign n3849 = ~n3847 & ~n3848;
  assign n3850 = n3846 & n3849;
  assign n3851 = ~n3843 & n3850;
  assign n3852 = n3843 & ~n3850;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = ~n3836 & n3853;
  assign n3855 = n3836 & ~n3853;
  assign n3856 = ~n3854 & ~n3855;
  assign n3857 = ~n3819 & n3856;
  assign n3858 = n3819 & ~n3856;
  assign n3859 = ~n3857 & ~n3858;
  assign n3860 = ~n3782 & n3859;
  assign n3861 = n3782 & ~n3859;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = pi1190 & ~n3862;
  assign n3864 = pi0384 & n3590;
  assign n3865 = pi0359 & n3594;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = pi0408 & n3599;
  assign n3868 = pi0432 & n3603;
  assign n3869 = ~n3867 & ~n3868;
  assign n3870 = n3866 & n3869;
  assign n3871 = pi0396 & n3599;
  assign n3872 = pi0322 & n3594;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = pi0421 & n3603;
  assign n3875 = pi0371 & n3590;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = n3873 & n3876;
  assign n3878 = pi0454 & n3603;
  assign n3879 = pi0349 & n3594;
  assign n3880 = pi0440 & n3590;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = pi0329 & n3599;
  assign n3883 = n3881 & ~n3882;
  assign n3884 = ~n3878 & n3883;
  assign n3885 = ~n3877 & n3884;
  assign n3886 = n3877 & ~n3884;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = pi0370 & n3590;
  assign n3889 = pi0347 & n3594;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = pi0395 & n3599;
  assign n3892 = pi0420 & n3603;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = n3890 & n3893;
  assign n3895 = pi0375 & n3590;
  assign n3896 = pi0316 & n3594;
  assign n3897 = ~n3895 & ~n3896;
  assign n3898 = pi0399 & n3599;
  assign n3899 = pi0424 & n3603;
  assign n3900 = ~n3898 & ~n3899;
  assign n3901 = n3897 & n3900;
  assign n3902 = ~n3894 & n3901;
  assign n3903 = n3894 & ~n3901;
  assign n3904 = ~n3902 & ~n3903;
  assign n3905 = ~n3887 & n3904;
  assign n3906 = n3887 & ~n3904;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = pi0374 & n3590;
  assign n3909 = pi0350 & n3594;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = pi0400 & n3599;
  assign n3912 = pi0425 & n3603;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = n3910 & n3913;
  assign n3915 = pi0369 & n3590;
  assign n3916 = pi0315 & n3594;
  assign n3917 = ~n3915 & ~n3916;
  assign n3918 = pi0394 & n3599;
  assign n3919 = pi0419 & n3603;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = n3917 & n3920;
  assign n3922 = ~n3914 & n3921;
  assign n3923 = n3914 & ~n3921;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = pi0442 & n3590;
  assign n3926 = pi0321 & n3594;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = pi0328 & n3599;
  assign n3929 = pi0459 & n3603;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = n3927 & n3930;
  assign n3932 = pi0423 & n3603;
  assign n3933 = pi0348 & n3594;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = pi0398 & n3599;
  assign n3936 = pi0373 & n3590;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = n3934 & n3937;
  assign n3939 = ~n3931 & n3938;
  assign n3940 = n3931 & ~n3938;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3924 & n3941;
  assign n3943 = n3924 & ~n3941;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~n3907 & n3944;
  assign n3946 = n3907 & ~n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = ~n3870 & n3947;
  assign n3949 = n3870 & ~n3947;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = pi1192 & ~n3950;
  assign n3952 = ~n3863 & ~n3951;
  assign n3953 = ~n3775 & n3952;
  assign n3954 = ~n3687 & n3953;
  assign n3955 = n3587 & ~n3954;
  assign n3956 = ~pi0098 & pi0567;
  assign n3957 = n2721 & ~n3956;
  assign n3958 = ~n3955 & ~n3957;
  assign n3959 = po0280 & n3958;
  assign n3960 = n3539 & n3959;
  assign n3961 = pi1155 & pi1156;
  assign n3962 = ~pi1157 & n3961;
  assign n3963 = ~n3539 & n3962;
  assign n3964 = ~pi0031 & n3963;
  assign n3965 = n2721 & n3964;
  assign po0189 = n3960 | n3965;
  assign n3967 = n2726 & n3540;
  assign n3968 = pi0032 & n2604;
  assign n3969 = n3967 & n3968;
  assign n3970 = ~n2749 & ~n2803;
  assign n3971 = ~pi0137 & ~n3540;
  assign n3972 = n3970 & n3971;
  assign n3973 = pi0683 & n2726;
  assign n3974 = n3540 & ~n3973;
  assign n3975 = ~n2749 & n3974;
  assign n3976 = pi0032 & n3975;
  assign n3977 = ~n2803 & n3976;
  assign n3978 = ~n3972 & ~n3977;
  assign n3979 = ~n2736 & ~n3978;
  assign n3980 = pi0032 & n2736;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = n2740 & ~n3981;
  assign n3983 = pi0032 & ~pi0314;
  assign n3984 = pi1044 & n3983;
  assign n3985 = n2619 & n3984;
  assign n3986 = pi0024 & pi0032;
  assign n3987 = n2591 & n3986;
  assign n3988 = ~n3985 & ~n3987;
  assign n3989 = ~pi0024 & n3102;
  assign n3990 = pi0032 & n3989;
  assign n3991 = ~n3986 & ~n3990;
  assign n3992 = n2563 & ~n3991;
  assign n3993 = n2795 & n3986;
  assign n3994 = ~n3992 & ~n3993;
  assign n3995 = pi0032 & pi0841;
  assign n3996 = n2644 & n3995;
  assign n3997 = ~n2583 & ~n2698;
  assign n3998 = ~n2747 & n3997;
  assign n3999 = n3995 & ~n3998;
  assign n4000 = ~n3996 & ~n3999;
  assign n4001 = n3994 & n4000;
  assign n4002 = n3988 & n4001;
  assign n4003 = ~po0740 & ~n3018;
  assign n4004 = n2651 & n4003;
  assign n4005 = pi0479 & n4004;
  assign n4006 = ~n3102 & n4005;
  assign n4007 = pi0032 & n4006;
  assign n4008 = pi0252 & po0740;
  assign n4009 = pi0314 & ~n4008;
  assign n4010 = n2614 & ~n4009;
  assign n4011 = n2614 & n4009;
  assign n4012 = pi0252 & pi0986;
  assign n4013 = n4011 & n4012;
  assign n4014 = ~n4010 & ~n4013;
  assign n4015 = pi0032 & ~n4014;
  assign n4016 = n3110 & n3986;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = pi0032 & po0740;
  assign n4019 = n2651 & n4018;
  assign n4020 = ~n3102 & n4019;
  assign n4021 = n4017 & ~n4020;
  assign n4022 = ~n4007 & n4021;
  assign n4023 = n4002 & n4022;
  assign n4024 = ~n3982 & n4023;
  assign n4025 = ~n3969 & n4024;
  assign n4026 = pi0252 & ~n3540;
  assign n4027 = n3042 & ~n4026;
  assign n4028 = n2716 & n3540;
  assign n4029 = ~po0840 & ~n4028;
  assign n4030 = n4027 & n4029;
  assign n4031 = ~pi0137 & n4030;
  assign n4032 = ~pi0024 & n4031;
  assign n4033 = n3042 & n3986;
  assign n4034 = ~n4032 & ~n4033;
  assign n4035 = pi0024 & ~pi0032;
  assign n4036 = n2913 & ~n4035;
  assign n4037 = n2533 & n3983;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = ~pi0137 & n3018;
  assign n4040 = pi0032 & ~n3553;
  assign n4041 = ~n4039 & ~n4040;
  assign n4042 = n2930 & ~n4041;
  assign n4043 = ~po0840 & ~n3577;
  assign n4044 = n4042 & ~n4043;
  assign n4045 = pi0032 & n4043;
  assign n4046 = n2930 & n4045;
  assign n4047 = ~n4044 & ~n4046;
  assign n4048 = n2936 & n3983;
  assign n4049 = n2917 & n3995;
  assign n4050 = ~n4048 & ~n4049;
  assign n4051 = n2544 & n3983;
  assign n4052 = n4050 & ~n4051;
  assign n4053 = n4047 & n4052;
  assign n4054 = n4038 & n4053;
  assign n4055 = pi0032 & ~pi1076;
  assign n4056 = n2926 & n4055;
  assign n4057 = n4054 & ~n4056;
  assign n4058 = ~pi0252 & n3540;
  assign n4059 = n2813 & n3540;
  assign n4060 = ~n4058 & n4059;
  assign n4061 = pi0252 & po0840;
  assign n4062 = n4060 & ~n4061;
  assign n4063 = pi0032 & n4062;
  assign n4064 = n2726 & n3577;
  assign n4065 = n2515 & ~n4064;
  assign n4066 = n2492 & n4065;
  assign n4067 = n2726 & n4066;
  assign n4068 = pi0032 & n4067;
  assign n4069 = n2910 & n3986;
  assign n4070 = ~n4068 & ~n4069;
  assign n4071 = n3033 & n3986;
  assign n4072 = n4070 & ~n4071;
  assign n4073 = ~n4063 & n4072;
  assign n4074 = n4057 & n4073;
  assign n4075 = n4034 & n4074;
  assign n4076 = n2681 & n3986;
  assign n4077 = ~n2770 & ~n2892;
  assign n4078 = n3995 & ~n4077;
  assign n4079 = ~n4076 & ~n4078;
  assign n4080 = n3057 & n3986;
  assign n4081 = pi0032 & ~n3057;
  assign n4082 = ~n4080 & ~n4081;
  assign n4083 = n2685 & ~n3053;
  assign n4084 = ~n4082 & n4083;
  assign n4085 = n2901 & n3983;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = n3406 & n3547;
  assign n4088 = ~pi1076 & ~n3397;
  assign n4089 = ~pi0786 & n4088;
  assign n4090 = pi0032 & n4089;
  assign n4091 = pi1076 & ~n3397;
  assign n4092 = pi0032 & n4091;
  assign n4093 = pi0032 & n3128;
  assign n4094 = pi0835 & ~po0740;
  assign n4095 = n4093 & ~n4094;
  assign n4096 = ~n3398 & ~n3402;
  assign n4097 = ~n2440 & n4096;
  assign n4098 = n4018 & ~n4097;
  assign n4099 = ~n4095 & ~n4098;
  assign n4100 = n3397 & ~n4099;
  assign n4101 = ~n4092 & ~n4100;
  assign n4102 = ~n4090 & n4101;
  assign n4103 = n4087 & ~n4102;
  assign n4104 = n4086 & ~n4103;
  assign n4105 = ~n2656 & ~n2662;
  assign n4106 = n3983 & ~n4105;
  assign n4107 = n2569 & n3986;
  assign n4108 = ~n4106 & ~n4107;
  assign n4109 = pi0032 & pi0993;
  assign n4110 = n2576 & n4109;
  assign n4111 = n2598 & n3986;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = n4108 & n4112;
  assign n4114 = n4104 & n4113;
  assign n4115 = n4079 & n4114;
  assign n4116 = ~n3072 & n3986;
  assign n4117 = n2847 & n3995;
  assign n4118 = n2834 & n3984;
  assign n4119 = ~n4117 & ~n4118;
  assign n4120 = n2858 & n3995;
  assign n4121 = pi0479 & n2856;
  assign n4122 = n2857 & n4121;
  assign n4123 = ~po0840 & n4122;
  assign n4124 = ~pi0841 & n4123;
  assign n4125 = pi0032 & n4124;
  assign n4126 = n2854 & n3986;
  assign n4127 = n2881 & n4018;
  assign n4128 = n2726 & n4127;
  assign n4129 = ~n4126 & ~n4128;
  assign n4130 = ~n4125 & n4129;
  assign n4131 = ~n4120 & n4130;
  assign n4132 = ~n2826 & ~n2831;
  assign n4133 = ~n2823 & n4132;
  assign n4134 = n3995 & ~n4133;
  assign n4135 = n4131 & ~n4134;
  assign n4136 = n2851 & n3983;
  assign n4137 = n3066 & n3986;
  assign n4138 = ~n4136 & ~n4137;
  assign n4139 = n4135 & n4138;
  assign n4140 = n4119 & n4139;
  assign n4141 = ~n4116 & n4140;
  assign n4142 = n4115 & n4141;
  assign n4143 = n4075 & n4142;
  assign po0190 = ~n4025 | ~n4143;
  assign n4145 = ~pi0979 & n3398;
  assign n4146 = ~n3403 & n4145;
  assign n4147 = n3397 & n4146;
  assign n4148 = n3102 & n4147;
  assign n4149 = ~n3405 & n4148;
  assign n4150 = n3547 & n4149;
  assign n4151 = n2619 & ~n2777;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = ~n3148 & ~n4152;
  assign n4154 = n2508 & ~n2823;
  assign n4155 = ~n3558 & ~n4154;
  assign n4156 = ~n3186 & ~n4155;
  assign n4157 = ~n2777 & n2834;
  assign n4158 = n3547 & n4146;
  assign n4159 = ~n3405 & n3468;
  assign n4160 = n3397 & n4159;
  assign n4161 = n4158 & n4160;
  assign n4162 = ~n4157 & ~n4161;
  assign n4163 = ~pi0075 & ~pi0100;
  assign n4164 = ~pi0183 & n2429;
  assign n4165 = ~pi0149 & ~n2429;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = n3481 & n4166;
  assign n4168 = ~pi0178 & n2429;
  assign n4169 = ~pi0157 & ~n2429;
  assign n4170 = ~n4168 & ~n4169;
  assign n4171 = n3481 & n4170;
  assign n4172 = ~n4167 & ~n4171;
  assign n4173 = n4167 & n4171;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = ~n4163 & ~n4174;
  assign n4176 = n4162 & ~n4175;
  assign n4177 = ~n2591 & ~n2854;
  assign n4178 = ~n2910 & n4177;
  assign n4179 = ~n2913 & n4178;
  assign n4180 = ~n2598 & n4179;
  assign n4181 = ~n2685 & ~n4180;
  assign n4182 = ~n3462 & ~n4181;
  assign n4183 = ~n3463 & n4182;
  assign n4184 = ~pi0038 & ~pi0059;
  assign n4185 = ~pi0057 & n4184;
  assign n4186 = ~pi0054 & n4185;
  assign n4187 = ~pi0079 & ~pi0118;
  assign n4188 = ~pi0033 & ~pi0139;
  assign n4189 = ~pi0034 & n4188;
  assign n4190 = n4187 & n4189;
  assign n4191 = ~pi0138 & n4190;
  assign n4192 = ~pi0195 & ~pi0196;
  assign po0997 = n4191 & n4192;
  assign n4194 = ~pi0954 & ~po0997;
  assign n4195 = pi0033 & n4194;
  assign n4196 = ~pi0033 & ~n4194;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = ~pi0040 & n2452;
  assign n4199 = ~n4197 & n4198;
  assign n4200 = n4186 & ~n4199;
  assign n4201 = ~pi0164 & ~n2429;
  assign n4202 = ~pi0186 & n2429;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = n3481 & n4203;
  assign n4205 = ~n4186 & ~n4204;
  assign n4206 = ~n4200 & ~n4205;
  assign n4207 = ~pi0074 & ~n4206;
  assign n4208 = n3254 & n3481;
  assign n4209 = pi0074 & ~n4208;
  assign n4210 = ~n4207 & ~n4209;
  assign n4211 = n4183 & ~n4210;
  assign n4212 = ~n4167 & ~n4182;
  assign n4213 = n3463 & n4182;
  assign n4214 = ~n3495 & n4213;
  assign n4215 = ~n4212 & ~n4214;
  assign n4216 = n4163 & n4215;
  assign n4217 = ~n4211 & n4216;
  assign n4218 = n4176 & ~n4217;
  assign n4219 = n2705 & n3481;
  assign n4220 = ~n4162 & ~n4219;
  assign n4221 = ~n4218 & ~n4220;
  assign n4222 = n4155 & ~n4221;
  assign n4223 = ~n4156 & ~n4222;
  assign n4224 = ~n3481 & ~n4155;
  assign n4225 = n4223 & ~n4224;
  assign n4226 = n4152 & ~n4225;
  assign n4227 = ~n4153 & ~n4226;
  assign n4228 = ~n3481 & ~n4152;
  assign po0191 = ~n4227 | n4228;
  assign n4230 = ~pi0177 & n2429;
  assign n4231 = ~pi0155 & ~n2429;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = ~n4152 & n4232;
  assign n4234 = ~n4163 & ~n4172;
  assign n4235 = ~pi0140 & n2429;
  assign n4236 = ~pi0162 & ~n2429;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = n3481 & n4237;
  assign n4239 = ~n3482 & ~n4238;
  assign n4240 = n3482 & n4238;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = n4234 & ~n4241;
  assign n4243 = ~n4163 & n4172;
  assign n4244 = n4241 & n4243;
  assign n4245 = ~n4242 & ~n4244;
  assign n4246 = n4162 & n4245;
  assign n4247 = ~pi0033 & ~pi0034;
  assign n4248 = pi0033 & pi0034;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = n4194 & ~n4249;
  assign n4251 = pi0034 & ~n4194;
  assign n4252 = ~n4250 & ~n4251;
  assign n4253 = n4198 & n4252;
  assign n4254 = n4186 & ~n4253;
  assign n4255 = ~pi0167 & ~n2429;
  assign n4256 = ~pi0188 & n2429;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = n3481 & n4257;
  assign n4259 = ~n4186 & ~n4258;
  assign n4260 = ~n4254 & ~n4259;
  assign n4261 = ~pi0074 & ~n4260;
  assign n4262 = n3237 & n3481;
  assign n4263 = pi0074 & ~n4262;
  assign n4264 = ~n4261 & ~n4263;
  assign n4265 = n4183 & ~n4264;
  assign n4266 = ~n4182 & ~n4238;
  assign n4267 = ~n3486 & n4213;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = n4163 & n4268;
  assign n4270 = ~n4265 & n4269;
  assign n4271 = n4246 & ~n4270;
  assign n4272 = n2710 & n3481;
  assign n4273 = ~n4162 & ~n4272;
  assign n4274 = ~n4271 & ~n4273;
  assign n4275 = n4155 & ~n4274;
  assign n4276 = ~n2702 & ~n4155;
  assign n4277 = ~n4151 & ~n4276;
  assign n4278 = ~n4150 & n4277;
  assign n4279 = ~n4224 & n4278;
  assign n4280 = ~n4275 & n4279;
  assign n4281 = ~n4233 & ~n4280;
  assign po0192 = n4228 | n4281;
  assign n4283 = pi0024 & pi0035;
  assign n4284 = n2681 & n4283;
  assign n4285 = pi0035 & pi0841;
  assign n4286 = ~n4077 & n4285;
  assign n4287 = ~n4284 & ~n4286;
  assign n4288 = pi0035 & ~pi0314;
  assign n4289 = n2901 & n4288;
  assign n4290 = pi0024 & ~pi0035;
  assign n4291 = n3057 & ~n4290;
  assign n4292 = pi0035 & ~n3057;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = n4083 & ~n4293;
  assign n4295 = ~n4289 & ~n4294;
  assign n4296 = pi0035 & n4089;
  assign n4297 = pi0035 & n4091;
  assign n4298 = pi0035 & n3128;
  assign n4299 = ~n4094 & n4298;
  assign n4300 = pi0035 & po0740;
  assign n4301 = ~n4097 & n4300;
  assign n4302 = ~n4299 & ~n4301;
  assign n4303 = n3397 & ~n4302;
  assign n4304 = ~n4297 & ~n4303;
  assign n4305 = ~n4296 & n4304;
  assign n4306 = n4087 & ~n4305;
  assign n4307 = n4295 & ~n4306;
  assign n4308 = ~n2823 & ~n2831;
  assign n4309 = n4285 & ~n4308;
  assign n4310 = n3066 & ~n4290;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = n2847 & n4285;
  assign n4313 = pi1044 & n4288;
  assign n4314 = n2834 & n4313;
  assign n4315 = ~n4312 & ~n4314;
  assign n4316 = n2858 & n4285;
  assign n4317 = pi0035 & n4124;
  assign n4318 = n2788 & ~n4290;
  assign n4319 = n2881 & n4300;
  assign n4320 = n2726 & n4319;
  assign n4321 = ~n4318 & ~n4320;
  assign n4322 = ~n4317 & n4321;
  assign n4323 = ~n4316 & n4322;
  assign n4324 = n2851 & n4288;
  assign n4325 = n4323 & ~n4324;
  assign n4326 = ~n2854 & ~n3071;
  assign n4327 = n4283 & ~n4326;
  assign n4328 = n4325 & ~n4327;
  assign n4329 = n4315 & n4328;
  assign n4330 = pi0035 & n2826;
  assign n4331 = n4329 & ~n4330;
  assign n4332 = ~n3414 & n4331;
  assign n4333 = n4311 & n4332;
  assign n4334 = n4307 & n4333;
  assign n4335 = n4287 & n4334;
  assign n4336 = n2604 & n3967;
  assign n4337 = pi0035 & n4336;
  assign n4338 = pi0035 & n3989;
  assign n4339 = ~n4283 & ~n4338;
  assign n4340 = n2563 & ~n4339;
  assign n4341 = n2795 & n4283;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = ~n2736 & n2749;
  assign n4344 = ~n2803 & ~n3971;
  assign n4345 = ~pi0035 & ~n3973;
  assign n4346 = n3540 & n4345;
  assign n4347 = ~n2736 & ~n4346;
  assign n4348 = n4344 & n4347;
  assign n4349 = ~n4343 & ~n4348;
  assign n4350 = pi0035 & n2736;
  assign n4351 = n4349 & ~n4350;
  assign n4352 = n2740 & ~n4351;
  assign n4353 = n4342 & ~n4352;
  assign n4354 = ~n3998 & n4285;
  assign n4355 = n4353 & ~n4354;
  assign n4356 = n3042 & n4283;
  assign n4357 = n3033 & n4283;
  assign n4358 = ~n4356 & ~n4357;
  assign n4359 = pi0035 & pi0993;
  assign n4360 = n2576 & n4359;
  assign n4361 = n2598 & n4283;
  assign n4362 = ~n4360 & ~n4361;
  assign n4363 = n4358 & n4362;
  assign n4364 = ~pi0035 & ~pi1076;
  assign n4365 = n2926 & ~n4364;
  assign n4366 = n4363 & ~n4365;
  assign n4367 = pi0137 & n4029;
  assign n4368 = ~n4026 & ~n4367;
  assign n4369 = ~pi0024 & n3042;
  assign n4370 = ~n4368 & n4369;
  assign n4371 = pi0035 & n4067;
  assign n4372 = n2910 & n4283;
  assign n4373 = ~n4371 & ~n4372;
  assign n4374 = ~n2508 & n4373;
  assign n4375 = ~n4370 & n4374;
  assign n4376 = n4366 & n4375;
  assign n4377 = n2917 & n4285;
  assign n4378 = n2913 & n4283;
  assign n4379 = ~n4377 & ~n4378;
  assign n4380 = n2936 & n4288;
  assign n4381 = n4379 & ~n4380;
  assign n4382 = n2619 & n4313;
  assign n4383 = n2644 & n4285;
  assign n4384 = ~n4382 & ~n4383;
  assign n4385 = pi0035 & n4006;
  assign n4386 = pi0035 & ~n4014;
  assign n4387 = n3110 & ~n4290;
  assign n4388 = ~n4386 & ~n4387;
  assign n4389 = n2651 & n4300;
  assign n4390 = ~n3102 & n4389;
  assign n4391 = n4388 & ~n4390;
  assign n4392 = ~n4385 & n4391;
  assign n4393 = n2591 & n4283;
  assign n4394 = n4392 & ~n4393;
  assign n4395 = pi0035 & n4043;
  assign n4396 = n2930 & n4395;
  assign n4397 = ~n4039 & ~n4043;
  assign n4398 = ~pi0035 & ~n3553;
  assign n4399 = n2930 & ~n4398;
  assign n4400 = n4397 & n4399;
  assign n4401 = ~n4396 & ~n4400;
  assign n4402 = ~n2533 & ~n2544;
  assign n4403 = n4288 & ~n4402;
  assign n4404 = n4401 & ~n4403;
  assign n4405 = n4394 & n4404;
  assign n4406 = n4384 & n4405;
  assign n4407 = n4381 & n4406;
  assign n4408 = n4376 & n4407;
  assign n4409 = n2569 & n4283;
  assign n4410 = pi0035 & n4062;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4105 & n4288;
  assign n4413 = n4411 & ~n4412;
  assign n4414 = n4408 & n4413;
  assign n4415 = n4355 & n4414;
  assign n4416 = ~n4337 & n4415;
  assign po0193 = ~n4335 | ~n4416;
  assign n4418 = pi0036 & ~pi0314;
  assign n4419 = ~n4105 & n4418;
  assign n4420 = pi0024 & pi0036;
  assign n4421 = n2569 & n4420;
  assign n4422 = ~n4419 & ~n4421;
  assign n4423 = pi0036 & pi0993;
  assign n4424 = n2576 & n4423;
  assign n4425 = n2598 & n4420;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = n4422 & n4426;
  assign n4428 = pi0036 & pi0841;
  assign n4429 = n2847 & n4428;
  assign n4430 = pi1044 & n4418;
  assign n4431 = n2834 & n4430;
  assign n4432 = ~n4429 & ~n4431;
  assign n4433 = ~n3072 & n4420;
  assign n4434 = n4432 & ~n4433;
  assign n4435 = n2851 & n4418;
  assign n4436 = n3066 & n4420;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438 = n2901 & n4418;
  assign n4439 = n2681 & n4420;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = ~n4077 & n4428;
  assign n4442 = n4440 & ~n4441;
  assign n4443 = n2858 & n4428;
  assign n4444 = pi0036 & n4124;
  assign n4445 = n2854 & n4420;
  assign n4446 = pi0036 & po0740;
  assign n4447 = n2881 & n4446;
  assign n4448 = n2726 & n4447;
  assign n4449 = ~n4445 & ~n4448;
  assign n4450 = ~n4444 & n4449;
  assign n4451 = ~n4443 & n4450;
  assign n4452 = ~n4133 & n4428;
  assign n4453 = n4451 & ~n4452;
  assign n4454 = n4442 & n4453;
  assign n4455 = n4437 & n4454;
  assign n4456 = n4434 & n4455;
  assign n4457 = pi0036 & n4091;
  assign n4458 = ~n4097 & n4446;
  assign n4459 = n3128 & ~n4094;
  assign n4460 = pi0036 & n4459;
  assign n4461 = ~n4458 & ~n4460;
  assign n4462 = n3397 & ~n4461;
  assign n4463 = pi0036 & ~pi0786;
  assign n4464 = n4088 & n4463;
  assign n4465 = ~n4462 & ~n4464;
  assign n4466 = ~n4457 & n4465;
  assign n4467 = n4087 & ~n4466;
  assign n4468 = po0740 & n2888;
  assign n4469 = n3057 & n4420;
  assign n4470 = pi0036 & ~n3057;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = n4083 & ~n4471;
  assign n4473 = ~n4468 & ~n4472;
  assign n4474 = ~n4467 & n4473;
  assign n4475 = n4456 & n4474;
  assign n4476 = pi0036 & n4006;
  assign n4477 = pi0036 & ~n4014;
  assign n4478 = n3110 & n4420;
  assign n4479 = ~n4477 & ~n4478;
  assign n4480 = n2651 & n4446;
  assign n4481 = ~n3102 & n4480;
  assign n4482 = n4479 & ~n4481;
  assign n4483 = ~n4476 & n4482;
  assign n4484 = n2591 & n4420;
  assign n4485 = n4483 & ~n4484;
  assign n4486 = n2619 & n4430;
  assign n4487 = n2644 & n4428;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = n2917 & n4428;
  assign n4490 = n2913 & n4420;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = n2936 & n4418;
  assign n4493 = n4491 & ~n4492;
  assign n4494 = pi0036 & n4043;
  assign n4495 = n2930 & n4494;
  assign n4496 = n2930 & ~n4039;
  assign n4497 = ~n4043 & n4496;
  assign n4498 = pi0036 & ~n3553;
  assign n4499 = n4497 & n4498;
  assign n4500 = ~n4495 & ~n4499;
  assign n4501 = ~n4402 & n4418;
  assign n4502 = n4500 & ~n4501;
  assign n4503 = n3042 & n4420;
  assign n4504 = ~pi1076 & n2926;
  assign n4505 = pi0036 & n4504;
  assign n4506 = ~n4503 & ~n4505;
  assign n4507 = n4502 & n4506;
  assign n4508 = n4493 & n4507;
  assign n4509 = n3033 & n4420;
  assign n4510 = n4508 & ~n4509;
  assign n4511 = n2910 & n4420;
  assign n4512 = pi0036 & n2726;
  assign n4513 = n4066 & n4512;
  assign n4514 = ~n4511 & ~n4513;
  assign n4515 = n4510 & n4514;
  assign n4516 = n4488 & n4515;
  assign n4517 = n4485 & n4516;
  assign n4518 = pi0036 & n2741;
  assign n4519 = n2795 & n4420;
  assign n4520 = n2740 & ~n2749;
  assign n4521 = ~n2736 & n4520;
  assign n4522 = ~n2803 & n4521;
  assign n4523 = n3540 & n4522;
  assign n4524 = pi0036 & n4523;
  assign n4525 = ~n3973 & n4524;
  assign n4526 = pi0036 & po0840;
  assign n4527 = ~po0740 & ~n4526;
  assign n4528 = n3552 & ~n4527;
  assign n4529 = n2563 & n4420;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = ~n4525 & n4530;
  assign n4532 = ~n4519 & n4531;
  assign n4533 = ~n4518 & n4532;
  assign n4534 = ~n3998 & n4428;
  assign n4535 = n4533 & ~n4534;
  assign n4536 = pi0036 & n4336;
  assign n4537 = pi0036 & n4062;
  assign n4538 = ~n4536 & ~n4537;
  assign n4539 = n4535 & n4538;
  assign n4540 = n4517 & n4539;
  assign n4541 = n4475 & n4540;
  assign po0194 = ~n4427 | ~n4541;
  assign n4543 = pi0038 & pi0841;
  assign n4544 = n2917 & n4543;
  assign n4545 = pi0024 & pi0038;
  assign n4546 = n2913 & n4545;
  assign n4547 = ~n4544 & ~n4546;
  assign n4548 = pi0038 & ~pi0314;
  assign n4549 = n2936 & n4548;
  assign n4550 = n4547 & ~n4549;
  assign n4551 = pi0038 & n4043;
  assign n4552 = n2930 & n4551;
  assign n4553 = pi0038 & ~n3553;
  assign n4554 = n4497 & n4553;
  assign n4555 = ~n4552 & ~n4554;
  assign n4556 = ~n4402 & n4548;
  assign n4557 = n4555 & ~n4556;
  assign n4558 = n3042 & n4545;
  assign n4559 = pi0038 & n4504;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = n4557 & n4560;
  assign n4562 = n4550 & n4561;
  assign n4563 = n3033 & n4545;
  assign n4564 = n4562 & ~n4563;
  assign n4565 = ~pi0038 & pi0841;
  assign n4566 = n2747 & ~n4565;
  assign n4567 = n2698 & n4543;
  assign n4568 = ~n4566 & ~n4567;
  assign n4569 = pi0038 & n2741;
  assign n4570 = pi0038 & n3989;
  assign n4571 = ~n4545 & ~n4570;
  assign n4572 = n2563 & ~n4571;
  assign n4573 = ~n4569 & ~n4572;
  assign n4574 = n4568 & n4573;
  assign n4575 = n2598 & n4545;
  assign n4576 = ~n4105 & n4548;
  assign n4577 = n2569 & n4545;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = pi0993 & n2576;
  assign n4580 = pi0038 & n4579;
  assign n4581 = n4578 & ~n4580;
  assign n4582 = ~n4575 & n4581;
  assign n4583 = n4574 & n4582;
  assign n4584 = n4564 & n4583;
  assign n4585 = ~n3973 & n4523;
  assign n4586 = pi0038 & n4585;
  assign n4587 = n2583 & n4543;
  assign n4588 = n2795 & n4545;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = pi1044 & n4548;
  assign n4591 = n2619 & n4590;
  assign n4592 = n2591 & n4545;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = n2910 & n4545;
  assign n4595 = pi0038 & n2726;
  assign n4596 = n4066 & n4595;
  assign n4597 = ~n4594 & ~n4596;
  assign n4598 = pi0038 & ~n4061;
  assign n4599 = n4060 & n4598;
  assign n4600 = n4597 & ~n4599;
  assign n4601 = n4593 & n4600;
  assign n4602 = n4589 & n4601;
  assign n4603 = pi0038 & n3967;
  assign n4604 = n2604 & n4603;
  assign n4605 = n4602 & ~n4604;
  assign n4606 = pi0038 & n4006;
  assign n4607 = pi0038 & ~n4014;
  assign n4608 = n2644 & n4543;
  assign n4609 = ~n4607 & ~n4608;
  assign n4610 = pi0038 & po0740;
  assign n4611 = n2651 & n4610;
  assign n4612 = ~n3102 & n4611;
  assign n4613 = n4609 & ~n4612;
  assign n4614 = ~n4606 & n4613;
  assign n4615 = n3110 & n4545;
  assign n4616 = n4614 & ~n4615;
  assign n4617 = n4605 & n4616;
  assign n4618 = ~n4586 & n4617;
  assign n4619 = n4584 & n4618;
  assign n4620 = n2726 & n4610;
  assign n4621 = n2881 & n4620;
  assign n4622 = n2847 & n4543;
  assign n4623 = ~n4621 & ~n4622;
  assign n4624 = n2858 & n4543;
  assign n4625 = pi0038 & ~pi0841;
  assign n4626 = n4123 & n4625;
  assign n4627 = ~n4624 & ~n4626;
  assign n4628 = n2831 & n4543;
  assign n4629 = n2851 & n4548;
  assign n4630 = ~n4628 & ~n4629;
  assign n4631 = n2788 & n4545;
  assign n4632 = n2834 & n4590;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = ~n4326 & n4545;
  assign n4635 = n4633 & ~n4634;
  assign n4636 = n4630 & n4635;
  assign n4637 = n4627 & n4636;
  assign n4638 = n4623 & n4637;
  assign n4639 = n2823 & n4543;
  assign n4640 = n4638 & ~n4639;
  assign n4641 = n2826 & n4543;
  assign n4642 = n3066 & n4545;
  assign n4643 = ~n4641 & ~n4642;
  assign n4644 = pi0038 & n4091;
  assign n4645 = ~n4097 & n4610;
  assign n4646 = pi0038 & n4459;
  assign n4647 = ~n4645 & ~n4646;
  assign n4648 = n3397 & ~n4647;
  assign n4649 = pi0038 & ~pi0786;
  assign n4650 = n4088 & n4649;
  assign n4651 = ~n4648 & ~n4650;
  assign n4652 = ~n4644 & n4651;
  assign n4653 = n3547 & ~n4652;
  assign n4654 = n3406 & n4653;
  assign n4655 = n3057 & n4545;
  assign n4656 = pi0038 & ~n3057;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = n4083 & ~n4657;
  assign n4659 = ~n4654 & ~n4658;
  assign n4660 = pi0332 & ~pi0841;
  assign n4661 = ~n4543 & ~n4660;
  assign n4662 = n2770 & ~n4661;
  assign n4663 = n4659 & ~n4662;
  assign n4664 = n2901 & n4548;
  assign n4665 = n4663 & ~n4664;
  assign n4666 = n2681 & n4545;
  assign n4667 = n2892 & n4543;
  assign n4668 = ~n4666 & ~n4667;
  assign n4669 = n4665 & n4668;
  assign n4670 = n4643 & n4669;
  assign n4671 = n4640 & n4670;
  assign po0196 = ~n4619 | ~n4671;
  assign n4673 = pi0024 & pi0039;
  assign n4674 = n3057 & n4673;
  assign n4675 = pi0039 & ~n3057;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = n2685 & ~n4676;
  assign n4678 = n2681 & n4673;
  assign n4679 = pi0039 & pi0841;
  assign n4680 = ~n4077 & n4679;
  assign n4681 = ~n4678 & ~n4680;
  assign n4682 = pi0039 & n4091;
  assign n4683 = pi0039 & po0740;
  assign n4684 = ~n4097 & n4683;
  assign n4685 = pi0039 & n4459;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = n3397 & ~n4686;
  assign n4688 = pi0039 & ~pi0786;
  assign n4689 = n4088 & n4688;
  assign n4690 = ~n4687 & ~n4689;
  assign n4691 = ~n4682 & n4690;
  assign n4692 = n3547 & ~n4691;
  assign n4693 = n3406 & n4692;
  assign n4694 = pi0039 & ~pi0314;
  assign n4695 = n2901 & n4694;
  assign n4696 = ~n4693 & ~n4695;
  assign n4697 = n4681 & n4696;
  assign n4698 = ~n3347 & n4697;
  assign n4699 = ~n4677 & n4698;
  assign n4700 = pi0039 & n2741;
  assign n4701 = ~n2583 & ~n2747;
  assign n4702 = n4679 & ~n4701;
  assign n4703 = n2795 & n4673;
  assign n4704 = ~n4702 & ~n4703;
  assign n4705 = ~n2736 & ~n2803;
  assign n4706 = ~n2749 & n4705;
  assign n4707 = n2740 & n4706;
  assign n4708 = n3540 & n4707;
  assign n4709 = pi0039 & n4708;
  assign n4710 = ~n3973 & n4709;
  assign n4711 = pi0039 & n3989;
  assign n4712 = ~n4673 & ~n4711;
  assign n4713 = n2563 & ~n4712;
  assign n4714 = ~pi0039 & pi0841;
  assign n4715 = n2698 & ~n4714;
  assign n4716 = ~n4713 & ~n4715;
  assign n4717 = ~n4710 & n4716;
  assign n4718 = n4704 & n4717;
  assign n4719 = ~n4700 & n4718;
  assign n4720 = n2591 & n4673;
  assign n4721 = n4719 & ~n4720;
  assign n4722 = pi0039 & ~n4009;
  assign n4723 = n2614 & n4722;
  assign n4724 = n3110 & n4673;
  assign n4725 = ~pi0039 & n4012;
  assign n4726 = n4011 & ~n4725;
  assign n4727 = ~n4724 & ~n4726;
  assign n4728 = ~n4723 & n4727;
  assign n4729 = ~n3102 & n4683;
  assign n4730 = n2651 & n4729;
  assign n4731 = pi0039 & ~n3102;
  assign n4732 = n4005 & n4731;
  assign n4733 = ~n4730 & ~n4732;
  assign n4734 = n4728 & n4733;
  assign n4735 = pi0039 & pi0993;
  assign n4736 = n2576 & n4735;
  assign n4737 = n2598 & n4673;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = pi1044 & n4694;
  assign n4740 = n2619 & n4739;
  assign n4741 = n2644 & n4679;
  assign n4742 = ~n4740 & ~n4741;
  assign n4743 = ~n2626 & n4742;
  assign n4744 = n4738 & n4743;
  assign n4745 = n4734 & n4744;
  assign n4746 = n4721 & n4745;
  assign n4747 = n4699 & n4746;
  assign n4748 = n2881 & n4683;
  assign n4749 = n2726 & n4748;
  assign n4750 = n2854 & n4673;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = pi0039 & n4124;
  assign n4753 = n2858 & n4679;
  assign n4754 = ~n4752 & ~n4753;
  assign n4755 = n4751 & n4754;
  assign n4756 = n2847 & n4679;
  assign n4757 = n2834 & n4739;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n3072 & n4673;
  assign n4760 = n4758 & ~n4759;
  assign n4761 = ~n2827 & n4679;
  assign n4762 = n3066 & n4673;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = n2831 & ~n4714;
  assign n4765 = n2851 & n4694;
  assign n4766 = ~n4764 & ~n4765;
  assign n4767 = n4763 & n4766;
  assign n4768 = n4760 & n4767;
  assign n4769 = n4755 & n4768;
  assign n4770 = n2913 & n4673;
  assign n4771 = pi0039 & n4043;
  assign n4772 = n2930 & n4771;
  assign n4773 = pi0039 & ~n3553;
  assign n4774 = n4497 & n4773;
  assign n4775 = ~n4772 & ~n4774;
  assign n4776 = ~n4770 & n4775;
  assign n4777 = n2917 & n4679;
  assign n4778 = pi0039 & n2926;
  assign n4779 = ~pi1076 & n4778;
  assign n4780 = n2936 & n4694;
  assign n4781 = ~n4402 & n4694;
  assign n4782 = ~n4780 & ~n4781;
  assign n4783 = ~n4779 & n4782;
  assign n4784 = n3042 & n4673;
  assign n4785 = n4783 & ~n4784;
  assign n4786 = ~n4777 & n4785;
  assign n4787 = n4776 & n4786;
  assign n4788 = n3033 & n4673;
  assign n4789 = n4787 & ~n4788;
  assign n4790 = n2910 & n4673;
  assign n4791 = pi0039 & n2726;
  assign n4792 = n4066 & n4791;
  assign n4793 = ~n4790 & ~n4792;
  assign n4794 = n2569 & n4673;
  assign n4795 = pi0039 & n4062;
  assign n4796 = ~n4794 & ~n4795;
  assign n4797 = ~n4105 & n4694;
  assign n4798 = n4796 & ~n4797;
  assign n4799 = pi0039 & n4336;
  assign n4800 = n4798 & ~n4799;
  assign n4801 = n4793 & n4800;
  assign n4802 = n4789 & n4801;
  assign n4803 = n4769 & n4802;
  assign po0197 = ~n4747 | ~n4803;
  assign n4805 = pi0040 & ~pi0314;
  assign n4806 = pi1044 & n4805;
  assign n4807 = n2619 & n4806;
  assign n4808 = pi0040 & pi0841;
  assign n4809 = n2644 & n4808;
  assign n4810 = ~n4807 & ~n4809;
  assign n4811 = pi0040 & n4062;
  assign n4812 = n2698 & n4808;
  assign n4813 = pi0024 & pi0040;
  assign n4814 = n2795 & n4813;
  assign n4815 = ~n4812 & ~n4814;
  assign n4816 = ~n4701 & n4808;
  assign n4817 = n4815 & ~n4816;
  assign n4818 = pi0040 & n2741;
  assign n4819 = pi0040 & n3102;
  assign n4820 = ~pi0024 & n4819;
  assign n4821 = ~n4813 & ~n4820;
  assign n4822 = n2563 & ~n4821;
  assign n4823 = ~n4818 & ~n4822;
  assign n4824 = n4817 & n4823;
  assign n4825 = ~n2679 & n4824;
  assign n4826 = pi0040 & n4579;
  assign n4827 = ~n4105 & n4805;
  assign n4828 = n2569 & n4813;
  assign n4829 = ~n4827 & ~n4828;
  assign n4830 = n2598 & n4813;
  assign n4831 = n4829 & ~n4830;
  assign n4832 = ~n4826 & n4831;
  assign n4833 = n4825 & n4832;
  assign n4834 = n2910 & n4813;
  assign n4835 = pi0040 & n2726;
  assign n4836 = n4066 & n4835;
  assign n4837 = ~n4834 & ~n4836;
  assign n4838 = n4833 & n4837;
  assign n4839 = ~n4811 & n4838;
  assign n4840 = n4810 & n4839;
  assign n4841 = pi0040 & n3967;
  assign n4842 = n2604 & n4841;
  assign n4843 = pi0040 & n4585;
  assign n4844 = n2917 & n4808;
  assign n4845 = n2913 & n4813;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = n2936 & n4805;
  assign n4848 = n4846 & ~n4847;
  assign n4849 = pi0040 & n4043;
  assign n4850 = n2930 & n4849;
  assign n4851 = pi0040 & ~n3553;
  assign n4852 = n4497 & n4851;
  assign n4853 = ~n4850 & ~n4852;
  assign n4854 = ~n4402 & n4805;
  assign n4855 = n4853 & ~n4854;
  assign n4856 = n3042 & n4813;
  assign n4857 = pi0040 & n4504;
  assign n4858 = ~n4856 & ~n4857;
  assign n4859 = n4855 & n4858;
  assign n4860 = n4848 & n4859;
  assign n4861 = n3033 & n4813;
  assign n4862 = n4860 & ~n4861;
  assign n4863 = pi0040 & n4006;
  assign n4864 = pi0040 & ~n4014;
  assign n4865 = n3110 & n4813;
  assign n4866 = ~n4864 & ~n4865;
  assign n4867 = pi0040 & po0740;
  assign n4868 = n2651 & n4867;
  assign n4869 = ~n3102 & n4868;
  assign n4870 = n4866 & ~n4869;
  assign n4871 = ~n4863 & n4870;
  assign n4872 = n2591 & n4813;
  assign n4873 = n4871 & ~n4872;
  assign n4874 = n4862 & n4873;
  assign n4875 = ~n4843 & n4874;
  assign n4876 = ~n4842 & n4875;
  assign n4877 = n4840 & n4876;
  assign n4878 = n3057 & n4813;
  assign n4879 = pi0040 & ~n3057;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = n4083 & ~n4880;
  assign n4882 = n2901 & n4805;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = n2681 & n4813;
  assign n4885 = ~n4077 & n4808;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = pi0040 & n4089;
  assign n4888 = pi0040 & n4091;
  assign n4889 = pi0040 & n3128;
  assign n4890 = ~n4094 & n4889;
  assign n4891 = ~n4097 & n4867;
  assign n4892 = ~n4890 & ~n4891;
  assign n4893 = n3397 & ~n4892;
  assign n4894 = ~n4888 & ~n4893;
  assign n4895 = ~n4887 & n4894;
  assign n4896 = n4087 & ~n4895;
  assign n4897 = n4886 & ~n4896;
  assign n4898 = n4883 & n4897;
  assign n4899 = ~n3072 & n4813;
  assign n4900 = n2847 & n4808;
  assign n4901 = n2834 & n4806;
  assign n4902 = ~n4900 & ~n4901;
  assign n4903 = n2858 & n4808;
  assign n4904 = pi0040 & n4124;
  assign n4905 = n2854 & n4813;
  assign n4906 = n2881 & n4867;
  assign n4907 = n2726 & n4906;
  assign n4908 = ~n4905 & ~n4907;
  assign n4909 = ~n4904 & n4908;
  assign n4910 = ~n4903 & n4909;
  assign n4911 = ~n4133 & n4808;
  assign n4912 = n4910 & ~n4911;
  assign n4913 = n2851 & n4805;
  assign n4914 = n3066 & n4813;
  assign n4915 = ~n4913 & ~n4914;
  assign n4916 = n4912 & n4915;
  assign n4917 = n4902 & n4916;
  assign n4918 = ~n4899 & n4917;
  assign n4919 = n4898 & n4918;
  assign po0198 = ~n4877 | ~n4919;
  assign n4921 = pi0039 & n4219;
  assign n4922 = n2714 & n3481;
  assign n4923 = ~n4272 & n4922;
  assign n4924 = n4921 & n4923;
  assign n4925 = ~pi0480 & pi0949;
  assign n4926 = n2604 & n4925;
  assign n4927 = ~pi0250 & pi0252;
  assign n4928 = ~pi0959 & n4927;
  assign n4929 = n2813 & n4928;
  assign n4930 = pi0901 & n4929;
  assign po0637 = n4926 | n4930;
  assign n4932 = ~pi0228 & ~po0637;
  assign n4933 = ~n3546 & ~n3555;
  assign n4934 = n3563 & n4933;
  assign n4935 = ~n3568 & n4934;
  assign n4936 = ~n3551 & ~n3570;
  assign n4937 = pi0228 & n4936;
  assign n4938 = n4935 & n4937;
  assign n4939 = ~n4932 & ~n4938;
  assign n4940 = ~pi0044 & ~pi0101;
  assign n4941 = ~pi0041 & n4940;
  assign n4942 = pi0041 & ~n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = n4939 & ~n4943;
  assign n4945 = pi0041 & ~n4939;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = ~pi0039 & ~n4946;
  assign n4948 = ~n4924 & ~n4947;
  assign po0199 = pi0072 | ~n4948;
  assign n4950 = pi0042 & ~n4939;
  assign n4951 = ~pi0114 & ~pi0115;
  assign n4952 = ~pi0113 & ~pi0116;
  assign n4953 = ~pi0099 & n4941;
  assign n4954 = n4952 & n4953;
  assign n4955 = n4951 & n4954;
  assign n4956 = pi0042 & n4955;
  assign n4957 = ~pi0042 & ~n4955;
  assign n4958 = ~n4956 & ~n4957;
  assign n4959 = n4939 & n4958;
  assign n4960 = ~n4950 & ~n4959;
  assign n4961 = ~pi0039 & ~n4960;
  assign n4962 = ~pi0219 & ~n2429;
  assign n4963 = ~pi0199 & n2429;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = pi0200 & n2429;
  assign n4966 = pi0211 & ~n2429;
  assign n4967 = ~n4965 & ~n4966;
  assign n4968 = ~pi0208 & n2429;
  assign n4969 = ~pi0212 & ~n2429;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = ~pi0207 & n2429;
  assign n4972 = ~pi0214 & ~n2429;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = n4970 & n4973;
  assign n4975 = ~n4967 & n4974;
  assign n4976 = ~n4964 & ~n4975;
  assign n4977 = pi0039 & ~n4922;
  assign n4978 = ~n4976 & n4977;
  assign n4979 = ~n4961 & ~n4978;
  assign po0200 = ~pi0072 & ~n4979;
  assign n4981 = ~n4922 & ~n4973;
  assign n4982 = ~n4967 & n4981;
  assign n4983 = ~n4964 & n4967;
  assign n4984 = n4974 & n4983;
  assign n4985 = ~n4967 & ~n4970;
  assign n4986 = ~n4984 & ~n4985;
  assign n4987 = ~n4922 & ~n4986;
  assign n4988 = ~n4982 & ~n4987;
  assign n4989 = pi0039 & ~n4988;
  assign n4990 = pi0043 & ~n4939;
  assign n4991 = ~pi0041 & ~pi0101;
  assign n4992 = n2752 & n4991;
  assign n4993 = ~pi0044 & n4992;
  assign n4994 = ~pi0042 & n4993;
  assign n4995 = n2751 & n4994;
  assign n4996 = ~pi0114 & n4995;
  assign n4997 = pi0043 & n4996;
  assign n4998 = ~pi0043 & ~n4996;
  assign n4999 = ~n4997 & ~n4998;
  assign n5000 = n4939 & n4999;
  assign n5001 = ~n4990 & ~n5000;
  assign n5002 = ~pi0039 & ~n5001;
  assign n5003 = ~n4989 & ~n5002;
  assign po0201 = ~pi0072 & ~n5003;
  assign n5005 = pi0044 & ~n4939;
  assign n5006 = ~pi0044 & n4939;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = ~pi0039 & ~n5007;
  assign n5009 = n4272 & n4922;
  assign n5010 = n4921 & n5009;
  assign n5011 = ~n5008 & ~n5010;
  assign po0202 = ~pi0072 & ~n5011;
  assign n5013 = pi0045 & pi0993;
  assign n5014 = n2576 & n5013;
  assign n5015 = pi0024 & pi0045;
  assign n5016 = n2598 & n5015;
  assign n5017 = ~n5014 & ~n5016;
  assign n5018 = pi0045 & n4062;
  assign n5019 = pi0045 & ~pi0314;
  assign n5020 = pi1044 & n5019;
  assign n5021 = n2619 & n5020;
  assign n5022 = pi0045 & pi0841;
  assign n5023 = n2644 & n5022;
  assign n5024 = ~n5021 & ~n5023;
  assign n5025 = ~n5018 & n5024;
  assign n5026 = pi0045 & n4336;
  assign n5027 = n5025 & ~n5026;
  assign n5028 = n5017 & n5027;
  assign n5029 = ~pi0287 & pi0979;
  assign n5030 = n2777 & n5029;
  assign n5031 = n2901 & n5019;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = pi0045 & n4089;
  assign n5034 = pi0045 & n4091;
  assign n5035 = pi0045 & n3128;
  assign n5036 = ~n4094 & n5035;
  assign n5037 = pi0045 & po0740;
  assign n5038 = ~n4097 & n5037;
  assign n5039 = ~n5036 & ~n5038;
  assign n5040 = n3397 & ~n5039;
  assign n5041 = ~n5034 & ~n5040;
  assign n5042 = ~n5033 & n5041;
  assign n5043 = n2777 & ~n5042;
  assign n5044 = n3466 & n5043;
  assign n5045 = ~pi0287 & n5044;
  assign n5046 = n2681 & n5015;
  assign n5047 = ~n4077 & n5022;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = n3057 & n5015;
  assign n5050 = pi0045 & ~n3057;
  assign n5051 = ~n5049 & ~n5050;
  assign n5052 = n4083 & ~n5051;
  assign n5053 = n5048 & ~n5052;
  assign n5054 = ~n5045 & n5053;
  assign n5055 = n5032 & n5054;
  assign n5056 = n5028 & n5055;
  assign n5057 = ~n3072 & n5015;
  assign n5058 = n2847 & n5022;
  assign n5059 = n2834 & n5020;
  assign n5060 = ~n5058 & ~n5059;
  assign n5061 = n2858 & n5022;
  assign n5062 = pi0045 & n4124;
  assign n5063 = n2854 & n5015;
  assign n5064 = n2881 & n5037;
  assign n5065 = n2726 & n5064;
  assign n5066 = ~n5063 & ~n5065;
  assign n5067 = ~n5062 & n5066;
  assign n5068 = ~n5061 & n5067;
  assign n5069 = ~n4133 & n5022;
  assign n5070 = n5068 & ~n5069;
  assign n5071 = n2851 & n5019;
  assign n5072 = n3066 & n5015;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = n5070 & n5073;
  assign n5075 = n5060 & n5074;
  assign n5076 = ~n5057 & n5075;
  assign n5077 = pi0045 & n4523;
  assign n5078 = ~n3973 & n5077;
  assign n5079 = pi0045 & n3989;
  assign n5080 = ~n5015 & ~n5079;
  assign n5081 = n2563 & ~n5080;
  assign n5082 = n2795 & n5015;
  assign n5083 = ~n5081 & ~n5082;
  assign n5084 = pi0045 & n2741;
  assign n5085 = n5083 & ~n5084;
  assign n5086 = ~n5078 & n5085;
  assign n5087 = ~n3998 & n5022;
  assign n5088 = n5086 & ~n5087;
  assign n5089 = n5076 & n5088;
  assign n5090 = n2910 & n5015;
  assign n5091 = pi0045 & n2726;
  assign n5092 = n4066 & n5091;
  assign n5093 = ~n5090 & ~n5092;
  assign n5094 = pi0045 & n4006;
  assign n5095 = pi0045 & ~n4014;
  assign n5096 = n3110 & n5015;
  assign n5097 = ~n5095 & ~n5096;
  assign n5098 = n2651 & n5037;
  assign n5099 = ~n3102 & n5098;
  assign n5100 = n5097 & ~n5099;
  assign n5101 = ~n5094 & n5100;
  assign n5102 = n2591 & n5015;
  assign n5103 = n5101 & ~n5102;
  assign n5104 = ~n4105 & n5019;
  assign n5105 = n2569 & n5015;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = n2917 & n5022;
  assign n5108 = n2913 & n5015;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = n2936 & n5019;
  assign n5111 = n5109 & ~n5110;
  assign n5112 = pi0045 & n4043;
  assign n5113 = n2930 & n5112;
  assign n5114 = pi0045 & ~n3553;
  assign n5115 = n4497 & n5114;
  assign n5116 = ~n5113 & ~n5115;
  assign n5117 = ~n4402 & n5019;
  assign n5118 = n5116 & ~n5117;
  assign n5119 = n3042 & n5015;
  assign n5120 = pi0045 & n4504;
  assign n5121 = ~n5119 & ~n5120;
  assign n5122 = n5118 & n5121;
  assign n5123 = n5111 & n5122;
  assign n5124 = n3033 & n5015;
  assign n5125 = n5123 & ~n5124;
  assign n5126 = n5106 & n5125;
  assign n5127 = n5103 & n5126;
  assign n5128 = n5093 & n5127;
  assign n5129 = n5089 & n5128;
  assign po0203 = ~n5056 | ~n5129;
  assign n5131 = pi0024 & pi0046;
  assign n5132 = n2910 & n5131;
  assign n5133 = pi0046 & n2726;
  assign n5134 = n4066 & n5133;
  assign n5135 = ~n5132 & ~n5134;
  assign n5136 = pi0046 & n4006;
  assign n5137 = pi0046 & ~n4014;
  assign n5138 = n3110 & n5131;
  assign n5139 = ~n5137 & ~n5138;
  assign n5140 = pi0046 & po0740;
  assign n5141 = n2651 & n5140;
  assign n5142 = ~n3102 & n5141;
  assign n5143 = n5139 & ~n5142;
  assign n5144 = ~n5136 & n5143;
  assign n5145 = n2591 & n5131;
  assign n5146 = n5144 & ~n5145;
  assign n5147 = pi0046 & ~pi0314;
  assign n5148 = ~n4105 & n5147;
  assign n5149 = n2569 & n5131;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = pi0046 & pi0841;
  assign n5152 = n2917 & n5151;
  assign n5153 = n2913 & n5131;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = n2936 & n5147;
  assign n5156 = n5154 & ~n5155;
  assign n5157 = pi0046 & n4043;
  assign n5158 = n2930 & n5157;
  assign n5159 = pi0046 & ~n3553;
  assign n5160 = n4497 & n5159;
  assign n5161 = ~n5158 & ~n5160;
  assign n5162 = ~n4402 & n5147;
  assign n5163 = n5161 & ~n5162;
  assign n5164 = n3042 & n5131;
  assign n5165 = pi0046 & n4504;
  assign n5166 = ~n5164 & ~n5165;
  assign n5167 = n5163 & n5166;
  assign n5168 = n5156 & n5167;
  assign n5169 = n3033 & n5131;
  assign n5170 = n5168 & ~n5169;
  assign n5171 = n5150 & n5170;
  assign n5172 = n5146 & n5171;
  assign n5173 = n5135 & n5172;
  assign n5174 = ~n3072 & n5131;
  assign n5175 = n2847 & n5151;
  assign n5176 = pi1044 & n5147;
  assign n5177 = n2834 & n5176;
  assign n5178 = ~n5175 & ~n5177;
  assign n5179 = n2858 & n5151;
  assign n5180 = pi0046 & n4124;
  assign n5181 = n2854 & n5131;
  assign n5182 = n2881 & n5140;
  assign n5183 = n2726 & n5182;
  assign n5184 = ~n5181 & ~n5183;
  assign n5185 = ~n5180 & n5184;
  assign n5186 = ~n5179 & n5185;
  assign n5187 = ~n4133 & n5151;
  assign n5188 = n5186 & ~n5187;
  assign n5189 = n2851 & n5147;
  assign n5190 = n3066 & n5131;
  assign n5191 = ~n5189 & ~n5190;
  assign n5192 = n5188 & n5191;
  assign n5193 = n5178 & n5192;
  assign n5194 = ~n5174 & n5193;
  assign n5195 = pi0046 & n4523;
  assign n5196 = ~n3973 & n5195;
  assign n5197 = pi0046 & n3989;
  assign n5198 = ~n5131 & ~n5197;
  assign n5199 = n2563 & ~n5198;
  assign n5200 = n2795 & n5131;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = pi0046 & n2741;
  assign n5203 = n5201 & ~n5202;
  assign n5204 = ~n5196 & n5203;
  assign n5205 = ~n3998 & n5151;
  assign n5206 = n5204 & ~n5205;
  assign n5207 = n5194 & n5206;
  assign n5208 = pi0046 & pi0993;
  assign n5209 = n2576 & n5208;
  assign n5210 = n2598 & n5131;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = pi0046 & n4062;
  assign n5213 = n2619 & n5176;
  assign n5214 = n2644 & n5151;
  assign n5215 = ~n5213 & ~n5214;
  assign n5216 = ~n5212 & n5215;
  assign n5217 = pi0046 & n4336;
  assign n5218 = n5216 & ~n5217;
  assign n5219 = n5211 & n5218;
  assign n5220 = n2770 & n5151;
  assign n5221 = pi0046 & n4089;
  assign n5222 = pi0046 & n4091;
  assign n5223 = pi0046 & n3128;
  assign n5224 = ~n4094 & n5223;
  assign n5225 = ~n4097 & n5140;
  assign n5226 = ~n5224 & ~n5225;
  assign n5227 = n3397 & ~n5226;
  assign n5228 = ~n5222 & ~n5227;
  assign n5229 = ~n5221 & n5228;
  assign n5230 = n4087 & ~n5229;
  assign n5231 = n3057 & ~n5131;
  assign n5232 = ~pi0046 & ~n3057;
  assign n5233 = ~n5231 & ~n5232;
  assign n5234 = n4083 & n5233;
  assign n5235 = ~pi0046 & pi0841;
  assign n5236 = n2892 & ~n5235;
  assign n5237 = ~n5234 & ~n5236;
  assign n5238 = ~n5230 & n5237;
  assign n5239 = n2901 & n5147;
  assign n5240 = n5238 & ~n5239;
  assign n5241 = n2681 & n5131;
  assign n5242 = n5240 & ~n5241;
  assign n5243 = ~n5220 & n5242;
  assign n5244 = n5219 & n5243;
  assign n5245 = n5207 & n5244;
  assign po0204 = ~n5173 | ~n5245;
  assign n5247 = pi0047 & ~pi0314;
  assign n5248 = ~n4105 & n5247;
  assign n5249 = pi0024 & pi0047;
  assign n5250 = n2569 & n5249;
  assign n5251 = ~n5248 & ~n5250;
  assign n5252 = pi0047 & pi0993;
  assign n5253 = n2576 & n5252;
  assign n5254 = n2598 & n5249;
  assign n5255 = ~n5253 & ~n5254;
  assign n5256 = n5251 & n5255;
  assign n5257 = pi0047 & pi0841;
  assign n5258 = n2847 & n5257;
  assign n5259 = pi1044 & n5247;
  assign n5260 = n2834 & n5259;
  assign n5261 = ~n5258 & ~n5260;
  assign n5262 = ~n3072 & n5249;
  assign n5263 = n5261 & ~n5262;
  assign n5264 = n2851 & n5247;
  assign n5265 = n3066 & n5249;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = n2901 & n5247;
  assign n5268 = n2681 & n5249;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = ~n4077 & n5257;
  assign n5271 = n5269 & ~n5270;
  assign n5272 = pi0047 & n4124;
  assign n5273 = pi0047 & po0740;
  assign n5274 = n2726 & ~n5273;
  assign n5275 = n2881 & ~n5274;
  assign n5276 = n2854 & n5249;
  assign n5277 = ~n5275 & ~n5276;
  assign n5278 = n2858 & n5257;
  assign n5279 = n5277 & ~n5278;
  assign n5280 = ~n5272 & n5279;
  assign n5281 = ~n4133 & n5257;
  assign n5282 = n5280 & ~n5281;
  assign n5283 = n5271 & n5282;
  assign n5284 = n5266 & n5283;
  assign n5285 = n5263 & n5284;
  assign n5286 = pi0047 & n4091;
  assign n5287 = ~n4097 & n5273;
  assign n5288 = pi0047 & n4459;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = n3397 & ~n5289;
  assign n5291 = pi0047 & ~pi0786;
  assign n5292 = n4088 & n5291;
  assign n5293 = ~n5290 & ~n5292;
  assign n5294 = ~n5286 & n5293;
  assign n5295 = n4087 & ~n5294;
  assign n5296 = n2888 & n3468;
  assign n5297 = n3057 & n5249;
  assign n5298 = pi0047 & ~n3057;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = n4083 & ~n5299;
  assign n5301 = ~n5296 & ~n5300;
  assign n5302 = ~n5295 & n5301;
  assign n5303 = n5285 & n5302;
  assign n5304 = n2619 & n5259;
  assign n5305 = n2644 & n5257;
  assign n5306 = ~n5304 & ~n5305;
  assign n5307 = n2917 & n5257;
  assign n5308 = n2913 & n5249;
  assign n5309 = ~n5307 & ~n5308;
  assign n5310 = n2936 & n5247;
  assign n5311 = n5309 & ~n5310;
  assign n5312 = ~n2726 & ~n4064;
  assign n5313 = pi0047 & ~n4064;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = n2516 & ~n5314;
  assign n5316 = pi0047 & n4043;
  assign n5317 = n2930 & n5316;
  assign n5318 = pi0047 & ~n3553;
  assign n5319 = n4497 & n5318;
  assign n5320 = ~n5317 & ~n5319;
  assign n5321 = ~n4402 & n5247;
  assign n5322 = n5320 & ~n5321;
  assign n5323 = pi0047 & n4504;
  assign n5324 = n5322 & ~n5323;
  assign n5325 = ~n5315 & n5324;
  assign n5326 = n5311 & n5325;
  assign n5327 = ~n2910 & ~n3033;
  assign n5328 = ~n3042 & n5327;
  assign n5329 = n5249 & ~n5328;
  assign n5330 = n5326 & ~n5329;
  assign n5331 = pi0047 & n4006;
  assign n5332 = pi0047 & ~n4014;
  assign n5333 = n3110 & n5249;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = n2651 & n5273;
  assign n5336 = ~n3102 & n5335;
  assign n5337 = n5334 & ~n5336;
  assign n5338 = ~n5331 & n5337;
  assign n5339 = n2591 & n5249;
  assign n5340 = n5338 & ~n5339;
  assign n5341 = n5330 & n5340;
  assign n5342 = n5306 & n5341;
  assign n5343 = pi0047 & n2741;
  assign n5344 = n2795 & n5249;
  assign n5345 = pi0047 & n4523;
  assign n5346 = ~n3973 & n5345;
  assign n5347 = pi0047 & ~po0740;
  assign n5348 = ~n3468 & ~n5347;
  assign n5349 = n3552 & ~n5348;
  assign n5350 = n2563 & n5249;
  assign n5351 = ~n5349 & ~n5350;
  assign n5352 = ~n5346 & n5351;
  assign n5353 = ~n5344 & n5352;
  assign n5354 = ~n5343 & n5353;
  assign n5355 = ~n3998 & n5257;
  assign n5356 = n5354 & ~n5355;
  assign n5357 = pi0047 & n4336;
  assign n5358 = pi0047 & n4062;
  assign n5359 = ~n5357 & ~n5358;
  assign n5360 = n5356 & n5359;
  assign n5361 = n5342 & n5360;
  assign n5362 = n5303 & n5361;
  assign po0205 = ~n5256 | ~n5362;
  assign n5364 = pi0048 & pi0841;
  assign n5365 = n2917 & n5364;
  assign n5366 = pi0024 & pi0048;
  assign n5367 = n2913 & n5366;
  assign n5368 = ~n5365 & ~n5367;
  assign n5369 = pi0048 & ~pi0314;
  assign n5370 = n2936 & n5369;
  assign n5371 = n5368 & ~n5370;
  assign n5372 = pi0048 & n4043;
  assign n5373 = n2930 & n5372;
  assign n5374 = pi0048 & ~n3553;
  assign n5375 = n4497 & n5374;
  assign n5376 = ~n5373 & ~n5375;
  assign n5377 = ~n4402 & n5369;
  assign n5378 = n5376 & ~n5377;
  assign n5379 = n3042 & n5366;
  assign n5380 = pi0048 & n4504;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = n5378 & n5381;
  assign n5383 = n5371 & n5382;
  assign n5384 = n3033 & n5366;
  assign n5385 = n5383 & ~n5384;
  assign n5386 = pi0048 & n4006;
  assign n5387 = pi0048 & ~n4014;
  assign n5388 = n3110 & n5366;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = pi0048 & po0740;
  assign n5391 = n2651 & n5390;
  assign n5392 = ~n3102 & n5391;
  assign n5393 = n5389 & ~n5392;
  assign n5394 = ~n5386 & n5393;
  assign n5395 = n2591 & n5366;
  assign n5396 = n5394 & ~n5395;
  assign n5397 = n2910 & n5366;
  assign n5398 = pi0048 & n2726;
  assign n5399 = n4066 & n5398;
  assign n5400 = ~n5397 & ~n5399;
  assign n5401 = n5396 & n5400;
  assign n5402 = n5385 & n5401;
  assign n5403 = ~n3072 & n5366;
  assign n5404 = n2847 & n5364;
  assign n5405 = pi1044 & n5369;
  assign n5406 = n2834 & n5405;
  assign n5407 = ~n5404 & ~n5406;
  assign n5408 = n2858 & n5364;
  assign n5409 = pi0048 & n4124;
  assign n5410 = n2854 & n5366;
  assign n5411 = n2881 & n5390;
  assign n5412 = n2726 & n5411;
  assign n5413 = ~n5410 & ~n5412;
  assign n5414 = ~n5409 & n5413;
  assign n5415 = ~n5408 & n5414;
  assign n5416 = ~n4133 & n5364;
  assign n5417 = n5415 & ~n5416;
  assign n5418 = n2851 & n5369;
  assign n5419 = n3066 & n5366;
  assign n5420 = ~n5418 & ~n5419;
  assign n5421 = n5417 & n5420;
  assign n5422 = n5407 & n5421;
  assign n5423 = ~n5403 & n5422;
  assign n5424 = n5402 & n5423;
  assign n5425 = pi0048 & pi0993;
  assign n5426 = n2576 & n5425;
  assign n5427 = n2598 & n5366;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = pi0048 & n4062;
  assign n5430 = n2619 & n5405;
  assign n5431 = n2644 & n5364;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = ~n5429 & n5432;
  assign n5434 = pi0048 & n4336;
  assign n5435 = n5433 & ~n5434;
  assign n5436 = n5428 & n5435;
  assign n5437 = n3057 & n5366;
  assign n5438 = pi0048 & ~n3057;
  assign n5439 = ~n5437 & ~n5438;
  assign n5440 = n4083 & ~n5439;
  assign n5441 = n2901 & n5369;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = n2681 & n5366;
  assign n5444 = ~n4077 & n5364;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = pi0048 & n4089;
  assign n5447 = pi0048 & n4091;
  assign n5448 = pi0048 & n3128;
  assign n5449 = ~n4094 & n5448;
  assign n5450 = ~n4097 & n5390;
  assign n5451 = ~n5449 & ~n5450;
  assign n5452 = n3397 & ~n5451;
  assign n5453 = ~n5447 & ~n5452;
  assign n5454 = ~n5446 & n5453;
  assign n5455 = n4087 & ~n5454;
  assign n5456 = n5445 & ~n5455;
  assign n5457 = n5442 & n5456;
  assign n5458 = n5436 & n5457;
  assign n5459 = pi0048 & n4523;
  assign n5460 = ~n3973 & n5459;
  assign n5461 = pi0048 & n3989;
  assign n5462 = ~n5366 & ~n5461;
  assign n5463 = n2563 & ~n5462;
  assign n5464 = n2795 & n5366;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = pi0048 & n2741;
  assign n5467 = n5465 & ~n5466;
  assign n5468 = ~n5460 & n5467;
  assign n5469 = ~n3998 & n5364;
  assign n5470 = n5468 & ~n5469;
  assign n5471 = ~n4105 & n5369;
  assign n5472 = n2569 & n5366;
  assign n5473 = ~n5471 & ~n5472;
  assign n5474 = n5470 & n5473;
  assign n5475 = n5458 & n5474;
  assign po0206 = ~n5424 | ~n5475;
  assign n5477 = pi0024 & pi0049;
  assign n5478 = n2910 & n5477;
  assign n5479 = pi0049 & n2726;
  assign n5480 = n4066 & n5479;
  assign n5481 = ~n5478 & ~n5480;
  assign n5482 = pi0049 & pi0841;
  assign n5483 = n2917 & n5482;
  assign n5484 = n2913 & n5477;
  assign n5485 = ~n5483 & ~n5484;
  assign n5486 = pi0049 & ~pi0314;
  assign n5487 = n2936 & n5486;
  assign n5488 = n5485 & ~n5487;
  assign n5489 = ~n3553 & n4497;
  assign n5490 = pi0049 & n5489;
  assign n5491 = n2930 & n4043;
  assign n5492 = pi0049 & n5491;
  assign n5493 = ~n5490 & ~n5492;
  assign n5494 = ~n4402 & n5486;
  assign n5495 = n5493 & ~n5494;
  assign n5496 = n3042 & n5477;
  assign n5497 = pi0049 & n4504;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = n5495 & n5498;
  assign n5500 = n5488 & n5499;
  assign n5501 = n3033 & n5477;
  assign n5502 = n5500 & ~n5501;
  assign n5503 = pi0049 & n4006;
  assign n5504 = pi0049 & ~n4014;
  assign n5505 = n3110 & n5477;
  assign n5506 = ~n5504 & ~n5505;
  assign n5507 = pi0049 & po0740;
  assign n5508 = n2651 & n5507;
  assign n5509 = ~n3102 & n5508;
  assign n5510 = n5506 & ~n5509;
  assign n5511 = ~n5503 & n5510;
  assign n5512 = n2591 & n5477;
  assign n5513 = n5511 & ~n5512;
  assign n5514 = n5502 & n5513;
  assign n5515 = n5481 & n5514;
  assign n5516 = pi1044 & n5486;
  assign n5517 = n2619 & n5516;
  assign n5518 = n2644 & n5482;
  assign n5519 = ~n5517 & ~n5518;
  assign n5520 = pi0049 & n4336;
  assign n5521 = pi0049 & n4062;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = n5519 & n5522;
  assign n5524 = n5515 & n5523;
  assign n5525 = pi0049 & n4523;
  assign n5526 = ~n3973 & n5525;
  assign n5527 = pi0049 & n3989;
  assign n5528 = ~n5477 & ~n5527;
  assign n5529 = n2563 & ~n5528;
  assign n5530 = n2795 & n5477;
  assign n5531 = ~n5529 & ~n5530;
  assign n5532 = pi0049 & n2741;
  assign n5533 = n5531 & ~n5532;
  assign n5534 = ~n5526 & n5533;
  assign n5535 = ~n3998 & n5482;
  assign n5536 = n5534 & ~n5535;
  assign n5537 = n3057 & n5477;
  assign n5538 = pi0049 & ~n3057;
  assign n5539 = ~n5537 & ~n5538;
  assign n5540 = n4083 & ~n5539;
  assign n5541 = n2901 & n5486;
  assign n5542 = ~n5540 & ~n5541;
  assign n5543 = n2681 & n5477;
  assign n5544 = ~n4077 & n5482;
  assign n5545 = ~n5543 & ~n5544;
  assign n5546 = pi0049 & n4089;
  assign n5547 = pi0049 & n4091;
  assign n5548 = pi0049 & n3128;
  assign n5549 = ~n4094 & n5548;
  assign n5550 = ~n4097 & n5507;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = n3397 & ~n5551;
  assign n5553 = ~n5547 & ~n5552;
  assign n5554 = ~n5546 & n5553;
  assign n5555 = n4087 & ~n5554;
  assign n5556 = n5545 & ~n5555;
  assign n5557 = n5542 & n5556;
  assign n5558 = ~n2788 & ~n2854;
  assign n5559 = n5477 & ~n5558;
  assign n5560 = n2847 & n5482;
  assign n5561 = n2834 & n5516;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = pi0024 & ~pi0049;
  assign n5564 = n3071 & ~n5563;
  assign n5565 = n2881 & n5507;
  assign n5566 = n2726 & n5565;
  assign n5567 = pi0049 & n4124;
  assign n5568 = n2858 & n5482;
  assign n5569 = ~n5567 & ~n5568;
  assign n5570 = ~n5566 & n5569;
  assign n5571 = ~n5564 & n5570;
  assign n5572 = ~n4133 & n5482;
  assign n5573 = n5571 & ~n5572;
  assign n5574 = n2851 & n5486;
  assign n5575 = n3066 & n5477;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = n5573 & n5576;
  assign n5578 = n5562 & n5577;
  assign n5579 = ~n5559 & n5578;
  assign n5580 = n5557 & n5579;
  assign n5581 = ~n4105 & n5486;
  assign n5582 = n2569 & n5477;
  assign n5583 = ~n5581 & ~n5582;
  assign n5584 = pi0049 & pi0993;
  assign n5585 = n2576 & n5584;
  assign n5586 = n2598 & n5477;
  assign n5587 = ~n5585 & ~n5586;
  assign n5588 = n5583 & n5587;
  assign n5589 = n5580 & n5588;
  assign n5590 = n5536 & n5589;
  assign po0207 = ~n5524 | ~n5590;
  assign n5592 = pi0050 & pi0841;
  assign n5593 = n2847 & n5592;
  assign n5594 = pi0050 & ~pi0314;
  assign n5595 = pi1044 & n5594;
  assign n5596 = n2834 & n5595;
  assign n5597 = ~n5593 & ~n5596;
  assign n5598 = pi0024 & pi0050;
  assign n5599 = ~n3072 & n5598;
  assign n5600 = n5597 & ~n5599;
  assign n5601 = n2851 & n5594;
  assign n5602 = n3066 & n5598;
  assign n5603 = ~n5601 & ~n5602;
  assign n5604 = ~n3998 & n5592;
  assign n5605 = n2598 & n5598;
  assign n5606 = pi0050 & pi0993;
  assign n5607 = n2576 & n5606;
  assign n5608 = ~n5605 & ~n5607;
  assign n5609 = ~n4105 & n5594;
  assign n5610 = n2569 & n5598;
  assign n5611 = ~n5609 & ~n5610;
  assign n5612 = pi0050 & n3989;
  assign n5613 = ~n5598 & ~n5612;
  assign n5614 = n2563 & ~n5613;
  assign n5615 = n2795 & n5598;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = n5611 & n5616;
  assign n5618 = n5608 & n5617;
  assign n5619 = ~n5604 & n5618;
  assign n5620 = pi0050 & n3540;
  assign n5621 = ~n4058 & ~n5620;
  assign n5622 = ~n4061 & n5621;
  assign n5623 = n2813 & ~n5622;
  assign n5624 = n5619 & ~n5623;
  assign n5625 = ~n2736 & n3540;
  assign n5626 = ~n3971 & n5625;
  assign n5627 = ~n2749 & ~n3973;
  assign n5628 = pi0050 & n5627;
  assign n5629 = n5626 & n5628;
  assign n5630 = pi0050 & n2736;
  assign n5631 = ~n5629 & ~n5630;
  assign n5632 = ~n3433 & n5631;
  assign n5633 = n2740 & ~n5632;
  assign n5634 = n5624 & ~n5633;
  assign n5635 = pi0050 & n4067;
  assign n5636 = n2910 & n5598;
  assign n5637 = ~n5635 & ~n5636;
  assign n5638 = n3033 & n5598;
  assign n5639 = n5637 & ~n5638;
  assign n5640 = ~pi0024 & n4027;
  assign n5641 = ~po0840 & n5640;
  assign n5642 = n4028 & n5641;
  assign n5643 = n3042 & n5598;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = n2936 & n5594;
  assign n5646 = n2913 & n5598;
  assign n5647 = n2917 & n5592;
  assign n5648 = ~n5646 & ~n5647;
  assign n5649 = pi0050 & n4504;
  assign n5650 = pi0050 & n4043;
  assign n5651 = n2930 & n5650;
  assign n5652 = pi0050 & ~n3553;
  assign n5653 = n4497 & n5652;
  assign n5654 = ~n5651 & ~n5653;
  assign n5655 = ~n4402 & n5594;
  assign n5656 = n5654 & ~n5655;
  assign n5657 = ~n5649 & n5656;
  assign n5658 = n5648 & n5657;
  assign n5659 = ~n5645 & n5658;
  assign n5660 = n5644 & n5659;
  assign n5661 = pi0050 & n4336;
  assign n5662 = pi0050 & n4006;
  assign n5663 = pi0050 & ~n4014;
  assign n5664 = n3110 & n5598;
  assign n5665 = ~n5663 & ~n5664;
  assign n5666 = pi0050 & po0740;
  assign n5667 = n2651 & n5666;
  assign n5668 = ~n3102 & n5667;
  assign n5669 = n5665 & ~n5668;
  assign n5670 = ~n5662 & n5669;
  assign n5671 = n2591 & n5598;
  assign n5672 = n5670 & ~n5671;
  assign n5673 = n2619 & n5595;
  assign n5674 = n2644 & n5592;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = n5672 & n5675;
  assign n5677 = ~n5661 & n5676;
  assign n5678 = n5660 & n5677;
  assign n5679 = n5639 & n5678;
  assign n5680 = n5634 & n5679;
  assign n5681 = pi0050 & n4089;
  assign n5682 = pi0050 & n4091;
  assign n5683 = pi0050 & n3128;
  assign n5684 = ~n4094 & n5683;
  assign n5685 = ~n4097 & n5666;
  assign n5686 = ~n5684 & ~n5685;
  assign n5687 = n3397 & ~n5686;
  assign n5688 = ~n5682 & ~n5687;
  assign n5689 = ~n5681 & n5688;
  assign n5690 = n4087 & ~n5689;
  assign n5691 = n3057 & n5598;
  assign n5692 = pi0050 & ~n3057;
  assign n5693 = ~n5691 & ~n5692;
  assign n5694 = n4083 & ~n5693;
  assign n5695 = n2901 & n5594;
  assign n5696 = ~n5694 & ~n5695;
  assign n5697 = n2881 & n5666;
  assign n5698 = n2726 & n5697;
  assign n5699 = n2854 & n5598;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = n2858 & n5592;
  assign n5702 = pi0050 & n4124;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = n5700 & n5703;
  assign n5705 = n2681 & n5598;
  assign n5706 = ~n4077 & n5592;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = n5704 & n5707;
  assign n5709 = n5696 & n5708;
  assign n5710 = ~n5690 & n5709;
  assign n5711 = ~n4133 & n5592;
  assign n5712 = n5710 & ~n5711;
  assign n5713 = n5680 & n5712;
  assign n5714 = n5603 & n5713;
  assign po0208 = ~n5600 | ~n5714;
  assign n5716 = pi0051 & n4006;
  assign n5717 = pi0051 & ~n4014;
  assign n5718 = pi0024 & pi0051;
  assign n5719 = n3110 & n5718;
  assign n5720 = ~n5717 & ~n5719;
  assign n5721 = pi0051 & po0740;
  assign n5722 = n2651 & n5721;
  assign n5723 = ~n3102 & n5722;
  assign n5724 = n5720 & ~n5723;
  assign n5725 = ~n5716 & n5724;
  assign n5726 = n2591 & n5718;
  assign n5727 = n5725 & ~n5726;
  assign n5728 = pi0051 & n4062;
  assign n5729 = n2910 & n5718;
  assign n5730 = pi0051 & n2726;
  assign n5731 = n4066 & n5730;
  assign n5732 = ~n5729 & ~n5731;
  assign n5733 = pi0051 & ~pi0314;
  assign n5734 = pi1044 & n5733;
  assign n5735 = n2619 & n5734;
  assign n5736 = pi0051 & pi0841;
  assign n5737 = n2644 & n5736;
  assign n5738 = ~n5735 & ~n5737;
  assign n5739 = n5732 & n5738;
  assign n5740 = ~n5728 & n5739;
  assign n5741 = pi0051 & n3967;
  assign n5742 = n2604 & n5741;
  assign n5743 = n5740 & ~n5742;
  assign n5744 = n2917 & n5736;
  assign n5745 = n2913 & n5718;
  assign n5746 = ~n5744 & ~n5745;
  assign n5747 = n2936 & n5733;
  assign n5748 = n5746 & ~n5747;
  assign n5749 = pi0051 & n4043;
  assign n5750 = n2930 & n5749;
  assign n5751 = pi0051 & ~n3553;
  assign n5752 = n4497 & n5751;
  assign n5753 = ~n5750 & ~n5752;
  assign n5754 = ~n4402 & n5733;
  assign n5755 = n5753 & ~n5754;
  assign n5756 = n3042 & n5718;
  assign n5757 = pi0051 & n4504;
  assign n5758 = ~n5756 & ~n5757;
  assign n5759 = n5755 & n5758;
  assign n5760 = n5748 & n5759;
  assign n5761 = n3033 & n5718;
  assign n5762 = n5760 & ~n5761;
  assign n5763 = n5743 & n5762;
  assign n5764 = n5727 & n5763;
  assign n5765 = pi0051 & n4708;
  assign n5766 = ~n3973 & n5765;
  assign n5767 = n2698 & n5736;
  assign n5768 = n2795 & n5718;
  assign n5769 = ~n5767 & ~n5768;
  assign n5770 = ~n4701 & n5736;
  assign n5771 = n5769 & ~n5770;
  assign n5772 = pi0051 & n2741;
  assign n5773 = pi0051 & n3102;
  assign n5774 = ~pi0024 & n5773;
  assign n5775 = ~n5718 & ~n5774;
  assign n5776 = n2563 & ~n5775;
  assign n5777 = ~n5772 & ~n5776;
  assign n5778 = n5771 & n5777;
  assign n5779 = ~n2694 & n5778;
  assign n5780 = pi0051 & n4579;
  assign n5781 = ~n4105 & n5733;
  assign n5782 = n2569 & n5718;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = n2598 & n5718;
  assign n5785 = n5783 & ~n5784;
  assign n5786 = ~n5780 & n5785;
  assign n5787 = n5779 & n5786;
  assign n5788 = ~n5766 & n5787;
  assign n5789 = n5764 & n5788;
  assign n5790 = n3057 & n5718;
  assign n5791 = pi0051 & ~n3057;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = n4083 & ~n5792;
  assign n5794 = n2901 & n5733;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = n2681 & n5718;
  assign n5797 = ~n4077 & n5736;
  assign n5798 = ~n5796 & ~n5797;
  assign n5799 = pi0051 & n4089;
  assign n5800 = pi0051 & n4091;
  assign n5801 = pi0051 & n3128;
  assign n5802 = ~n4094 & n5801;
  assign n5803 = ~n4097 & n5721;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = n3397 & ~n5804;
  assign n5806 = ~n5800 & ~n5805;
  assign n5807 = ~n5799 & n5806;
  assign n5808 = n4087 & ~n5807;
  assign n5809 = n5798 & ~n5808;
  assign n5810 = n5795 & n5809;
  assign n5811 = ~n3072 & n5718;
  assign n5812 = n2847 & n5736;
  assign n5813 = n2834 & n5734;
  assign n5814 = ~n5812 & ~n5813;
  assign n5815 = n2858 & n5736;
  assign n5816 = pi0051 & n4124;
  assign n5817 = n2854 & n5718;
  assign n5818 = n2881 & n5721;
  assign n5819 = n2726 & n5818;
  assign n5820 = ~n5817 & ~n5819;
  assign n5821 = ~n5816 & n5820;
  assign n5822 = ~n5815 & n5821;
  assign n5823 = ~n4133 & n5736;
  assign n5824 = n5822 & ~n5823;
  assign n5825 = n2851 & n5733;
  assign n5826 = n3066 & n5718;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = n5824 & n5827;
  assign n5829 = n5814 & n5828;
  assign n5830 = ~n5811 & n5829;
  assign n5831 = n5810 & n5830;
  assign po0209 = ~n5789 | ~n5831;
  assign n5833 = ~n4974 & n4977;
  assign n5834 = n4983 & n5833;
  assign n5835 = ~pi0052 & ~n4939;
  assign n5836 = ~pi0116 & n2752;
  assign n5837 = n4941 & n5836;
  assign n5838 = n4951 & n5837;
  assign n5839 = n2755 & n5838;
  assign n5840 = ~pi0052 & n5839;
  assign n5841 = pi0052 & ~n5839;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = n4939 & n5842;
  assign n5844 = ~pi0039 & ~n5843;
  assign n5845 = ~n5835 & n5844;
  assign n5846 = ~n5834 & ~n5845;
  assign po0210 = ~pi0072 & ~n5846;
  assign n5848 = pi0024 & pi0053;
  assign n5849 = n2910 & n5848;
  assign n5850 = pi0053 & n2726;
  assign n5851 = n4066 & n5850;
  assign n5852 = ~n5849 & ~n5851;
  assign n5853 = pi0053 & n4006;
  assign n5854 = pi0053 & ~n4014;
  assign n5855 = n3110 & n5848;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = pi0053 & po0740;
  assign n5858 = n2651 & n5857;
  assign n5859 = ~n3102 & n5858;
  assign n5860 = n5856 & ~n5859;
  assign n5861 = ~n5853 & n5860;
  assign n5862 = n2591 & n5848;
  assign n5863 = n5861 & ~n5862;
  assign n5864 = pi0053 & ~pi0314;
  assign n5865 = ~n4105 & n5864;
  assign n5866 = n2569 & n5848;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = pi0053 & pi0841;
  assign n5869 = n2917 & n5868;
  assign n5870 = n2913 & n5848;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = n2936 & n5864;
  assign n5873 = n5871 & ~n5872;
  assign n5874 = pi0053 & n4043;
  assign n5875 = n2930 & n5874;
  assign n5876 = pi0053 & ~n3553;
  assign n5877 = n4497 & n5876;
  assign n5878 = ~n5875 & ~n5877;
  assign n5879 = ~n4402 & n5864;
  assign n5880 = n5878 & ~n5879;
  assign n5881 = n3042 & n5848;
  assign n5882 = pi0053 & n4504;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = n5880 & n5883;
  assign n5885 = n5873 & n5884;
  assign n5886 = n3033 & n5848;
  assign n5887 = n5885 & ~n5886;
  assign n5888 = n5867 & n5887;
  assign n5889 = n5863 & n5888;
  assign n5890 = n5852 & n5889;
  assign n5891 = n3403 & n3464;
  assign n5892 = n2777 & n5891;
  assign n5893 = n2901 & n5864;
  assign n5894 = ~n5892 & ~n5893;
  assign n5895 = pi0053 & n3128;
  assign n5896 = ~n4094 & n5895;
  assign n5897 = ~n4097 & n5857;
  assign n5898 = ~n5896 & ~n5897;
  assign n5899 = n3397 & ~n3405;
  assign n5900 = ~n5898 & n5899;
  assign n5901 = ~n4089 & ~n4091;
  assign n5902 = ~n3405 & ~n5901;
  assign n5903 = pi0053 & n5902;
  assign n5904 = ~n5900 & ~n5903;
  assign n5905 = n3465 & ~n5904;
  assign n5906 = n2681 & n5848;
  assign n5907 = ~n4077 & n5868;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = n3057 & n5848;
  assign n5910 = pi0053 & ~n3057;
  assign n5911 = ~n5909 & ~n5910;
  assign n5912 = n4083 & ~n5911;
  assign n5913 = n5908 & ~n5912;
  assign n5914 = ~n5905 & n5913;
  assign n5915 = n5894 & n5914;
  assign n5916 = pi0053 & n4708;
  assign n5917 = ~n3973 & n5916;
  assign n5918 = pi0053 & n3989;
  assign n5919 = ~n5848 & ~n5918;
  assign n5920 = n2563 & ~n5919;
  assign n5921 = n2795 & n5848;
  assign n5922 = ~n5920 & ~n5921;
  assign n5923 = pi0053 & n2741;
  assign n5924 = n5922 & ~n5923;
  assign n5925 = ~n5917 & n5924;
  assign n5926 = ~n3998 & n5868;
  assign n5927 = n5925 & ~n5926;
  assign n5928 = n5915 & n5927;
  assign n5929 = pi1044 & n5864;
  assign n5930 = n2619 & n5929;
  assign n5931 = n2644 & n5868;
  assign n5932 = ~n5930 & ~n5931;
  assign n5933 = pi0053 & pi0993;
  assign n5934 = n2576 & n5933;
  assign n5935 = n2598 & n5848;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = pi0053 & n4336;
  assign n5938 = pi0053 & n4062;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = n5936 & n5939;
  assign n5941 = n5932 & n5940;
  assign n5942 = ~n3072 & n5848;
  assign n5943 = n2847 & n5868;
  assign n5944 = n2834 & n5929;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = n2858 & n5868;
  assign n5947 = pi0053 & n4124;
  assign n5948 = n2854 & n5848;
  assign n5949 = n2881 & n5857;
  assign n5950 = n2726 & n5949;
  assign n5951 = ~n5948 & ~n5950;
  assign n5952 = ~n5947 & n5951;
  assign n5953 = ~n5946 & n5952;
  assign n5954 = ~n4133 & n5868;
  assign n5955 = n5953 & ~n5954;
  assign n5956 = n2851 & n5864;
  assign n5957 = n3066 & n5848;
  assign n5958 = ~n5956 & ~n5957;
  assign n5959 = n5955 & n5958;
  assign n5960 = n5945 & n5959;
  assign n5961 = ~n5942 & n5960;
  assign n5962 = n5941 & n5961;
  assign n5963 = n5928 & n5962;
  assign po0211 = ~n5890 | ~n5963;
  assign n5965 = ~n3973 & n4708;
  assign n5966 = pi0054 & n5965;
  assign n5967 = pi0024 & pi0054;
  assign n5968 = pi0054 & n3989;
  assign n5969 = ~n5967 & ~n5968;
  assign n5970 = n2563 & ~n5969;
  assign n5971 = n2795 & n5967;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = pi0054 & n2741;
  assign n5974 = n5972 & ~n5973;
  assign n5975 = ~n5966 & n5974;
  assign n5976 = pi0054 & pi0841;
  assign n5977 = ~n3998 & n5976;
  assign n5978 = n5975 & ~n5977;
  assign n5979 = pi0054 & ~pi0314;
  assign n5980 = pi1044 & n5979;
  assign n5981 = n2619 & n5980;
  assign n5982 = n2591 & n5967;
  assign n5983 = ~n5981 & ~n5982;
  assign n5984 = pi0054 & n4336;
  assign n5985 = pi0054 & n4062;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = n5983 & n5986;
  assign n5988 = ~n3072 & n5967;
  assign n5989 = n2847 & n5976;
  assign n5990 = n2834 & n5980;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = n2858 & n5976;
  assign n5993 = pi0054 & n4124;
  assign n5994 = n2854 & n5967;
  assign n5995 = pi0054 & po0740;
  assign n5996 = n2881 & n5995;
  assign n5997 = n2726 & n5996;
  assign n5998 = ~n5994 & ~n5997;
  assign n5999 = ~n5993 & n5998;
  assign n6000 = ~n5992 & n5999;
  assign n6001 = ~n4133 & n5976;
  assign n6002 = n6000 & ~n6001;
  assign n6003 = n2851 & n5979;
  assign n6004 = n3066 & n5967;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = n6002 & n6005;
  assign n6007 = n5991 & n6006;
  assign n6008 = ~n5988 & n6007;
  assign n6009 = n5987 & n6008;
  assign n6010 = n2910 & n5967;
  assign n6011 = pi0054 & n2726;
  assign n6012 = n4066 & n6011;
  assign n6013 = ~n6010 & ~n6012;
  assign n6014 = n2917 & n5976;
  assign n6015 = n2913 & n5967;
  assign n6016 = ~n6014 & ~n6015;
  assign n6017 = n2936 & n5979;
  assign n6018 = n6016 & ~n6017;
  assign n6019 = n3042 & n5967;
  assign n6020 = pi0054 & n4043;
  assign n6021 = n2930 & n6020;
  assign n6022 = pi0054 & ~n3553;
  assign n6023 = n4497 & n6022;
  assign n6024 = ~n6021 & ~n6023;
  assign n6025 = ~n4402 & n5979;
  assign n6026 = n6024 & ~n6025;
  assign n6027 = pi0054 & n4504;
  assign n6028 = n6026 & ~n6027;
  assign n6029 = ~n6019 & n6028;
  assign n6030 = n6018 & n6029;
  assign n6031 = n3033 & n5967;
  assign n6032 = n6030 & ~n6031;
  assign n6033 = n2651 & n5995;
  assign n6034 = ~n3102 & n6033;
  assign n6035 = pi0054 & n4006;
  assign n6036 = pi0054 & ~n4014;
  assign n6037 = ~pi0054 & pi0841;
  assign n6038 = n2644 & ~n6037;
  assign n6039 = ~n6036 & ~n6038;
  assign n6040 = ~n6035 & n6039;
  assign n6041 = ~n6034 & n6040;
  assign n6042 = n3110 & n5967;
  assign n6043 = n6041 & ~n6042;
  assign n6044 = n6032 & n6043;
  assign n6045 = n6013 & n6044;
  assign n6046 = ~n4105 & n5979;
  assign n6047 = n2569 & n5967;
  assign n6048 = ~n6046 & ~n6047;
  assign n6049 = pi0054 & pi0993;
  assign n6050 = n2576 & n6049;
  assign n6051 = n2598 & n5967;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = n6048 & n6052;
  assign n6054 = n6045 & n6053;
  assign n6055 = n3057 & n5967;
  assign n6056 = pi0054 & ~n3057;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = n4083 & ~n6057;
  assign n6059 = n2901 & n5979;
  assign n6060 = ~n6058 & ~n6059;
  assign n6061 = n2681 & n5967;
  assign n6062 = ~n4077 & n5976;
  assign n6063 = ~n6061 & ~n6062;
  assign n6064 = pi0054 & n4089;
  assign n6065 = pi0054 & n4091;
  assign n6066 = pi0054 & n3128;
  assign n6067 = ~n4094 & n6066;
  assign n6068 = ~n4097 & n5995;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = n3397 & ~n6069;
  assign n6071 = ~n6065 & ~n6070;
  assign n6072 = ~n6064 & n6071;
  assign n6073 = n4087 & ~n6072;
  assign n6074 = n6063 & ~n6073;
  assign n6075 = n6060 & n6074;
  assign n6076 = n6054 & n6075;
  assign n6077 = n6009 & n6076;
  assign po0212 = ~n5978 | ~n6077;
  assign n6079 = pi0024 & pi0055;
  assign n6080 = n2910 & n6079;
  assign n6081 = pi0055 & n2726;
  assign n6082 = n4066 & n6081;
  assign n6083 = ~n6080 & ~n6082;
  assign n6084 = pi0055 & pi0993;
  assign n6085 = n2576 & n6084;
  assign n6086 = n2598 & n6079;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = pi0055 & n4043;
  assign n6089 = n2930 & n6088;
  assign n6090 = pi0055 & ~n3553;
  assign n6091 = n4497 & n6090;
  assign n6092 = ~n6089 & ~n6091;
  assign n6093 = pi0055 & ~pi0314;
  assign n6094 = ~n4402 & n6093;
  assign n6095 = n6092 & ~n6094;
  assign n6096 = pi0055 & pi0841;
  assign n6097 = n2917 & n6096;
  assign n6098 = n2913 & n6079;
  assign n6099 = ~n6097 & ~n6098;
  assign n6100 = n2936 & n6093;
  assign n6101 = n6099 & ~n6100;
  assign n6102 = n3042 & n6079;
  assign n6103 = pi0055 & n4504;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = n6101 & n6104;
  assign n6106 = n6095 & n6105;
  assign n6107 = n3033 & n6079;
  assign n6108 = n6106 & ~n6107;
  assign n6109 = pi0055 & n4006;
  assign n6110 = pi0055 & ~n4014;
  assign n6111 = n3110 & n6079;
  assign n6112 = ~n6110 & ~n6111;
  assign n6113 = pi0055 & po0740;
  assign n6114 = n2651 & n6113;
  assign n6115 = ~n3102 & n6114;
  assign n6116 = n6112 & ~n6115;
  assign n6117 = ~n6109 & n6116;
  assign n6118 = n2591 & n6079;
  assign n6119 = n6117 & ~n6118;
  assign n6120 = n6108 & n6119;
  assign n6121 = n6087 & n6120;
  assign n6122 = n6083 & n6121;
  assign n6123 = pi1044 & n6093;
  assign n6124 = n2619 & n6123;
  assign n6125 = n2644 & n6096;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = pi0055 & n4336;
  assign n6128 = pi0055 & n4062;
  assign n6129 = ~n6127 & ~n6128;
  assign n6130 = n6126 & n6129;
  assign n6131 = ~n3072 & n6079;
  assign n6132 = n2847 & n6096;
  assign n6133 = n2834 & n6123;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = n2881 & n6113;
  assign n6136 = n2726 & n6135;
  assign n6137 = n2858 & n6096;
  assign n6138 = pi0055 & n4124;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = ~n2841 & n6139;
  assign n6141 = n2854 & n6079;
  assign n6142 = n6140 & ~n6141;
  assign n6143 = ~n6136 & n6142;
  assign n6144 = ~n4133 & n6096;
  assign n6145 = n6143 & ~n6144;
  assign n6146 = n2851 & n6093;
  assign n6147 = n3066 & n6079;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = n6145 & n6148;
  assign n6150 = n6134 & n6149;
  assign n6151 = ~n6131 & n6150;
  assign n6152 = n6130 & n6151;
  assign n6153 = ~n4105 & n6093;
  assign n6154 = n2569 & n6079;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = pi0055 & n4708;
  assign n6157 = ~n3973 & n6156;
  assign n6158 = pi0055 & n3989;
  assign n6159 = ~n6079 & ~n6158;
  assign n6160 = n2563 & ~n6159;
  assign n6161 = n2795 & n6079;
  assign n6162 = ~n6160 & ~n6161;
  assign n6163 = pi0055 & n2741;
  assign n6164 = n6162 & ~n6163;
  assign n6165 = ~n6157 & n6164;
  assign n6166 = ~n3998 & n6096;
  assign n6167 = n6165 & ~n6166;
  assign n6168 = n6155 & n6167;
  assign n6169 = n3057 & n6079;
  assign n6170 = pi0055 & ~n3057;
  assign n6171 = ~n6169 & ~n6170;
  assign n6172 = n4083 & ~n6171;
  assign n6173 = n2901 & n6093;
  assign n6174 = ~n6172 & ~n6173;
  assign n6175 = n2681 & n6079;
  assign n6176 = ~n4077 & n6096;
  assign n6177 = ~n6175 & ~n6176;
  assign n6178 = pi0055 & n4089;
  assign n6179 = pi0055 & n4091;
  assign n6180 = pi0055 & n3128;
  assign n6181 = ~n4094 & n6180;
  assign n6182 = ~n4097 & n6113;
  assign n6183 = ~n6181 & ~n6182;
  assign n6184 = n3397 & ~n6183;
  assign n6185 = ~n6179 & ~n6184;
  assign n6186 = ~n6178 & n6185;
  assign n6187 = n4087 & ~n6186;
  assign n6188 = n6177 & ~n6187;
  assign n6189 = n6174 & n6188;
  assign n6190 = n6168 & n6189;
  assign n6191 = n6152 & n6190;
  assign po0213 = ~n6122 | ~n6191;
  assign n6193 = pi0056 & ~pi0314;
  assign n6194 = pi1044 & n6193;
  assign n6195 = n2619 & n6194;
  assign n6196 = pi0056 & pi0841;
  assign n6197 = n2644 & n6196;
  assign n6198 = ~n6195 & ~n6197;
  assign n6199 = pi0056 & pi0993;
  assign n6200 = n2576 & n6199;
  assign n6201 = pi0024 & pi0056;
  assign n6202 = n2598 & n6201;
  assign n6203 = ~n6200 & ~n6202;
  assign n6204 = pi0056 & n4336;
  assign n6205 = pi0056 & n4062;
  assign n6206 = ~n6204 & ~n6205;
  assign n6207 = n6203 & n6206;
  assign n6208 = n6198 & n6207;
  assign n6209 = n3057 & n6201;
  assign n6210 = pi0056 & ~n3057;
  assign n6211 = ~n6209 & ~n6210;
  assign n6212 = n4083 & ~n6211;
  assign n6213 = n2901 & n6193;
  assign n6214 = ~n6212 & ~n6213;
  assign n6215 = n2681 & n6201;
  assign n6216 = ~n4077 & n6196;
  assign n6217 = ~n6215 & ~n6216;
  assign n6218 = pi0056 & n4089;
  assign n6219 = pi0056 & n4091;
  assign n6220 = pi0056 & n3128;
  assign n6221 = ~n4094 & n6220;
  assign n6222 = pi0056 & po0740;
  assign n6223 = ~n4097 & n6222;
  assign n6224 = ~n6221 & ~n6223;
  assign n6225 = n3397 & ~n6224;
  assign n6226 = ~n6219 & ~n6225;
  assign n6227 = ~n6218 & n6226;
  assign n6228 = n4087 & ~n6227;
  assign n6229 = n6217 & ~n6228;
  assign n6230 = n6214 & n6229;
  assign n6231 = n2917 & n6196;
  assign n6232 = n2913 & n6201;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = n2936 & n6193;
  assign n6235 = n6233 & ~n6234;
  assign n6236 = pi0056 & n4043;
  assign n6237 = n2930 & n6236;
  assign n6238 = pi0056 & ~n3553;
  assign n6239 = n4497 & n6238;
  assign n6240 = ~n6237 & ~n6239;
  assign n6241 = ~n4402 & n6193;
  assign n6242 = n6240 & ~n6241;
  assign n6243 = n3042 & n6201;
  assign n6244 = pi0056 & n4504;
  assign n6245 = ~n6243 & ~n6244;
  assign n6246 = n6242 & n6245;
  assign n6247 = n6235 & n6246;
  assign n6248 = n3033 & n6201;
  assign n6249 = n6247 & ~n6248;
  assign n6250 = n2651 & n6222;
  assign n6251 = ~n3102 & n6250;
  assign n6252 = pi0056 & n4006;
  assign n6253 = pi0056 & ~n4014;
  assign n6254 = pi0024 & ~pi0056;
  assign n6255 = n2591 & ~n6254;
  assign n6256 = ~n6253 & ~n6255;
  assign n6257 = ~n6252 & n6256;
  assign n6258 = ~n6251 & n6257;
  assign n6259 = n3110 & n6201;
  assign n6260 = n6258 & ~n6259;
  assign n6261 = n2910 & n6201;
  assign n6262 = pi0056 & n2726;
  assign n6263 = n4066 & n6262;
  assign n6264 = ~n6261 & ~n6263;
  assign n6265 = n6260 & n6264;
  assign n6266 = n6249 & n6265;
  assign n6267 = ~n3072 & n6201;
  assign n6268 = n2847 & n6196;
  assign n6269 = n2834 & n6194;
  assign n6270 = ~n6268 & ~n6269;
  assign n6271 = n2858 & n6196;
  assign n6272 = pi0056 & n4124;
  assign n6273 = n2854 & n6201;
  assign n6274 = n2881 & n6222;
  assign n6275 = n2726 & n6274;
  assign n6276 = ~n6273 & ~n6275;
  assign n6277 = ~n6272 & n6276;
  assign n6278 = ~n6271 & n6277;
  assign n6279 = ~n4133 & n6196;
  assign n6280 = n6278 & ~n6279;
  assign n6281 = n2851 & n6193;
  assign n6282 = n3066 & n6201;
  assign n6283 = ~n6281 & ~n6282;
  assign n6284 = n6280 & n6283;
  assign n6285 = n6270 & n6284;
  assign n6286 = ~n6267 & n6285;
  assign n6287 = n6266 & n6286;
  assign n6288 = pi0056 & n4708;
  assign n6289 = ~n3973 & n6288;
  assign n6290 = pi0056 & n3989;
  assign n6291 = ~n6201 & ~n6290;
  assign n6292 = n2563 & ~n6291;
  assign n6293 = n2795 & n6201;
  assign n6294 = ~n6292 & ~n6293;
  assign n6295 = pi0056 & n2741;
  assign n6296 = n6294 & ~n6295;
  assign n6297 = ~n6289 & n6296;
  assign n6298 = ~n3998 & n6196;
  assign n6299 = n6297 & ~n6298;
  assign n6300 = ~n4105 & n6193;
  assign n6301 = n2569 & n6201;
  assign n6302 = ~n6300 & ~n6301;
  assign n6303 = n6299 & n6302;
  assign n6304 = n6287 & n6303;
  assign n6305 = n6230 & n6304;
  assign po0214 = ~n6208 | ~n6305;
  assign n6307 = pi0057 & ~pi0314;
  assign n6308 = ~n4105 & n6307;
  assign n6309 = pi0024 & pi0057;
  assign n6310 = n2569 & n6309;
  assign n6311 = ~n6308 & ~n6310;
  assign n6312 = pi0057 & pi0993;
  assign n6313 = n2576 & n6312;
  assign n6314 = n2598 & n6309;
  assign n6315 = ~n6313 & ~n6314;
  assign n6316 = n6311 & n6315;
  assign n6317 = n3057 & n6309;
  assign n6318 = pi0057 & ~n3057;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = n4083 & ~n6319;
  assign n6321 = n2901 & n6307;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = n2681 & n6309;
  assign n6324 = pi0057 & pi0841;
  assign n6325 = ~n4077 & n6324;
  assign n6326 = ~n6323 & ~n6325;
  assign n6327 = pi0057 & n4089;
  assign n6328 = pi0057 & n4091;
  assign n6329 = pi0057 & n3128;
  assign n6330 = ~n4094 & n6329;
  assign n6331 = pi0057 & po0740;
  assign n6332 = ~n4097 & n6331;
  assign n6333 = ~n6330 & ~n6332;
  assign n6334 = n3397 & ~n6333;
  assign n6335 = ~n6328 & ~n6334;
  assign n6336 = ~n6327 & n6335;
  assign n6337 = n4087 & ~n6336;
  assign n6338 = n6326 & ~n6337;
  assign n6339 = n6322 & n6338;
  assign n6340 = ~n3072 & n6309;
  assign n6341 = n2847 & n6324;
  assign n6342 = pi1044 & n6307;
  assign n6343 = n2834 & n6342;
  assign n6344 = ~n6341 & ~n6343;
  assign n6345 = n2858 & n6324;
  assign n6346 = pi0057 & n4124;
  assign n6347 = n2854 & n6309;
  assign n6348 = n2881 & n6331;
  assign n6349 = n2726 & n6348;
  assign n6350 = ~n6347 & ~n6349;
  assign n6351 = ~n6346 & n6350;
  assign n6352 = ~n6345 & n6351;
  assign n6353 = ~n4133 & n6324;
  assign n6354 = n6352 & ~n6353;
  assign n6355 = n2851 & n6307;
  assign n6356 = n3066 & n6309;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = n6354 & n6357;
  assign n6359 = n6344 & n6358;
  assign n6360 = ~n6340 & n6359;
  assign n6361 = n6339 & n6360;
  assign n6362 = pi0057 & n4006;
  assign n6363 = pi0057 & ~n4014;
  assign n6364 = n3110 & n6309;
  assign n6365 = ~n6363 & ~n6364;
  assign n6366 = n2651 & n6331;
  assign n6367 = ~n3102 & n6366;
  assign n6368 = n6365 & ~n6367;
  assign n6369 = ~n6362 & n6368;
  assign n6370 = n2591 & n6309;
  assign n6371 = n6369 & ~n6370;
  assign n6372 = n2619 & n6342;
  assign n6373 = n2644 & n6324;
  assign n6374 = ~n6372 & ~n6373;
  assign n6375 = pi0057 & n4043;
  assign n6376 = n2930 & n6375;
  assign n6377 = pi0057 & ~n3553;
  assign n6378 = n4497 & n6377;
  assign n6379 = ~n6376 & ~n6378;
  assign n6380 = n2913 & n6309;
  assign n6381 = n6379 & ~n6380;
  assign n6382 = n2936 & n6307;
  assign n6383 = n2544 & n6307;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = n2533 & n6307;
  assign n6386 = ~pi0841 & ~pi0924;
  assign n6387 = ~n6324 & ~n6386;
  assign n6388 = n2917 & ~n6387;
  assign n6389 = n3042 & n6309;
  assign n6390 = pi0057 & ~pi1076;
  assign n6391 = n2926 & n6390;
  assign n6392 = ~n6389 & ~n6391;
  assign n6393 = ~n6388 & n6392;
  assign n6394 = ~n6385 & n6393;
  assign n6395 = n6384 & n6394;
  assign n6396 = n6381 & n6395;
  assign n6397 = n3033 & n6309;
  assign n6398 = n6396 & ~n6397;
  assign n6399 = n2910 & n6309;
  assign n6400 = pi0057 & n2726;
  assign n6401 = n4066 & n6400;
  assign n6402 = ~n6399 & ~n6401;
  assign n6403 = n6398 & n6402;
  assign n6404 = n6374 & n6403;
  assign n6405 = n6371 & n6404;
  assign n6406 = pi0057 & n4336;
  assign n6407 = pi0057 & n2741;
  assign n6408 = pi0057 & n4708;
  assign n6409 = ~n3973 & n6408;
  assign n6410 = ~n2698 & ~n2747;
  assign n6411 = n6324 & ~n6410;
  assign n6412 = n2795 & n6309;
  assign n6413 = ~n6411 & ~n6412;
  assign n6414 = pi0057 & n3989;
  assign n6415 = ~n6309 & ~n6414;
  assign n6416 = n2563 & ~n6415;
  assign n6417 = ~pi0057 & pi0841;
  assign n6418 = n2583 & ~n6417;
  assign n6419 = ~n6416 & ~n6418;
  assign n6420 = n6413 & n6419;
  assign n6421 = ~n6409 & n6420;
  assign n6422 = ~n6407 & n6421;
  assign n6423 = pi0057 & ~n4061;
  assign n6424 = n4060 & n6423;
  assign n6425 = n6422 & ~n6424;
  assign n6426 = ~n6406 & n6425;
  assign n6427 = n6405 & n6426;
  assign n6428 = n6361 & n6427;
  assign po0215 = ~n6316 | ~n6428;
  assign n6430 = pi0058 & po0740;
  assign n6431 = n2651 & n6430;
  assign n6432 = ~n3102 & n6431;
  assign n6433 = pi0058 & n4006;
  assign n6434 = ~n6432 & ~n6433;
  assign n6435 = pi0058 & ~n4014;
  assign n6436 = pi0024 & pi0058;
  assign n6437 = n3110 & n6436;
  assign n6438 = ~n6435 & ~n6437;
  assign n6439 = n6434 & n6438;
  assign n6440 = pi0058 & ~n4061;
  assign n6441 = n4060 & n6440;
  assign n6442 = n6439 & ~n6441;
  assign n6443 = pi0058 & n4067;
  assign n6444 = n2591 & n6436;
  assign n6445 = ~n6443 & ~n6444;
  assign n6446 = pi0058 & ~pi0314;
  assign n6447 = pi1044 & n6446;
  assign n6448 = n2619 & n6447;
  assign n6449 = pi0058 & pi0841;
  assign n6450 = n2644 & n6449;
  assign n6451 = ~n6448 & ~n6450;
  assign n6452 = n2910 & n6436;
  assign n6453 = n6451 & ~n6452;
  assign n6454 = n6445 & n6453;
  assign n6455 = ~n3558 & n6454;
  assign n6456 = n2847 & n6449;
  assign n6457 = n2834 & n6447;
  assign n6458 = ~n6456 & ~n6457;
  assign n6459 = n2858 & n6449;
  assign n6460 = pi0058 & n4124;
  assign n6461 = n2854 & n6436;
  assign n6462 = n2881 & n6430;
  assign n6463 = n2726 & n6462;
  assign n6464 = ~n6461 & ~n6463;
  assign n6465 = ~n6460 & n6464;
  assign n6466 = ~n6459 & n6465;
  assign n6467 = n2851 & n6446;
  assign n6468 = n6466 & ~n6467;
  assign n6469 = ~n3072 & n6436;
  assign n6470 = n6468 & ~n6469;
  assign n6471 = n6458 & n6470;
  assign n6472 = pi0058 & n2823;
  assign n6473 = n6471 & ~n6472;
  assign n6474 = ~n4132 & n6449;
  assign n6475 = n3066 & n6436;
  assign n6476 = ~n6474 & ~n6475;
  assign n6477 = n6473 & n6476;
  assign n6478 = n6455 & n6477;
  assign n6479 = pi0058 & n2741;
  assign n6480 = pi0058 & n4523;
  assign n6481 = ~n3973 & n6480;
  assign n6482 = ~n3998 & n6449;
  assign n6483 = pi0058 & n3989;
  assign n6484 = ~n6436 & ~n6483;
  assign n6485 = n2563 & ~n6484;
  assign n6486 = n2795 & n6436;
  assign n6487 = ~n6485 & ~n6486;
  assign n6488 = ~n6482 & n6487;
  assign n6489 = ~n6481 & n6488;
  assign n6490 = ~n6479 & n6489;
  assign n6491 = n2917 & n6449;
  assign n6492 = n2913 & n6436;
  assign n6493 = ~n6491 & ~n6492;
  assign n6494 = n2936 & n6446;
  assign n6495 = n6493 & ~n6494;
  assign n6496 = pi0058 & n4043;
  assign n6497 = n2930 & n6496;
  assign n6498 = pi0058 & ~n3553;
  assign n6499 = n4497 & n6498;
  assign n6500 = ~n6497 & ~n6499;
  assign n6501 = ~n4402 & n6446;
  assign n6502 = n6500 & ~n6501;
  assign n6503 = n3042 & n6436;
  assign n6504 = pi0058 & n4504;
  assign n6505 = ~n6503 & ~n6504;
  assign n6506 = n6502 & n6505;
  assign n6507 = n6495 & n6506;
  assign n6508 = n3033 & n6436;
  assign n6509 = n6507 & ~n6508;
  assign n6510 = n6490 & n6509;
  assign n6511 = pi0058 & n4336;
  assign n6512 = n6510 & ~n6511;
  assign n6513 = n6478 & n6512;
  assign n6514 = n6442 & n6513;
  assign n6515 = n2681 & n6436;
  assign n6516 = ~n4077 & n6449;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = n2901 & n6446;
  assign n6519 = n3057 & n6436;
  assign n6520 = pi0058 & ~n3057;
  assign n6521 = ~n6519 & ~n6520;
  assign n6522 = n4083 & ~n6521;
  assign n6523 = ~n6518 & ~n6522;
  assign n6524 = pi0058 & n4089;
  assign n6525 = pi0058 & n4091;
  assign n6526 = pi0058 & n3128;
  assign n6527 = ~n4094 & n6526;
  assign n6528 = ~n4097 & n6430;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = n3397 & ~n6529;
  assign n6531 = ~n6525 & ~n6530;
  assign n6532 = ~n6524 & n6531;
  assign n6533 = n4087 & ~n6532;
  assign n6534 = n6523 & ~n6533;
  assign n6535 = ~n4105 & n6446;
  assign n6536 = n2569 & n6436;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = pi0058 & pi0993;
  assign n6539 = n2576 & n6538;
  assign n6540 = n2598 & n6436;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = n6537 & n6541;
  assign n6543 = n6534 & n6542;
  assign n6544 = n6517 & n6543;
  assign po0216 = ~n6514 | ~n6544;
  assign n6546 = pi0059 & n4043;
  assign n6547 = n2930 & n6546;
  assign n6548 = pi0059 & ~n3553;
  assign n6549 = n4497 & n6548;
  assign n6550 = ~n6547 & ~n6549;
  assign n6551 = pi0059 & ~pi0314;
  assign n6552 = n2533 & n6551;
  assign n6553 = n6550 & ~n6552;
  assign n6554 = pi0059 & pi0841;
  assign n6555 = ~pi0841 & pi0924;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = n2917 & ~n6556;
  assign n6558 = pi0059 & ~pi1076;
  assign n6559 = n2926 & n6558;
  assign n6560 = pi0024 & pi0059;
  assign n6561 = n3042 & n6560;
  assign n6562 = ~n6559 & ~n6561;
  assign n6563 = n2936 & n6551;
  assign n6564 = n2913 & n6560;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = n2544 & n6551;
  assign n6567 = n6565 & ~n6566;
  assign n6568 = n6562 & n6567;
  assign n6569 = ~n6557 & n6568;
  assign n6570 = n6553 & n6569;
  assign n6571 = n3033 & n6560;
  assign n6572 = n6570 & ~n6571;
  assign n6573 = pi0059 & n4006;
  assign n6574 = pi0059 & ~n4014;
  assign n6575 = n3110 & n6560;
  assign n6576 = ~n6574 & ~n6575;
  assign n6577 = pi0059 & po0740;
  assign n6578 = n2651 & n6577;
  assign n6579 = ~n3102 & n6578;
  assign n6580 = n6576 & ~n6579;
  assign n6581 = ~n6573 & n6580;
  assign n6582 = n2591 & n6560;
  assign n6583 = n6581 & ~n6582;
  assign n6584 = n2910 & n6560;
  assign n6585 = pi0059 & n2726;
  assign n6586 = n4066 & n6585;
  assign n6587 = ~n6584 & ~n6586;
  assign n6588 = n6583 & n6587;
  assign n6589 = n6572 & n6588;
  assign n6590 = ~n3072 & n6560;
  assign n6591 = n2847 & n6554;
  assign n6592 = pi1044 & n6551;
  assign n6593 = n2834 & n6592;
  assign n6594 = ~n6591 & ~n6593;
  assign n6595 = n2858 & n6554;
  assign n6596 = pi0059 & n4124;
  assign n6597 = n2854 & n6560;
  assign n6598 = n2881 & n6577;
  assign n6599 = n2726 & n6598;
  assign n6600 = ~n6597 & ~n6599;
  assign n6601 = ~n6596 & n6600;
  assign n6602 = ~n6595 & n6601;
  assign n6603 = ~n4133 & n6554;
  assign n6604 = n6602 & ~n6603;
  assign n6605 = n2851 & n6551;
  assign n6606 = n3066 & n6560;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6604 & n6607;
  assign n6609 = n6594 & n6608;
  assign n6610 = ~n6590 & n6609;
  assign n6611 = n6589 & n6610;
  assign n6612 = pi0059 & pi0993;
  assign n6613 = n2576 & n6612;
  assign n6614 = n2598 & n6560;
  assign n6615 = ~n6613 & ~n6614;
  assign n6616 = pi0059 & n4062;
  assign n6617 = n2619 & n6592;
  assign n6618 = n2644 & n6554;
  assign n6619 = ~n6617 & ~n6618;
  assign n6620 = ~n6616 & n6619;
  assign n6621 = pi0059 & n4336;
  assign n6622 = n6620 & ~n6621;
  assign n6623 = n6615 & n6622;
  assign n6624 = n3057 & n6560;
  assign n6625 = pi0059 & ~n3057;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = n4083 & ~n6626;
  assign n6628 = n2901 & n6551;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = n2681 & n6560;
  assign n6631 = ~n4077 & n6554;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = pi0059 & n4089;
  assign n6634 = pi0059 & n4091;
  assign n6635 = pi0059 & n3128;
  assign n6636 = ~n4094 & n6635;
  assign n6637 = ~n4097 & n6577;
  assign n6638 = ~n6636 & ~n6637;
  assign n6639 = n3397 & ~n6638;
  assign n6640 = ~n6634 & ~n6639;
  assign n6641 = ~n6633 & n6640;
  assign n6642 = n4087 & ~n6641;
  assign n6643 = n6632 & ~n6642;
  assign n6644 = n6629 & n6643;
  assign n6645 = n6623 & n6644;
  assign n6646 = ~n4105 & n6551;
  assign n6647 = n2569 & n6560;
  assign n6648 = ~n6646 & ~n6647;
  assign n6649 = pi0059 & n4708;
  assign n6650 = ~n3973 & n6649;
  assign n6651 = pi0059 & n3989;
  assign n6652 = ~n6560 & ~n6651;
  assign n6653 = n2563 & ~n6652;
  assign n6654 = n2795 & n6560;
  assign n6655 = ~n6653 & ~n6654;
  assign n6656 = pi0059 & n2741;
  assign n6657 = n6655 & ~n6656;
  assign n6658 = ~n6650 & n6657;
  assign n6659 = ~n3998 & n6554;
  assign n6660 = n6658 & ~n6659;
  assign n6661 = n6648 & n6660;
  assign n6662 = n6645 & n6661;
  assign po0217 = ~n6611 | ~n6662;
  assign n6664 = pi0060 & pi0841;
  assign n6665 = n2917 & n6664;
  assign n6666 = pi0024 & pi0060;
  assign n6667 = n2913 & n6666;
  assign n6668 = ~n6665 & ~n6667;
  assign n6669 = pi0060 & ~pi0314;
  assign n6670 = n2936 & n6669;
  assign n6671 = n6668 & ~n6670;
  assign n6672 = pi0060 & n4043;
  assign n6673 = n2930 & n6672;
  assign n6674 = pi0060 & ~n3553;
  assign n6675 = n4497 & n6674;
  assign n6676 = ~n6673 & ~n6675;
  assign n6677 = ~n4402 & n6669;
  assign n6678 = n6676 & ~n6677;
  assign n6679 = n3042 & n6666;
  assign n6680 = pi0060 & n4504;
  assign n6681 = ~n6679 & ~n6680;
  assign n6682 = n6678 & n6681;
  assign n6683 = n6671 & n6682;
  assign n6684 = n3033 & n6666;
  assign n6685 = n6683 & ~n6684;
  assign n6686 = pi0060 & n4006;
  assign n6687 = pi0060 & ~n4014;
  assign n6688 = n3110 & n6666;
  assign n6689 = ~n6687 & ~n6688;
  assign n6690 = pi0060 & po0740;
  assign n6691 = n2651 & n6690;
  assign n6692 = ~n3102 & n6691;
  assign n6693 = n6689 & ~n6692;
  assign n6694 = ~n6686 & n6693;
  assign n6695 = n2591 & n6666;
  assign n6696 = n6694 & ~n6695;
  assign n6697 = n2910 & n6666;
  assign n6698 = pi0060 & n2726;
  assign n6699 = n4066 & n6698;
  assign n6700 = ~n6697 & ~n6699;
  assign n6701 = n6696 & n6700;
  assign n6702 = n6685 & n6701;
  assign n6703 = ~n3072 & n6666;
  assign n6704 = n2847 & n6664;
  assign n6705 = pi1044 & n6669;
  assign n6706 = n2834 & n6705;
  assign n6707 = ~n6704 & ~n6706;
  assign n6708 = n2858 & n6664;
  assign n6709 = pi0060 & n4124;
  assign n6710 = n2854 & n6666;
  assign n6711 = n2881 & n6690;
  assign n6712 = n2726 & n6711;
  assign n6713 = ~n6710 & ~n6712;
  assign n6714 = ~n6709 & n6713;
  assign n6715 = ~n6708 & n6714;
  assign n6716 = ~n4133 & n6664;
  assign n6717 = n6715 & ~n6716;
  assign n6718 = n2851 & n6669;
  assign n6719 = n3066 & n6666;
  assign n6720 = ~n6718 & ~n6719;
  assign n6721 = n6717 & n6720;
  assign n6722 = n6707 & n6721;
  assign n6723 = ~n6703 & n6722;
  assign n6724 = n6702 & n6723;
  assign n6725 = pi0060 & pi0993;
  assign n6726 = n2576 & n6725;
  assign n6727 = n2598 & n6666;
  assign n6728 = ~n6726 & ~n6727;
  assign n6729 = pi0060 & n4062;
  assign n6730 = n2619 & n6705;
  assign n6731 = n2644 & n6664;
  assign n6732 = ~n6730 & ~n6731;
  assign n6733 = ~n6729 & n6732;
  assign n6734 = pi0060 & n4336;
  assign n6735 = n6733 & ~n6734;
  assign n6736 = n6728 & n6735;
  assign n6737 = n3397 & ~n3403;
  assign n6738 = ~n4097 & n6690;
  assign n6739 = pi0060 & n4459;
  assign n6740 = ~n6738 & ~n6739;
  assign n6741 = n6737 & ~n6740;
  assign n6742 = ~n3403 & ~n5901;
  assign n6743 = pi0060 & n6742;
  assign n6744 = ~n6741 & ~n6743;
  assign n6745 = ~n3403 & n3405;
  assign n6746 = n6744 & ~n6745;
  assign n6747 = n2777 & ~n6746;
  assign n6748 = n3464 & n6747;
  assign n6749 = n2681 & n6666;
  assign n6750 = ~n4077 & n6664;
  assign n6751 = ~n6749 & ~n6750;
  assign n6752 = n3057 & n6666;
  assign n6753 = pi0060 & ~n3057;
  assign n6754 = ~n6752 & ~n6753;
  assign n6755 = n4083 & ~n6754;
  assign n6756 = n2901 & n6669;
  assign n6757 = ~n6755 & ~n6756;
  assign n6758 = n6751 & n6757;
  assign n6759 = ~n6748 & n6758;
  assign n6760 = n6736 & n6759;
  assign n6761 = ~n4105 & n6669;
  assign n6762 = n2569 & n6666;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = pi0060 & n4708;
  assign n6765 = ~n3973 & n6764;
  assign n6766 = pi0060 & n3989;
  assign n6767 = ~n6666 & ~n6766;
  assign n6768 = n2563 & ~n6767;
  assign n6769 = n2795 & n6666;
  assign n6770 = ~n6768 & ~n6769;
  assign n6771 = pi0060 & n2741;
  assign n6772 = n6770 & ~n6771;
  assign n6773 = ~n6765 & n6772;
  assign n6774 = ~n3998 & n6664;
  assign n6775 = n6773 & ~n6774;
  assign n6776 = n6763 & n6775;
  assign n6777 = n6760 & n6776;
  assign po0218 = ~n6724 | ~n6777;
  assign n6779 = pi0061 & pi0993;
  assign n6780 = n2576 & n6779;
  assign n6781 = pi0024 & pi0061;
  assign n6782 = n2598 & n6781;
  assign n6783 = ~n6780 & ~n6782;
  assign n6784 = pi0061 & n4067;
  assign n6785 = n3033 & n6781;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = n3042 & n6781;
  assign n6788 = n6786 & ~n6787;
  assign n6789 = pi0024 & ~pi0061;
  assign n6790 = n2910 & ~n6789;
  assign n6791 = pi0061 & ~pi0314;
  assign n6792 = n2936 & n6791;
  assign n6793 = n2913 & n6781;
  assign n6794 = pi0061 & pi0841;
  assign n6795 = n2917 & n6794;
  assign n6796 = ~n6793 & ~n6795;
  assign n6797 = pi0061 & n4504;
  assign n6798 = pi0061 & n4043;
  assign n6799 = n2930 & n6798;
  assign n6800 = pi0061 & ~n3553;
  assign n6801 = n4497 & n6800;
  assign n6802 = ~n6799 & ~n6801;
  assign n6803 = ~n4402 & n6791;
  assign n6804 = n6802 & ~n6803;
  assign n6805 = ~n6797 & n6804;
  assign n6806 = n6796 & n6805;
  assign n6807 = ~n6792 & n6806;
  assign n6808 = ~n6790 & n6807;
  assign n6809 = pi0061 & n4006;
  assign n6810 = pi0061 & ~n4014;
  assign n6811 = n3110 & n6781;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = pi0061 & po0740;
  assign n6814 = n2651 & n6813;
  assign n6815 = ~n3102 & n6814;
  assign n6816 = n6812 & ~n6815;
  assign n6817 = ~n6809 & n6816;
  assign n6818 = n2591 & n6781;
  assign n6819 = n6817 & ~n6818;
  assign n6820 = n6808 & n6819;
  assign n6821 = n6788 & n6820;
  assign n6822 = n6783 & n6821;
  assign n6823 = pi1044 & n6791;
  assign n6824 = n2619 & n6823;
  assign n6825 = n2644 & n6794;
  assign n6826 = ~n6824 & ~n6825;
  assign n6827 = pi0061 & n4336;
  assign n6828 = pi0061 & n4062;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = n6826 & n6829;
  assign n6831 = ~n3072 & n6781;
  assign n6832 = n2847 & n6794;
  assign n6833 = n2834 & n6823;
  assign n6834 = ~n6832 & ~n6833;
  assign n6835 = n2858 & n6794;
  assign n6836 = pi0061 & n4124;
  assign n6837 = n2854 & n6781;
  assign n6838 = n2881 & n6813;
  assign n6839 = n2726 & n6838;
  assign n6840 = ~n6837 & ~n6839;
  assign n6841 = ~n6836 & n6840;
  assign n6842 = ~n6835 & n6841;
  assign n6843 = ~n4133 & n6794;
  assign n6844 = n6842 & ~n6843;
  assign n6845 = n2851 & n6791;
  assign n6846 = n3066 & n6781;
  assign n6847 = ~n6845 & ~n6846;
  assign n6848 = n6844 & n6847;
  assign n6849 = n6834 & n6848;
  assign n6850 = ~n6831 & n6849;
  assign n6851 = n6830 & n6850;
  assign n6852 = ~n4105 & n6791;
  assign n6853 = n2569 & n6781;
  assign n6854 = ~n6852 & ~n6853;
  assign n6855 = pi0061 & n4708;
  assign n6856 = ~n3973 & n6855;
  assign n6857 = pi0061 & n3989;
  assign n6858 = ~n6781 & ~n6857;
  assign n6859 = n2563 & ~n6858;
  assign n6860 = n2795 & n6781;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = pi0061 & n2741;
  assign n6863 = n6861 & ~n6862;
  assign n6864 = ~n6856 & n6863;
  assign n6865 = ~n3998 & n6794;
  assign n6866 = n6864 & ~n6865;
  assign n6867 = n6854 & n6866;
  assign n6868 = n3057 & n6781;
  assign n6869 = pi0061 & ~n3057;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = n4083 & ~n6870;
  assign n6872 = n2901 & n6791;
  assign n6873 = ~n6871 & ~n6872;
  assign n6874 = n2681 & n6781;
  assign n6875 = ~n4077 & n6794;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = pi0061 & n4089;
  assign n6878 = pi0061 & n4091;
  assign n6879 = pi0061 & n3128;
  assign n6880 = ~n4094 & n6879;
  assign n6881 = ~n4097 & n6813;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = n3397 & ~n6882;
  assign n6884 = ~n6878 & ~n6883;
  assign n6885 = ~n6877 & n6884;
  assign n6886 = n4087 & ~n6885;
  assign n6887 = n6876 & ~n6886;
  assign n6888 = n6873 & n6887;
  assign n6889 = n6867 & n6888;
  assign n6890 = n6851 & n6889;
  assign po0219 = ~n6822 | ~n6890;
  assign n6892 = ~pi0024 & n3033;
  assign n6893 = pi0062 & pi0993;
  assign n6894 = n2576 & n6893;
  assign n6895 = pi0024 & pi0062;
  assign n6896 = n2598 & n6895;
  assign n6897 = ~n6894 & ~n6896;
  assign n6898 = pi0062 & n4336;
  assign n6899 = pi0062 & n4062;
  assign n6900 = ~n6898 & ~n6899;
  assign n6901 = n6897 & n6900;
  assign n6902 = ~n6892 & n6901;
  assign n6903 = pi0062 & n4067;
  assign n6904 = n2910 & n6895;
  assign n6905 = ~n6903 & ~n6904;
  assign n6906 = n3042 & n6895;
  assign n6907 = n6905 & ~n6906;
  assign n6908 = pi0062 & n4006;
  assign n6909 = pi0062 & ~n4014;
  assign n6910 = n3110 & n6895;
  assign n6911 = ~n6909 & ~n6910;
  assign n6912 = pi0062 & po0740;
  assign n6913 = n2651 & n6912;
  assign n6914 = ~n3102 & n6913;
  assign n6915 = n6911 & ~n6914;
  assign n6916 = ~n6908 & n6915;
  assign n6917 = n2591 & n6895;
  assign n6918 = n6916 & ~n6917;
  assign n6919 = pi0062 & ~pi0314;
  assign n6920 = pi1044 & n6919;
  assign n6921 = n2619 & n6920;
  assign n6922 = pi0062 & pi0841;
  assign n6923 = n2644 & n6922;
  assign n6924 = ~n6921 & ~n6923;
  assign n6925 = n6918 & n6924;
  assign n6926 = n2936 & n6919;
  assign n6927 = n2913 & n6895;
  assign n6928 = n2917 & n6922;
  assign n6929 = ~n6927 & ~n6928;
  assign n6930 = pi0062 & n4504;
  assign n6931 = pi0062 & n4043;
  assign n6932 = n2930 & n6931;
  assign n6933 = pi0062 & ~n3553;
  assign n6934 = n4497 & n6933;
  assign n6935 = ~n6932 & ~n6934;
  assign n6936 = ~n4402 & n6919;
  assign n6937 = n6935 & ~n6936;
  assign n6938 = ~n6930 & n6937;
  assign n6939 = n6929 & n6938;
  assign n6940 = ~n6926 & n6939;
  assign n6941 = pi0062 & n3033;
  assign n6942 = n6940 & ~n6941;
  assign n6943 = n6925 & n6942;
  assign n6944 = n6907 & n6943;
  assign n6945 = ~n3072 & n6895;
  assign n6946 = n2847 & n6922;
  assign n6947 = n2834 & n6920;
  assign n6948 = ~n6946 & ~n6947;
  assign n6949 = n2858 & n6922;
  assign n6950 = pi0062 & n4124;
  assign n6951 = n2854 & n6895;
  assign n6952 = n2881 & n6912;
  assign n6953 = n2726 & n6952;
  assign n6954 = ~n6951 & ~n6953;
  assign n6955 = ~n6950 & n6954;
  assign n6956 = ~n6949 & n6955;
  assign n6957 = ~n4133 & n6922;
  assign n6958 = n6956 & ~n6957;
  assign n6959 = n2851 & n6919;
  assign n6960 = n3066 & n6895;
  assign n6961 = ~n6959 & ~n6960;
  assign n6962 = n6958 & n6961;
  assign n6963 = n6948 & n6962;
  assign n6964 = ~n6945 & n6963;
  assign n6965 = n6944 & n6964;
  assign n6966 = ~n4105 & n6919;
  assign n6967 = n2569 & n6895;
  assign n6968 = ~n6966 & ~n6967;
  assign n6969 = pi0062 & n4708;
  assign n6970 = ~n3973 & n6969;
  assign n6971 = pi0062 & n3989;
  assign n6972 = ~n6895 & ~n6971;
  assign n6973 = n2563 & ~n6972;
  assign n6974 = n2795 & n6895;
  assign n6975 = ~n6973 & ~n6974;
  assign n6976 = pi0062 & n2741;
  assign n6977 = n6975 & ~n6976;
  assign n6978 = ~n6970 & n6977;
  assign n6979 = ~n3998 & n6922;
  assign n6980 = n6978 & ~n6979;
  assign n6981 = n6968 & n6980;
  assign n6982 = n3057 & n6895;
  assign n6983 = pi0062 & ~n3057;
  assign n6984 = ~n6982 & ~n6983;
  assign n6985 = n4083 & ~n6984;
  assign n6986 = n2901 & n6919;
  assign n6987 = ~n6985 & ~n6986;
  assign n6988 = n2681 & n6895;
  assign n6989 = ~n4077 & n6922;
  assign n6990 = ~n6988 & ~n6989;
  assign n6991 = pi0062 & n4089;
  assign n6992 = pi0062 & n4091;
  assign n6993 = pi0062 & n3128;
  assign n6994 = ~n4094 & n6993;
  assign n6995 = ~n4097 & n6912;
  assign n6996 = ~n6994 & ~n6995;
  assign n6997 = n3397 & ~n6996;
  assign n6998 = ~n6992 & ~n6997;
  assign n6999 = ~n6991 & n6998;
  assign n7000 = n4087 & ~n6999;
  assign n7001 = n6990 & ~n7000;
  assign n7002 = n6987 & n7001;
  assign n7003 = n6981 & n7002;
  assign n7004 = n6965 & n7003;
  assign po0220 = ~n6902 | ~n7004;
  assign n7006 = pi0063 & ~pi0314;
  assign n7007 = pi1044 & n7006;
  assign n7008 = n2619 & n7007;
  assign n7009 = pi0063 & pi0841;
  assign n7010 = n2644 & n7009;
  assign n7011 = ~n7008 & ~n7010;
  assign n7012 = pi0063 & pi0993;
  assign n7013 = n2576 & n7012;
  assign n7014 = pi0024 & pi0063;
  assign n7015 = n2598 & n7014;
  assign n7016 = ~n7013 & ~n7015;
  assign n7017 = pi0063 & n4336;
  assign n7018 = pi0063 & n4062;
  assign n7019 = ~n7017 & ~n7018;
  assign n7020 = n7016 & n7019;
  assign n7021 = n7011 & n7020;
  assign n7022 = pi0063 & n4006;
  assign n7023 = pi0063 & ~n4014;
  assign n7024 = n3110 & n7014;
  assign n7025 = ~n7023 & ~n7024;
  assign n7026 = pi0063 & po0740;
  assign n7027 = n2651 & n7026;
  assign n7028 = ~n3102 & n7027;
  assign n7029 = n7025 & ~n7028;
  assign n7030 = ~n7022 & n7029;
  assign n7031 = n2591 & n7014;
  assign n7032 = n7030 & ~n7031;
  assign n7033 = n2910 & n7014;
  assign n7034 = pi0063 & n2726;
  assign n7035 = n4066 & n7034;
  assign n7036 = ~n7033 & ~n7035;
  assign n7037 = n7032 & n7036;
  assign n7038 = n2917 & n7009;
  assign n7039 = n2913 & n7014;
  assign n7040 = ~n7038 & ~n7039;
  assign n7041 = n2936 & n7006;
  assign n7042 = n7040 & ~n7041;
  assign n7043 = pi0063 & n4043;
  assign n7044 = n2930 & n7043;
  assign n7045 = pi0063 & ~n3553;
  assign n7046 = n4497 & n7045;
  assign n7047 = ~n7044 & ~n7046;
  assign n7048 = ~n4402 & n7006;
  assign n7049 = n7047 & ~n7048;
  assign n7050 = n3042 & n7014;
  assign n7051 = pi0063 & n4504;
  assign n7052 = ~n7050 & ~n7051;
  assign n7053 = n7049 & n7052;
  assign n7054 = n7042 & n7053;
  assign n7055 = n3033 & n7014;
  assign n7056 = n7054 & ~n7055;
  assign n7057 = n7037 & n7056;
  assign n7058 = ~n3072 & n7014;
  assign n7059 = n2847 & n7009;
  assign n7060 = n2834 & n7007;
  assign n7061 = ~n7059 & ~n7060;
  assign n7062 = n2858 & n7009;
  assign n7063 = pi0063 & n4124;
  assign n7064 = n2854 & n7014;
  assign n7065 = n2881 & n7026;
  assign n7066 = n2726 & n7065;
  assign n7067 = ~n7064 & ~n7066;
  assign n7068 = ~n7063 & n7067;
  assign n7069 = ~n7062 & n7068;
  assign n7070 = ~n4133 & n7009;
  assign n7071 = n7069 & ~n7070;
  assign n7072 = n2851 & n7006;
  assign n7073 = n3066 & n7014;
  assign n7074 = ~n7072 & ~n7073;
  assign n7075 = n7071 & n7074;
  assign n7076 = n7061 & n7075;
  assign n7077 = ~n7058 & n7076;
  assign n7078 = n7057 & n7077;
  assign n7079 = ~n4105 & n7006;
  assign n7080 = n2569 & n7014;
  assign n7081 = ~n7079 & ~n7080;
  assign n7082 = pi0063 & n4708;
  assign n7083 = ~n3973 & n7082;
  assign n7084 = pi0063 & n3989;
  assign n7085 = ~n7014 & ~n7084;
  assign n7086 = n2563 & ~n7085;
  assign n7087 = pi0024 & ~pi0063;
  assign n7088 = n2795 & ~n7087;
  assign n7089 = ~n7086 & ~n7088;
  assign n7090 = pi0063 & n2741;
  assign n7091 = n7089 & ~n7090;
  assign n7092 = ~n7083 & n7091;
  assign n7093 = ~n3998 & n7009;
  assign n7094 = n7092 & ~n7093;
  assign n7095 = n7081 & n7094;
  assign n7096 = n3057 & n7014;
  assign n7097 = pi0063 & ~n3057;
  assign n7098 = ~n7096 & ~n7097;
  assign n7099 = n4083 & ~n7098;
  assign n7100 = n2901 & n7006;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = n2681 & n7014;
  assign n7103 = ~n4077 & n7009;
  assign n7104 = ~n7102 & ~n7103;
  assign n7105 = pi0063 & n4089;
  assign n7106 = pi0063 & n4091;
  assign n7107 = pi0063 & n3128;
  assign n7108 = ~n4094 & n7107;
  assign n7109 = ~n4097 & n7026;
  assign n7110 = ~n7108 & ~n7109;
  assign n7111 = n3397 & ~n7110;
  assign n7112 = ~n7106 & ~n7111;
  assign n7113 = ~n7105 & n7112;
  assign n7114 = n4087 & ~n7113;
  assign n7115 = n7104 & ~n7114;
  assign n7116 = n7101 & n7115;
  assign n7117 = n7095 & n7116;
  assign n7118 = n7078 & n7117;
  assign po0221 = ~n7021 | ~n7118;
  assign n7120 = pi0064 & ~pi0314;
  assign n7121 = pi1044 & n7120;
  assign n7122 = n2619 & n7121;
  assign n7123 = pi0064 & pi0841;
  assign n7124 = n2644 & n7123;
  assign n7125 = ~n7122 & ~n7124;
  assign n7126 = pi0064 & pi0993;
  assign n7127 = n2576 & n7126;
  assign n7128 = pi0024 & pi0064;
  assign n7129 = n2598 & n7128;
  assign n7130 = ~n7127 & ~n7129;
  assign n7131 = pi0064 & n4336;
  assign n7132 = pi0064 & n4062;
  assign n7133 = ~n7131 & ~n7132;
  assign n7134 = n7130 & n7133;
  assign n7135 = n7125 & n7134;
  assign n7136 = n2901 & n7120;
  assign n7137 = n2681 & n7128;
  assign n7138 = ~n7136 & ~n7137;
  assign n7139 = ~n4077 & n7123;
  assign n7140 = n7138 & ~n7139;
  assign n7141 = pi0064 & n4091;
  assign n7142 = pi0064 & po0740;
  assign n7143 = ~n4097 & n7142;
  assign n7144 = pi0064 & n4459;
  assign n7145 = ~n7143 & ~n7144;
  assign n7146 = n3397 & ~n7145;
  assign n7147 = pi0064 & ~pi0786;
  assign n7148 = n4088 & n7147;
  assign n7149 = ~n7146 & ~n7148;
  assign n7150 = ~n7141 & n7149;
  assign n7151 = n3547 & ~n7150;
  assign n7152 = n3406 & n7151;
  assign n7153 = n3057 & n7128;
  assign n7154 = pi0064 & ~n3057;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = n4083 & ~n7155;
  assign n7157 = ~n7152 & ~n7156;
  assign n7158 = n7140 & n7157;
  assign n7159 = ~n2895 & n7158;
  assign n7160 = n2917 & n7123;
  assign n7161 = n2913 & n7128;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = n2936 & n7120;
  assign n7164 = n7162 & ~n7163;
  assign n7165 = pi0064 & n4043;
  assign n7166 = n2930 & n7165;
  assign n7167 = pi0064 & ~n3553;
  assign n7168 = n4497 & n7167;
  assign n7169 = ~n7166 & ~n7168;
  assign n7170 = ~n4402 & n7120;
  assign n7171 = n7169 & ~n7170;
  assign n7172 = n3042 & n7128;
  assign n7173 = pi0064 & n4504;
  assign n7174 = ~n7172 & ~n7173;
  assign n7175 = n7171 & n7174;
  assign n7176 = n7164 & n7175;
  assign n7177 = n3033 & n7128;
  assign n7178 = n7176 & ~n7177;
  assign n7179 = pi0064 & n4006;
  assign n7180 = pi0064 & ~n4014;
  assign n7181 = n3110 & n7128;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = n2651 & n7142;
  assign n7184 = ~n3102 & n7183;
  assign n7185 = n7182 & ~n7184;
  assign n7186 = ~n7179 & n7185;
  assign n7187 = n2591 & n7128;
  assign n7188 = n7186 & ~n7187;
  assign n7189 = n2910 & n7128;
  assign n7190 = pi0064 & n2726;
  assign n7191 = n4066 & n7190;
  assign n7192 = ~n7189 & ~n7191;
  assign n7193 = n7188 & n7192;
  assign n7194 = n7178 & n7193;
  assign n7195 = n7159 & n7194;
  assign n7196 = ~n4105 & n7120;
  assign n7197 = n2569 & n7128;
  assign n7198 = ~n7196 & ~n7197;
  assign n7199 = pi0064 & n4708;
  assign n7200 = ~n3973 & n7199;
  assign n7201 = pi0064 & n3989;
  assign n7202 = ~n7128 & ~n7201;
  assign n7203 = n2563 & ~n7202;
  assign n7204 = n2795 & n7128;
  assign n7205 = ~n7203 & ~n7204;
  assign n7206 = pi0064 & n2741;
  assign n7207 = n7205 & ~n7206;
  assign n7208 = ~n7200 & n7207;
  assign n7209 = ~n3998 & n7123;
  assign n7210 = n7208 & ~n7209;
  assign n7211 = n7198 & n7210;
  assign n7212 = ~n3072 & n7128;
  assign n7213 = n2847 & n7123;
  assign n7214 = n2834 & n7121;
  assign n7215 = ~n7213 & ~n7214;
  assign n7216 = n2858 & n7123;
  assign n7217 = pi0064 & n4124;
  assign n7218 = n2854 & n7128;
  assign n7219 = n2881 & n7142;
  assign n7220 = n2726 & n7219;
  assign n7221 = ~n7218 & ~n7220;
  assign n7222 = ~n7217 & n7221;
  assign n7223 = ~n7216 & n7222;
  assign n7224 = ~n4133 & n7123;
  assign n7225 = n7223 & ~n7224;
  assign n7226 = n2851 & n7120;
  assign n7227 = n3066 & n7128;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = n7225 & n7228;
  assign n7230 = n7215 & n7229;
  assign n7231 = ~n7212 & n7230;
  assign n7232 = n7211 & n7231;
  assign n7233 = n7195 & n7232;
  assign po0222 = ~n7135 | ~n7233;
  assign n7235 = pi0065 & pi0841;
  assign n7236 = n2917 & n7235;
  assign n7237 = pi0024 & pi0065;
  assign n7238 = n2913 & n7237;
  assign n7239 = ~n7236 & ~n7238;
  assign n7240 = pi0065 & ~pi0314;
  assign n7241 = n2936 & n7240;
  assign n7242 = n7239 & ~n7241;
  assign n7243 = pi0065 & n4043;
  assign n7244 = n2930 & n7243;
  assign n7245 = pi0065 & ~n3553;
  assign n7246 = n4497 & n7245;
  assign n7247 = ~n7244 & ~n7246;
  assign n7248 = ~n4402 & n7240;
  assign n7249 = n7247 & ~n7248;
  assign n7250 = n3042 & n7237;
  assign n7251 = pi0065 & n4504;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = n7249 & n7252;
  assign n7254 = n7242 & n7253;
  assign n7255 = n3033 & n7237;
  assign n7256 = n7254 & ~n7255;
  assign n7257 = pi0065 & n4006;
  assign n7258 = pi0065 & ~n4014;
  assign n7259 = n3110 & n7237;
  assign n7260 = ~n7258 & ~n7259;
  assign n7261 = pi0065 & po0740;
  assign n7262 = n2651 & n7261;
  assign n7263 = ~n3102 & n7262;
  assign n7264 = n7260 & ~n7263;
  assign n7265 = ~n7257 & n7264;
  assign n7266 = n2591 & n7237;
  assign n7267 = n7265 & ~n7266;
  assign n7268 = n2910 & n7237;
  assign n7269 = pi0065 & n2726;
  assign n7270 = n4066 & n7269;
  assign n7271 = ~n7268 & ~n7270;
  assign n7272 = n7267 & n7271;
  assign n7273 = n7256 & n7272;
  assign n7274 = ~n3072 & n7237;
  assign n7275 = n2847 & n7235;
  assign n7276 = pi1044 & n7240;
  assign n7277 = n2834 & n7276;
  assign n7278 = ~n7275 & ~n7277;
  assign n7279 = n2858 & n7235;
  assign n7280 = pi0065 & n4124;
  assign n7281 = n2854 & n7237;
  assign n7282 = n2881 & n7261;
  assign n7283 = n2726 & n7282;
  assign n7284 = ~n7281 & ~n7283;
  assign n7285 = ~n7280 & n7284;
  assign n7286 = ~n7279 & n7285;
  assign n7287 = ~n4133 & n7235;
  assign n7288 = n7286 & ~n7287;
  assign n7289 = n2851 & n7240;
  assign n7290 = n3066 & n7237;
  assign n7291 = ~n7289 & ~n7290;
  assign n7292 = n7288 & n7291;
  assign n7293 = n7278 & n7292;
  assign n7294 = ~n7274 & n7293;
  assign n7295 = n7273 & n7294;
  assign n7296 = n2619 & n7276;
  assign n7297 = n2644 & n7235;
  assign n7298 = ~n7296 & ~n7297;
  assign n7299 = pi0065 & pi0993;
  assign n7300 = n2576 & n7299;
  assign n7301 = n2598 & n7237;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = pi0065 & n4336;
  assign n7304 = pi0065 & n4062;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = n7302 & n7305;
  assign n7307 = n7298 & n7306;
  assign n7308 = n7295 & n7307;
  assign n7309 = n3057 & n7237;
  assign n7310 = pi0065 & ~n3057;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = n4083 & ~n7311;
  assign n7313 = n2901 & n7240;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = n2681 & n7237;
  assign n7316 = ~n4077 & n7235;
  assign n7317 = ~n7315 & ~n7316;
  assign n7318 = pi0065 & n4091;
  assign n7319 = ~n4097 & n7261;
  assign n7320 = pi0065 & n4459;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = n3397 & ~n7321;
  assign n7323 = ~pi0065 & ~pi0786;
  assign n7324 = n4088 & ~n7323;
  assign n7325 = ~n7322 & ~n7324;
  assign n7326 = ~n7318 & n7325;
  assign n7327 = n4087 & ~n7326;
  assign n7328 = n7317 & ~n7327;
  assign n7329 = n7314 & n7328;
  assign n7330 = ~n4105 & n7240;
  assign n7331 = n2569 & n7237;
  assign n7332 = ~n7330 & ~n7331;
  assign n7333 = pi0065 & n4708;
  assign n7334 = ~n3973 & n7333;
  assign n7335 = pi0065 & n3989;
  assign n7336 = ~n7237 & ~n7335;
  assign n7337 = n2563 & ~n7336;
  assign n7338 = n2795 & n7237;
  assign n7339 = ~n7337 & ~n7338;
  assign n7340 = pi0065 & n2741;
  assign n7341 = n7339 & ~n7340;
  assign n7342 = ~n7334 & n7341;
  assign n7343 = ~n3998 & n7235;
  assign n7344 = n7342 & ~n7343;
  assign n7345 = n7332 & n7344;
  assign n7346 = n7329 & n7345;
  assign po0223 = ~n7308 | ~n7346;
  assign n7348 = pi0066 & ~pi0314;
  assign n7349 = pi1044 & n7348;
  assign n7350 = n2619 & n7349;
  assign n7351 = pi0066 & pi0841;
  assign n7352 = n2644 & n7351;
  assign n7353 = ~n7350 & ~n7352;
  assign n7354 = pi0066 & pi0993;
  assign n7355 = n2576 & n7354;
  assign n7356 = pi0024 & pi0066;
  assign n7357 = n2598 & n7356;
  assign n7358 = ~n7355 & ~n7357;
  assign n7359 = pi0066 & n4336;
  assign n7360 = pi0066 & n4062;
  assign n7361 = ~n7359 & ~n7360;
  assign n7362 = n7358 & n7361;
  assign n7363 = n7353 & n7362;
  assign n7364 = n2917 & n7351;
  assign n7365 = n2913 & n7356;
  assign n7366 = ~n7364 & ~n7365;
  assign n7367 = n2936 & n7348;
  assign n7368 = n7366 & ~n7367;
  assign n7369 = pi0066 & n4043;
  assign n7370 = n2930 & n7369;
  assign n7371 = pi0066 & ~n3553;
  assign n7372 = n4497 & n7371;
  assign n7373 = ~n7370 & ~n7372;
  assign n7374 = ~n4402 & n7348;
  assign n7375 = n7373 & ~n7374;
  assign n7376 = n3042 & n7356;
  assign n7377 = pi0066 & n4504;
  assign n7378 = ~n7376 & ~n7377;
  assign n7379 = n7375 & n7378;
  assign n7380 = n7368 & n7379;
  assign n7381 = n3033 & n7356;
  assign n7382 = n7380 & ~n7381;
  assign n7383 = pi0066 & n4006;
  assign n7384 = pi0066 & ~n4014;
  assign n7385 = n3110 & n7356;
  assign n7386 = ~n7384 & ~n7385;
  assign n7387 = pi0066 & po0740;
  assign n7388 = n2651 & n7387;
  assign n7389 = ~n3102 & n7388;
  assign n7390 = n7386 & ~n7389;
  assign n7391 = ~n7383 & n7390;
  assign n7392 = n2591 & n7356;
  assign n7393 = n7391 & ~n7392;
  assign n7394 = n2910 & n7356;
  assign n7395 = pi0066 & n2726;
  assign n7396 = n4066 & n7395;
  assign n7397 = ~n7394 & ~n7396;
  assign n7398 = n7393 & n7397;
  assign n7399 = n7382 & n7398;
  assign n7400 = ~n4964 & ~n4967;
  assign n7401 = pi0314 & ~n4983;
  assign n7402 = ~n7400 & n7401;
  assign n7403 = ~n7348 & ~n7402;
  assign n7404 = n2901 & ~n7403;
  assign n7405 = n2681 & n7356;
  assign n7406 = ~n4077 & n7351;
  assign n7407 = ~n7405 & ~n7406;
  assign n7408 = pi0066 & n4091;
  assign n7409 = ~n4097 & n7387;
  assign n7410 = pi0066 & n4459;
  assign n7411 = ~n7409 & ~n7410;
  assign n7412 = n3397 & ~n7411;
  assign n7413 = pi0066 & ~pi0786;
  assign n7414 = n4088 & n7413;
  assign n7415 = ~n7412 & ~n7414;
  assign n7416 = ~n7408 & n7415;
  assign n7417 = n3547 & ~n7416;
  assign n7418 = n3406 & n7417;
  assign n7419 = n3057 & n7356;
  assign n7420 = pi0066 & ~n3057;
  assign n7421 = ~n7419 & ~n7420;
  assign n7422 = n4083 & ~n7421;
  assign n7423 = ~n7418 & ~n7422;
  assign n7424 = n7407 & n7423;
  assign n7425 = ~n7404 & n7424;
  assign n7426 = n7399 & n7425;
  assign n7427 = ~n4105 & n7348;
  assign n7428 = n2569 & n7356;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 = pi0066 & n4708;
  assign n7431 = ~n3973 & n7430;
  assign n7432 = pi0066 & n3989;
  assign n7433 = ~n7356 & ~n7432;
  assign n7434 = n2563 & ~n7433;
  assign n7435 = n2795 & n7356;
  assign n7436 = ~n7434 & ~n7435;
  assign n7437 = pi0066 & n2741;
  assign n7438 = n7436 & ~n7437;
  assign n7439 = ~n7431 & n7438;
  assign n7440 = ~n3998 & n7351;
  assign n7441 = n7439 & ~n7440;
  assign n7442 = n7429 & n7441;
  assign n7443 = ~n3072 & n7356;
  assign n7444 = n2847 & n7351;
  assign n7445 = n2834 & n7349;
  assign n7446 = ~n7444 & ~n7445;
  assign n7447 = n2858 & n7351;
  assign n7448 = pi0066 & n4124;
  assign n7449 = n2854 & n7356;
  assign n7450 = n2881 & n7387;
  assign n7451 = n2726 & n7450;
  assign n7452 = ~n7449 & ~n7451;
  assign n7453 = ~n7448 & n7452;
  assign n7454 = ~n7447 & n7453;
  assign n7455 = ~n4133 & n7351;
  assign n7456 = n7454 & ~n7455;
  assign n7457 = n2851 & n7348;
  assign n7458 = n3066 & n7356;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = n7456 & n7459;
  assign n7461 = n7446 & n7460;
  assign n7462 = ~n7443 & n7461;
  assign n7463 = n7442 & n7462;
  assign n7464 = n7426 & n7463;
  assign po0224 = ~n7363 | ~n7464;
  assign n7466 = pi0067 & n4336;
  assign n7467 = pi0067 & n2741;
  assign n7468 = pi0067 & n4523;
  assign n7469 = ~n3973 & n7468;
  assign n7470 = pi0067 & pi0841;
  assign n7471 = ~n3998 & n7470;
  assign n7472 = pi0024 & pi0067;
  assign n7473 = pi0067 & n3989;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = n2563 & ~n7474;
  assign n7476 = n2795 & n7472;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~n7471 & n7477;
  assign n7479 = ~n7469 & n7478;
  assign n7480 = ~n7467 & n7479;
  assign n7481 = pi0067 & ~n4061;
  assign n7482 = n4060 & n7481;
  assign n7483 = n7480 & ~n7482;
  assign n7484 = pi0067 & ~pi0314;
  assign n7485 = ~n4105 & n7484;
  assign n7486 = n2569 & n7472;
  assign n7487 = ~n7485 & ~n7486;
  assign n7488 = pi0067 & pi0993;
  assign n7489 = n2576 & n7488;
  assign n7490 = n2598 & n7472;
  assign n7491 = ~n7489 & ~n7490;
  assign n7492 = n7487 & n7491;
  assign n7493 = pi0067 & n4067;
  assign n7494 = n3042 & n7472;
  assign n7495 = n2913 & n7472;
  assign n7496 = n2917 & n7470;
  assign n7497 = ~n7495 & ~n7496;
  assign n7498 = pi0067 & ~n3553;
  assign n7499 = n4497 & n7498;
  assign n7500 = ~pi0067 & ~pi0314;
  assign n7501 = n2533 & ~n7500;
  assign n7502 = n2544 & n7484;
  assign n7503 = ~n7501 & ~n7502;
  assign n7504 = pi0067 & n5491;
  assign n7505 = n7503 & ~n7504;
  assign n7506 = ~n7499 & n7505;
  assign n7507 = n2936 & n7484;
  assign n7508 = n7506 & ~n7507;
  assign n7509 = pi0067 & n4504;
  assign n7510 = n7508 & ~n7509;
  assign n7511 = n7497 & n7510;
  assign n7512 = ~n7494 & n7511;
  assign n7513 = n3033 & n7472;
  assign n7514 = n7512 & ~n7513;
  assign n7515 = n2910 & n7472;
  assign n7516 = n7514 & ~n7515;
  assign n7517 = ~n7493 & n7516;
  assign n7518 = pi0067 & ~n4014;
  assign n7519 = n3110 & n7472;
  assign n7520 = ~n7518 & ~n7519;
  assign n7521 = pi0067 & po0740;
  assign n7522 = n2651 & n7521;
  assign n7523 = ~n3102 & n7522;
  assign n7524 = pi0067 & n4006;
  assign n7525 = ~n7523 & ~n7524;
  assign n7526 = pi1044 & n7484;
  assign n7527 = n2619 & n7526;
  assign n7528 = n2644 & n7470;
  assign n7529 = ~n7527 & ~n7528;
  assign n7530 = n2591 & n7472;
  assign n7531 = n7529 & ~n7530;
  assign n7532 = n7525 & n7531;
  assign n7533 = n7520 & n7532;
  assign n7534 = n7517 & n7533;
  assign n7535 = n7492 & n7534;
  assign n7536 = n7483 & n7535;
  assign n7537 = ~n7466 & n7536;
  assign n7538 = pi0067 & n4089;
  assign n7539 = pi0067 & n4091;
  assign n7540 = pi0067 & n3128;
  assign n7541 = ~n4094 & n7540;
  assign n7542 = ~n4097 & n7521;
  assign n7543 = ~n7541 & ~n7542;
  assign n7544 = n3397 & ~n7543;
  assign n7545 = ~n7539 & ~n7544;
  assign n7546 = ~n7538 & n7545;
  assign n7547 = n4087 & ~n7546;
  assign n7548 = n3057 & n7472;
  assign n7549 = pi0067 & ~n3057;
  assign n7550 = ~n7548 & ~n7549;
  assign n7551 = n4083 & ~n7550;
  assign n7552 = n2901 & n7484;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n3072 & n7472;
  assign n7555 = n2847 & n7470;
  assign n7556 = n2834 & n7526;
  assign n7557 = ~n7555 & ~n7556;
  assign n7558 = n2858 & n7470;
  assign n7559 = pi0067 & n4124;
  assign n7560 = n2854 & n7472;
  assign n7561 = n2881 & n7521;
  assign n7562 = n2726 & n7561;
  assign n7563 = ~n7560 & ~n7562;
  assign n7564 = ~n7559 & n7563;
  assign n7565 = ~n7558 & n7564;
  assign n7566 = ~n4133 & n7470;
  assign n7567 = n7565 & ~n7566;
  assign n7568 = n2851 & n7484;
  assign n7569 = n3066 & n7472;
  assign n7570 = ~n7568 & ~n7569;
  assign n7571 = n7567 & n7570;
  assign n7572 = n7557 & n7571;
  assign n7573 = ~n7554 & n7572;
  assign n7574 = n2681 & n7472;
  assign n7575 = ~n4077 & n7470;
  assign n7576 = ~n7574 & ~n7575;
  assign n7577 = n7573 & n7576;
  assign n7578 = n7553 & n7577;
  assign n7579 = ~n7547 & n7578;
  assign po0225 = ~n7537 | ~n7579;
  assign n7581 = pi0068 & pi0841;
  assign n7582 = n2917 & n7581;
  assign n7583 = pi0024 & pi0068;
  assign n7584 = n2913 & n7583;
  assign n7585 = ~n7582 & ~n7584;
  assign n7586 = pi0068 & ~pi0314;
  assign n7587 = n2936 & n7586;
  assign n7588 = n7585 & ~n7587;
  assign n7589 = pi0068 & n4043;
  assign n7590 = n2930 & n7589;
  assign n7591 = pi0068 & ~n3553;
  assign n7592 = n4497 & n7591;
  assign n7593 = ~n7590 & ~n7592;
  assign n7594 = ~n4402 & n7586;
  assign n7595 = n7593 & ~n7594;
  assign n7596 = n3042 & n7583;
  assign n7597 = pi0068 & n4504;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = n7595 & n7598;
  assign n7600 = n7588 & n7599;
  assign n7601 = n3033 & n7583;
  assign n7602 = n7600 & ~n7601;
  assign n7603 = pi0068 & n4006;
  assign n7604 = pi0068 & ~n4014;
  assign n7605 = n3110 & n7583;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = pi0068 & po0740;
  assign n7608 = n2651 & n7607;
  assign n7609 = ~n3102 & n7608;
  assign n7610 = n7606 & ~n7609;
  assign n7611 = ~n7603 & n7610;
  assign n7612 = n2591 & n7583;
  assign n7613 = n7611 & ~n7612;
  assign n7614 = n2910 & n7583;
  assign n7615 = pi0068 & n2726;
  assign n7616 = n4066 & n7615;
  assign n7617 = ~n7614 & ~n7616;
  assign n7618 = n7613 & n7617;
  assign n7619 = n7602 & n7618;
  assign n7620 = ~n3072 & n7583;
  assign n7621 = n2847 & n7581;
  assign n7622 = pi1044 & n7586;
  assign n7623 = n2834 & n7622;
  assign n7624 = ~n7621 & ~n7623;
  assign n7625 = n2858 & n7581;
  assign n7626 = pi0068 & n4124;
  assign n7627 = n2854 & n7583;
  assign n7628 = n2881 & n7607;
  assign n7629 = n2726 & n7628;
  assign n7630 = ~n7627 & ~n7629;
  assign n7631 = ~n7626 & n7630;
  assign n7632 = ~n7625 & n7631;
  assign n7633 = ~n4133 & n7581;
  assign n7634 = n7632 & ~n7633;
  assign n7635 = n2851 & n7586;
  assign n7636 = n3066 & n7583;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = n7634 & n7637;
  assign n7639 = n7624 & n7638;
  assign n7640 = ~n7620 & n7639;
  assign n7641 = n7619 & n7640;
  assign n7642 = n2619 & n7622;
  assign n7643 = n2644 & n7581;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = pi0068 & pi0993;
  assign n7646 = n2576 & n7645;
  assign n7647 = n2598 & n7583;
  assign n7648 = ~n7646 & ~n7647;
  assign n7649 = pi0068 & n4336;
  assign n7650 = pi0068 & n4062;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = n7648 & n7651;
  assign n7653 = n7644 & n7652;
  assign n7654 = n7641 & n7653;
  assign n7655 = n3057 & n7583;
  assign n7656 = pi0068 & ~n3057;
  assign n7657 = ~n7655 & ~n7656;
  assign n7658 = n4083 & ~n7657;
  assign n7659 = n2901 & n7586;
  assign n7660 = ~n7658 & ~n7659;
  assign n7661 = n2681 & n7583;
  assign n7662 = ~n4077 & n7581;
  assign n7663 = ~n7661 & ~n7662;
  assign n7664 = pi0068 & n4091;
  assign n7665 = pi0068 & n4459;
  assign n7666 = ~n4097 & n7607;
  assign n7667 = n2440 & n3468;
  assign n7668 = ~n7666 & ~n7667;
  assign n7669 = ~n7665 & n7668;
  assign n7670 = n3397 & ~n7669;
  assign n7671 = pi0068 & ~pi0786;
  assign n7672 = n4088 & n7671;
  assign n7673 = ~n7670 & ~n7672;
  assign n7674 = ~n7664 & n7673;
  assign n7675 = n4087 & ~n7674;
  assign n7676 = n7663 & ~n7675;
  assign n7677 = n7660 & n7676;
  assign n7678 = ~n4105 & n7586;
  assign n7679 = n2569 & n7583;
  assign n7680 = ~n7678 & ~n7679;
  assign n7681 = pi0068 & n4708;
  assign n7682 = ~n3973 & n7681;
  assign n7683 = pi0068 & n3989;
  assign n7684 = ~n7583 & ~n7683;
  assign n7685 = n2563 & ~n7684;
  assign n7686 = n2795 & n7583;
  assign n7687 = ~n7685 & ~n7686;
  assign n7688 = pi0068 & n2741;
  assign n7689 = n7687 & ~n7688;
  assign n7690 = ~n7682 & n7689;
  assign n7691 = ~n3998 & n7581;
  assign n7692 = n7690 & ~n7691;
  assign n7693 = n7680 & n7692;
  assign n7694 = n7677 & n7693;
  assign po0226 = ~n7654 | ~n7694;
  assign n7696 = pi0069 & n2741;
  assign n7697 = pi0069 & n4523;
  assign n7698 = ~n3973 & n7697;
  assign n7699 = pi0069 & pi0841;
  assign n7700 = ~n3998 & n7699;
  assign n7701 = pi0024 & pi0069;
  assign n7702 = pi0069 & n3989;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = n2563 & ~n7703;
  assign n7705 = n2795 & n7701;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = ~n7700 & n7706;
  assign n7708 = ~n7698 & n7707;
  assign n7709 = ~n7696 & n7708;
  assign n7710 = pi0069 & po0740;
  assign n7711 = n2651 & n7710;
  assign n7712 = ~n3102 & n7711;
  assign n7713 = pi0069 & n4006;
  assign n7714 = ~n7712 & ~n7713;
  assign n7715 = pi0069 & n4336;
  assign n7716 = pi0069 & ~pi0314;
  assign n7717 = ~n4105 & n7716;
  assign n7718 = n2569 & n7701;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = pi0069 & pi0993;
  assign n7721 = n2576 & n7720;
  assign n7722 = n2598 & n7701;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = n7719 & n7723;
  assign n7725 = n2591 & n7701;
  assign n7726 = pi0069 & ~n4014;
  assign n7727 = n3110 & n7701;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = pi1044 & n7716;
  assign n7730 = n2619 & n7729;
  assign n7731 = n2644 & n7699;
  assign n7732 = ~n7730 & ~n7731;
  assign n7733 = n7728 & n7732;
  assign n7734 = ~n7725 & n7733;
  assign n7735 = n7724 & n7734;
  assign n7736 = ~n7715 & n7735;
  assign n7737 = n7714 & n7736;
  assign n7738 = n7709 & n7737;
  assign n7739 = pi0069 & n4067;
  assign n7740 = n2533 & n7716;
  assign n7741 = ~n2537 & ~n7740;
  assign n7742 = pi0069 & ~n3553;
  assign n7743 = n4497 & n7742;
  assign n7744 = pi0069 & n4043;
  assign n7745 = n2930 & n7744;
  assign n7746 = ~n7743 & ~n7745;
  assign n7747 = pi0069 & n4504;
  assign n7748 = n3042 & n7701;
  assign n7749 = ~n7747 & ~n7748;
  assign n7750 = ~n3455 & n7716;
  assign n7751 = n7749 & ~n7750;
  assign n7752 = n2913 & n7701;
  assign n7753 = n2917 & n7699;
  assign n7754 = ~n7752 & ~n7753;
  assign n7755 = n7751 & n7754;
  assign n7756 = n7746 & n7755;
  assign n7757 = n7741 & n7756;
  assign n7758 = n3033 & n7701;
  assign n7759 = n7757 & ~n7758;
  assign n7760 = n2910 & n7701;
  assign n7761 = n7759 & ~n7760;
  assign n7762 = ~n7739 & n7761;
  assign n7763 = pi0069 & ~n4061;
  assign n7764 = n4060 & n7763;
  assign n7765 = n7762 & ~n7764;
  assign n7766 = n7738 & n7765;
  assign n7767 = pi0069 & n4089;
  assign n7768 = pi0069 & n4091;
  assign n7769 = pi0069 & n3128;
  assign n7770 = ~n4094 & n7769;
  assign n7771 = ~n4097 & n7710;
  assign n7772 = ~n7770 & ~n7771;
  assign n7773 = n3397 & ~n7772;
  assign n7774 = ~n7768 & ~n7773;
  assign n7775 = ~n7767 & n7774;
  assign n7776 = n4087 & ~n7775;
  assign n7777 = n3057 & n7701;
  assign n7778 = pi0069 & ~n3057;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = n4083 & ~n7779;
  assign n7781 = n2901 & n7716;
  assign n7782 = ~n7780 & ~n7781;
  assign n7783 = ~n3072 & n7701;
  assign n7784 = n2847 & n7699;
  assign n7785 = n2834 & n7729;
  assign n7786 = ~n7784 & ~n7785;
  assign n7787 = n2858 & n7699;
  assign n7788 = pi0069 & n4124;
  assign n7789 = n2854 & n7701;
  assign n7790 = n2881 & n7710;
  assign n7791 = n2726 & n7790;
  assign n7792 = ~n7789 & ~n7791;
  assign n7793 = ~n7788 & n7792;
  assign n7794 = ~n7787 & n7793;
  assign n7795 = ~n4133 & n7699;
  assign n7796 = n7794 & ~n7795;
  assign n7797 = n2851 & n7716;
  assign n7798 = n3066 & n7701;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = n7796 & n7799;
  assign n7801 = n7786 & n7800;
  assign n7802 = ~n7783 & n7801;
  assign n7803 = n2681 & n7701;
  assign n7804 = ~n4077 & n7699;
  assign n7805 = ~n7803 & ~n7804;
  assign n7806 = n7802 & n7805;
  assign n7807 = n7782 & n7806;
  assign n7808 = ~n7776 & n7807;
  assign po0227 = ~n7766 | ~n7808;
  assign n7810 = pi0070 & ~pi0314;
  assign n7811 = pi1044 & n7810;
  assign n7812 = n2619 & n7811;
  assign n7813 = pi0070 & pi0841;
  assign n7814 = n2644 & n7813;
  assign n7815 = ~n7812 & ~n7814;
  assign n7816 = pi0070 & n4336;
  assign n7817 = pi0070 & n4062;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = n7815 & n7818;
  assign n7820 = pi0024 & pi0070;
  assign n7821 = n2910 & n7820;
  assign n7822 = pi0070 & n2726;
  assign n7823 = n4066 & n7822;
  assign n7824 = ~n7821 & ~n7823;
  assign n7825 = n2917 & n7813;
  assign n7826 = n2913 & n7820;
  assign n7827 = ~n7825 & ~n7826;
  assign n7828 = n2936 & n7810;
  assign n7829 = n7827 & ~n7828;
  assign n7830 = pi0070 & n4043;
  assign n7831 = n2930 & n7830;
  assign n7832 = pi0070 & ~n3553;
  assign n7833 = n4497 & n7832;
  assign n7834 = ~n7831 & ~n7833;
  assign n7835 = ~n4402 & n7810;
  assign n7836 = n7834 & ~n7835;
  assign n7837 = n3042 & n7820;
  assign n7838 = pi0070 & n4504;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = n7836 & n7839;
  assign n7841 = n7829 & n7840;
  assign n7842 = n3033 & n7820;
  assign n7843 = n7841 & ~n7842;
  assign n7844 = pi0070 & n4006;
  assign n7845 = pi0070 & ~n4014;
  assign n7846 = n3110 & n7820;
  assign n7847 = ~n7845 & ~n7846;
  assign n7848 = pi0070 & po0740;
  assign n7849 = n2651 & n7848;
  assign n7850 = ~n3102 & n7849;
  assign n7851 = n7847 & ~n7850;
  assign n7852 = ~n7844 & n7851;
  assign n7853 = n2591 & n7820;
  assign n7854 = n7852 & ~n7853;
  assign n7855 = n7843 & n7854;
  assign n7856 = n7824 & n7855;
  assign n7857 = n7819 & n7856;
  assign n7858 = pi0070 & pi0993;
  assign n7859 = n2576 & n7858;
  assign n7860 = n2598 & n7820;
  assign n7861 = ~n7859 & ~n7860;
  assign n7862 = pi0070 & n4708;
  assign n7863 = ~n3973 & n7862;
  assign n7864 = pi0070 & n3989;
  assign n7865 = ~n7820 & ~n7864;
  assign n7866 = n2563 & ~n7865;
  assign n7867 = n2795 & n7820;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = pi0070 & n2741;
  assign n7870 = n7868 & ~n7869;
  assign n7871 = ~n7863 & n7870;
  assign n7872 = ~n3998 & n7813;
  assign n7873 = n7871 & ~n7872;
  assign n7874 = ~n4105 & n7810;
  assign n7875 = n2569 & n7820;
  assign n7876 = ~n7874 & ~n7875;
  assign n7877 = n7873 & n7876;
  assign n7878 = n7861 & n7877;
  assign n7879 = ~n3072 & n7820;
  assign n7880 = n2847 & n7813;
  assign n7881 = n2834 & n7811;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = n2858 & n7813;
  assign n7884 = pi0070 & n4124;
  assign n7885 = n2854 & n7820;
  assign n7886 = n2881 & n7848;
  assign n7887 = n2726 & n7886;
  assign n7888 = ~n7885 & ~n7887;
  assign n7889 = ~n7884 & n7888;
  assign n7890 = ~n7883 & n7889;
  assign n7891 = ~n4133 & n7813;
  assign n7892 = n7890 & ~n7891;
  assign n7893 = n2851 & n7810;
  assign n7894 = n3066 & n7820;
  assign n7895 = ~n7893 & ~n7894;
  assign n7896 = n7892 & n7895;
  assign n7897 = n7882 & n7896;
  assign n7898 = ~n7879 & n7897;
  assign n7899 = pi0589 & ~n3018;
  assign n7900 = pi0593 & n7899;
  assign n7901 = n7899 & ~n7900;
  assign n7902 = n4094 & ~n7901;
  assign n7903 = ~pi0070 & ~n4094;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = n3128 & n7904;
  assign n7906 = ~n4097 & n7848;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = n3397 & ~n7907;
  assign n7909 = pi0070 & n4091;
  assign n7910 = pi0070 & n4089;
  assign n7911 = ~n7909 & ~n7910;
  assign n7912 = ~n7908 & n7911;
  assign n7913 = n2777 & ~n7912;
  assign n7914 = n3406 & n7913;
  assign n7915 = n3057 & n7820;
  assign n7916 = pi0070 & ~n3057;
  assign n7917 = ~n7915 & ~n7916;
  assign n7918 = n4083 & ~n7917;
  assign n7919 = n2901 & n7810;
  assign n7920 = ~n7918 & ~n7919;
  assign n7921 = n2681 & n7820;
  assign n7922 = ~n4077 & n7813;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = ~n3350 & n7923;
  assign n7925 = n7920 & n7924;
  assign n7926 = ~n7914 & n7925;
  assign n7927 = n7898 & n7926;
  assign n7928 = n7878 & n7927;
  assign po0228 = ~n7857 | ~n7928;
  assign n7930 = pi0071 & ~pi0314;
  assign n7931 = ~n4105 & n7930;
  assign n7932 = pi0024 & pi0071;
  assign n7933 = n2569 & n7932;
  assign n7934 = ~n7931 & ~n7933;
  assign n7935 = pi0071 & pi0993;
  assign n7936 = n2576 & n7935;
  assign n7937 = n2598 & n7932;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = n7934 & n7938;
  assign n7940 = pi0071 & n2741;
  assign n7941 = pi0071 & n4523;
  assign n7942 = ~n3973 & n7941;
  assign n7943 = pi0071 & pi0841;
  assign n7944 = ~n3998 & n7943;
  assign n7945 = pi0071 & n3989;
  assign n7946 = ~n7932 & ~n7945;
  assign n7947 = n2563 & ~n7946;
  assign n7948 = n2795 & n7932;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = ~n7944 & n7949;
  assign n7951 = ~n7942 & n7950;
  assign n7952 = ~n7940 & n7951;
  assign n7953 = pi0071 & ~n4061;
  assign n7954 = n4060 & n7953;
  assign n7955 = n7952 & ~n7954;
  assign n7956 = pi0071 & n4336;
  assign n7957 = pi0071 & n4067;
  assign n7958 = n3042 & n7932;
  assign n7959 = n2913 & n7932;
  assign n7960 = n2917 & n7943;
  assign n7961 = ~n7959 & ~n7960;
  assign n7962 = pi0071 & ~n3553;
  assign n7963 = n4497 & n7962;
  assign n7964 = ~pi0071 & ~pi0314;
  assign n7965 = n2544 & ~n7964;
  assign n7966 = n2533 & n7930;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = pi0071 & n5491;
  assign n7969 = n7967 & ~n7968;
  assign n7970 = ~n7963 & n7969;
  assign n7971 = n2936 & n7930;
  assign n7972 = n7970 & ~n7971;
  assign n7973 = pi0071 & n4504;
  assign n7974 = n7972 & ~n7973;
  assign n7975 = n7961 & n7974;
  assign n7976 = ~n7958 & n7975;
  assign n7977 = n3033 & n7932;
  assign n7978 = n7976 & ~n7977;
  assign n7979 = n2910 & n7932;
  assign n7980 = n7978 & ~n7979;
  assign n7981 = ~n7957 & n7980;
  assign n7982 = pi0071 & ~n4014;
  assign n7983 = n3110 & n7932;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = pi0071 & po0740;
  assign n7986 = n2651 & n7985;
  assign n7987 = ~n3102 & n7986;
  assign n7988 = pi0071 & n4006;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = pi1044 & n7930;
  assign n7991 = n2619 & n7990;
  assign n7992 = n2644 & n7943;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = n2591 & n7932;
  assign n7995 = n7993 & ~n7994;
  assign n7996 = n7989 & n7995;
  assign n7997 = n7984 & n7996;
  assign n7998 = n7981 & n7997;
  assign n7999 = ~n7956 & n7998;
  assign n8000 = n7955 & n7999;
  assign n8001 = n7939 & n8000;
  assign n8002 = pi0071 & n4091;
  assign n8003 = ~n4097 & n7985;
  assign n8004 = pi0071 & n4459;
  assign n8005 = ~n8003 & ~n8004;
  assign n8006 = n3397 & ~n8005;
  assign n8007 = pi0071 & ~pi0786;
  assign n8008 = n4088 & n8007;
  assign n8009 = ~n8006 & ~n8008;
  assign n8010 = ~n8002 & n8009;
  assign n8011 = n3547 & ~n8010;
  assign n8012 = n3406 & n8011;
  assign n8013 = n3057 & n7932;
  assign n8014 = pi0071 & ~n3057;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = n4083 & ~n8015;
  assign n8017 = ~n8012 & ~n8016;
  assign n8018 = n7400 & n7401;
  assign n8019 = ~n7930 & ~n8018;
  assign n8020 = n2901 & ~n8019;
  assign n8021 = ~n3072 & n7932;
  assign n8022 = n2847 & n7943;
  assign n8023 = n2834 & n7990;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = n2858 & n7943;
  assign n8026 = pi0071 & n4124;
  assign n8027 = n2854 & n7932;
  assign n8028 = n2881 & n7985;
  assign n8029 = n2726 & n8028;
  assign n8030 = ~n8027 & ~n8029;
  assign n8031 = ~n8026 & n8030;
  assign n8032 = ~n8025 & n8031;
  assign n8033 = ~n4133 & n7943;
  assign n8034 = n8032 & ~n8033;
  assign n8035 = n2851 & n7930;
  assign n8036 = n3066 & n7932;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = n8034 & n8037;
  assign n8039 = n8024 & n8038;
  assign n8040 = ~n8021 & n8039;
  assign n8041 = n2681 & n7932;
  assign n8042 = ~n4077 & n7943;
  assign n8043 = ~n8041 & ~n8042;
  assign n8044 = n8040 & n8043;
  assign n8045 = ~n8020 & n8044;
  assign n8046 = n8017 & n8045;
  assign po0229 = ~n8001 | ~n8046;
  assign n8048 = pi0072 & n4336;
  assign n8049 = pi0072 & n2741;
  assign n8050 = pi0072 & n4585;
  assign n8051 = pi0072 & pi0841;
  assign n8052 = ~n3998 & n8051;
  assign n8053 = pi0024 & pi0072;
  assign n8054 = pi0072 & n3989;
  assign n8055 = ~n8053 & ~n8054;
  assign n8056 = n2563 & ~n8055;
  assign n8057 = n2795 & n8053;
  assign n8058 = ~n8056 & ~n8057;
  assign n8059 = ~n8052 & n8058;
  assign n8060 = ~n8050 & n8059;
  assign n8061 = ~n8049 & n8060;
  assign n8062 = pi0072 & ~n4061;
  assign n8063 = n4060 & n8062;
  assign n8064 = n8061 & ~n8063;
  assign n8065 = pi0072 & ~pi0314;
  assign n8066 = ~n4105 & n8065;
  assign n8067 = n2569 & n8053;
  assign n8068 = ~n8066 & ~n8067;
  assign n8069 = pi0072 & pi0993;
  assign n8070 = n2576 & n8069;
  assign n8071 = n2598 & n8053;
  assign n8072 = ~n8070 & ~n8071;
  assign n8073 = n8068 & n8072;
  assign n8074 = pi0072 & n4006;
  assign n8075 = pi0072 & ~n4014;
  assign n8076 = n3110 & n8053;
  assign n8077 = ~n8075 & ~n8076;
  assign n8078 = pi0072 & po0740;
  assign n8079 = n2651 & n8078;
  assign n8080 = ~n3102 & n8079;
  assign n8081 = n8077 & ~n8080;
  assign n8082 = ~n8074 & n8081;
  assign n8083 = n2591 & n8053;
  assign n8084 = n8082 & ~n8083;
  assign n8085 = pi1044 & n8065;
  assign n8086 = n2619 & n8085;
  assign n8087 = n2644 & n8051;
  assign n8088 = ~n8086 & ~n8087;
  assign n8089 = n2917 & n8051;
  assign n8090 = n2913 & n8053;
  assign n8091 = ~n8089 & ~n8090;
  assign n8092 = n2936 & n8065;
  assign n8093 = n8091 & ~n8092;
  assign n8094 = pi0072 & n4043;
  assign n8095 = n2930 & n8094;
  assign n8096 = pi0072 & ~n3553;
  assign n8097 = n4497 & n8096;
  assign n8098 = ~n8095 & ~n8097;
  assign n8099 = ~n4402 & n8065;
  assign n8100 = n8098 & ~n8099;
  assign n8101 = n3042 & n8053;
  assign n8102 = pi0072 & n4504;
  assign n8103 = ~n8101 & ~n8102;
  assign n8104 = n8100 & n8103;
  assign n8105 = n8093 & n8104;
  assign n8106 = n3033 & n8053;
  assign n8107 = n8105 & ~n8106;
  assign n8108 = n2910 & n8053;
  assign n8109 = pi0072 & n2726;
  assign n8110 = n4066 & n8109;
  assign n8111 = ~n8108 & ~n8110;
  assign n8112 = n8107 & n8111;
  assign n8113 = n8088 & n8112;
  assign n8114 = n8084 & n8113;
  assign n8115 = n8073 & n8114;
  assign n8116 = n8064 & n8115;
  assign n8117 = ~n8048 & n8116;
  assign n8118 = pi0072 & n4091;
  assign n8119 = pi0072 & n4459;
  assign n8120 = ~n4097 & n8078;
  assign n8121 = ~n3469 & ~n8120;
  assign n8122 = ~n8119 & n8121;
  assign n8123 = n3397 & ~n8122;
  assign n8124 = pi0072 & ~pi0786;
  assign n8125 = n4088 & n8124;
  assign n8126 = ~n8123 & ~n8125;
  assign n8127 = ~n8118 & n8126;
  assign n8128 = n4087 & ~n8127;
  assign n8129 = n3057 & n8053;
  assign n8130 = pi0072 & ~n3057;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = n4083 & ~n8131;
  assign n8133 = n2901 & n8065;
  assign n8134 = ~n8132 & ~n8133;
  assign n8135 = ~n3072 & n8053;
  assign n8136 = n2847 & n8051;
  assign n8137 = n2834 & n8085;
  assign n8138 = ~n8136 & ~n8137;
  assign n8139 = n2858 & n8051;
  assign n8140 = pi0072 & n4124;
  assign n8141 = n2854 & n8053;
  assign n8142 = n2881 & n8109;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~po0740 & n2881;
  assign n8145 = n2726 & n8144;
  assign n8146 = n8143 & ~n8145;
  assign n8147 = ~n8140 & n8146;
  assign n8148 = ~n8139 & n8147;
  assign n8149 = ~n4133 & n8051;
  assign n8150 = n8148 & ~n8149;
  assign n8151 = n2851 & n8065;
  assign n8152 = n3066 & n8053;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = n8150 & n8153;
  assign n8155 = n8138 & n8154;
  assign n8156 = ~n8135 & n8155;
  assign n8157 = n2681 & n8053;
  assign n8158 = ~n4077 & n8051;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = n8156 & n8159;
  assign n8161 = n8134 & n8160;
  assign n8162 = ~n8128 & n8161;
  assign po0230 = ~n8117 | ~n8162;
  assign n8164 = pi0073 & n4336;
  assign n8165 = pi0073 & n2741;
  assign n8166 = pi0073 & n4523;
  assign n8167 = ~n3973 & n8166;
  assign n8168 = pi0073 & pi0841;
  assign n8169 = ~n3998 & n8168;
  assign n8170 = pi0024 & pi0073;
  assign n8171 = pi0073 & n3989;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = n2563 & ~n8172;
  assign n8174 = n2795 & n8170;
  assign n8175 = ~n8173 & ~n8174;
  assign n8176 = ~n8169 & n8175;
  assign n8177 = ~n8167 & n8176;
  assign n8178 = ~n8165 & n8177;
  assign n8179 = pi0073 & ~n4061;
  assign n8180 = n4060 & n8179;
  assign n8181 = n8178 & ~n8180;
  assign n8182 = pi0073 & ~pi0314;
  assign n8183 = ~n4105 & n8182;
  assign n8184 = n2569 & n8170;
  assign n8185 = ~n8183 & ~n8184;
  assign n8186 = pi0073 & pi0993;
  assign n8187 = n2576 & n8186;
  assign n8188 = n2598 & n8170;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = n8185 & n8189;
  assign n8191 = pi0073 & n4067;
  assign n8192 = n2917 & n8168;
  assign n8193 = n2913 & n8170;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = n2936 & n8182;
  assign n8196 = n8194 & ~n8195;
  assign n8197 = pi0073 & n4043;
  assign n8198 = n2930 & n8197;
  assign n8199 = pi0073 & ~n3553;
  assign n8200 = n4497 & n8199;
  assign n8201 = ~n8198 & ~n8200;
  assign n8202 = ~n4402 & n8182;
  assign n8203 = n8201 & ~n8202;
  assign n8204 = n3042 & n8170;
  assign n8205 = pi0073 & n4504;
  assign n8206 = ~n8204 & ~n8205;
  assign n8207 = n8203 & n8206;
  assign n8208 = n8196 & n8207;
  assign n8209 = n3033 & n8170;
  assign n8210 = n8208 & ~n8209;
  assign n8211 = n2910 & n8170;
  assign n8212 = n8210 & ~n8211;
  assign n8213 = ~n8191 & n8212;
  assign n8214 = pi0073 & ~n4014;
  assign n8215 = n3110 & n8170;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = pi0073 & po0740;
  assign n8218 = n2651 & n8217;
  assign n8219 = ~n3102 & n8218;
  assign n8220 = pi0073 & n4006;
  assign n8221 = ~n8219 & ~n8220;
  assign n8222 = pi1044 & n8182;
  assign n8223 = n2619 & n8222;
  assign n8224 = n2644 & n8168;
  assign n8225 = ~n8223 & ~n8224;
  assign n8226 = n2591 & n8170;
  assign n8227 = n8225 & ~n8226;
  assign n8228 = n8221 & n8227;
  assign n8229 = n8216 & n8228;
  assign n8230 = n8213 & n8229;
  assign n8231 = n8190 & n8230;
  assign n8232 = n8181 & n8231;
  assign n8233 = ~n8164 & n8232;
  assign n8234 = pi0073 & n4091;
  assign n8235 = pi0073 & n4459;
  assign n8236 = n3398 & n3468;
  assign n8237 = ~n4097 & n8217;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~n8235 & n8238;
  assign n8240 = n3397 & ~n8239;
  assign n8241 = pi0073 & ~pi0786;
  assign n8242 = n4088 & n8241;
  assign n8243 = ~n8240 & ~n8242;
  assign n8244 = ~n8234 & n8243;
  assign n8245 = n4087 & ~n8244;
  assign n8246 = n3057 & n8170;
  assign n8247 = pi0073 & ~n3057;
  assign n8248 = ~n8246 & ~n8247;
  assign n8249 = n4083 & ~n8248;
  assign n8250 = n2901 & n8182;
  assign n8251 = ~n8249 & ~n8250;
  assign n8252 = ~n3072 & n8170;
  assign n8253 = n2847 & n8168;
  assign n8254 = n2834 & n8222;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = n2858 & n8168;
  assign n8257 = pi0073 & n4124;
  assign n8258 = n2854 & n8170;
  assign n8259 = n2881 & n8217;
  assign n8260 = n2726 & n8259;
  assign n8261 = ~n8258 & ~n8260;
  assign n8262 = ~n8257 & n8261;
  assign n8263 = ~n8256 & n8262;
  assign n8264 = ~n4133 & n8168;
  assign n8265 = n8263 & ~n8264;
  assign n8266 = n2851 & n8182;
  assign n8267 = n3066 & n8170;
  assign n8268 = ~n8266 & ~n8267;
  assign n8269 = n8265 & n8268;
  assign n8270 = n8255 & n8269;
  assign n8271 = ~n8252 & n8270;
  assign n8272 = n2681 & n8170;
  assign n8273 = ~n4077 & n8168;
  assign n8274 = ~n8272 & ~n8273;
  assign n8275 = n8271 & n8274;
  assign n8276 = n8251 & n8275;
  assign n8277 = ~n8245 & n8276;
  assign po0231 = ~n8233 | ~n8277;
  assign n8279 = pi0024 & pi0074;
  assign n8280 = ~n3072 & n8279;
  assign n8281 = pi0074 & pi0841;
  assign n8282 = n2847 & n8281;
  assign n8283 = pi0074 & ~pi0314;
  assign n8284 = pi1044 & n8283;
  assign n8285 = n2834 & n8284;
  assign n8286 = ~n8282 & ~n8285;
  assign n8287 = n2851 & n8283;
  assign n8288 = n3066 & n8279;
  assign n8289 = ~n8287 & ~n8288;
  assign n8290 = ~pi0074 & pi0479;
  assign n8291 = ~po0840 & ~n8290;
  assign n8292 = ~pi0841 & n8291;
  assign n8293 = ~n8281 & ~n8292;
  assign n8294 = n2858 & ~n8293;
  assign n8295 = pi0074 & po0740;
  assign n8296 = n2881 & n8295;
  assign n8297 = n2726 & n8296;
  assign n8298 = n2854 & n8279;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = ~n8294 & n8299;
  assign n8301 = n8289 & n8300;
  assign n8302 = n8286 & n8301;
  assign n8303 = ~n8280 & n8302;
  assign n8304 = n3057 & n8279;
  assign n8305 = pi0074 & ~n3057;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = n4083 & ~n8306;
  assign n8308 = n2901 & n8283;
  assign n8309 = ~n8307 & ~n8308;
  assign n8310 = n2681 & n8279;
  assign n8311 = ~n4077 & n8281;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = pi0074 & n4089;
  assign n8314 = pi0074 & n4091;
  assign n8315 = pi0074 & n3128;
  assign n8316 = ~n4094 & n8315;
  assign n8317 = ~n4097 & n8295;
  assign n8318 = ~n8316 & ~n8317;
  assign n8319 = n3397 & ~n8318;
  assign n8320 = ~n8314 & ~n8319;
  assign n8321 = ~n8313 & n8320;
  assign n8322 = n4087 & ~n8321;
  assign n8323 = n8312 & ~n8322;
  assign n8324 = n8309 & n8323;
  assign n8325 = n8303 & n8324;
  assign n8326 = n2651 & ~n3102;
  assign n8327 = ~n3018 & n8290;
  assign n8328 = ~po0740 & ~n8327;
  assign n8329 = ~n8295 & ~n8328;
  assign n8330 = n8326 & ~n8329;
  assign n8331 = n3110 & n8279;
  assign n8332 = ~n8330 & ~n8331;
  assign n8333 = pi0074 & ~n4014;
  assign n8334 = n8332 & ~n8333;
  assign n8335 = n2591 & n8279;
  assign n8336 = n8334 & ~n8335;
  assign n8337 = n2619 & n8284;
  assign n8338 = n2644 & n8281;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = n2917 & n8281;
  assign n8341 = n2913 & n8279;
  assign n8342 = ~n8340 & ~n8341;
  assign n8343 = n2936 & n8283;
  assign n8344 = n8342 & ~n8343;
  assign n8345 = pi0074 & n4043;
  assign n8346 = n2930 & n8345;
  assign n8347 = pi0074 & ~n3553;
  assign n8348 = n4497 & n8347;
  assign n8349 = ~n8346 & ~n8348;
  assign n8350 = ~n4402 & n8283;
  assign n8351 = n8349 & ~n8350;
  assign n8352 = n3042 & n8279;
  assign n8353 = pi0074 & n4504;
  assign n8354 = ~n8352 & ~n8353;
  assign n8355 = n8351 & n8354;
  assign n8356 = n8344 & n8355;
  assign n8357 = n3033 & n8279;
  assign n8358 = n8356 & ~n8357;
  assign n8359 = n2910 & n8279;
  assign n8360 = pi0074 & n2726;
  assign n8361 = n4066 & n8360;
  assign n8362 = ~n8359 & ~n8361;
  assign n8363 = n8358 & n8362;
  assign n8364 = n8339 & n8363;
  assign n8365 = n8336 & n8364;
  assign n8366 = pi0074 & n4523;
  assign n8367 = ~n3973 & n8366;
  assign n8368 = pi0074 & n3989;
  assign n8369 = ~n8279 & ~n8368;
  assign n8370 = n2563 & ~n8369;
  assign n8371 = n2795 & n8279;
  assign n8372 = ~n8370 & ~n8371;
  assign n8373 = pi0074 & n2741;
  assign n8374 = n8372 & ~n8373;
  assign n8375 = ~n8367 & n8374;
  assign n8376 = ~n3998 & n8281;
  assign n8377 = n8375 & ~n8376;
  assign n8378 = pi0074 & n4336;
  assign n8379 = pi0074 & n4062;
  assign n8380 = ~n8378 & ~n8379;
  assign n8381 = n8377 & n8380;
  assign n8382 = n8365 & n8381;
  assign n8383 = pi0074 & n4579;
  assign n8384 = ~n4105 & n8283;
  assign n8385 = n2569 & n8279;
  assign n8386 = ~n8384 & ~n8385;
  assign n8387 = n2598 & n8279;
  assign n8388 = n8386 & ~n8387;
  assign n8389 = ~n8383 & n8388;
  assign n8390 = ~n4133 & n8281;
  assign n8391 = n8389 & ~n8390;
  assign n8392 = n8382 & n8391;
  assign po0232 = ~n8325 | ~n8392;
  assign n8394 = pi0075 & pi0993;
  assign n8395 = n2576 & n8394;
  assign n8396 = pi0024 & pi0075;
  assign n8397 = n2598 & n8396;
  assign n8398 = ~n8395 & ~n8397;
  assign n8399 = pi0075 & n4062;
  assign n8400 = pi0075 & ~pi0314;
  assign n8401 = pi1044 & n8400;
  assign n8402 = n2619 & n8401;
  assign n8403 = pi0075 & pi0841;
  assign n8404 = n2644 & n8403;
  assign n8405 = ~n8402 & ~n8404;
  assign n8406 = ~n8399 & n8405;
  assign n8407 = pi0075 & n4336;
  assign n8408 = n8406 & ~n8407;
  assign n8409 = n8398 & n8408;
  assign n8410 = ~n3072 & n8396;
  assign n8411 = n2847 & n8403;
  assign n8412 = n2834 & n8401;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = pi0075 & po0740;
  assign n8415 = n2881 & n8414;
  assign n8416 = n2726 & n8415;
  assign n8417 = n2854 & n8396;
  assign n8418 = ~n8416 & ~n8417;
  assign n8419 = pi0075 & pi0479;
  assign n8420 = ~po0840 & ~n8419;
  assign n8421 = ~pi0841 & ~n8420;
  assign n8422 = ~n8403 & ~n8421;
  assign n8423 = n2858 & ~n8422;
  assign n8424 = n8418 & ~n8423;
  assign n8425 = ~n4133 & n8403;
  assign n8426 = n8424 & ~n8425;
  assign n8427 = n2851 & n8400;
  assign n8428 = n3066 & n8396;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = n8426 & n8429;
  assign n8431 = n8413 & n8430;
  assign n8432 = ~n8410 & n8431;
  assign n8433 = n8409 & n8432;
  assign n8434 = n3057 & n8396;
  assign n8435 = pi0075 & ~n3057;
  assign n8436 = ~n8434 & ~n8435;
  assign n8437 = n4083 & ~n8436;
  assign n8438 = n2901 & n8400;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = n2681 & n8396;
  assign n8441 = ~n4077 & n8403;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = pi0075 & n4089;
  assign n8444 = pi0075 & n4091;
  assign n8445 = pi0075 & n3128;
  assign n8446 = ~n4094 & n8445;
  assign n8447 = ~n4097 & n8414;
  assign n8448 = ~n8446 & ~n8447;
  assign n8449 = n3397 & ~n8448;
  assign n8450 = ~n8444 & ~n8449;
  assign n8451 = ~n8443 & n8450;
  assign n8452 = n4087 & ~n8451;
  assign n8453 = n8442 & ~n8452;
  assign n8454 = n8439 & n8453;
  assign n8455 = pi0075 & n4708;
  assign n8456 = ~n3973 & n8455;
  assign n8457 = pi0075 & n3989;
  assign n8458 = ~n8396 & ~n8457;
  assign n8459 = n2563 & ~n8458;
  assign n8460 = n2795 & n8396;
  assign n8461 = ~n8459 & ~n8460;
  assign n8462 = pi0075 & n2741;
  assign n8463 = n8461 & ~n8462;
  assign n8464 = ~n8456 & n8463;
  assign n8465 = ~n3998 & n8403;
  assign n8466 = n8464 & ~n8465;
  assign n8467 = n8454 & n8466;
  assign n8468 = n2910 & n8396;
  assign n8469 = pi0075 & n2726;
  assign n8470 = n4066 & n8469;
  assign n8471 = ~n8468 & ~n8470;
  assign n8472 = n2651 & n3102;
  assign n8473 = pi0075 & ~n4014;
  assign n8474 = n3110 & n8396;
  assign n8475 = ~n8473 & ~n8474;
  assign n8476 = n4003 & n8419;
  assign n8477 = ~n8414 & ~n8476;
  assign n8478 = n2651 & ~n8477;
  assign n8479 = n8475 & ~n8478;
  assign n8480 = ~n8472 & n8479;
  assign n8481 = n2591 & n8396;
  assign n8482 = n8480 & ~n8481;
  assign n8483 = ~n4105 & n8400;
  assign n8484 = n2569 & n8396;
  assign n8485 = ~n8483 & ~n8484;
  assign n8486 = n2917 & n8403;
  assign n8487 = n2913 & n8396;
  assign n8488 = ~n8486 & ~n8487;
  assign n8489 = n2936 & n8400;
  assign n8490 = n8488 & ~n8489;
  assign n8491 = pi0075 & n4043;
  assign n8492 = n2930 & n8491;
  assign n8493 = pi0075 & ~n3553;
  assign n8494 = n4497 & n8493;
  assign n8495 = ~n8492 & ~n8494;
  assign n8496 = ~n4402 & n8400;
  assign n8497 = n8495 & ~n8496;
  assign n8498 = n3042 & n8396;
  assign n8499 = pi0075 & n4504;
  assign n8500 = ~n8498 & ~n8499;
  assign n8501 = n8497 & n8500;
  assign n8502 = n8490 & n8501;
  assign n8503 = n3033 & n8396;
  assign n8504 = n8502 & ~n8503;
  assign n8505 = n8485 & n8504;
  assign n8506 = n8482 & n8505;
  assign n8507 = n8471 & n8506;
  assign n8508 = n8467 & n8507;
  assign po0233 = ~n8433 | ~n8508;
  assign n8510 = pi0076 & ~pi0314;
  assign n8511 = pi1044 & n8510;
  assign n8512 = n2619 & n8511;
  assign n8513 = pi0076 & pi0841;
  assign n8514 = n2644 & n8513;
  assign n8515 = ~n8512 & ~n8514;
  assign n8516 = pi0076 & pi0993;
  assign n8517 = n2576 & n8516;
  assign n8518 = pi0024 & pi0076;
  assign n8519 = n2598 & n8518;
  assign n8520 = ~n8517 & ~n8519;
  assign n8521 = pi0076 & n4336;
  assign n8522 = ~pi0076 & n3540;
  assign n8523 = n2813 & ~n8522;
  assign n8524 = ~n4058 & n8523;
  assign n8525 = ~n4061 & n8524;
  assign n8526 = ~n8521 & ~n8525;
  assign n8527 = n8520 & n8526;
  assign n8528 = n8515 & n8527;
  assign n8529 = n3057 & n8518;
  assign n8530 = pi0076 & ~n3057;
  assign n8531 = ~n8529 & ~n8530;
  assign n8532 = n4083 & ~n8531;
  assign n8533 = n2901 & n8510;
  assign n8534 = ~n8532 & ~n8533;
  assign n8535 = pi0076 & n4089;
  assign n8536 = pi0076 & n4091;
  assign n8537 = pi0076 & n3128;
  assign n8538 = ~n4094 & n8537;
  assign n8539 = pi0076 & po0740;
  assign n8540 = ~n4097 & n8539;
  assign n8541 = ~n8538 & ~n8540;
  assign n8542 = n3397 & ~n8541;
  assign n8543 = ~n8536 & ~n8542;
  assign n8544 = ~n8535 & n8543;
  assign n8545 = n4087 & ~n8544;
  assign n8546 = pi0076 & n4006;
  assign n8547 = pi0076 & ~n4014;
  assign n8548 = n3110 & n8518;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = n2651 & n8539;
  assign n8551 = ~n3102 & n8550;
  assign n8552 = n8549 & ~n8551;
  assign n8553 = ~n8546 & n8552;
  assign n8554 = n2591 & n8518;
  assign n8555 = n8553 & ~n8554;
  assign n8556 = n2910 & n8518;
  assign n8557 = pi0076 & n2726;
  assign n8558 = n4066 & n8557;
  assign n8559 = ~n8556 & ~n8558;
  assign n8560 = n8555 & n8559;
  assign n8561 = n2917 & n8513;
  assign n8562 = n2913 & n8518;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = n2936 & n8510;
  assign n8565 = n8563 & ~n8564;
  assign n8566 = pi0076 & n4043;
  assign n8567 = n2930 & n8566;
  assign n8568 = pi0076 & ~n3553;
  assign n8569 = n4497 & n8568;
  assign n8570 = ~n8567 & ~n8569;
  assign n8571 = ~n4402 & n8510;
  assign n8572 = n8570 & ~n8571;
  assign n8573 = n3042 & n8518;
  assign n8574 = pi0076 & n4504;
  assign n8575 = ~n8573 & ~n8574;
  assign n8576 = n8572 & n8575;
  assign n8577 = n8565 & n8576;
  assign n8578 = n3033 & n8518;
  assign n8579 = n8577 & ~n8578;
  assign n8580 = n8560 & n8579;
  assign n8581 = ~n8545 & n8580;
  assign n8582 = n8534 & n8581;
  assign n8583 = n8528 & n8582;
  assign n8584 = n2681 & n8518;
  assign n8585 = ~n4077 & n8513;
  assign n8586 = ~n8584 & ~n8585;
  assign n8587 = ~n4105 & n8510;
  assign n8588 = n2569 & n8518;
  assign n8589 = ~n8587 & ~n8588;
  assign n8590 = n8586 & n8589;
  assign n8591 = n2847 & n8513;
  assign n8592 = n2834 & n8511;
  assign n8593 = ~n8591 & ~n8592;
  assign n8594 = n2851 & n8510;
  assign n8595 = n3066 & n8518;
  assign n8596 = ~n8594 & ~n8595;
  assign n8597 = ~n3072 & n8518;
  assign n8598 = n8596 & ~n8597;
  assign n8599 = n8593 & n8598;
  assign n8600 = n8590 & n8599;
  assign n8601 = n2858 & n8513;
  assign n8602 = pi0076 & n4124;
  assign n8603 = n2854 & n8518;
  assign n8604 = n2881 & n8539;
  assign n8605 = n2726 & n8604;
  assign n8606 = ~n8603 & ~n8605;
  assign n8607 = ~n8602 & n8606;
  assign n8608 = ~n8601 & n8607;
  assign n8609 = ~n4133 & n8513;
  assign n8610 = n8608 & ~n8609;
  assign n8611 = pi0076 & n4708;
  assign n8612 = ~n3973 & n8611;
  assign n8613 = pi0076 & n3989;
  assign n8614 = ~n8518 & ~n8613;
  assign n8615 = n2563 & ~n8614;
  assign n8616 = n2795 & n8518;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = pi0076 & n2741;
  assign n8619 = n8617 & ~n8618;
  assign n8620 = ~n8612 & n8619;
  assign n8621 = ~n3998 & n8513;
  assign n8622 = n8620 & ~n8621;
  assign n8623 = n8610 & n8622;
  assign n8624 = n8600 & n8623;
  assign po0234 = ~n8583 | ~n8624;
  assign n8626 = pi0077 & n4585;
  assign n8627 = pi0024 & pi0077;
  assign n8628 = pi0077 & n3989;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = n2563 & ~n8629;
  assign n8631 = n2795 & n8627;
  assign n8632 = ~n8630 & ~n8631;
  assign n8633 = pi0077 & n2741;
  assign n8634 = n8632 & ~n8633;
  assign n8635 = ~n8626 & n8634;
  assign n8636 = pi0077 & pi0841;
  assign n8637 = ~n3998 & n8636;
  assign n8638 = n8635 & ~n8637;
  assign n8639 = pi0077 & n4062;
  assign n8640 = n2569 & n8627;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = pi0077 & ~pi0314;
  assign n8643 = ~n4105 & n8642;
  assign n8644 = n8641 & ~n8643;
  assign n8645 = pi0077 & n4336;
  assign n8646 = n8644 & ~n8645;
  assign n8647 = n8638 & n8646;
  assign n8648 = ~n3072 & n8627;
  assign n8649 = n2847 & n8636;
  assign n8650 = pi1044 & n8642;
  assign n8651 = n2834 & n8650;
  assign n8652 = ~n8649 & ~n8651;
  assign n8653 = n2858 & n8636;
  assign n8654 = pi0077 & n4124;
  assign n8655 = n2854 & n8627;
  assign n8656 = pi0077 & po0740;
  assign n8657 = n2881 & n8656;
  assign n8658 = n2726 & n8657;
  assign n8659 = ~n8655 & ~n8658;
  assign n8660 = ~n8654 & n8659;
  assign n8661 = ~n8653 & n8660;
  assign n8662 = ~n4133 & n8636;
  assign n8663 = n8661 & ~n8662;
  assign n8664 = n2851 & n8642;
  assign n8665 = n3066 & n8627;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = n8663 & n8666;
  assign n8668 = n8652 & n8667;
  assign n8669 = ~n8648 & n8668;
  assign n8670 = n3057 & n8627;
  assign n8671 = pi0077 & ~n3057;
  assign n8672 = ~n8670 & ~n8671;
  assign n8673 = n4083 & ~n8672;
  assign n8674 = n2901 & n8642;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = n2681 & n8627;
  assign n8677 = ~n4077 & n8636;
  assign n8678 = ~n8676 & ~n8677;
  assign n8679 = pi0077 & n4089;
  assign n8680 = pi0077 & n4091;
  assign n8681 = ~n4097 & n8656;
  assign n8682 = pi0077 & n3128;
  assign n8683 = ~n4094 & n8682;
  assign n8684 = ~n8681 & ~n8683;
  assign n8685 = n3397 & ~n8684;
  assign n8686 = ~n8680 & ~n8685;
  assign n8687 = ~n8679 & n8686;
  assign n8688 = n4087 & ~n8687;
  assign n8689 = n8678 & ~n8688;
  assign n8690 = n8675 & n8689;
  assign n8691 = pi0077 & ~n4014;
  assign n8692 = n3110 & n8627;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = ~n3102 & n8656;
  assign n8695 = n2651 & n8694;
  assign n8696 = pi0077 & ~n3102;
  assign n8697 = n4005 & n8696;
  assign n8698 = ~n8695 & ~n8697;
  assign n8699 = n8693 & n8698;
  assign n8700 = n2619 & n8650;
  assign n8701 = n2644 & n8636;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = pi0077 & pi0993;
  assign n8704 = n2576 & n8703;
  assign n8705 = n2598 & n8627;
  assign n8706 = ~n8704 & ~n8705;
  assign n8707 = n2910 & n8627;
  assign n8708 = pi0077 & n4067;
  assign n8709 = pi0077 & n5491;
  assign n8710 = pi0077 & ~n3553;
  assign n8711 = n4497 & n8710;
  assign n8712 = n2917 & n8636;
  assign n8713 = n2913 & n8627;
  assign n8714 = ~n8712 & ~n8713;
  assign n8715 = n2936 & n8642;
  assign n8716 = n8714 & ~n8715;
  assign n8717 = ~n4402 & n8642;
  assign n8718 = n8716 & ~n8717;
  assign n8719 = ~n8711 & n8718;
  assign n8720 = ~n8709 & n8719;
  assign n8721 = ~n2941 & n8720;
  assign n8722 = pi0077 & n4504;
  assign n8723 = n3042 & n8627;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = n3033 & n8627;
  assign n8726 = n8724 & ~n8725;
  assign n8727 = n8721 & n8726;
  assign n8728 = ~n8708 & n8727;
  assign n8729 = ~n8707 & n8728;
  assign n8730 = n2591 & n8627;
  assign n8731 = n8729 & ~n8730;
  assign n8732 = n8706 & n8731;
  assign n8733 = n8702 & n8732;
  assign n8734 = n8699 & n8733;
  assign n8735 = n8690 & n8734;
  assign n8736 = n8669 & n8735;
  assign po0235 = ~n8647 | ~n8736;
  assign n8738 = pi0232 & ~pi0468;
  assign po0236 = pi0119 & n8738;
  assign n8740 = ~pi0179 & n2429;
  assign n8741 = ~pi0156 & ~n2429;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = ~n4152 & n8742;
  assign n8744 = ~n4162 & ~n4922;
  assign n8745 = ~pi0184 & n2429;
  assign n8746 = ~pi0163 & ~n2429;
  assign n8747 = ~n8745 & ~n8746;
  assign n8748 = n3481 & n8747;
  assign n8749 = ~n4182 & ~n8748;
  assign n8750 = ~n3491 & n4213;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~pi0074 & ~n3463;
  assign n8753 = n4182 & n8752;
  assign n8754 = ~pi0187 & n2429;
  assign n8755 = ~pi0147 & ~n2429;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = n3481 & n8756;
  assign n8758 = ~n4186 & ~n8757;
  assign n8759 = ~pi0040 & n4186;
  assign n8760 = ~pi0079 & n4247;
  assign n8761 = pi0079 & ~n4247;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = n4194 & ~n8762;
  assign n8764 = pi0079 & ~n4194;
  assign n8765 = ~n8763 & ~n8764;
  assign n8766 = n2452 & n8765;
  assign n8767 = n8759 & ~n8766;
  assign n8768 = ~n8758 & ~n8767;
  assign n8769 = n8753 & ~n8768;
  assign n8770 = n8751 & ~n8769;
  assign n8771 = n4163 & ~n8770;
  assign n8772 = ~n4166 & ~n4170;
  assign n8773 = n3481 & ~n8772;
  assign n8774 = ~n4240 & ~n8773;
  assign n8775 = ~n4239 & ~n8774;
  assign n8776 = n8748 & ~n8775;
  assign n8777 = ~n8748 & n8775;
  assign n8778 = ~n8776 & ~n8777;
  assign n8779 = ~n4163 & ~n8778;
  assign n8780 = ~n8771 & ~n8779;
  assign n8781 = n4162 & ~n8780;
  assign n8782 = ~n8744 & ~n8781;
  assign n8783 = n4155 & n8782;
  assign n8784 = n2444 & ~n4155;
  assign n8785 = ~n8783 & ~n8784;
  assign n8786 = n4152 & ~n4224;
  assign n8787 = ~n8785 & n8786;
  assign n8788 = ~n8743 & ~n8787;
  assign po0237 = n4228 | n8788;
  assign n8790 = ~pi0080 & n3539;
  assign po0238 = ~n3958 & n8790;
  assign n8792 = pi0081 & pi0841;
  assign n8793 = ~n3998 & n8792;
  assign n8794 = pi0081 & ~pi0314;
  assign n8795 = pi1044 & n8794;
  assign n8796 = n2619 & n8795;
  assign n8797 = n2644 & n8792;
  assign n8798 = ~n8796 & ~n8797;
  assign n8799 = n2851 & n8794;
  assign n8800 = pi0024 & pi0081;
  assign n8801 = n3066 & n8800;
  assign n8802 = ~n8799 & ~n8801;
  assign n8803 = ~n4105 & n8794;
  assign n8804 = n2569 & n8800;
  assign n8805 = ~n8803 & ~n8804;
  assign n8806 = n2598 & n8800;
  assign n8807 = n8805 & ~n8806;
  assign n8808 = n8802 & n8807;
  assign n8809 = ~n2878 & n8808;
  assign n8810 = pi0081 & n4060;
  assign n8811 = ~n4061 & n8810;
  assign n8812 = n8809 & ~n8811;
  assign n8813 = n8798 & n8812;
  assign n8814 = ~n8793 & n8813;
  assign n8815 = pi0081 & n2604;
  assign n8816 = n3967 & n8815;
  assign n8817 = n8814 & ~n8816;
  assign n8818 = pi0081 & n4708;
  assign n8819 = ~n3973 & n8818;
  assign n8820 = pi0081 & n3989;
  assign n8821 = ~n8800 & ~n8820;
  assign n8822 = n2563 & ~n8821;
  assign n8823 = n2795 & n8800;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = pi0081 & n2741;
  assign n8826 = n8824 & ~n8825;
  assign n8827 = ~n8819 & n8826;
  assign n8828 = ~n4077 & n8792;
  assign n8829 = n2681 & n8800;
  assign n8830 = ~n8828 & ~n8829;
  assign n8831 = pi0081 & n4091;
  assign n8832 = pi0081 & po0740;
  assign n8833 = ~n4097 & n8832;
  assign n8834 = pi0081 & n4459;
  assign n8835 = ~n8833 & ~n8834;
  assign n8836 = n3397 & ~n8835;
  assign n8837 = pi0081 & ~pi0786;
  assign n8838 = n4088 & n8837;
  assign n8839 = ~n8836 & ~n8838;
  assign n8840 = ~n8831 & n8839;
  assign n8841 = n4087 & ~n8840;
  assign n8842 = n2901 & n8794;
  assign n8843 = n3057 & n8800;
  assign n8844 = pi0081 & ~n3057;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = n4083 & ~n8845;
  assign n8847 = ~n8842 & ~n8846;
  assign n8848 = ~n8841 & n8847;
  assign n8849 = n8830 & n8848;
  assign n8850 = n8827 & n8849;
  assign n8851 = n2910 & n8800;
  assign n8852 = pi0081 & n2726;
  assign n8853 = n4066 & n8852;
  assign n8854 = ~n8851 & ~n8853;
  assign n8855 = pi0081 & n4579;
  assign n8856 = n2858 & n8792;
  assign n8857 = pi0081 & n4124;
  assign n8858 = n2854 & n8800;
  assign n8859 = n2881 & n8832;
  assign n8860 = n2726 & n8859;
  assign n8861 = ~n8858 & ~n8860;
  assign n8862 = ~n8857 & n8861;
  assign n8863 = ~n8856 & n8862;
  assign n8864 = ~n3072 & n8800;
  assign n8865 = n8863 & ~n8864;
  assign n8866 = n2847 & n8792;
  assign n8867 = n2834 & n8795;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = n8865 & n8868;
  assign n8870 = ~n4133 & n8792;
  assign n8871 = n8869 & ~n8870;
  assign n8872 = pi0081 & n4006;
  assign n8873 = pi0081 & ~n4014;
  assign n8874 = n3110 & n8800;
  assign n8875 = ~n8873 & ~n8874;
  assign n8876 = n2651 & n8832;
  assign n8877 = ~n3102 & n8876;
  assign n8878 = n8875 & ~n8877;
  assign n8879 = ~n8872 & n8878;
  assign n8880 = n2591 & n8800;
  assign n8881 = n8879 & ~n8880;
  assign n8882 = n8871 & n8881;
  assign n8883 = ~n8855 & n8882;
  assign n8884 = n8854 & n8883;
  assign n8885 = n2917 & n8792;
  assign n8886 = n2913 & n8800;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = n2936 & n8794;
  assign n8889 = n8887 & ~n8888;
  assign n8890 = pi0081 & n4043;
  assign n8891 = n2930 & n8890;
  assign n8892 = pi0081 & ~n3553;
  assign n8893 = n4497 & n8892;
  assign n8894 = ~n8891 & ~n8893;
  assign n8895 = ~n4402 & n8794;
  assign n8896 = n8894 & ~n8895;
  assign n8897 = n3042 & n8800;
  assign n8898 = pi0081 & n4504;
  assign n8899 = ~n8897 & ~n8898;
  assign n8900 = n8896 & n8899;
  assign n8901 = n8889 & n8900;
  assign n8902 = n3033 & n8800;
  assign n8903 = n8901 & ~n8902;
  assign n8904 = n8884 & n8903;
  assign n8905 = n8850 & n8904;
  assign po0239 = ~n8817 | ~n8905;
  assign n8907 = pi0024 & pi0082;
  assign n8908 = n2913 & n8907;
  assign n8909 = pi0082 & pi0841;
  assign n8910 = n2917 & n8909;
  assign n8911 = ~n8908 & ~n8910;
  assign n8912 = pi0082 & n4336;
  assign n8913 = ~n3998 & n8909;
  assign n8914 = ~n8912 & ~n8913;
  assign n8915 = pi0082 & n4062;
  assign n8916 = n8914 & ~n8915;
  assign n8917 = n8911 & n8916;
  assign n8918 = ~n4077 & n8909;
  assign n8919 = n2681 & n8907;
  assign n8920 = ~n8918 & ~n8919;
  assign n8921 = pi0082 & n4091;
  assign n8922 = pi0082 & po0740;
  assign n8923 = ~n4097 & n8922;
  assign n8924 = pi0082 & n4459;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = n3397 & ~n8925;
  assign n8927 = pi0082 & ~pi0786;
  assign n8928 = n4088 & n8927;
  assign n8929 = ~n8926 & ~n8928;
  assign n8930 = ~n8921 & n8929;
  assign n8931 = n4087 & ~n8930;
  assign n8932 = pi0082 & ~pi0314;
  assign n8933 = n2901 & n8932;
  assign n8934 = n3057 & n8907;
  assign n8935 = pi0082 & ~n3057;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = n4083 & ~n8936;
  assign n8938 = ~n8933 & ~n8937;
  assign n8939 = ~n8931 & n8938;
  assign n8940 = n8920 & n8939;
  assign n8941 = n2858 & n8909;
  assign n8942 = pi0082 & n4124;
  assign n8943 = n2854 & n8907;
  assign n8944 = n2881 & n8922;
  assign n8945 = n2726 & n8944;
  assign n8946 = ~n8943 & ~n8945;
  assign n8947 = ~n8942 & n8946;
  assign n8948 = ~n8941 & n8947;
  assign n8949 = ~n3072 & n8907;
  assign n8950 = n8948 & ~n8949;
  assign n8951 = n2847 & n8909;
  assign n8952 = pi1044 & n8932;
  assign n8953 = n2834 & n8952;
  assign n8954 = ~n8951 & ~n8953;
  assign n8955 = n8950 & n8954;
  assign n8956 = ~n4133 & n8909;
  assign n8957 = n8955 & ~n8956;
  assign n8958 = pi0082 & n4708;
  assign n8959 = ~n3973 & n8958;
  assign n8960 = pi0082 & n3989;
  assign n8961 = ~n8907 & ~n8960;
  assign n8962 = n2563 & ~n8961;
  assign n8963 = n2795 & n8907;
  assign n8964 = ~n8962 & ~n8963;
  assign n8965 = pi0082 & n2741;
  assign n8966 = n8964 & ~n8965;
  assign n8967 = ~n8959 & n8966;
  assign n8968 = n8957 & n8967;
  assign n8969 = n8940 & n8968;
  assign n8970 = n8917 & n8969;
  assign n8971 = pi0082 & n4504;
  assign n8972 = n2619 & n8952;
  assign n8973 = n3042 & n8907;
  assign n8974 = pi0082 & n2726;
  assign n8975 = n4066 & n8974;
  assign n8976 = n2591 & n8907;
  assign n8977 = ~n8975 & ~n8976;
  assign n8978 = n2644 & n8909;
  assign n8979 = n8977 & ~n8978;
  assign n8980 = ~n8973 & n8979;
  assign n8981 = ~n8972 & n8980;
  assign n8982 = ~n8971 & n8981;
  assign n8983 = n2910 & n8907;
  assign n8984 = pi0082 & n4006;
  assign n8985 = pi0082 & ~n4014;
  assign n8986 = n3110 & n8907;
  assign n8987 = ~n8985 & ~n8986;
  assign n8988 = n2651 & n8922;
  assign n8989 = ~n3102 & n8988;
  assign n8990 = n8987 & ~n8989;
  assign n8991 = ~n8984 & n8990;
  assign n8992 = ~n8983 & n8991;
  assign n8993 = n8982 & n8992;
  assign n8994 = n2598 & n8907;
  assign n8995 = ~n4105 & n8932;
  assign n8996 = n2569 & n8907;
  assign n8997 = ~n8995 & ~n8996;
  assign n8998 = n2851 & n8932;
  assign n8999 = n3066 & n8907;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = n8997 & n9000;
  assign n9002 = ~n8994 & n9001;
  assign n9003 = ~n2872 & n9002;
  assign n9004 = n3033 & n8907;
  assign n9005 = pi0082 & ~n3553;
  assign n9006 = n4497 & n9005;
  assign n9007 = ~pi0082 & ~pi0314;
  assign n9008 = n2936 & ~n9007;
  assign n9009 = n2533 & n8932;
  assign n9010 = ~n9008 & ~n9009;
  assign n9011 = pi0082 & n5491;
  assign n9012 = n9010 & ~n9011;
  assign n9013 = ~n9006 & n9012;
  assign n9014 = n2544 & n8932;
  assign n9015 = n9013 & ~n9014;
  assign n9016 = pi0082 & n4579;
  assign n9017 = n9015 & ~n9016;
  assign n9018 = ~n9004 & n9017;
  assign n9019 = n9003 & n9018;
  assign n9020 = n8993 & n9019;
  assign po0240 = ~n8970 | ~n9020;
  assign n9022 = pi0083 & n4067;
  assign n9023 = pi0083 & pi0841;
  assign n9024 = n2917 & n9023;
  assign n9025 = pi0024 & pi0083;
  assign n9026 = n2913 & n9025;
  assign n9027 = ~n9024 & ~n9026;
  assign n9028 = pi0083 & ~pi0314;
  assign n9029 = n2936 & n9028;
  assign n9030 = n9027 & ~n9029;
  assign n9031 = n3042 & n9025;
  assign n9032 = pi0083 & n4043;
  assign n9033 = n2930 & n9032;
  assign n9034 = pi0083 & ~n3553;
  assign n9035 = n4497 & n9034;
  assign n9036 = ~n9033 & ~n9035;
  assign n9037 = ~n4402 & n9028;
  assign n9038 = n9036 & ~n9037;
  assign n9039 = pi0083 & n4504;
  assign n9040 = n9038 & ~n9039;
  assign n9041 = ~n9031 & n9040;
  assign n9042 = n9030 & n9041;
  assign n9043 = n3033 & n9025;
  assign n9044 = n9042 & ~n9043;
  assign n9045 = n2910 & n9025;
  assign n9046 = n9044 & ~n9045;
  assign n9047 = ~n9022 & n9046;
  assign n9048 = ~n4105 & n9028;
  assign n9049 = n2569 & n9025;
  assign n9050 = ~n9048 & ~n9049;
  assign n9051 = pi0083 & pi0993;
  assign n9052 = n2576 & n9051;
  assign n9053 = n2598 & n9025;
  assign n9054 = ~n9052 & ~n9053;
  assign n9055 = n9050 & n9054;
  assign n9056 = pi0083 & ~n4014;
  assign n9057 = n3110 & n9025;
  assign n9058 = ~n9056 & ~n9057;
  assign n9059 = pi0083 & po0740;
  assign n9060 = n2651 & n9059;
  assign n9061 = ~n3102 & n9060;
  assign n9062 = pi0083 & n4006;
  assign n9063 = ~n9061 & ~n9062;
  assign n9064 = pi1044 & n9028;
  assign n9065 = n2619 & n9064;
  assign n9066 = n2644 & n9023;
  assign n9067 = ~n9065 & ~n9066;
  assign n9068 = n2591 & n9025;
  assign n9069 = n9067 & ~n9068;
  assign n9070 = n9063 & n9069;
  assign n9071 = n9058 & n9070;
  assign n9072 = n9055 & n9071;
  assign n9073 = pi0083 & n3967;
  assign n9074 = n2604 & n9073;
  assign n9075 = pi0083 & ~n4061;
  assign n9076 = n4060 & n9075;
  assign n9077 = ~n9074 & ~n9076;
  assign n9078 = pi0083 & n2741;
  assign n9079 = ~n3998 & n9023;
  assign n9080 = pi0083 & n4708;
  assign n9081 = ~n3973 & n9080;
  assign n9082 = pi0083 & n3989;
  assign n9083 = ~n9025 & ~n9082;
  assign n9084 = n2563 & ~n9083;
  assign n9085 = n2795 & n9025;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = ~n9081 & n9086;
  assign n9088 = ~n9079 & n9087;
  assign n9089 = ~n9078 & n9088;
  assign n9090 = n9077 & n9089;
  assign n9091 = n9072 & n9090;
  assign n9092 = n9047 & n9091;
  assign n9093 = n2851 & n9028;
  assign n9094 = n3066 & n9025;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = ~n4077 & n9023;
  assign n9097 = n2681 & n9025;
  assign n9098 = ~n9096 & ~n9097;
  assign n9099 = pi0083 & n4091;
  assign n9100 = ~n4097 & n9059;
  assign n9101 = pi0083 & n4459;
  assign n9102 = ~n9100 & ~n9101;
  assign n9103 = n3397 & ~n9102;
  assign n9104 = pi0083 & ~pi0786;
  assign n9105 = n4088 & n9104;
  assign n9106 = ~n9103 & ~n9105;
  assign n9107 = ~n9099 & n9106;
  assign n9108 = n4087 & ~n9107;
  assign n9109 = n2901 & n9028;
  assign n9110 = n3057 & n9025;
  assign n9111 = pi0083 & ~n3057;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = n4083 & ~n9112;
  assign n9114 = ~n9109 & ~n9113;
  assign n9115 = ~n9108 & n9114;
  assign n9116 = n9098 & n9115;
  assign n9117 = n2858 & n9023;
  assign n9118 = pi0083 & n4124;
  assign n9119 = n2854 & n9025;
  assign n9120 = n2881 & n9059;
  assign n9121 = n2726 & n9120;
  assign n9122 = ~n9119 & ~n9121;
  assign n9123 = ~n9118 & n9122;
  assign n9124 = ~n9117 & n9123;
  assign n9125 = ~n3072 & n9025;
  assign n9126 = n9124 & ~n9125;
  assign n9127 = n2847 & n9023;
  assign n9128 = n2834 & n9064;
  assign n9129 = ~n9127 & ~n9128;
  assign n9130 = n9126 & n9129;
  assign n9131 = ~n4133 & n9023;
  assign n9132 = n9130 & ~n9131;
  assign n9133 = n9116 & n9132;
  assign n9134 = n9095 & n9133;
  assign n9135 = ~n2867 & n9134;
  assign po0241 = ~n9092 | ~n9135;
  assign n9137 = pi0084 & pi0993;
  assign n9138 = n2576 & n9137;
  assign n9139 = pi0024 & pi0084;
  assign n9140 = n2598 & n9139;
  assign n9141 = ~n9138 & ~n9140;
  assign n9142 = pi0084 & ~pi0314;
  assign n9143 = ~n4105 & n9142;
  assign n9144 = n2569 & n9139;
  assign n9145 = ~n9143 & ~n9144;
  assign n9146 = pi0084 & ~n4014;
  assign n9147 = n3110 & n9139;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = pi0084 & po0740;
  assign n9150 = n2651 & n9149;
  assign n9151 = ~n3102 & n9150;
  assign n9152 = pi0084 & n4006;
  assign n9153 = ~n9151 & ~n9152;
  assign n9154 = n9148 & n9153;
  assign n9155 = n9145 & n9154;
  assign n9156 = n9141 & n9155;
  assign n9157 = pi0084 & n2741;
  assign n9158 = pi0084 & n4708;
  assign n9159 = ~n3973 & n9158;
  assign n9160 = pi0084 & pi0841;
  assign n9161 = ~n3998 & n9160;
  assign n9162 = pi0084 & n3989;
  assign n9163 = ~n9139 & ~n9162;
  assign n9164 = n2563 & ~n9163;
  assign n9165 = n2795 & n9139;
  assign n9166 = ~n9164 & ~n9165;
  assign n9167 = ~n9161 & n9166;
  assign n9168 = ~n9159 & n9167;
  assign n9169 = ~n9157 & n9168;
  assign n9170 = n9156 & n9169;
  assign n9171 = n2591 & n9139;
  assign n9172 = pi1044 & n9142;
  assign n9173 = n2619 & n9172;
  assign n9174 = n2644 & n9160;
  assign n9175 = ~n9173 & ~n9174;
  assign n9176 = n2917 & n9160;
  assign n9177 = n2913 & n9139;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = n2936 & n9142;
  assign n9180 = n9178 & ~n9179;
  assign n9181 = pi0084 & n4043;
  assign n9182 = n2930 & n9181;
  assign n9183 = pi0084 & ~n3553;
  assign n9184 = n4497 & n9183;
  assign n9185 = ~n9182 & ~n9184;
  assign n9186 = ~n4402 & n9142;
  assign n9187 = n9185 & ~n9186;
  assign n9188 = n3042 & n9139;
  assign n9189 = pi0084 & n4504;
  assign n9190 = ~n9188 & ~n9189;
  assign n9191 = n9187 & n9190;
  assign n9192 = n9180 & n9191;
  assign n9193 = n3033 & n9139;
  assign n9194 = n9192 & ~n9193;
  assign n9195 = n2910 & n9139;
  assign n9196 = pi0084 & n4067;
  assign n9197 = ~n9195 & ~n9196;
  assign n9198 = n9194 & n9197;
  assign n9199 = n9175 & n9198;
  assign n9200 = ~n9171 & n9199;
  assign n9201 = pi0084 & ~n4061;
  assign n9202 = n4060 & n9201;
  assign n9203 = n9200 & ~n9202;
  assign n9204 = pi0084 & n2604;
  assign n9205 = n3967 & n9204;
  assign n9206 = n9203 & ~n9205;
  assign n9207 = n9170 & n9206;
  assign n9208 = pi0084 & n4091;
  assign n9209 = ~n4097 & n9149;
  assign n9210 = pi0084 & n4459;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = n3397 & ~n9211;
  assign n9213 = pi0084 & ~pi0786;
  assign n9214 = n4088 & n9213;
  assign n9215 = ~n9212 & ~n9214;
  assign n9216 = ~n9208 & n9215;
  assign n9217 = n3547 & ~n9216;
  assign n9218 = n3406 & n9217;
  assign n9219 = n3057 & n9139;
  assign n9220 = pi0084 & ~n3057;
  assign n9221 = ~n9219 & ~n9220;
  assign n9222 = n4083 & ~n9221;
  assign n9223 = ~n9218 & ~n9222;
  assign n9224 = pi0314 & n4983;
  assign n9225 = ~n9142 & ~n9224;
  assign n9226 = n2901 & ~n9225;
  assign n9227 = ~n3072 & n9139;
  assign n9228 = n2847 & n9160;
  assign n9229 = n2834 & n9172;
  assign n9230 = ~n9228 & ~n9229;
  assign n9231 = n2858 & n9160;
  assign n9232 = pi0084 & n4124;
  assign n9233 = n2854 & n9139;
  assign n9234 = n2881 & n9149;
  assign n9235 = n2726 & n9234;
  assign n9236 = ~n9233 & ~n9235;
  assign n9237 = ~n9232 & n9236;
  assign n9238 = ~n9231 & n9237;
  assign n9239 = ~n4133 & n9160;
  assign n9240 = n9238 & ~n9239;
  assign n9241 = n2851 & n9142;
  assign n9242 = n3066 & n9139;
  assign n9243 = ~n9241 & ~n9242;
  assign n9244 = n9240 & n9243;
  assign n9245 = n9230 & n9244;
  assign n9246 = ~n9227 & n9245;
  assign n9247 = n2681 & n9139;
  assign n9248 = ~n4077 & n9160;
  assign n9249 = ~n9247 & ~n9248;
  assign n9250 = n9246 & n9249;
  assign n9251 = ~n9226 & n9250;
  assign n9252 = n9223 & n9251;
  assign po0242 = ~n9207 | ~n9252;
  assign n9254 = pi0085 & n4336;
  assign n9255 = pi0085 & n2741;
  assign n9256 = pi0085 & n5965;
  assign n9257 = pi0085 & pi0841;
  assign n9258 = ~n3998 & n9257;
  assign n9259 = pi0024 & pi0085;
  assign n9260 = pi0085 & n3989;
  assign n9261 = ~n9259 & ~n9260;
  assign n9262 = n2563 & ~n9261;
  assign n9263 = n2795 & n9259;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = ~n9258 & n9264;
  assign n9266 = ~n9256 & n9265;
  assign n9267 = ~n9255 & n9266;
  assign n9268 = pi0085 & ~n4061;
  assign n9269 = n4060 & n9268;
  assign n9270 = n9267 & ~n9269;
  assign n9271 = pi0085 & n4067;
  assign n9272 = pi0085 & ~n3553;
  assign n9273 = n4497 & n9272;
  assign n9274 = n2917 & n9257;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = n2913 & n9259;
  assign n9277 = pi0085 & n4504;
  assign n9278 = n3042 & n9259;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = pi0085 & ~pi0314;
  assign n9281 = n2533 & n9280;
  assign n9282 = pi0085 & n4043;
  assign n9283 = n2930 & n9282;
  assign n9284 = ~n9281 & ~n9283;
  assign n9285 = ~n2527 & n9284;
  assign n9286 = n9279 & n9285;
  assign n9287 = ~n9276 & n9286;
  assign n9288 = ~n3455 & n9280;
  assign n9289 = n9287 & ~n9288;
  assign n9290 = n9275 & n9289;
  assign n9291 = n3033 & n9259;
  assign n9292 = n9290 & ~n9291;
  assign n9293 = n2910 & n9259;
  assign n9294 = n9292 & ~n9293;
  assign n9295 = ~n9271 & n9294;
  assign n9296 = pi0085 & ~n4014;
  assign n9297 = n3110 & n9259;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = pi0085 & po0740;
  assign n9300 = n2651 & n9299;
  assign n9301 = ~n3102 & n9300;
  assign n9302 = pi0085 & n4006;
  assign n9303 = ~n9301 & ~n9302;
  assign n9304 = pi1044 & n9280;
  assign n9305 = n2619 & n9304;
  assign n9306 = n2644 & n9257;
  assign n9307 = ~n9305 & ~n9306;
  assign n9308 = n2591 & n9259;
  assign n9309 = n9307 & ~n9308;
  assign n9310 = n9303 & n9309;
  assign n9311 = n9298 & n9310;
  assign n9312 = n9295 & n9311;
  assign n9313 = ~n4105 & n9280;
  assign n9314 = n2569 & n9259;
  assign n9315 = ~n9313 & ~n9314;
  assign n9316 = pi0085 & pi0993;
  assign n9317 = n2576 & n9316;
  assign n9318 = n2598 & n9259;
  assign n9319 = ~n9317 & ~n9318;
  assign n9320 = n9315 & n9319;
  assign n9321 = n9312 & n9320;
  assign n9322 = n9270 & n9321;
  assign n9323 = ~n9254 & n9322;
  assign n9324 = pi0085 & n4089;
  assign n9325 = pi0085 & n4091;
  assign n9326 = pi0085 & n3128;
  assign n9327 = ~n4094 & n9326;
  assign n9328 = ~n4097 & n9299;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = n3397 & ~n9329;
  assign n9331 = ~n9325 & ~n9330;
  assign n9332 = ~n9324 & n9331;
  assign n9333 = n4087 & ~n9332;
  assign n9334 = n3057 & n9259;
  assign n9335 = pi0085 & ~n3057;
  assign n9336 = ~n9334 & ~n9335;
  assign n9337 = n4083 & ~n9336;
  assign n9338 = n2901 & n9280;
  assign n9339 = ~n9337 & ~n9338;
  assign n9340 = ~n3072 & n9259;
  assign n9341 = n2847 & n9257;
  assign n9342 = n2834 & n9304;
  assign n9343 = ~n9341 & ~n9342;
  assign n9344 = n2858 & n9257;
  assign n9345 = pi0085 & n4124;
  assign n9346 = n2854 & n9259;
  assign n9347 = n2881 & n9299;
  assign n9348 = n2726 & n9347;
  assign n9349 = ~n9346 & ~n9348;
  assign n9350 = ~n9345 & n9349;
  assign n9351 = ~n9344 & n9350;
  assign n9352 = ~n4133 & n9257;
  assign n9353 = n9351 & ~n9352;
  assign n9354 = n2851 & n9280;
  assign n9355 = n3066 & n9259;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = n9353 & n9356;
  assign n9358 = n9343 & n9357;
  assign n9359 = ~n9340 & n9358;
  assign n9360 = n2681 & n9259;
  assign n9361 = ~n4077 & n9257;
  assign n9362 = ~n9360 & ~n9361;
  assign n9363 = n9359 & n9362;
  assign n9364 = n9339 & n9363;
  assign n9365 = ~n9333 & n9364;
  assign po0243 = ~n9323 | ~n9365;
  assign n9367 = pi0086 & ~n4061;
  assign n9368 = n4060 & n9367;
  assign n9369 = pi0086 & pi0841;
  assign n9370 = n2917 & n9369;
  assign n9371 = pi0024 & pi0086;
  assign n9372 = n2913 & n9371;
  assign n9373 = ~n9370 & ~n9372;
  assign n9374 = pi0086 & ~pi0314;
  assign n9375 = n2936 & n9374;
  assign n9376 = n9373 & ~n9375;
  assign n9377 = pi0086 & n4043;
  assign n9378 = n2930 & n9377;
  assign n9379 = pi0086 & ~n3553;
  assign n9380 = n4497 & n9379;
  assign n9381 = ~n9378 & ~n9380;
  assign n9382 = ~n4402 & n9374;
  assign n9383 = n9381 & ~n9382;
  assign n9384 = n3042 & n9371;
  assign n9385 = pi0086 & n4504;
  assign n9386 = ~n9384 & ~n9385;
  assign n9387 = n9383 & n9386;
  assign n9388 = n9376 & n9387;
  assign n9389 = n3033 & n9371;
  assign n9390 = n9388 & ~n9389;
  assign n9391 = n2591 & n9371;
  assign n9392 = pi0086 & n4067;
  assign n9393 = pi1044 & n9374;
  assign n9394 = n2619 & n9393;
  assign n9395 = n2644 & n9369;
  assign n9396 = ~n9394 & ~n9395;
  assign n9397 = n2910 & n9371;
  assign n9398 = n9396 & ~n9397;
  assign n9399 = ~n9392 & n9398;
  assign n9400 = ~n9391 & n9399;
  assign n9401 = pi0086 & pi0993;
  assign n9402 = n2576 & n9401;
  assign n9403 = n2598 & n9371;
  assign n9404 = ~n9402 & ~n9403;
  assign n9405 = pi0086 & po0740;
  assign n9406 = n2651 & n9405;
  assign n9407 = ~n3102 & n9406;
  assign n9408 = pi0086 & n4006;
  assign n9409 = ~n9407 & ~n9408;
  assign n9410 = ~n4105 & n9374;
  assign n9411 = n2569 & n9371;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = pi0086 & ~n4014;
  assign n9414 = n3110 & n9371;
  assign n9415 = ~n9413 & ~n9414;
  assign n9416 = n9412 & n9415;
  assign n9417 = n9409 & n9416;
  assign n9418 = n9404 & n9417;
  assign n9419 = n9400 & n9418;
  assign n9420 = pi0086 & n2741;
  assign n9421 = pi0086 & n4708;
  assign n9422 = ~n3973 & n9421;
  assign n9423 = ~n3998 & n9369;
  assign n9424 = pi0086 & n3989;
  assign n9425 = ~n9371 & ~n9424;
  assign n9426 = n2563 & ~n9425;
  assign n9427 = n2795 & n9371;
  assign n9428 = ~n9426 & ~n9427;
  assign n9429 = ~n9423 & n9428;
  assign n9430 = ~n9422 & n9429;
  assign n9431 = ~n9420 & n9430;
  assign n9432 = n9419 & n9431;
  assign n9433 = pi0086 & n2604;
  assign n9434 = n3967 & n9433;
  assign n9435 = n9432 & ~n9434;
  assign n9436 = n9390 & n9435;
  assign n9437 = ~n9368 & n9436;
  assign n9438 = pi0086 & n4091;
  assign n9439 = pi0086 & n4459;
  assign n9440 = n2440 & n3102;
  assign n9441 = ~n4097 & n9405;
  assign n9442 = ~n9440 & ~n9441;
  assign n9443 = ~n9439 & n9442;
  assign n9444 = n3397 & ~n9443;
  assign n9445 = pi0086 & ~pi0786;
  assign n9446 = n4088 & n9445;
  assign n9447 = ~n9444 & ~n9446;
  assign n9448 = ~n9438 & n9447;
  assign n9449 = n4087 & ~n9448;
  assign n9450 = n3057 & n9371;
  assign n9451 = pi0086 & ~n3057;
  assign n9452 = ~n9450 & ~n9451;
  assign n9453 = n4083 & ~n9452;
  assign n9454 = n2901 & n9374;
  assign n9455 = ~n9453 & ~n9454;
  assign n9456 = ~n3072 & n9371;
  assign n9457 = n2847 & n9369;
  assign n9458 = n2834 & n9393;
  assign n9459 = ~n9457 & ~n9458;
  assign n9460 = n2858 & n9369;
  assign n9461 = pi0086 & n4124;
  assign n9462 = n2854 & n9371;
  assign n9463 = n2881 & n9405;
  assign n9464 = n2726 & n9463;
  assign n9465 = ~n9462 & ~n9464;
  assign n9466 = ~n9461 & n9465;
  assign n9467 = ~n9460 & n9466;
  assign n9468 = ~n4133 & n9369;
  assign n9469 = n9467 & ~n9468;
  assign n9470 = n2851 & n9374;
  assign n9471 = n3066 & n9371;
  assign n9472 = ~n9470 & ~n9471;
  assign n9473 = n9469 & n9472;
  assign n9474 = n9459 & n9473;
  assign n9475 = ~n9456 & n9474;
  assign n9476 = n2681 & n9371;
  assign n9477 = ~n4077 & n9369;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = n9475 & n9478;
  assign n9480 = n9455 & n9479;
  assign n9481 = ~n9449 & n9480;
  assign po0244 = ~n9437 | ~n9481;
  assign n9483 = pi0024 & pi0087;
  assign n9484 = n3057 & n9483;
  assign n9485 = pi0087 & ~n3057;
  assign n9486 = ~n9484 & ~n9485;
  assign n9487 = n4083 & ~n9486;
  assign n9488 = pi0087 & ~pi0314;
  assign n9489 = n2901 & n9488;
  assign n9490 = ~n9487 & ~n9489;
  assign n9491 = n2681 & n9483;
  assign n9492 = pi0087 & pi0841;
  assign n9493 = ~n4077 & n9492;
  assign n9494 = ~n9491 & ~n9493;
  assign n9495 = pi0087 & n4089;
  assign n9496 = pi0087 & n4091;
  assign n9497 = pi0087 & n3128;
  assign n9498 = ~n4094 & n9497;
  assign n9499 = pi0087 & po0740;
  assign n9500 = ~n4097 & n9499;
  assign n9501 = ~n9498 & ~n9500;
  assign n9502 = n3397 & ~n9501;
  assign n9503 = ~n9496 & ~n9502;
  assign n9504 = ~n9495 & n9503;
  assign n9505 = n4087 & ~n9504;
  assign n9506 = n9494 & ~n9505;
  assign n9507 = n9490 & n9506;
  assign n9508 = ~n3072 & n9483;
  assign n9509 = n2847 & n9492;
  assign n9510 = pi1044 & n9488;
  assign n9511 = n2834 & n9510;
  assign n9512 = ~n9509 & ~n9511;
  assign n9513 = ~pi0087 & ~pi0314;
  assign n9514 = n2851 & ~n9513;
  assign n9515 = n2858 & n9492;
  assign n9516 = pi0087 & n4124;
  assign n9517 = n2854 & n9483;
  assign n9518 = n2881 & n9499;
  assign n9519 = n2726 & n9518;
  assign n9520 = ~n9517 & ~n9519;
  assign n9521 = ~n9516 & n9520;
  assign n9522 = ~n9515 & n9521;
  assign n9523 = n3066 & n9483;
  assign n9524 = n9522 & ~n9523;
  assign n9525 = ~n9514 & n9524;
  assign n9526 = n9512 & n9525;
  assign n9527 = ~n9508 & n9526;
  assign n9528 = n9507 & n9527;
  assign n9529 = ~n4105 & n9488;
  assign n9530 = n2569 & n9483;
  assign n9531 = ~n9529 & ~n9530;
  assign n9532 = pi0087 & pi0993;
  assign n9533 = n2576 & n9532;
  assign n9534 = n2598 & n9483;
  assign n9535 = ~n9533 & ~n9534;
  assign n9536 = n9531 & n9535;
  assign n9537 = pi0087 & n4006;
  assign n9538 = pi0087 & ~n4014;
  assign n9539 = n3110 & n9483;
  assign n9540 = ~n9538 & ~n9539;
  assign n9541 = n2651 & n9499;
  assign n9542 = ~n3102 & n9541;
  assign n9543 = n9540 & ~n9542;
  assign n9544 = ~n9537 & n9543;
  assign n9545 = n2591 & n9483;
  assign n9546 = n9544 & ~n9545;
  assign n9547 = n2619 & n9510;
  assign n9548 = n2644 & n9492;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = n2917 & n9492;
  assign n9551 = n2913 & n9483;
  assign n9552 = ~n9550 & ~n9551;
  assign n9553 = n2936 & n9488;
  assign n9554 = n9552 & ~n9553;
  assign n9555 = n3042 & n9483;
  assign n9556 = pi0087 & n4043;
  assign n9557 = n2930 & n9556;
  assign n9558 = pi0087 & ~n3553;
  assign n9559 = n4497 & n9558;
  assign n9560 = ~n9557 & ~n9559;
  assign n9561 = ~n4402 & n9488;
  assign n9562 = n9560 & ~n9561;
  assign n9563 = pi0087 & n4504;
  assign n9564 = n9562 & ~n9563;
  assign n9565 = ~n9555 & n9564;
  assign n9566 = n9554 & n9565;
  assign n9567 = n3033 & n9483;
  assign n9568 = n9566 & ~n9567;
  assign n9569 = n2910 & n9483;
  assign n9570 = pi0087 & n2726;
  assign n9571 = n4066 & n9570;
  assign n9572 = ~n9569 & ~n9571;
  assign n9573 = n9568 & n9572;
  assign n9574 = n9549 & n9573;
  assign n9575 = n9546 & n9574;
  assign n9576 = pi0087 & n4585;
  assign n9577 = pi0087 & n3989;
  assign n9578 = ~n9483 & ~n9577;
  assign n9579 = n2563 & ~n9578;
  assign n9580 = n2795 & n9483;
  assign n9581 = ~n9579 & ~n9580;
  assign n9582 = pi0087 & n2741;
  assign n9583 = n9581 & ~n9582;
  assign n9584 = ~n9576 & n9583;
  assign n9585 = ~n3998 & n9492;
  assign n9586 = n9584 & ~n9585;
  assign n9587 = pi0087 & n4336;
  assign n9588 = pi0087 & n4062;
  assign n9589 = ~n9587 & ~n9588;
  assign n9590 = n9586 & n9589;
  assign n9591 = n9575 & n9590;
  assign n9592 = ~n4133 & n9492;
  assign n9593 = n9591 & ~n9592;
  assign n9594 = n9536 & n9593;
  assign po0245 = ~n9528 | ~n9594;
  assign n9596 = pi0088 & pi0993;
  assign n9597 = n2576 & n9596;
  assign n9598 = pi0024 & pi0088;
  assign n9599 = n2598 & n9598;
  assign n9600 = ~n9597 & ~n9599;
  assign n9601 = pi0088 & ~pi0314;
  assign n9602 = ~n4105 & n9601;
  assign n9603 = n2569 & n9598;
  assign n9604 = ~n9602 & ~n9603;
  assign n9605 = pi0088 & n4336;
  assign n9606 = pi0088 & ~n4061;
  assign n9607 = n4060 & n9606;
  assign n9608 = ~n9605 & ~n9607;
  assign n9609 = n9604 & n9608;
  assign n9610 = n9600 & n9609;
  assign n9611 = pi0088 & n2741;
  assign n9612 = pi0088 & n4523;
  assign n9613 = ~n3973 & n9612;
  assign n9614 = pi0088 & pi0841;
  assign n9615 = ~n3998 & n9614;
  assign n9616 = pi0088 & n3989;
  assign n9617 = ~n9598 & ~n9616;
  assign n9618 = n2563 & ~n9617;
  assign n9619 = n2795 & n9598;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = ~n9615 & n9620;
  assign n9622 = ~n9613 & n9621;
  assign n9623 = ~n9611 & n9622;
  assign n9624 = n9610 & n9623;
  assign n9625 = ~n3072 & n9598;
  assign n9626 = n2847 & n9614;
  assign n9627 = pi1044 & n9601;
  assign n9628 = n2834 & n9627;
  assign n9629 = ~n9626 & ~n9628;
  assign n9630 = n2858 & n9614;
  assign n9631 = pi0088 & n4124;
  assign n9632 = n2854 & n9598;
  assign n9633 = pi0088 & po0740;
  assign n9634 = n2881 & n9633;
  assign n9635 = n2726 & n9634;
  assign n9636 = ~n9632 & ~n9635;
  assign n9637 = ~n9631 & n9636;
  assign n9638 = ~n9630 & n9637;
  assign n9639 = ~n4133 & n9614;
  assign n9640 = n9638 & ~n9639;
  assign n9641 = n2851 & n9601;
  assign n9642 = n3066 & n9598;
  assign n9643 = ~n9641 & ~n9642;
  assign n9644 = n9640 & n9643;
  assign n9645 = n9629 & n9644;
  assign n9646 = ~n9625 & n9645;
  assign n9647 = n2619 & n9627;
  assign n9648 = n2644 & n9614;
  assign n9649 = ~n9647 & ~n9648;
  assign n9650 = n2917 & n9614;
  assign n9651 = n2913 & n9598;
  assign n9652 = ~n9650 & ~n9651;
  assign n9653 = n2936 & n9601;
  assign n9654 = n9652 & ~n9653;
  assign n9655 = pi0088 & n4043;
  assign n9656 = n2930 & n9655;
  assign n9657 = pi0088 & ~n3553;
  assign n9658 = n4497 & n9657;
  assign n9659 = ~n9656 & ~n9658;
  assign n9660 = ~n4402 & n9601;
  assign n9661 = n9659 & ~n9660;
  assign n9662 = pi0088 & n2726;
  assign n9663 = ~n4064 & ~n9662;
  assign n9664 = n2516 & ~n9663;
  assign n9665 = pi0088 & n4504;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = n9661 & n9666;
  assign n9668 = n9654 & n9667;
  assign n9669 = ~n5328 & n9598;
  assign n9670 = n9668 & ~n9669;
  assign n9671 = pi0088 & n4006;
  assign n9672 = pi0088 & ~n4014;
  assign n9673 = n3110 & n9598;
  assign n9674 = ~n9672 & ~n9673;
  assign n9675 = n2651 & n9633;
  assign n9676 = ~n3102 & n9675;
  assign n9677 = n9674 & ~n9676;
  assign n9678 = ~n9671 & n9677;
  assign n9679 = n2591 & n9598;
  assign n9680 = n9678 & ~n9679;
  assign n9681 = n9670 & n9680;
  assign n9682 = n9649 & n9681;
  assign n9683 = n2681 & n9598;
  assign n9684 = ~n4077 & n9614;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = pi0088 & n4089;
  assign n9687 = pi0088 & n4091;
  assign n9688 = pi0088 & n3128;
  assign n9689 = ~n4094 & n9688;
  assign n9690 = ~n4097 & n9633;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = n3397 & ~n9691;
  assign n9693 = ~n9687 & ~n9692;
  assign n9694 = ~n9686 & n9693;
  assign n9695 = n4087 & ~n9694;
  assign n9696 = n3057 & n9598;
  assign n9697 = pi0088 & ~n3057;
  assign n9698 = ~n9696 & ~n9697;
  assign n9699 = n4083 & ~n9698;
  assign n9700 = n2901 & n9601;
  assign n9701 = ~n9699 & ~n9700;
  assign n9702 = ~n9695 & n9701;
  assign n9703 = n9685 & n9702;
  assign n9704 = n9682 & n9703;
  assign n9705 = n9646 & n9704;
  assign po0246 = ~n9624 | ~n9705;
  assign n9707 = pi0089 & ~pi0314;
  assign n9708 = ~n4105 & n9707;
  assign n9709 = pi0024 & pi0089;
  assign n9710 = n2569 & n9709;
  assign n9711 = ~n9708 & ~n9710;
  assign n9712 = pi0089 & pi0993;
  assign n9713 = n2576 & n9712;
  assign n9714 = n2598 & n9709;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = n9711 & n9715;
  assign n9717 = pi0089 & n4067;
  assign n9718 = pi0089 & ~n4014;
  assign n9719 = n3110 & n9709;
  assign n9720 = ~n9718 & ~n9719;
  assign n9721 = n2910 & n9709;
  assign n9722 = n9720 & ~n9721;
  assign n9723 = ~n9717 & n9722;
  assign n9724 = n9716 & n9723;
  assign n9725 = pi0089 & n2604;
  assign n9726 = n3967 & n9725;
  assign n9727 = n2591 & n9709;
  assign n9728 = pi1044 & n9707;
  assign n9729 = n2619 & n9728;
  assign n9730 = pi0089 & pi0841;
  assign n9731 = n2644 & n9730;
  assign n9732 = ~n9729 & ~n9731;
  assign n9733 = pi0089 & ~n4061;
  assign n9734 = n4060 & n9733;
  assign n9735 = pi0089 & po0740;
  assign n9736 = n2651 & n9735;
  assign n9737 = ~n3102 & n9736;
  assign n9738 = pi0089 & n4006;
  assign n9739 = ~n9737 & ~n9738;
  assign n9740 = ~n9734 & n9739;
  assign n9741 = n9732 & n9740;
  assign n9742 = ~n9727 & n9741;
  assign n9743 = pi0089 & n2741;
  assign n9744 = pi0089 & n4523;
  assign n9745 = ~n3973 & n9744;
  assign n9746 = ~n3998 & n9730;
  assign n9747 = pi0089 & n3989;
  assign n9748 = ~n9709 & ~n9747;
  assign n9749 = n2563 & ~n9748;
  assign n9750 = n2795 & n9709;
  assign n9751 = ~n9749 & ~n9750;
  assign n9752 = ~n9746 & n9751;
  assign n9753 = ~n9745 & n9752;
  assign n9754 = ~n9743 & n9753;
  assign n9755 = n9742 & n9754;
  assign n9756 = n2917 & n9730;
  assign n9757 = n2913 & n9709;
  assign n9758 = ~n9756 & ~n9757;
  assign n9759 = n2936 & n9707;
  assign n9760 = n9758 & ~n9759;
  assign n9761 = pi0089 & n4043;
  assign n9762 = n2930 & n9761;
  assign n9763 = pi0089 & ~n3553;
  assign n9764 = n4497 & n9763;
  assign n9765 = ~n9762 & ~n9764;
  assign n9766 = ~n4402 & n9707;
  assign n9767 = n9765 & ~n9766;
  assign n9768 = n3042 & n9709;
  assign n9769 = pi0089 & n4504;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = n9767 & n9770;
  assign n9772 = n9760 & n9771;
  assign n9773 = n3033 & n9709;
  assign n9774 = n9772 & ~n9773;
  assign n9775 = n9755 & n9774;
  assign n9776 = ~n9726 & n9775;
  assign n9777 = n9724 & n9776;
  assign n9778 = pi0089 & n4089;
  assign n9779 = pi0089 & n4091;
  assign n9780 = pi0089 & n3128;
  assign n9781 = ~n4094 & n9780;
  assign n9782 = ~n4097 & n9735;
  assign n9783 = ~n9781 & ~n9782;
  assign n9784 = n3397 & ~n9783;
  assign n9785 = ~n9779 & ~n9784;
  assign n9786 = ~n9778 & n9785;
  assign n9787 = n4087 & ~n9786;
  assign n9788 = n3057 & n9709;
  assign n9789 = pi0089 & ~n3057;
  assign n9790 = ~n9788 & ~n9789;
  assign n9791 = n4083 & ~n9790;
  assign n9792 = n2901 & n9707;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = ~n3072 & n9709;
  assign n9795 = n2847 & n9730;
  assign n9796 = n2834 & n9728;
  assign n9797 = ~n9795 & ~n9796;
  assign n9798 = pi0024 & ~pi0089;
  assign n9799 = n2854 & ~n9798;
  assign n9800 = n2881 & n9735;
  assign n9801 = n2726 & n9800;
  assign n9802 = pi0089 & n4124;
  assign n9803 = n2858 & n9730;
  assign n9804 = ~n9802 & ~n9803;
  assign n9805 = ~n9801 & n9804;
  assign n9806 = ~n9799 & n9805;
  assign n9807 = ~n4133 & n9730;
  assign n9808 = n9806 & ~n9807;
  assign n9809 = n2851 & n9707;
  assign n9810 = n3066 & n9709;
  assign n9811 = ~n9809 & ~n9810;
  assign n9812 = n9808 & n9811;
  assign n9813 = n9797 & n9812;
  assign n9814 = ~n9794 & n9813;
  assign n9815 = n2681 & n9709;
  assign n9816 = ~n4077 & n9730;
  assign n9817 = ~n9815 & ~n9816;
  assign n9818 = n9814 & n9817;
  assign n9819 = n9793 & n9818;
  assign n9820 = ~n9787 & n9819;
  assign po0247 = ~n9777 | ~n9820;
  assign n9822 = pi0090 & n4336;
  assign n9823 = pi0090 & n2741;
  assign n9824 = pi0090 & n4523;
  assign n9825 = ~n3973 & n9824;
  assign n9826 = pi0090 & pi0841;
  assign n9827 = ~n3998 & n9826;
  assign n9828 = pi0024 & pi0090;
  assign n9829 = pi0090 & n3989;
  assign n9830 = ~n9828 & ~n9829;
  assign n9831 = n2563 & ~n9830;
  assign n9832 = n2795 & n9828;
  assign n9833 = ~n9831 & ~n9832;
  assign n9834 = ~n9827 & n9833;
  assign n9835 = ~n9825 & n9834;
  assign n9836 = ~n9823 & n9835;
  assign n9837 = pi0090 & ~n4061;
  assign n9838 = n4060 & n9837;
  assign n9839 = n9836 & ~n9838;
  assign n9840 = pi0090 & ~pi0314;
  assign n9841 = ~n4105 & n9840;
  assign n9842 = n2569 & n9828;
  assign n9843 = ~n9841 & ~n9842;
  assign n9844 = pi0090 & pi0993;
  assign n9845 = n2576 & n9844;
  assign n9846 = n2598 & n9828;
  assign n9847 = ~n9845 & ~n9846;
  assign n9848 = n9843 & n9847;
  assign n9849 = pi0090 & n4067;
  assign n9850 = ~n4402 & n9840;
  assign n9851 = pi0090 & n2926;
  assign n9852 = ~pi1076 & n9851;
  assign n9853 = n3042 & n9828;
  assign n9854 = n2936 & n9840;
  assign n9855 = ~n9853 & ~n9854;
  assign n9856 = ~n9852 & n9855;
  assign n9857 = ~n9850 & n9856;
  assign n9858 = n2917 & n9826;
  assign n9859 = n2913 & n9828;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = n9857 & n9860;
  assign n9862 = pi0090 & n4043;
  assign n9863 = n2930 & n9862;
  assign n9864 = pi0090 & ~n3553;
  assign n9865 = n4497 & n9864;
  assign n9866 = ~n9863 & ~n9865;
  assign n9867 = n9861 & n9866;
  assign n9868 = n3033 & n9828;
  assign n9869 = n9867 & ~n9868;
  assign n9870 = n2910 & n9828;
  assign n9871 = n9869 & ~n9870;
  assign n9872 = ~n9849 & n9871;
  assign n9873 = pi0090 & po0740;
  assign n9874 = n2651 & n9873;
  assign n9875 = ~n3102 & n9874;
  assign n9876 = pi0090 & n4006;
  assign n9877 = n2644 & n9826;
  assign n9878 = n2619 & n9840;
  assign n9879 = pi1044 & n9878;
  assign n9880 = ~n9877 & ~n9879;
  assign n9881 = n2591 & n9828;
  assign n9882 = n9880 & ~n9881;
  assign n9883 = pi0090 & ~n4014;
  assign n9884 = n3110 & n9828;
  assign n9885 = ~n9883 & ~n9884;
  assign n9886 = n9882 & n9885;
  assign n9887 = ~n9876 & n9886;
  assign n9888 = ~n9875 & n9887;
  assign n9889 = n9872 & n9888;
  assign n9890 = n9848 & n9889;
  assign n9891 = n9839 & n9890;
  assign n9892 = ~n9822 & n9891;
  assign n9893 = n2847 & n9826;
  assign n9894 = n2788 & n9828;
  assign n9895 = ~n9893 & ~n9894;
  assign n9896 = ~n4326 & n9828;
  assign n9897 = n9895 & ~n9896;
  assign n9898 = n2851 & n9840;
  assign n9899 = n3066 & n9828;
  assign n9900 = ~n9898 & ~n9899;
  assign n9901 = ~n4077 & n9826;
  assign n9902 = n2681 & n9828;
  assign n9903 = ~n9901 & ~n9902;
  assign n9904 = pi0090 & n4091;
  assign n9905 = ~n4097 & n9873;
  assign n9906 = pi0090 & n4459;
  assign n9907 = ~n9905 & ~n9906;
  assign n9908 = n3397 & ~n9907;
  assign n9909 = pi0090 & ~pi0786;
  assign n9910 = n4088 & n9909;
  assign n9911 = ~n9908 & ~n9910;
  assign n9912 = ~n9904 & n9911;
  assign n9913 = n4087 & ~n9912;
  assign n9914 = n2901 & n9840;
  assign n9915 = n3057 & n9828;
  assign n9916 = pi0090 & ~n3057;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 = n4083 & ~n9917;
  assign n9919 = ~n9914 & ~n9918;
  assign n9920 = ~n9913 & n9919;
  assign n9921 = n9903 & n9920;
  assign n9922 = pi1044 & ~n9840;
  assign n9923 = n2834 & ~n9922;
  assign n9924 = n2881 & n9873;
  assign n9925 = n2726 & n9924;
  assign n9926 = pi0090 & n4124;
  assign n9927 = n2858 & n9826;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = ~n9925 & n9928;
  assign n9930 = ~n9923 & n9929;
  assign n9931 = ~n4133 & n9826;
  assign n9932 = n9930 & ~n9931;
  assign n9933 = n9921 & n9932;
  assign n9934 = n9900 & n9933;
  assign n9935 = n9897 & n9934;
  assign po0248 = ~n9892 | ~n9935;
  assign n9937 = pi0091 & n4336;
  assign n9938 = pi0091 & n2741;
  assign n9939 = pi0091 & n4708;
  assign n9940 = ~n3973 & n9939;
  assign n9941 = pi0091 & pi0841;
  assign n9942 = ~n3998 & n9941;
  assign n9943 = pi0024 & pi0091;
  assign n9944 = pi0091 & n3989;
  assign n9945 = ~n9943 & ~n9944;
  assign n9946 = n2563 & ~n9945;
  assign n9947 = n2795 & n9943;
  assign n9948 = ~n9946 & ~n9947;
  assign n9949 = ~n9942 & n9948;
  assign n9950 = ~n9940 & n9949;
  assign n9951 = ~n9938 & n9950;
  assign n9952 = pi0091 & ~n4061;
  assign n9953 = n4060 & n9952;
  assign n9954 = n9951 & ~n9953;
  assign n9955 = pi0091 & ~pi0314;
  assign n9956 = ~n4105 & n9955;
  assign n9957 = n2569 & n9943;
  assign n9958 = ~n9956 & ~n9957;
  assign n9959 = pi0091 & pi0993;
  assign n9960 = n2576 & n9959;
  assign n9961 = n2598 & n9943;
  assign n9962 = ~n9960 & ~n9961;
  assign n9963 = n9958 & n9962;
  assign n9964 = pi0091 & n4067;
  assign n9965 = n2917 & n9941;
  assign n9966 = n2913 & n9943;
  assign n9967 = ~n9965 & ~n9966;
  assign n9968 = n2936 & n9955;
  assign n9969 = n9967 & ~n9968;
  assign n9970 = pi0091 & n4043;
  assign n9971 = n2930 & n9970;
  assign n9972 = pi0091 & ~n3553;
  assign n9973 = n4497 & n9972;
  assign n9974 = ~n9971 & ~n9973;
  assign n9975 = ~n4402 & n9955;
  assign n9976 = n9974 & ~n9975;
  assign n9977 = n3042 & n9943;
  assign n9978 = pi0091 & n4504;
  assign n9979 = ~n9977 & ~n9978;
  assign n9980 = n9976 & n9979;
  assign n9981 = n9969 & n9980;
  assign n9982 = n3033 & n9943;
  assign n9983 = n9981 & ~n9982;
  assign n9984 = n2910 & n9943;
  assign n9985 = n9983 & ~n9984;
  assign n9986 = ~n9964 & n9985;
  assign n9987 = pi0091 & ~n4014;
  assign n9988 = n3110 & n9943;
  assign n9989 = ~n9987 & ~n9988;
  assign n9990 = pi0091 & po0740;
  assign n9991 = n2651 & n9990;
  assign n9992 = ~n3102 & n9991;
  assign n9993 = pi0091 & n4006;
  assign n9994 = ~n9992 & ~n9993;
  assign n9995 = pi1044 & n9955;
  assign n9996 = n2619 & n9995;
  assign n9997 = n2644 & n9941;
  assign n9998 = ~n9996 & ~n9997;
  assign n9999 = n2591 & n9943;
  assign n10000 = n9998 & ~n9999;
  assign n10001 = n9994 & n10000;
  assign n10002 = n9989 & n10001;
  assign n10003 = n9986 & n10002;
  assign n10004 = n9963 & n10003;
  assign n10005 = n9954 & n10004;
  assign n10006 = ~n9937 & n10005;
  assign n10007 = pi0091 & n4091;
  assign n10008 = pi0091 & n4459;
  assign n10009 = ~n4097 & n9990;
  assign n10010 = ~n3549 & ~n10009;
  assign n10011 = ~n10008 & n10010;
  assign n10012 = n3397 & ~n10011;
  assign n10013 = pi0091 & ~pi0786;
  assign n10014 = n4088 & n10013;
  assign n10015 = ~n10012 & ~n10014;
  assign n10016 = ~n10007 & n10015;
  assign n10017 = n3547 & ~n10016;
  assign n10018 = n3406 & n10017;
  assign n10019 = n3057 & n9943;
  assign n10020 = pi0091 & ~n3057;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = n4083 & ~n10021;
  assign n10023 = ~n10018 & ~n10022;
  assign n10024 = n2888 & n3102;
  assign n10025 = ~n3072 & n9943;
  assign n10026 = n2847 & n9941;
  assign n10027 = n2834 & n9995;
  assign n10028 = ~n10026 & ~n10027;
  assign n10029 = n2858 & n9941;
  assign n10030 = pi0091 & n4124;
  assign n10031 = n2854 & n9943;
  assign n10032 = n2881 & n9990;
  assign n10033 = n2726 & n10032;
  assign n10034 = ~n10031 & ~n10033;
  assign n10035 = ~n10030 & n10034;
  assign n10036 = ~n10029 & n10035;
  assign n10037 = ~n4133 & n9941;
  assign n10038 = n10036 & ~n10037;
  assign n10039 = n2851 & n9955;
  assign n10040 = n3066 & n9943;
  assign n10041 = ~n10039 & ~n10040;
  assign n10042 = n10038 & n10041;
  assign n10043 = n10028 & n10042;
  assign n10044 = ~n10025 & n10043;
  assign n10045 = n2901 & n9955;
  assign n10046 = n2681 & n9943;
  assign n10047 = ~n10045 & ~n10046;
  assign n10048 = ~n4077 & n9941;
  assign n10049 = n10047 & ~n10048;
  assign n10050 = n10044 & n10049;
  assign n10051 = ~n10024 & n10050;
  assign n10052 = n10023 & n10051;
  assign po0249 = ~n10006 | ~n10052;
  assign n10054 = pi0092 & ~pi0314;
  assign n10055 = ~n4105 & n10054;
  assign n10056 = pi0024 & pi0092;
  assign n10057 = n2569 & n10056;
  assign n10058 = ~n10055 & ~n10057;
  assign n10059 = pi0092 & pi0993;
  assign n10060 = n2576 & n10059;
  assign n10061 = n2598 & n10056;
  assign n10062 = ~n10060 & ~n10061;
  assign n10063 = n10058 & n10062;
  assign n10064 = pi0092 & n4067;
  assign n10065 = pi0092 & ~n4014;
  assign n10066 = n3110 & n10056;
  assign n10067 = ~n10065 & ~n10066;
  assign n10068 = n2910 & n10056;
  assign n10069 = n10067 & ~n10068;
  assign n10070 = ~n10064 & n10069;
  assign n10071 = n10063 & n10070;
  assign n10072 = pi0092 & n2604;
  assign n10073 = n3967 & n10072;
  assign n10074 = n2591 & n10056;
  assign n10075 = pi1044 & n10054;
  assign n10076 = n2619 & n10075;
  assign n10077 = pi0092 & pi0841;
  assign n10078 = n2644 & n10077;
  assign n10079 = ~n10076 & ~n10078;
  assign n10080 = pi0092 & ~n4061;
  assign n10081 = n4060 & n10080;
  assign n10082 = pi0092 & po0740;
  assign n10083 = n2651 & n10082;
  assign n10084 = ~n3102 & n10083;
  assign n10085 = pi0092 & n4006;
  assign n10086 = ~n10084 & ~n10085;
  assign n10087 = ~n10081 & n10086;
  assign n10088 = n10079 & n10087;
  assign n10089 = ~n10074 & n10088;
  assign n10090 = pi0092 & n2741;
  assign n10091 = pi0092 & n4708;
  assign n10092 = ~n3973 & n10091;
  assign n10093 = ~n3998 & n10077;
  assign n10094 = pi0092 & n3989;
  assign n10095 = ~n10056 & ~n10094;
  assign n10096 = n2563 & ~n10095;
  assign n10097 = n2795 & n10056;
  assign n10098 = ~n10096 & ~n10097;
  assign n10099 = ~n10093 & n10098;
  assign n10100 = ~n10092 & n10099;
  assign n10101 = ~n10090 & n10100;
  assign n10102 = n10089 & n10101;
  assign n10103 = n2917 & n10077;
  assign n10104 = n2913 & n10056;
  assign n10105 = ~n10103 & ~n10104;
  assign n10106 = n2936 & n10054;
  assign n10107 = n10105 & ~n10106;
  assign n10108 = pi0092 & n4043;
  assign n10109 = n2930 & n10108;
  assign n10110 = pi0092 & ~n3553;
  assign n10111 = n4497 & n10110;
  assign n10112 = ~n10109 & ~n10111;
  assign n10113 = ~n4402 & n10054;
  assign n10114 = n10112 & ~n10113;
  assign n10115 = n3042 & n10056;
  assign n10116 = pi0092 & n4504;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = n10114 & n10117;
  assign n10119 = n10107 & n10118;
  assign n10120 = n3033 & n10056;
  assign n10121 = n10119 & ~n10120;
  assign n10122 = n10102 & n10121;
  assign n10123 = ~n10073 & n10122;
  assign n10124 = n10071 & n10123;
  assign n10125 = pi0092 & n4091;
  assign n10126 = pi0092 & n4459;
  assign n10127 = n3102 & n3398;
  assign n10128 = ~n4097 & n10082;
  assign n10129 = ~n10127 & ~n10128;
  assign n10130 = ~n10126 & n10129;
  assign n10131 = n3397 & ~n10130;
  assign n10132 = pi0092 & ~pi0786;
  assign n10133 = n4088 & n10132;
  assign n10134 = ~n10131 & ~n10133;
  assign n10135 = ~n10125 & n10134;
  assign n10136 = n4087 & ~n10135;
  assign n10137 = n3057 & n10056;
  assign n10138 = pi0092 & ~n3057;
  assign n10139 = ~n10137 & ~n10138;
  assign n10140 = n4083 & ~n10139;
  assign n10141 = n2901 & n10054;
  assign n10142 = ~n10140 & ~n10141;
  assign n10143 = ~n3072 & n10056;
  assign n10144 = n2847 & n10077;
  assign n10145 = n2834 & n10075;
  assign n10146 = ~n10144 & ~n10145;
  assign n10147 = n2858 & n10077;
  assign n10148 = pi0092 & n4124;
  assign n10149 = n2854 & n10056;
  assign n10150 = n2881 & n10082;
  assign n10151 = n2726 & n10150;
  assign n10152 = ~n10149 & ~n10151;
  assign n10153 = ~n10148 & n10152;
  assign n10154 = ~n10147 & n10153;
  assign n10155 = ~n4133 & n10077;
  assign n10156 = n10154 & ~n10155;
  assign n10157 = n2851 & n10054;
  assign n10158 = n3066 & n10056;
  assign n10159 = ~n10157 & ~n10158;
  assign n10160 = n10156 & n10159;
  assign n10161 = n10146 & n10160;
  assign n10162 = ~n10143 & n10161;
  assign n10163 = n2681 & n10056;
  assign n10164 = ~n4077 & n10077;
  assign n10165 = ~n10163 & ~n10164;
  assign n10166 = n10162 & n10165;
  assign n10167 = n10142 & n10166;
  assign n10168 = ~n10136 & n10167;
  assign po0250 = ~n10124 | ~n10168;
  assign n10170 = pi0093 & n4336;
  assign n10171 = pi0093 & n2741;
  assign n10172 = pi0093 & n4708;
  assign n10173 = ~n3973 & n10172;
  assign n10174 = pi0093 & pi0841;
  assign n10175 = ~n3998 & n10174;
  assign n10176 = pi0024 & pi0093;
  assign n10177 = pi0093 & n3989;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = n2563 & ~n10178;
  assign n10180 = n2795 & n10176;
  assign n10181 = ~n10179 & ~n10180;
  assign n10182 = ~n10175 & n10181;
  assign n10183 = ~n10173 & n10182;
  assign n10184 = ~n10171 & n10183;
  assign n10185 = pi0093 & ~n4061;
  assign n10186 = n4060 & n10185;
  assign n10187 = n10184 & ~n10186;
  assign n10188 = pi0093 & ~pi0314;
  assign n10189 = ~n4105 & n10188;
  assign n10190 = n2569 & n10176;
  assign n10191 = ~n10189 & ~n10190;
  assign n10192 = pi0093 & pi0993;
  assign n10193 = n2576 & n10192;
  assign n10194 = n2598 & n10176;
  assign n10195 = ~n10193 & ~n10194;
  assign n10196 = n10191 & n10195;
  assign n10197 = pi0093 & n4067;
  assign n10198 = n2917 & n10174;
  assign n10199 = n2913 & n10176;
  assign n10200 = ~n10198 & ~n10199;
  assign n10201 = n2936 & n10188;
  assign n10202 = n10200 & ~n10201;
  assign n10203 = pi0093 & n4043;
  assign n10204 = n2930 & n10203;
  assign n10205 = pi0093 & ~n3553;
  assign n10206 = n4497 & n10205;
  assign n10207 = ~n10204 & ~n10206;
  assign n10208 = ~n4402 & n10188;
  assign n10209 = n10207 & ~n10208;
  assign n10210 = n3042 & n10176;
  assign n10211 = pi0093 & n4504;
  assign n10212 = ~n10210 & ~n10211;
  assign n10213 = n10209 & n10212;
  assign n10214 = n10202 & n10213;
  assign n10215 = n3033 & n10176;
  assign n10216 = n10214 & ~n10215;
  assign n10217 = n2910 & n10176;
  assign n10218 = n10216 & ~n10217;
  assign n10219 = ~n10197 & n10218;
  assign n10220 = pi0093 & ~n4014;
  assign n10221 = pi1044 & ~n10188;
  assign n10222 = n2619 & ~n10221;
  assign n10223 = pi0093 & po0740;
  assign n10224 = ~n3102 & n10223;
  assign n10225 = n2651 & n10224;
  assign n10226 = pi0093 & ~n3102;
  assign n10227 = n4005 & n10226;
  assign n10228 = ~n10225 & ~n10227;
  assign n10229 = ~n10222 & n10228;
  assign n10230 = n2644 & n10174;
  assign n10231 = n2591 & n10176;
  assign n10232 = ~n10230 & ~n10231;
  assign n10233 = n3110 & n10176;
  assign n10234 = n10232 & ~n10233;
  assign n10235 = n10229 & n10234;
  assign n10236 = ~n10220 & n10235;
  assign n10237 = n10219 & n10236;
  assign n10238 = n10196 & n10237;
  assign n10239 = n10187 & n10238;
  assign n10240 = ~n10170 & n10239;
  assign n10241 = n2847 & n10174;
  assign n10242 = n2834 & n10188;
  assign n10243 = pi1044 & n10242;
  assign n10244 = ~n10241 & ~n10243;
  assign n10245 = ~n3072 & n10176;
  assign n10246 = n10244 & ~n10245;
  assign n10247 = n2851 & n10188;
  assign n10248 = n3066 & n10176;
  assign n10249 = ~n10247 & ~n10248;
  assign n10250 = ~n4077 & n10174;
  assign n10251 = n2681 & n10176;
  assign n10252 = ~n10250 & ~n10251;
  assign n10253 = pi0093 & n4091;
  assign n10254 = ~n4097 & n10223;
  assign n10255 = pi0093 & n4459;
  assign n10256 = ~n10254 & ~n10255;
  assign n10257 = n3397 & ~n10256;
  assign n10258 = pi0093 & ~pi0786;
  assign n10259 = n4088 & n10258;
  assign n10260 = ~n10257 & ~n10259;
  assign n10261 = ~n10253 & n10260;
  assign n10262 = n4087 & ~n10261;
  assign n10263 = n2901 & n10188;
  assign n10264 = n3057 & n10176;
  assign n10265 = pi0093 & ~n3057;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = n4083 & ~n10266;
  assign n10268 = ~n10263 & ~n10267;
  assign n10269 = ~n10262 & n10268;
  assign n10270 = n10252 & n10269;
  assign n10271 = n2858 & n10174;
  assign n10272 = pi0093 & n4124;
  assign n10273 = n2854 & n10176;
  assign n10274 = n2881 & n10223;
  assign n10275 = n2726 & n10274;
  assign n10276 = ~n10273 & ~n10275;
  assign n10277 = ~n10272 & n10276;
  assign n10278 = ~n10271 & n10277;
  assign n10279 = ~n4133 & n10174;
  assign n10280 = n10278 & ~n10279;
  assign n10281 = n10270 & n10280;
  assign n10282 = n10249 & n10281;
  assign n10283 = n10246 & n10282;
  assign po0251 = ~n10240 | ~n10283;
  assign n10285 = pi0094 & n4043;
  assign n10286 = n2930 & n10285;
  assign n10287 = pi0094 & ~n3553;
  assign n10288 = n4497 & n10287;
  assign n10289 = ~n10286 & ~n10288;
  assign n10290 = pi0094 & ~pi0314;
  assign n10291 = ~n4402 & n10290;
  assign n10292 = n10289 & ~n10291;
  assign n10293 = pi0094 & n2726;
  assign n10294 = n4066 & n10293;
  assign n10295 = pi0024 & pi0094;
  assign n10296 = n2591 & n10295;
  assign n10297 = ~n10294 & ~n10296;
  assign n10298 = pi0094 & pi0841;
  assign n10299 = n2644 & n10298;
  assign n10300 = n2910 & n10295;
  assign n10301 = n3033 & n10295;
  assign n10302 = pi1044 & n10290;
  assign n10303 = n2619 & n10302;
  assign n10304 = pi0094 & n4504;
  assign n10305 = ~n10303 & ~n10304;
  assign n10306 = ~n10301 & n10305;
  assign n10307 = ~n10300 & n10306;
  assign n10308 = n3042 & n10295;
  assign n10309 = n10307 & ~n10308;
  assign n10310 = ~n10299 & n10309;
  assign n10311 = n10297 & n10310;
  assign n10312 = pi0094 & n4006;
  assign n10313 = pi0094 & ~n4014;
  assign n10314 = n3110 & n10295;
  assign n10315 = ~n10313 & ~n10314;
  assign n10316 = pi0094 & po0740;
  assign n10317 = n2651 & n10316;
  assign n10318 = ~n3102 & n10317;
  assign n10319 = n10315 & ~n10318;
  assign n10320 = ~n10312 & n10319;
  assign n10321 = n10311 & n10320;
  assign n10322 = n2917 & n10298;
  assign n10323 = n2913 & n10295;
  assign n10324 = ~n10322 & ~n10323;
  assign n10325 = n2936 & n10290;
  assign n10326 = n10324 & ~n10325;
  assign n10327 = n10321 & n10326;
  assign n10328 = n10292 & n10327;
  assign n10329 = ~n3998 & n10298;
  assign n10330 = pi0094 & n4336;
  assign n10331 = pi0094 & n4062;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = ~n10329 & n10332;
  assign n10334 = pi0094 & n4708;
  assign n10335 = ~n3973 & n10334;
  assign n10336 = pi0094 & n3989;
  assign n10337 = ~n10295 & ~n10336;
  assign n10338 = n2563 & ~n10337;
  assign n10339 = n2795 & n10295;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = pi0094 & n2741;
  assign n10342 = n10340 & ~n10341;
  assign n10343 = ~n10335 & n10342;
  assign n10344 = n10333 & n10343;
  assign n10345 = n2788 & n10295;
  assign n10346 = n2834 & n10302;
  assign n10347 = ~n10345 & ~n10346;
  assign n10348 = ~n4326 & n10295;
  assign n10349 = n10347 & ~n10348;
  assign n10350 = n2851 & n10290;
  assign n10351 = n3066 & n10295;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = ~n4077 & n10298;
  assign n10354 = n2681 & n10295;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356 = pi0094 & n4091;
  assign n10357 = ~n4097 & n10316;
  assign n10358 = pi0094 & n4459;
  assign n10359 = ~n10357 & ~n10358;
  assign n10360 = n3397 & ~n10359;
  assign n10361 = pi0094 & ~pi0786;
  assign n10362 = n4088 & n10361;
  assign n10363 = ~n10360 & ~n10362;
  assign n10364 = ~n10356 & n10363;
  assign n10365 = n4087 & ~n10364;
  assign n10366 = n2901 & n10290;
  assign n10367 = n3057 & n10295;
  assign n10368 = pi0094 & ~n3057;
  assign n10369 = ~n10367 & ~n10368;
  assign n10370 = n4083 & ~n10369;
  assign n10371 = ~n10366 & ~n10370;
  assign n10372 = ~n10365 & n10371;
  assign n10373 = n10355 & n10372;
  assign n10374 = ~pi0094 & pi0841;
  assign n10375 = n2847 & ~n10374;
  assign n10376 = n2881 & n10316;
  assign n10377 = n2726 & n10376;
  assign n10378 = pi0094 & n4124;
  assign n10379 = n2858 & n10298;
  assign n10380 = ~n10378 & ~n10379;
  assign n10381 = ~n10377 & n10380;
  assign n10382 = ~n10375 & n10381;
  assign n10383 = ~n4133 & n10298;
  assign n10384 = n10382 & ~n10383;
  assign n10385 = n10373 & n10384;
  assign n10386 = n10352 & n10385;
  assign n10387 = n10349 & n10386;
  assign n10388 = pi0094 & n4579;
  assign n10389 = ~n4105 & n10290;
  assign n10390 = n2569 & n10295;
  assign n10391 = ~n10389 & ~n10390;
  assign n10392 = n2598 & n10295;
  assign n10393 = n10391 & ~n10392;
  assign n10394 = ~n10388 & n10393;
  assign n10395 = n10387 & n10394;
  assign n10396 = n10344 & n10395;
  assign po0252 = ~n10328 | ~n10396;
  assign n10398 = pi0095 & n4091;
  assign n10399 = ~n7899 & ~n7900;
  assign n10400 = n4094 & ~n10399;
  assign n10401 = ~pi0095 & ~n4094;
  assign n10402 = ~n10400 & ~n10401;
  assign n10403 = n3128 & n10402;
  assign n10404 = pi0095 & po0740;
  assign n10405 = ~n4097 & n10404;
  assign n10406 = ~n10403 & ~n10405;
  assign n10407 = n3397 & ~n10406;
  assign n10408 = pi0095 & ~pi0786;
  assign n10409 = n4088 & n10408;
  assign n10410 = ~n10407 & ~n10409;
  assign n10411 = ~n10398 & n10410;
  assign n10412 = n3547 & ~n10411;
  assign n10413 = n3406 & n10412;
  assign n10414 = pi0024 & pi0095;
  assign n10415 = n3057 & n10414;
  assign n10416 = pi0095 & ~n3057;
  assign n10417 = ~n10415 & ~n10416;
  assign n10418 = n4083 & ~n10417;
  assign n10419 = ~n10413 & ~n10418;
  assign n10420 = pi0095 & pi0841;
  assign n10421 = ~pi0332 & ~pi0841;
  assign n10422 = ~n10420 & ~n10421;
  assign n10423 = n2770 & ~n10422;
  assign n10424 = n10419 & ~n10423;
  assign n10425 = pi0095 & ~pi0314;
  assign n10426 = n2901 & n10425;
  assign n10427 = n10424 & ~n10426;
  assign n10428 = n2681 & n10414;
  assign n10429 = n2892 & n10420;
  assign n10430 = ~n10428 & ~n10429;
  assign n10431 = n2858 & n10420;
  assign n10432 = pi0095 & n4124;
  assign n10433 = n2854 & n10414;
  assign n10434 = n2881 & n10404;
  assign n10435 = n2726 & n10434;
  assign n10436 = ~n10433 & ~n10435;
  assign n10437 = ~n10432 & n10436;
  assign n10438 = ~n10431 & n10437;
  assign n10439 = ~n4133 & n10420;
  assign n10440 = n10438 & ~n10439;
  assign n10441 = n2847 & n10420;
  assign n10442 = pi1044 & n10425;
  assign n10443 = n2834 & n10442;
  assign n10444 = ~n10441 & ~n10443;
  assign n10445 = ~n3072 & n10414;
  assign n10446 = n10444 & ~n10445;
  assign n10447 = n2851 & n10425;
  assign n10448 = n3066 & n10414;
  assign n10449 = ~n10447 & ~n10448;
  assign n10450 = n10446 & n10449;
  assign n10451 = n10440 & n10450;
  assign n10452 = n10430 & n10451;
  assign n10453 = n10427 & n10452;
  assign n10454 = pi0095 & n4067;
  assign n10455 = n2910 & n10414;
  assign n10456 = n2651 & n10404;
  assign n10457 = ~n3102 & n10456;
  assign n10458 = pi0095 & n4006;
  assign n10459 = ~n10457 & ~n10458;
  assign n10460 = pi0095 & ~n4014;
  assign n10461 = n3110 & n10414;
  assign n10462 = ~n10460 & ~n10461;
  assign n10463 = n10459 & n10462;
  assign n10464 = ~n10455 & n10463;
  assign n10465 = ~n10454 & n10464;
  assign n10466 = n2917 & n10420;
  assign n10467 = n2913 & n10414;
  assign n10468 = ~n10466 & ~n10467;
  assign n10469 = n2936 & n10425;
  assign n10470 = n10468 & ~n10469;
  assign n10471 = pi0095 & n4043;
  assign n10472 = n2930 & n10471;
  assign n10473 = pi0095 & ~n3553;
  assign n10474 = n4497 & n10473;
  assign n10475 = ~n10472 & ~n10474;
  assign n10476 = ~n4402 & n10425;
  assign n10477 = n10475 & ~n10476;
  assign n10478 = n3042 & n10414;
  assign n10479 = pi0095 & n4504;
  assign n10480 = ~n10478 & ~n10479;
  assign n10481 = n10477 & n10480;
  assign n10482 = n10470 & n10481;
  assign n10483 = n3033 & n10414;
  assign n10484 = n10482 & ~n10483;
  assign n10485 = n2591 & n10414;
  assign n10486 = pi0095 & pi0993;
  assign n10487 = n2576 & n10486;
  assign n10488 = n2598 & n10414;
  assign n10489 = ~n10487 & ~n10488;
  assign n10490 = ~n4105 & n10425;
  assign n10491 = n2569 & n10414;
  assign n10492 = ~n10490 & ~n10491;
  assign n10493 = n2619 & n10442;
  assign n10494 = n2644 & n10420;
  assign n10495 = ~n10493 & ~n10494;
  assign n10496 = n10492 & n10495;
  assign n10497 = n10489 & n10496;
  assign n10498 = ~n10485 & n10497;
  assign n10499 = pi0095 & ~n4061;
  assign n10500 = n4060 & n10499;
  assign n10501 = n10498 & ~n10500;
  assign n10502 = pi0095 & n2741;
  assign n10503 = pi0095 & n4708;
  assign n10504 = ~n3973 & n10503;
  assign n10505 = ~n3998 & n10420;
  assign n10506 = pi0095 & n3989;
  assign n10507 = ~n10414 & ~n10506;
  assign n10508 = n2563 & ~n10507;
  assign n10509 = n2795 & n10414;
  assign n10510 = ~n10508 & ~n10509;
  assign n10511 = ~n10505 & n10510;
  assign n10512 = ~n10504 & n10511;
  assign n10513 = ~n10502 & n10512;
  assign n10514 = n10501 & n10513;
  assign n10515 = pi0095 & n2604;
  assign n10516 = n3967 & n10515;
  assign n10517 = n10514 & ~n10516;
  assign n10518 = n10484 & n10517;
  assign n10519 = n10465 & n10518;
  assign po0253 = ~n10453 | ~n10519;
  assign n10521 = pi0096 & n4336;
  assign n10522 = pi0096 & n2741;
  assign n10523 = pi0096 & n4708;
  assign n10524 = ~n3973 & n10523;
  assign n10525 = pi0096 & pi0841;
  assign n10526 = ~n3998 & n10525;
  assign n10527 = pi0024 & pi0096;
  assign n10528 = pi0096 & n3989;
  assign n10529 = ~n10527 & ~n10528;
  assign n10530 = n2563 & ~n10529;
  assign n10531 = n2795 & n10527;
  assign n10532 = ~n10530 & ~n10531;
  assign n10533 = ~n10526 & n10532;
  assign n10534 = ~n10524 & n10533;
  assign n10535 = ~n10522 & n10534;
  assign n10536 = pi0096 & ~n4061;
  assign n10537 = n4060 & n10536;
  assign n10538 = n10535 & ~n10537;
  assign n10539 = pi0096 & ~pi0314;
  assign n10540 = ~n4105 & n10539;
  assign n10541 = n2569 & n10527;
  assign n10542 = ~n10540 & ~n10541;
  assign n10543 = pi0096 & pi0993;
  assign n10544 = n2576 & n10543;
  assign n10545 = n2598 & n10527;
  assign n10546 = ~n10544 & ~n10545;
  assign n10547 = n10542 & n10546;
  assign n10548 = pi0096 & n4067;
  assign n10549 = n2917 & n10525;
  assign n10550 = n2913 & n10527;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = n2936 & n10539;
  assign n10553 = n10551 & ~n10552;
  assign n10554 = pi0096 & n4043;
  assign n10555 = n2930 & n10554;
  assign n10556 = pi0096 & ~n3553;
  assign n10557 = n4497 & n10556;
  assign n10558 = ~n10555 & ~n10557;
  assign n10559 = ~n4402 & n10539;
  assign n10560 = n10558 & ~n10559;
  assign n10561 = n3042 & n10527;
  assign n10562 = pi0096 & n4504;
  assign n10563 = ~n10561 & ~n10562;
  assign n10564 = n10560 & n10563;
  assign n10565 = n10553 & n10564;
  assign n10566 = n3033 & n10527;
  assign n10567 = n10565 & ~n10566;
  assign n10568 = n2910 & n10527;
  assign n10569 = n10567 & ~n10568;
  assign n10570 = ~n10548 & n10569;
  assign n10571 = pi0096 & ~n3018;
  assign n10572 = ~po0740 & n10571;
  assign n10573 = pi0479 & n10572;
  assign n10574 = pi0096 & po0740;
  assign n10575 = ~n10573 & ~n10574;
  assign n10576 = n8326 & ~n10575;
  assign n10577 = n3110 & n10527;
  assign n10578 = ~n10576 & ~n10577;
  assign n10579 = pi0096 & ~n4014;
  assign n10580 = pi1044 & n10539;
  assign n10581 = n2619 & n10580;
  assign n10582 = n2644 & n10525;
  assign n10583 = ~n10581 & ~n10582;
  assign n10584 = n2591 & n10527;
  assign n10585 = n10583 & ~n10584;
  assign n10586 = ~n10579 & n10585;
  assign n10587 = n10578 & n10586;
  assign n10588 = n10570 & n10587;
  assign n10589 = n10547 & n10588;
  assign n10590 = n10538 & n10589;
  assign n10591 = ~n10521 & n10590;
  assign n10592 = pi0096 & n4089;
  assign n10593 = pi0096 & n4091;
  assign n10594 = pi0096 & n3128;
  assign n10595 = ~n4094 & n10594;
  assign n10596 = ~n4097 & n10574;
  assign n10597 = ~n10595 & ~n10596;
  assign n10598 = n3397 & ~n10597;
  assign n10599 = ~n10593 & ~n10598;
  assign n10600 = ~n10592 & n10599;
  assign n10601 = n4087 & ~n10600;
  assign n10602 = pi0024 & ~pi0096;
  assign n10603 = n2681 & ~n10602;
  assign n10604 = n3057 & ~n10527;
  assign n10605 = ~pi0096 & ~n3057;
  assign n10606 = ~n10604 & ~n10605;
  assign n10607 = n4083 & n10606;
  assign n10608 = ~n10603 & ~n10607;
  assign n10609 = ~n3072 & n10527;
  assign n10610 = n2847 & n10525;
  assign n10611 = n2834 & n10580;
  assign n10612 = ~n10610 & ~n10611;
  assign n10613 = n2858 & n10525;
  assign n10614 = pi0096 & n4124;
  assign n10615 = n2854 & n10527;
  assign n10616 = n2881 & n10574;
  assign n10617 = n2726 & n10616;
  assign n10618 = ~n10615 & ~n10617;
  assign n10619 = ~n10614 & n10618;
  assign n10620 = ~n10613 & n10619;
  assign n10621 = ~n4133 & n10525;
  assign n10622 = n10620 & ~n10621;
  assign n10623 = n2851 & n10539;
  assign n10624 = n3066 & n10527;
  assign n10625 = ~n10623 & ~n10624;
  assign n10626 = n10622 & n10625;
  assign n10627 = n10612 & n10626;
  assign n10628 = ~n10609 & n10627;
  assign n10629 = ~n4077 & n10525;
  assign n10630 = n2901 & n10539;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = n10628 & n10631;
  assign n10633 = n10608 & n10632;
  assign n10634 = ~n10601 & n10633;
  assign po0254 = ~n10591 | ~n10634;
  assign n10636 = pi0097 & n4336;
  assign n10637 = pi0097 & n2741;
  assign n10638 = pi0097 & n4708;
  assign n10639 = ~n3973 & n10638;
  assign n10640 = pi0097 & pi0841;
  assign n10641 = ~n3998 & n10640;
  assign n10642 = pi0024 & pi0097;
  assign n10643 = pi0097 & n3989;
  assign n10644 = ~n10642 & ~n10643;
  assign n10645 = n2563 & ~n10644;
  assign n10646 = n2795 & n10642;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = ~n10641 & n10647;
  assign n10649 = ~n10639 & n10648;
  assign n10650 = ~n10637 & n10649;
  assign n10651 = pi0097 & ~n4061;
  assign n10652 = n4060 & n10651;
  assign n10653 = n10650 & ~n10652;
  assign n10654 = pi0097 & ~pi0314;
  assign n10655 = ~n4105 & n10654;
  assign n10656 = n2569 & n10642;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = pi0097 & pi0993;
  assign n10659 = n2576 & n10658;
  assign n10660 = n2598 & n10642;
  assign n10661 = ~n10659 & ~n10660;
  assign n10662 = n10657 & n10661;
  assign n10663 = pi0097 & n4067;
  assign n10664 = pi0097 & n4043;
  assign n10665 = n2930 & n10664;
  assign n10666 = pi0097 & ~n3553;
  assign n10667 = n4497 & n10666;
  assign n10668 = ~n10665 & ~n10667;
  assign n10669 = n2917 & n10640;
  assign n10670 = n2913 & n10642;
  assign n10671 = ~n10669 & ~n10670;
  assign n10672 = n3042 & n10642;
  assign n10673 = pi0097 & ~pi1076;
  assign n10674 = n2926 & n10673;
  assign n10675 = ~n10672 & ~n10674;
  assign n10676 = n2936 & n10654;
  assign n10677 = ~n4402 & n10654;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = n10675 & n10678;
  assign n10680 = n10671 & n10679;
  assign n10681 = n10668 & n10680;
  assign n10682 = n3033 & n10642;
  assign n10683 = n10681 & ~n10682;
  assign n10684 = n2910 & n10642;
  assign n10685 = n10683 & ~n10684;
  assign n10686 = ~n10663 & n10685;
  assign n10687 = pi0097 & ~n4014;
  assign n10688 = n3110 & n10642;
  assign n10689 = ~n10687 & ~n10688;
  assign n10690 = pi0097 & po0740;
  assign n10691 = n2651 & n10690;
  assign n10692 = ~n3102 & n10691;
  assign n10693 = pi0097 & n4006;
  assign n10694 = ~n10692 & ~n10693;
  assign n10695 = pi1044 & n10654;
  assign n10696 = n2619 & n10695;
  assign n10697 = n2644 & n10640;
  assign n10698 = ~n10696 & ~n10697;
  assign n10699 = n2591 & n10642;
  assign n10700 = n10698 & ~n10699;
  assign n10701 = n10694 & n10700;
  assign n10702 = n10689 & n10701;
  assign n10703 = n10686 & n10702;
  assign n10704 = n10662 & n10703;
  assign n10705 = n10653 & n10704;
  assign n10706 = ~n10636 & n10705;
  assign n10707 = pi0097 & n4089;
  assign n10708 = pi0097 & n4091;
  assign n10709 = ~n4097 & n10690;
  assign n10710 = pi0097 & ~n4094;
  assign n10711 = n4094 & n7900;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = n3128 & ~n10712;
  assign n10714 = ~n10709 & ~n10713;
  assign n10715 = n3397 & ~n10714;
  assign n10716 = ~n10708 & ~n10715;
  assign n10717 = ~n10707 & n10716;
  assign n10718 = n4087 & ~n10717;
  assign n10719 = n3057 & n10642;
  assign n10720 = pi0097 & ~n3057;
  assign n10721 = ~n10719 & ~n10720;
  assign n10722 = n4083 & ~n10721;
  assign n10723 = n2901 & n10654;
  assign n10724 = ~n10722 & ~n10723;
  assign n10725 = ~n3072 & n10642;
  assign n10726 = n2847 & n10640;
  assign n10727 = n2834 & n10695;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = n2858 & n10640;
  assign n10730 = pi0097 & n4124;
  assign n10731 = n2854 & n10642;
  assign n10732 = n2881 & n10690;
  assign n10733 = n2726 & n10732;
  assign n10734 = ~n10731 & ~n10733;
  assign n10735 = ~n10730 & n10734;
  assign n10736 = ~n10729 & n10735;
  assign n10737 = ~n4133 & n10640;
  assign n10738 = n10736 & ~n10737;
  assign n10739 = n2851 & n10654;
  assign n10740 = n3066 & n10642;
  assign n10741 = ~n10739 & ~n10740;
  assign n10742 = n10738 & n10741;
  assign n10743 = n10728 & n10742;
  assign n10744 = ~n10725 & n10743;
  assign n10745 = n2681 & n10642;
  assign n10746 = ~n4077 & n10640;
  assign n10747 = ~n10745 & ~n10746;
  assign n10748 = n10744 & n10747;
  assign n10749 = n10724 & n10748;
  assign n10750 = ~n10718 & n10749;
  assign po0255 = ~n10706 | ~n10750;
  assign n10752 = pi0098 & ~pi0314;
  assign n10753 = ~n4105 & n10752;
  assign n10754 = pi0024 & pi0098;
  assign n10755 = n2569 & n10754;
  assign n10756 = ~n10753 & ~n10755;
  assign n10757 = pi0098 & pi0993;
  assign n10758 = n2576 & n10757;
  assign n10759 = n2598 & n10754;
  assign n10760 = ~n10758 & ~n10759;
  assign n10761 = n10756 & n10760;
  assign n10762 = pi0098 & n4060;
  assign n10763 = ~n4061 & n10762;
  assign n10764 = pi0098 & n4523;
  assign n10765 = ~n3973 & n10764;
  assign n10766 = pi0098 & n2741;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = ~n10763 & n10767;
  assign n10769 = pi0098 & pi0841;
  assign n10770 = ~n3998 & n10769;
  assign n10771 = pi0098 & n3989;
  assign n10772 = ~n10754 & ~n10771;
  assign n10773 = n2563 & ~n10772;
  assign n10774 = n2795 & n10754;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = ~n10770 & n10775;
  assign n10777 = pi0098 & n2604;
  assign n10778 = n3967 & n10777;
  assign n10779 = n10776 & ~n10778;
  assign n10780 = pi0098 & n4067;
  assign n10781 = pi0098 & n4043;
  assign n10782 = n2930 & n10781;
  assign n10783 = pi0098 & ~n3553;
  assign n10784 = n4497 & n10783;
  assign n10785 = ~n10782 & ~n10784;
  assign n10786 = n2917 & n10769;
  assign n10787 = n2913 & n10754;
  assign n10788 = ~n10786 & ~n10787;
  assign n10789 = n3042 & n10754;
  assign n10790 = pi0098 & ~pi1076;
  assign n10791 = n2926 & n10790;
  assign n10792 = ~n10789 & ~n10791;
  assign n10793 = n2936 & n10752;
  assign n10794 = ~n4402 & n10752;
  assign n10795 = ~n10793 & ~n10794;
  assign n10796 = n10792 & n10795;
  assign n10797 = n10788 & n10796;
  assign n10798 = n10785 & n10797;
  assign n10799 = n3033 & n10754;
  assign n10800 = n10798 & ~n10799;
  assign n10801 = n2910 & n10754;
  assign n10802 = n10800 & ~n10801;
  assign n10803 = ~n10780 & n10802;
  assign n10804 = ~pi0098 & ~pi0314;
  assign n10805 = pi1044 & ~n10804;
  assign n10806 = n2619 & n10805;
  assign n10807 = pi0098 & ~n4014;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = pi0098 & po0740;
  assign n10810 = n2651 & n10809;
  assign n10811 = ~n3102 & n10810;
  assign n10812 = pi0098 & n4006;
  assign n10813 = ~n10811 & ~n10812;
  assign n10814 = n2644 & n10769;
  assign n10815 = n2591 & n10754;
  assign n10816 = ~n10814 & ~n10815;
  assign n10817 = n3110 & n10754;
  assign n10818 = n10816 & ~n10817;
  assign n10819 = n10813 & n10818;
  assign n10820 = n10808 & n10819;
  assign n10821 = n10803 & n10820;
  assign n10822 = n10779 & n10821;
  assign n10823 = n10768 & n10822;
  assign n10824 = n10761 & n10823;
  assign n10825 = n2847 & n10769;
  assign n10826 = n2788 & n10754;
  assign n10827 = ~n10825 & ~n10826;
  assign n10828 = ~n4326 & n10754;
  assign n10829 = n10827 & ~n10828;
  assign n10830 = n2851 & n10752;
  assign n10831 = n3066 & n10754;
  assign n10832 = ~n10830 & ~n10831;
  assign n10833 = ~n4077 & n10769;
  assign n10834 = n2681 & n10754;
  assign n10835 = ~n10833 & ~n10834;
  assign n10836 = pi0098 & n4091;
  assign n10837 = ~n4097 & n10809;
  assign n10838 = pi0098 & n4459;
  assign n10839 = ~n10837 & ~n10838;
  assign n10840 = n3397 & ~n10839;
  assign n10841 = pi0098 & ~pi0786;
  assign n10842 = n4088 & n10841;
  assign n10843 = ~n10840 & ~n10842;
  assign n10844 = ~n10836 & n10843;
  assign n10845 = n4087 & ~n10844;
  assign n10846 = n2901 & n10752;
  assign n10847 = n3057 & n10754;
  assign n10848 = pi0098 & ~n3057;
  assign n10849 = ~n10847 & ~n10848;
  assign n10850 = n4083 & ~n10849;
  assign n10851 = ~n10846 & ~n10850;
  assign n10852 = ~n10845 & n10851;
  assign n10853 = n10835 & n10852;
  assign n10854 = n2858 & n10769;
  assign n10855 = pi0098 & n4124;
  assign n10856 = n2834 & n10805;
  assign n10857 = n2881 & n10809;
  assign n10858 = n2726 & n10857;
  assign n10859 = ~n10856 & ~n10858;
  assign n10860 = ~n10855 & n10859;
  assign n10861 = ~n10854 & n10860;
  assign n10862 = ~n4133 & n10769;
  assign n10863 = n10861 & ~n10862;
  assign n10864 = n10853 & n10863;
  assign n10865 = n10832 & n10864;
  assign n10866 = n10829 & n10865;
  assign po0256 = ~n10824 | ~n10866;
  assign n10868 = pi0099 & ~n4941;
  assign n10869 = ~n4953 & ~n10868;
  assign n10870 = n4939 & ~n10869;
  assign n10871 = pi0099 & ~n4939;
  assign n10872 = ~n10870 & ~n10871;
  assign n10873 = ~pi0039 & ~pi0072;
  assign n10874 = ~n10872 & n10873;
  assign n10875 = ~pi0072 & ~n4219;
  assign n10876 = pi0039 & n10875;
  assign n10877 = n4923 & n10876;
  assign po0257 = n10874 | n10877;
  assign n10879 = pi0100 & n4006;
  assign n10880 = pi0100 & ~n4014;
  assign n10881 = pi0024 & pi0100;
  assign n10882 = n3110 & n10881;
  assign n10883 = ~n10880 & ~n10882;
  assign n10884 = pi0100 & po0740;
  assign n10885 = n2651 & n10884;
  assign n10886 = ~n3102 & n10885;
  assign n10887 = n10883 & ~n10886;
  assign n10888 = ~n10879 & n10887;
  assign n10889 = n2591 & n10881;
  assign n10890 = n10888 & ~n10889;
  assign n10891 = pi0100 & ~pi0314;
  assign n10892 = pi1044 & n10891;
  assign n10893 = n2619 & n10892;
  assign n10894 = pi0100 & pi0841;
  assign n10895 = n2644 & n10894;
  assign n10896 = ~n10893 & ~n10895;
  assign n10897 = pi0100 & n4523;
  assign n10898 = ~n3973 & n10897;
  assign n10899 = pi0100 & n3989;
  assign n10900 = ~n10881 & ~n10899;
  assign n10901 = n2563 & ~n10900;
  assign n10902 = n2795 & n10881;
  assign n10903 = ~n10901 & ~n10902;
  assign n10904 = pi0100 & n2741;
  assign n10905 = n10903 & ~n10904;
  assign n10906 = ~n10898 & n10905;
  assign n10907 = ~n3998 & n10894;
  assign n10908 = n10906 & ~n10907;
  assign n10909 = pi0100 & n4336;
  assign n10910 = n10908 & ~n10909;
  assign n10911 = n10896 & n10910;
  assign n10912 = n10890 & n10911;
  assign n10913 = n2910 & n10881;
  assign n10914 = pi0100 & n4067;
  assign n10915 = pi0100 & n4062;
  assign n10916 = n2936 & n10891;
  assign n10917 = n2913 & n10881;
  assign n10918 = n2917 & n10894;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = ~pi0024 & ~n4026;
  assign n10921 = po0840 & n10920;
  assign n10922 = ~n10881 & ~n10921;
  assign n10923 = n3042 & ~n10922;
  assign n10924 = pi0100 & ~pi1076;
  assign n10925 = n2926 & n10924;
  assign n10926 = ~n10923 & ~n10925;
  assign n10927 = pi0100 & n4043;
  assign n10928 = n2930 & n10927;
  assign n10929 = pi0100 & ~n3553;
  assign n10930 = n4497 & n10929;
  assign n10931 = ~n10928 & ~n10930;
  assign n10932 = ~n4402 & n10891;
  assign n10933 = n10931 & ~n10932;
  assign n10934 = n10926 & n10933;
  assign n10935 = n10919 & n10934;
  assign n10936 = ~n10916 & n10935;
  assign n10937 = n3033 & n10881;
  assign n10938 = n10936 & ~n10937;
  assign n10939 = ~n10915 & n10938;
  assign n10940 = ~n10914 & n10939;
  assign n10941 = ~n10913 & n10940;
  assign n10942 = n2681 & n10881;
  assign n10943 = ~n4077 & n10894;
  assign n10944 = ~n10942 & ~n10943;
  assign n10945 = n2901 & n10891;
  assign n10946 = n3057 & n10881;
  assign n10947 = pi0100 & ~n3057;
  assign n10948 = ~n10946 & ~n10947;
  assign n10949 = n4083 & ~n10948;
  assign n10950 = ~n10945 & ~n10949;
  assign n10951 = pi0100 & n4089;
  assign n10952 = pi0100 & n4091;
  assign n10953 = pi0100 & n3128;
  assign n10954 = ~n4094 & n10953;
  assign n10955 = ~n4097 & n10884;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = n3397 & ~n10956;
  assign n10958 = ~n10952 & ~n10957;
  assign n10959 = ~n10951 & n10958;
  assign n10960 = n4087 & ~n10959;
  assign n10961 = n10950 & ~n10960;
  assign n10962 = ~n4105 & n10891;
  assign n10963 = n2569 & n10881;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = pi0100 & pi0993;
  assign n10966 = n2576 & n10965;
  assign n10967 = n2598 & n10881;
  assign n10968 = ~n10966 & ~n10967;
  assign n10969 = n10964 & n10968;
  assign n10970 = n10961 & n10969;
  assign n10971 = n10944 & n10970;
  assign n10972 = ~n3072 & n10881;
  assign n10973 = n2847 & n10894;
  assign n10974 = n2834 & n10892;
  assign n10975 = ~n10973 & ~n10974;
  assign n10976 = n2858 & n10894;
  assign n10977 = pi0100 & n4124;
  assign n10978 = n2854 & n10881;
  assign n10979 = n2881 & n10884;
  assign n10980 = n2726 & n10979;
  assign n10981 = ~n10978 & ~n10980;
  assign n10982 = ~n10977 & n10981;
  assign n10983 = ~n10976 & n10982;
  assign n10984 = ~n4133 & n10894;
  assign n10985 = n10983 & ~n10984;
  assign n10986 = n2851 & n10891;
  assign n10987 = n3066 & n10881;
  assign n10988 = ~n10986 & ~n10987;
  assign n10989 = n10985 & n10988;
  assign n10990 = n10975 & n10989;
  assign n10991 = ~n10972 & n10990;
  assign n10992 = n10971 & n10991;
  assign n10993 = n10941 & n10992;
  assign po0258 = ~n10912 | ~n10993;
  assign n10995 = pi0044 & pi0101;
  assign n10996 = ~n4940 & ~n10995;
  assign n10997 = n4939 & ~n10996;
  assign n10998 = pi0101 & ~n4939;
  assign n10999 = ~n10997 & ~n10998;
  assign n11000 = n10873 & ~n10999;
  assign n11001 = n5009 & n10876;
  assign po0259 = n11000 | n11001;
  assign n11003 = pi0102 & n4062;
  assign n11004 = pi0024 & pi0102;
  assign n11005 = n2569 & n11004;
  assign n11006 = ~n11003 & ~n11005;
  assign n11007 = pi0102 & ~pi0314;
  assign n11008 = ~n4105 & n11007;
  assign n11009 = n11006 & ~n11008;
  assign n11010 = pi1044 & n11007;
  assign n11011 = n2619 & n11010;
  assign n11012 = pi0102 & pi0841;
  assign n11013 = n2644 & n11012;
  assign n11014 = ~n11011 & ~n11013;
  assign n11015 = pi0102 & n4006;
  assign n11016 = pi0102 & ~n4014;
  assign n11017 = n3110 & n11004;
  assign n11018 = ~n11016 & ~n11017;
  assign n11019 = pi0102 & po0740;
  assign n11020 = n2651 & n11019;
  assign n11021 = ~n3102 & n11020;
  assign n11022 = n11018 & ~n11021;
  assign n11023 = ~n11015 & n11022;
  assign n11024 = n2591 & n11004;
  assign n11025 = n11023 & ~n11024;
  assign n11026 = ~n2556 & n11025;
  assign n11027 = n11014 & n11026;
  assign n11028 = pi0102 & n4089;
  assign n11029 = pi0102 & n4091;
  assign n11030 = pi0102 & n3128;
  assign n11031 = ~n4094 & n11030;
  assign n11032 = ~n4097 & n11019;
  assign n11033 = ~n11031 & ~n11032;
  assign n11034 = n3397 & ~n11033;
  assign n11035 = ~n11029 & ~n11034;
  assign n11036 = ~n11028 & n11035;
  assign n11037 = n4087 & ~n11036;
  assign n11038 = n11027 & ~n11037;
  assign n11039 = pi0102 & n3989;
  assign n11040 = ~n11004 & ~n11039;
  assign n11041 = n2563 & ~n11040;
  assign n11042 = n2795 & n11004;
  assign n11043 = ~n11041 & ~n11042;
  assign n11044 = pi0102 & n4708;
  assign n11045 = ~n3973 & n11044;
  assign n11046 = pi0102 & n2741;
  assign n11047 = ~n11045 & ~n11046;
  assign n11048 = n11043 & n11047;
  assign n11049 = ~n3998 & n11012;
  assign n11050 = n11048 & ~n11049;
  assign n11051 = pi0102 & pi0993;
  assign n11052 = n2576 & n11051;
  assign n11053 = n2598 & n11004;
  assign n11054 = ~n11052 & ~n11053;
  assign n11055 = n11050 & n11054;
  assign n11056 = n2910 & n11004;
  assign n11057 = pi0102 & n2726;
  assign n11058 = n4066 & n11057;
  assign n11059 = ~n11056 & ~n11058;
  assign n11060 = n2851 & n11007;
  assign n11061 = n3066 & n11004;
  assign n11062 = ~n11060 & ~n11061;
  assign n11063 = n2858 & n11012;
  assign n11064 = pi0102 & n4124;
  assign n11065 = n2854 & n11004;
  assign n11066 = n2881 & n11019;
  assign n11067 = n2726 & n11066;
  assign n11068 = ~n11065 & ~n11067;
  assign n11069 = ~n11064 & n11068;
  assign n11070 = ~n11063 & n11069;
  assign n11071 = ~n4133 & n11012;
  assign n11072 = n11070 & ~n11071;
  assign n11073 = n2917 & n11012;
  assign n11074 = n2913 & n11004;
  assign n11075 = ~n11073 & ~n11074;
  assign n11076 = n2936 & n11007;
  assign n11077 = n11075 & ~n11076;
  assign n11078 = pi0102 & n4043;
  assign n11079 = n2930 & n11078;
  assign n11080 = pi0102 & ~n3553;
  assign n11081 = n4497 & n11080;
  assign n11082 = ~n11079 & ~n11081;
  assign n11083 = ~n4402 & n11007;
  assign n11084 = n11082 & ~n11083;
  assign n11085 = n3042 & n11004;
  assign n11086 = pi0102 & n4504;
  assign n11087 = ~n11085 & ~n11086;
  assign n11088 = n11084 & n11087;
  assign n11089 = n11077 & n11088;
  assign n11090 = n3033 & n11004;
  assign n11091 = n11089 & ~n11090;
  assign n11092 = n11072 & n11091;
  assign n11093 = n11062 & n11092;
  assign n11094 = n11059 & n11093;
  assign n11095 = n11055 & n11094;
  assign n11096 = ~n4077 & n11012;
  assign n11097 = ~n3072 & n11004;
  assign n11098 = n2681 & n11004;
  assign n11099 = n2847 & n11012;
  assign n11100 = n2834 & n11010;
  assign n11101 = ~n11099 & ~n11100;
  assign n11102 = ~n11098 & n11101;
  assign n11103 = ~n11097 & n11102;
  assign n11104 = ~n11096 & n11103;
  assign n11105 = n2901 & n11007;
  assign n11106 = n3057 & n11004;
  assign n11107 = pi0102 & ~n3057;
  assign n11108 = ~n11106 & ~n11107;
  assign n11109 = n4083 & ~n11108;
  assign n11110 = ~n11105 & ~n11109;
  assign n11111 = n11104 & n11110;
  assign n11112 = pi0102 & n4336;
  assign n11113 = n11111 & ~n11112;
  assign n11114 = n11095 & n11113;
  assign n11115 = n11038 & n11114;
  assign po0260 = ~n11009 | ~n11115;
  assign n11117 = pi0103 & n4062;
  assign n11118 = pi0024 & pi0103;
  assign n11119 = n2569 & n11118;
  assign n11120 = ~n11117 & ~n11119;
  assign n11121 = pi0103 & ~pi0314;
  assign n11122 = ~n4105 & n11121;
  assign n11123 = n11120 & ~n11122;
  assign n11124 = pi1044 & n11121;
  assign n11125 = n2619 & n11124;
  assign n11126 = pi0103 & pi0841;
  assign n11127 = n2644 & n11126;
  assign n11128 = ~n11125 & ~n11127;
  assign n11129 = pi0103 & n4006;
  assign n11130 = pi0103 & ~n4014;
  assign n11131 = n3110 & n11118;
  assign n11132 = ~n11130 & ~n11131;
  assign n11133 = pi0103 & po0740;
  assign n11134 = n2651 & n11133;
  assign n11135 = ~n3102 & n11134;
  assign n11136 = n11132 & ~n11135;
  assign n11137 = ~n11129 & n11136;
  assign n11138 = n2591 & n11118;
  assign n11139 = n11137 & ~n11138;
  assign n11140 = ~n2637 & n11139;
  assign n11141 = n11128 & n11140;
  assign n11142 = pi0103 & n4089;
  assign n11143 = pi0103 & n4091;
  assign n11144 = pi0103 & n3128;
  assign n11145 = ~n4094 & n11144;
  assign n11146 = ~n4097 & n11133;
  assign n11147 = ~n11145 & ~n11146;
  assign n11148 = n3397 & ~n11147;
  assign n11149 = ~n11143 & ~n11148;
  assign n11150 = ~n11142 & n11149;
  assign n11151 = n4087 & ~n11150;
  assign n11152 = n11141 & ~n11151;
  assign n11153 = pi0103 & n3989;
  assign n11154 = ~n11118 & ~n11153;
  assign n11155 = n2563 & ~n11154;
  assign n11156 = n2795 & n11118;
  assign n11157 = ~n11155 & ~n11156;
  assign n11158 = pi0103 & n4708;
  assign n11159 = ~n3973 & n11158;
  assign n11160 = pi0103 & n2741;
  assign n11161 = ~n11159 & ~n11160;
  assign n11162 = n11157 & n11161;
  assign n11163 = ~n3998 & n11126;
  assign n11164 = n11162 & ~n11163;
  assign n11165 = pi0103 & pi0993;
  assign n11166 = n2576 & n11165;
  assign n11167 = n2598 & n11118;
  assign n11168 = ~n11166 & ~n11167;
  assign n11169 = n11164 & n11168;
  assign n11170 = n2910 & n11118;
  assign n11171 = pi0103 & n2726;
  assign n11172 = n4066 & n11171;
  assign n11173 = ~n11170 & ~n11172;
  assign n11174 = n2851 & n11121;
  assign n11175 = n3066 & n11118;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = n2858 & n11126;
  assign n11178 = pi0103 & n4124;
  assign n11179 = n2854 & n11118;
  assign n11180 = n2881 & n11133;
  assign n11181 = n2726 & n11180;
  assign n11182 = ~n11179 & ~n11181;
  assign n11183 = ~n11178 & n11182;
  assign n11184 = ~n11177 & n11183;
  assign n11185 = ~n4133 & n11126;
  assign n11186 = n11184 & ~n11185;
  assign n11187 = n2917 & n11126;
  assign n11188 = n2913 & n11118;
  assign n11189 = ~n11187 & ~n11188;
  assign n11190 = n2936 & n11121;
  assign n11191 = n11189 & ~n11190;
  assign n11192 = pi0103 & n4043;
  assign n11193 = n2930 & n11192;
  assign n11194 = pi0103 & ~n3553;
  assign n11195 = n4497 & n11194;
  assign n11196 = ~n11193 & ~n11195;
  assign n11197 = ~n4402 & n11121;
  assign n11198 = n11196 & ~n11197;
  assign n11199 = n3042 & n11118;
  assign n11200 = pi0103 & n4504;
  assign n11201 = ~n11199 & ~n11200;
  assign n11202 = n11198 & n11201;
  assign n11203 = n11191 & n11202;
  assign n11204 = n3033 & n11118;
  assign n11205 = n11203 & ~n11204;
  assign n11206 = n11186 & n11205;
  assign n11207 = n11176 & n11206;
  assign n11208 = n11173 & n11207;
  assign n11209 = n11169 & n11208;
  assign n11210 = ~n4077 & n11126;
  assign n11211 = ~n3072 & n11118;
  assign n11212 = n2681 & n11118;
  assign n11213 = n2847 & n11126;
  assign n11214 = n2834 & n11124;
  assign n11215 = ~n11213 & ~n11214;
  assign n11216 = ~n11212 & n11215;
  assign n11217 = ~n11211 & n11216;
  assign n11218 = ~n11210 & n11217;
  assign n11219 = n2901 & n11121;
  assign n11220 = n3057 & n11118;
  assign n11221 = pi0103 & ~n3057;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = n4083 & ~n11222;
  assign n11224 = ~n11219 & ~n11223;
  assign n11225 = n11218 & n11224;
  assign n11226 = pi0103 & n4336;
  assign n11227 = n11225 & ~n11226;
  assign n11228 = n11209 & n11227;
  assign n11229 = n11152 & n11228;
  assign po0261 = ~n11123 | ~n11229;
  assign n11231 = pi0104 & n4062;
  assign n11232 = pi0104 & n4523;
  assign n11233 = ~n3973 & n11232;
  assign n11234 = pi0024 & pi0104;
  assign n11235 = pi0104 & n3989;
  assign n11236 = ~n11234 & ~n11235;
  assign n11237 = n2563 & ~n11236;
  assign n11238 = n2795 & n11234;
  assign n11239 = ~n11237 & ~n11238;
  assign n11240 = pi0104 & n2741;
  assign n11241 = n11239 & ~n11240;
  assign n11242 = ~n11233 & n11241;
  assign n11243 = pi0104 & pi0841;
  assign n11244 = ~n3998 & n11243;
  assign n11245 = n11242 & ~n11244;
  assign n11246 = ~pi0104 & n3967;
  assign n11247 = n2604 & ~n11246;
  assign n11248 = n11245 & ~n11247;
  assign n11249 = ~n11231 & n11248;
  assign n11250 = pi0104 & n4006;
  assign n11251 = pi0104 & ~n4014;
  assign n11252 = n3110 & n11234;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = pi0104 & po0740;
  assign n11255 = n2651 & n11254;
  assign n11256 = ~n3102 & n11255;
  assign n11257 = n11253 & ~n11256;
  assign n11258 = ~n11250 & n11257;
  assign n11259 = n2591 & n11234;
  assign n11260 = n11258 & ~n11259;
  assign n11261 = pi0104 & ~pi0314;
  assign n11262 = pi1044 & n11261;
  assign n11263 = n2619 & n11262;
  assign n11264 = n2644 & n11243;
  assign n11265 = ~n11263 & ~n11264;
  assign n11266 = n2917 & n11243;
  assign n11267 = n2913 & n11234;
  assign n11268 = ~n11266 & ~n11267;
  assign n11269 = n2936 & n11261;
  assign n11270 = n11268 & ~n11269;
  assign n11271 = n3042 & n11234;
  assign n11272 = pi0104 & n4043;
  assign n11273 = n2930 & n11272;
  assign n11274 = pi0104 & ~n3553;
  assign n11275 = n4497 & n11274;
  assign n11276 = ~n11273 & ~n11275;
  assign n11277 = ~n4402 & n11261;
  assign n11278 = n11276 & ~n11277;
  assign n11279 = pi0104 & n4504;
  assign n11280 = n11278 & ~n11279;
  assign n11281 = ~n11271 & n11280;
  assign n11282 = n11270 & n11281;
  assign n11283 = n3033 & n11234;
  assign n11284 = n11282 & ~n11283;
  assign n11285 = n2910 & n11234;
  assign n11286 = pi0104 & n2726;
  assign n11287 = n4066 & n11286;
  assign n11288 = ~n11285 & ~n11287;
  assign n11289 = n11284 & n11288;
  assign n11290 = n11265 & n11289;
  assign n11291 = n11260 & n11290;
  assign n11292 = n2681 & n11234;
  assign n11293 = ~n4077 & n11243;
  assign n11294 = ~n11292 & ~n11293;
  assign n11295 = n2901 & n11261;
  assign n11296 = n3057 & n11234;
  assign n11297 = pi0104 & ~n3057;
  assign n11298 = ~n11296 & ~n11297;
  assign n11299 = n4083 & ~n11298;
  assign n11300 = ~n11295 & ~n11299;
  assign n11301 = pi0104 & n4089;
  assign n11302 = pi0104 & n4091;
  assign n11303 = pi0104 & n3128;
  assign n11304 = ~n4094 & n11303;
  assign n11305 = ~n4097 & n11254;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = n3397 & ~n11306;
  assign n11308 = ~n11302 & ~n11307;
  assign n11309 = ~n11301 & n11308;
  assign n11310 = n4087 & ~n11309;
  assign n11311 = n11300 & ~n11310;
  assign n11312 = ~n4105 & n11261;
  assign n11313 = n2569 & n11234;
  assign n11314 = ~n11312 & ~n11313;
  assign n11315 = pi0104 & pi0993;
  assign n11316 = n2576 & n11315;
  assign n11317 = n2598 & n11234;
  assign n11318 = ~n11316 & ~n11317;
  assign n11319 = n11314 & n11318;
  assign n11320 = n11311 & n11319;
  assign n11321 = n11294 & n11320;
  assign n11322 = ~n3072 & n11234;
  assign n11323 = n2847 & n11243;
  assign n11324 = n2834 & n11262;
  assign n11325 = ~n11323 & ~n11324;
  assign n11326 = n2858 & n11243;
  assign n11327 = pi0104 & n4124;
  assign n11328 = n2854 & n11234;
  assign n11329 = n2881 & n11254;
  assign n11330 = n2726 & n11329;
  assign n11331 = ~n11328 & ~n11330;
  assign n11332 = ~n11327 & n11331;
  assign n11333 = ~n11326 & n11332;
  assign n11334 = ~n4133 & n11243;
  assign n11335 = n11333 & ~n11334;
  assign n11336 = n2851 & n11261;
  assign n11337 = n3066 & n11234;
  assign n11338 = ~n11336 & ~n11337;
  assign n11339 = n11335 & n11338;
  assign n11340 = n11325 & n11339;
  assign n11341 = ~n11322 & n11340;
  assign n11342 = n11321 & n11341;
  assign n11343 = n11291 & n11342;
  assign po0262 = ~n11249 | ~n11343;
  assign n11345 = pi0106 & pi0841;
  assign n11346 = n2847 & n11345;
  assign n11347 = pi0106 & ~pi0314;
  assign n11348 = pi1044 & n11347;
  assign n11349 = n2834 & n11348;
  assign n11350 = ~n11346 & ~n11349;
  assign n11351 = pi0024 & pi0106;
  assign n11352 = ~n3072 & n11351;
  assign n11353 = n11350 & ~n11352;
  assign n11354 = n2851 & n11347;
  assign n11355 = n3066 & n11351;
  assign n11356 = ~n11354 & ~n11355;
  assign n11357 = pi0106 & n2741;
  assign n11358 = pi0106 & n4523;
  assign n11359 = ~n3973 & n11358;
  assign n11360 = ~n3998 & n11345;
  assign n11361 = pi0106 & n3989;
  assign n11362 = ~n11351 & ~n11361;
  assign n11363 = n2563 & ~n11362;
  assign n11364 = n2795 & n11351;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 = ~n11360 & n11365;
  assign n11367 = ~n11359 & n11366;
  assign n11368 = ~n11357 & n11367;
  assign n11369 = n2619 & n11348;
  assign n11370 = n2644 & n11345;
  assign n11371 = ~n11369 & ~n11370;
  assign n11372 = pi0106 & n4336;
  assign n11373 = pi0106 & n4006;
  assign n11374 = pi0106 & ~n4014;
  assign n11375 = n3110 & n11351;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = pi0106 & po0740;
  assign n11378 = n2651 & n11377;
  assign n11379 = ~n3102 & n11378;
  assign n11380 = n11376 & ~n11379;
  assign n11381 = ~n11373 & n11380;
  assign n11382 = n2591 & n11351;
  assign n11383 = n11381 & ~n11382;
  assign n11384 = ~n11372 & n11383;
  assign n11385 = n11371 & n11384;
  assign n11386 = n11368 & n11385;
  assign n11387 = pi0024 & ~pi0106;
  assign n11388 = n2598 & ~n11387;
  assign n11389 = pi0106 & n4062;
  assign n11390 = n2910 & n11351;
  assign n11391 = pi0106 & n4067;
  assign n11392 = n2662 & n11347;
  assign n11393 = n3033 & n11351;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = pi0106 & n4504;
  assign n11396 = n3042 & n11351;
  assign n11397 = ~n11395 & ~n11396;
  assign n11398 = pi0106 & n5491;
  assign n11399 = pi0106 & ~n3553;
  assign n11400 = n4497 & n11399;
  assign n11401 = n2917 & n11345;
  assign n11402 = n2913 & n11351;
  assign n11403 = ~n11401 & ~n11402;
  assign n11404 = n2936 & n11347;
  assign n11405 = n11403 & ~n11404;
  assign n11406 = ~n4402 & n11347;
  assign n11407 = n11405 & ~n11406;
  assign n11408 = ~n11400 & n11407;
  assign n11409 = ~n11398 & n11408;
  assign n11410 = n11397 & n11409;
  assign n11411 = n11394 & n11410;
  assign n11412 = ~n11391 & n11411;
  assign n11413 = ~n11390 & n11412;
  assign n11414 = n2656 & n11347;
  assign n11415 = n11413 & ~n11414;
  assign n11416 = pi0106 & pi0993;
  assign n11417 = n2576 & n11416;
  assign n11418 = n2569 & n11351;
  assign n11419 = ~n11417 & ~n11418;
  assign n11420 = n11415 & n11419;
  assign n11421 = ~n11389 & n11420;
  assign n11422 = ~n11388 & n11421;
  assign n11423 = n11386 & n11422;
  assign n11424 = pi0106 & n4089;
  assign n11425 = pi0106 & n4091;
  assign n11426 = pi0106 & n3128;
  assign n11427 = ~n4094 & n11426;
  assign n11428 = ~n4097 & n11377;
  assign n11429 = ~n11427 & ~n11428;
  assign n11430 = n3397 & ~n11429;
  assign n11431 = ~n11425 & ~n11430;
  assign n11432 = ~n11424 & n11431;
  assign n11433 = n4087 & ~n11432;
  assign n11434 = n3057 & n11351;
  assign n11435 = pi0106 & ~n3057;
  assign n11436 = ~n11434 & ~n11435;
  assign n11437 = n4083 & ~n11436;
  assign n11438 = n2901 & n11347;
  assign n11439 = ~n11437 & ~n11438;
  assign n11440 = n2881 & n11377;
  assign n11441 = n2726 & n11440;
  assign n11442 = n2854 & n11351;
  assign n11443 = ~n11441 & ~n11442;
  assign n11444 = n2858 & n11345;
  assign n11445 = pi0106 & n4124;
  assign n11446 = ~n11444 & ~n11445;
  assign n11447 = n11443 & n11446;
  assign n11448 = n2681 & n11351;
  assign n11449 = ~n4077 & n11345;
  assign n11450 = ~n11448 & ~n11449;
  assign n11451 = n11447 & n11450;
  assign n11452 = n11439 & n11451;
  assign n11453 = ~n11433 & n11452;
  assign n11454 = ~n4133 & n11345;
  assign n11455 = n11453 & ~n11454;
  assign n11456 = n11423 & n11455;
  assign n11457 = n11356 & n11456;
  assign po0264 = ~n11353 | ~n11457;
  assign n11459 = pi0107 & pi0841;
  assign n11460 = n2847 & n11459;
  assign n11461 = pi0107 & ~pi0314;
  assign n11462 = pi1044 & n11461;
  assign n11463 = n2834 & n11462;
  assign n11464 = ~n11460 & ~n11463;
  assign n11465 = pi0024 & pi0107;
  assign n11466 = ~n3072 & n11465;
  assign n11467 = n11464 & ~n11466;
  assign n11468 = n2851 & n11461;
  assign n11469 = n3066 & n11465;
  assign n11470 = ~n11468 & ~n11469;
  assign n11471 = pi0107 & n2741;
  assign n11472 = pi0107 & n4523;
  assign n11473 = ~n3973 & n11472;
  assign n11474 = ~n3998 & n11459;
  assign n11475 = pi0107 & n3989;
  assign n11476 = ~n11465 & ~n11475;
  assign n11477 = n2563 & ~n11476;
  assign n11478 = n2795 & n11465;
  assign n11479 = ~n11477 & ~n11478;
  assign n11480 = ~n11474 & n11479;
  assign n11481 = ~n11473 & n11480;
  assign n11482 = ~n11471 & n11481;
  assign n11483 = n2662 & n11461;
  assign n11484 = n3033 & n11465;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486 = ~n2569 & ~n2598;
  assign n11487 = n11465 & ~n11486;
  assign n11488 = n2656 & n11461;
  assign n11489 = ~n11487 & ~n11488;
  assign n11490 = n2917 & n11459;
  assign n11491 = n2913 & n11465;
  assign n11492 = ~n11490 & ~n11491;
  assign n11493 = n2936 & n11461;
  assign n11494 = n11492 & ~n11493;
  assign n11495 = pi0107 & n4043;
  assign n11496 = n2930 & n11495;
  assign n11497 = pi0107 & ~n3553;
  assign n11498 = n4497 & n11497;
  assign n11499 = ~n11496 & ~n11498;
  assign n11500 = ~n4402 & n11461;
  assign n11501 = n11499 & ~n11500;
  assign n11502 = n3042 & n11465;
  assign n11503 = pi0107 & n4504;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = n11501 & n11504;
  assign n11506 = n11494 & n11505;
  assign n11507 = pi0107 & n4067;
  assign n11508 = n2910 & n11465;
  assign n11509 = ~n11507 & ~n11508;
  assign n11510 = n11506 & n11509;
  assign n11511 = n11489 & n11510;
  assign n11512 = n11485 & n11511;
  assign n11513 = n11482 & n11512;
  assign n11514 = ~pi0107 & pi0993;
  assign n11515 = n2576 & ~n11514;
  assign n11516 = pi0107 & n4062;
  assign n11517 = pi0107 & n4336;
  assign n11518 = pi0107 & n4006;
  assign n11519 = pi0107 & ~n4014;
  assign n11520 = n3110 & n11465;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = pi0107 & po0740;
  assign n11523 = n2651 & n11522;
  assign n11524 = ~n3102 & n11523;
  assign n11525 = n11521 & ~n11524;
  assign n11526 = ~n11518 & n11525;
  assign n11527 = n2591 & n11465;
  assign n11528 = n11526 & ~n11527;
  assign n11529 = n2619 & n11462;
  assign n11530 = n2644 & n11459;
  assign n11531 = ~n11529 & ~n11530;
  assign n11532 = n11528 & n11531;
  assign n11533 = ~n11517 & n11532;
  assign n11534 = ~n11516 & n11533;
  assign n11535 = ~n11515 & n11534;
  assign n11536 = n11513 & n11535;
  assign n11537 = pi0107 & n4089;
  assign n11538 = pi0107 & n4091;
  assign n11539 = pi0107 & n3128;
  assign n11540 = ~n4094 & n11539;
  assign n11541 = ~n4097 & n11522;
  assign n11542 = ~n11540 & ~n11541;
  assign n11543 = n3397 & ~n11542;
  assign n11544 = ~n11538 & ~n11543;
  assign n11545 = ~n11537 & n11544;
  assign n11546 = n4087 & ~n11545;
  assign n11547 = n3057 & n11465;
  assign n11548 = pi0107 & ~n3057;
  assign n11549 = ~n11547 & ~n11548;
  assign n11550 = n4083 & ~n11549;
  assign n11551 = n2901 & n11461;
  assign n11552 = ~n11550 & ~n11551;
  assign n11553 = n2881 & n11522;
  assign n11554 = n2726 & n11553;
  assign n11555 = n2854 & n11465;
  assign n11556 = ~n11554 & ~n11555;
  assign n11557 = n2858 & n11459;
  assign n11558 = pi0107 & n4124;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = n11556 & n11559;
  assign n11561 = n2681 & n11465;
  assign n11562 = ~n4077 & n11459;
  assign n11563 = ~n11561 & ~n11562;
  assign n11564 = n11560 & n11563;
  assign n11565 = n11552 & n11564;
  assign n11566 = ~n11546 & n11565;
  assign n11567 = ~n4133 & n11459;
  assign n11568 = n11566 & ~n11567;
  assign n11569 = n11536 & n11568;
  assign n11570 = n11470 & n11569;
  assign po0265 = ~n11467 | ~n11570;
  assign n11572 = pi0108 & n2741;
  assign n11573 = pi0108 & n4523;
  assign n11574 = ~n3973 & n11573;
  assign n11575 = pi0108 & pi0841;
  assign n11576 = ~n3998 & n11575;
  assign n11577 = pi0024 & pi0108;
  assign n11578 = pi0108 & n3989;
  assign n11579 = ~n11577 & ~n11578;
  assign n11580 = n2563 & ~n11579;
  assign n11581 = n2795 & n11577;
  assign n11582 = ~n11580 & ~n11581;
  assign n11583 = ~n11576 & n11582;
  assign n11584 = ~n11574 & n11583;
  assign n11585 = ~n11572 & n11584;
  assign n11586 = n2910 & n11577;
  assign n11587 = pi0108 & n4067;
  assign n11588 = pi0108 & n4504;
  assign n11589 = n3042 & n11577;
  assign n11590 = ~n11588 & ~n11589;
  assign n11591 = n3033 & n11577;
  assign n11592 = n11590 & ~n11591;
  assign n11593 = ~n2922 & n11592;
  assign n11594 = ~n11587 & n11593;
  assign n11595 = ~n11586 & n11594;
  assign n11596 = pi0108 & ~n4061;
  assign n11597 = n4060 & n11596;
  assign n11598 = n11595 & ~n11597;
  assign n11599 = ~n3072 & n11577;
  assign n11600 = n2847 & n11575;
  assign n11601 = pi0108 & ~pi0314;
  assign n11602 = pi1044 & n11601;
  assign n11603 = n2834 & n11602;
  assign n11604 = ~n11600 & ~n11603;
  assign n11605 = n2858 & n11575;
  assign n11606 = pi0108 & n4124;
  assign n11607 = n2854 & n11577;
  assign n11608 = pi0108 & po0740;
  assign n11609 = n2881 & n11608;
  assign n11610 = n2726 & n11609;
  assign n11611 = ~n11607 & ~n11610;
  assign n11612 = ~n11606 & n11611;
  assign n11613 = ~n11605 & n11612;
  assign n11614 = ~n4133 & n11575;
  assign n11615 = n11613 & ~n11614;
  assign n11616 = n2851 & n11601;
  assign n11617 = n3066 & n11577;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = n11615 & n11618;
  assign n11620 = n11604 & n11619;
  assign n11621 = ~n11599 & n11620;
  assign n11622 = pi0108 & n5491;
  assign n11623 = pi0108 & ~n3553;
  assign n11624 = n4497 & n11623;
  assign n11625 = n2917 & n11575;
  assign n11626 = n2913 & n11577;
  assign n11627 = ~n11625 & ~n11626;
  assign n11628 = n2936 & n11601;
  assign n11629 = n11627 & ~n11628;
  assign n11630 = ~n4402 & n11601;
  assign n11631 = n11629 & ~n11630;
  assign n11632 = ~n11624 & n11631;
  assign n11633 = ~n11622 & n11632;
  assign n11634 = pi0108 & n4579;
  assign n11635 = n2569 & n11577;
  assign n11636 = ~n11634 & ~n11635;
  assign n11637 = n11633 & n11636;
  assign n11638 = n11621 & n11637;
  assign n11639 = n2901 & n11601;
  assign n11640 = n3057 & n11577;
  assign n11641 = pi0108 & ~n3057;
  assign n11642 = ~n11640 & ~n11641;
  assign n11643 = n4083 & ~n11642;
  assign n11644 = ~n11639 & ~n11643;
  assign n11645 = pi0108 & n4089;
  assign n11646 = pi0108 & n4091;
  assign n11647 = pi0108 & n3128;
  assign n11648 = ~n4094 & n11647;
  assign n11649 = ~n4097 & n11608;
  assign n11650 = ~n11648 & ~n11649;
  assign n11651 = n3397 & ~n11650;
  assign n11652 = ~n11646 & ~n11651;
  assign n11653 = ~n11645 & n11652;
  assign n11654 = n4087 & ~n11653;
  assign n11655 = n11644 & ~n11654;
  assign n11656 = pi0108 & ~n4014;
  assign n11657 = n3110 & n11577;
  assign n11658 = ~n11656 & ~n11657;
  assign n11659 = n2651 & n11608;
  assign n11660 = ~n3102 & n11659;
  assign n11661 = pi0108 & n4006;
  assign n11662 = ~n11660 & ~n11661;
  assign n11663 = n2619 & n11602;
  assign n11664 = n2644 & n11575;
  assign n11665 = ~n11663 & ~n11664;
  assign n11666 = n2591 & n11577;
  assign n11667 = n11665 & ~n11666;
  assign n11668 = n11662 & n11667;
  assign n11669 = n11658 & n11668;
  assign n11670 = n2662 & n11601;
  assign n11671 = n11669 & ~n11670;
  assign n11672 = n11655 & n11671;
  assign n11673 = n2681 & n11577;
  assign n11674 = ~n4077 & n11575;
  assign n11675 = ~n11673 & ~n11674;
  assign n11676 = n2656 & n11601;
  assign n11677 = n2598 & n11577;
  assign n11678 = ~n11676 & ~n11677;
  assign n11679 = n11675 & n11678;
  assign n11680 = ~n2632 & n11679;
  assign n11681 = ~n2667 & n11680;
  assign n11682 = pi0108 & n4336;
  assign n11683 = n11681 & ~n11682;
  assign n11684 = n11672 & n11683;
  assign n11685 = n11638 & n11684;
  assign n11686 = n11598 & n11685;
  assign po0266 = ~n11585 | ~n11686;
  assign n11688 = pi0109 & pi0841;
  assign n11689 = n2847 & n11688;
  assign n11690 = pi0109 & ~pi0314;
  assign n11691 = pi1044 & n11690;
  assign n11692 = n2834 & n11691;
  assign n11693 = ~n11689 & ~n11692;
  assign n11694 = pi0024 & pi0109;
  assign n11695 = ~n3072 & n11694;
  assign n11696 = n11693 & ~n11695;
  assign n11697 = n2851 & n11690;
  assign n11698 = n3066 & n11694;
  assign n11699 = ~n11697 & ~n11698;
  assign n11700 = pi0109 & n2741;
  assign n11701 = pi0109 & n4523;
  assign n11702 = ~n3973 & n11701;
  assign n11703 = ~n3998 & n11688;
  assign n11704 = pi0109 & n3989;
  assign n11705 = ~n11694 & ~n11704;
  assign n11706 = n2563 & ~n11705;
  assign n11707 = n2795 & n11694;
  assign n11708 = ~n11706 & ~n11707;
  assign n11709 = ~n11703 & n11708;
  assign n11710 = ~n11702 & n11709;
  assign n11711 = ~n11700 & n11710;
  assign n11712 = n2619 & n11691;
  assign n11713 = n2644 & n11688;
  assign n11714 = ~n11712 & ~n11713;
  assign n11715 = pi0109 & n4336;
  assign n11716 = pi0109 & n4006;
  assign n11717 = pi0109 & ~n4014;
  assign n11718 = n3110 & n11694;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = pi0109 & po0740;
  assign n11721 = n2651 & n11720;
  assign n11722 = ~n3102 & n11721;
  assign n11723 = n11719 & ~n11722;
  assign n11724 = ~n11716 & n11723;
  assign n11725 = n2591 & n11694;
  assign n11726 = n11724 & ~n11725;
  assign n11727 = ~n11715 & n11726;
  assign n11728 = n11714 & n11727;
  assign n11729 = n11711 & n11728;
  assign n11730 = pi0109 & ~n4061;
  assign n11731 = n4060 & n11730;
  assign n11732 = pi0109 & n2656;
  assign n11733 = ~n11731 & ~n11732;
  assign n11734 = pi0314 & n2656;
  assign n11735 = n2910 & n11694;
  assign n11736 = pi0109 & n4067;
  assign n11737 = n2662 & n11690;
  assign n11738 = n3033 & n11694;
  assign n11739 = ~n11737 & ~n11738;
  assign n11740 = pi0109 & n4504;
  assign n11741 = n3042 & n11694;
  assign n11742 = ~n11740 & ~n11741;
  assign n11743 = pi0109 & n5491;
  assign n11744 = pi0109 & ~n3553;
  assign n11745 = n4497 & n11744;
  assign n11746 = n2917 & n11688;
  assign n11747 = n2913 & n11694;
  assign n11748 = ~n11746 & ~n11747;
  assign n11749 = n2936 & n11690;
  assign n11750 = n11748 & ~n11749;
  assign n11751 = ~n4402 & n11690;
  assign n11752 = n11750 & ~n11751;
  assign n11753 = ~n11745 & n11752;
  assign n11754 = ~n11743 & n11753;
  assign n11755 = n11742 & n11754;
  assign n11756 = n11739 & n11755;
  assign n11757 = ~n11736 & n11756;
  assign n11758 = ~n11735 & n11757;
  assign n11759 = n2569 & n11694;
  assign n11760 = n11758 & ~n11759;
  assign n11761 = pi0109 & pi0993;
  assign n11762 = n2576 & n11761;
  assign n11763 = n2598 & n11694;
  assign n11764 = ~n11762 & ~n11763;
  assign n11765 = n11760 & n11764;
  assign n11766 = ~n11734 & n11765;
  assign n11767 = n11733 & n11766;
  assign n11768 = n11729 & n11767;
  assign n11769 = pi0109 & n4089;
  assign n11770 = pi0109 & n4091;
  assign n11771 = pi0109 & n3128;
  assign n11772 = ~n4094 & n11771;
  assign n11773 = ~n4097 & n11720;
  assign n11774 = ~n11772 & ~n11773;
  assign n11775 = n3397 & ~n11774;
  assign n11776 = ~n11770 & ~n11775;
  assign n11777 = ~n11769 & n11776;
  assign n11778 = n4087 & ~n11777;
  assign n11779 = n3057 & n11694;
  assign n11780 = pi0109 & ~n3057;
  assign n11781 = ~n11779 & ~n11780;
  assign n11782 = n4083 & ~n11781;
  assign n11783 = n2901 & n11690;
  assign n11784 = ~n11782 & ~n11783;
  assign n11785 = n2881 & n11720;
  assign n11786 = n2726 & n11785;
  assign n11787 = n2854 & n11694;
  assign n11788 = ~n11786 & ~n11787;
  assign n11789 = n2858 & n11688;
  assign n11790 = pi0109 & n4124;
  assign n11791 = ~n11789 & ~n11790;
  assign n11792 = n11788 & n11791;
  assign n11793 = n2681 & n11694;
  assign n11794 = ~n4077 & n11688;
  assign n11795 = ~n11793 & ~n11794;
  assign n11796 = n11792 & n11795;
  assign n11797 = n11784 & n11796;
  assign n11798 = ~n11778 & n11797;
  assign n11799 = ~n4133 & n11688;
  assign n11800 = n11798 & ~n11799;
  assign n11801 = n11768 & n11800;
  assign n11802 = n11699 & n11801;
  assign po0267 = ~n11696 | ~n11802;
  assign n11804 = pi0110 & pi0841;
  assign n11805 = n2847 & n11804;
  assign n11806 = pi0110 & ~pi0314;
  assign n11807 = pi1044 & n11806;
  assign n11808 = n2834 & n11807;
  assign n11809 = ~n11805 & ~n11808;
  assign n11810 = pi0024 & pi0110;
  assign n11811 = ~n3072 & n11810;
  assign n11812 = n11809 & ~n11811;
  assign n11813 = n2851 & n11806;
  assign n11814 = n3066 & n11810;
  assign n11815 = ~n11813 & ~n11814;
  assign n11816 = pi0110 & n2741;
  assign n11817 = pi0110 & n5965;
  assign n11818 = ~n3998 & n11804;
  assign n11819 = pi0110 & n3989;
  assign n11820 = ~n11810 & ~n11819;
  assign n11821 = n2563 & ~n11820;
  assign n11822 = n2795 & n11810;
  assign n11823 = ~n11821 & ~n11822;
  assign n11824 = ~n11818 & n11823;
  assign n11825 = ~n11817 & n11824;
  assign n11826 = ~n11816 & n11825;
  assign n11827 = n2619 & n11807;
  assign n11828 = n2644 & n11804;
  assign n11829 = ~n11827 & ~n11828;
  assign n11830 = pi0110 & n4336;
  assign n11831 = pi0110 & n4006;
  assign n11832 = pi0110 & ~n4014;
  assign n11833 = n3110 & n11810;
  assign n11834 = ~n11832 & ~n11833;
  assign n11835 = pi0110 & po0740;
  assign n11836 = n2651 & n11835;
  assign n11837 = ~n3102 & n11836;
  assign n11838 = n11834 & ~n11837;
  assign n11839 = ~n11831 & n11838;
  assign n11840 = n2591 & n11810;
  assign n11841 = n11839 & ~n11840;
  assign n11842 = ~n11830 & n11841;
  assign n11843 = n11829 & n11842;
  assign n11844 = n11826 & n11843;
  assign n11845 = ~pi0110 & ~pi0314;
  assign n11846 = n2662 & ~n11845;
  assign n11847 = pi0110 & n4062;
  assign n11848 = n2910 & n11810;
  assign n11849 = pi0110 & n4067;
  assign n11850 = n2656 & n11806;
  assign n11851 = n3033 & n11810;
  assign n11852 = ~n11850 & ~n11851;
  assign n11853 = pi0110 & n4504;
  assign n11854 = n3042 & n11810;
  assign n11855 = ~n11853 & ~n11854;
  assign n11856 = pi0110 & n5491;
  assign n11857 = pi0110 & ~n3553;
  assign n11858 = n4497 & n11857;
  assign n11859 = n2917 & n11804;
  assign n11860 = n2913 & n11810;
  assign n11861 = ~n11859 & ~n11860;
  assign n11862 = n2936 & n11806;
  assign n11863 = n11861 & ~n11862;
  assign n11864 = ~n4402 & n11806;
  assign n11865 = n11863 & ~n11864;
  assign n11866 = ~n11858 & n11865;
  assign n11867 = ~n11856 & n11866;
  assign n11868 = n11855 & n11867;
  assign n11869 = n11852 & n11868;
  assign n11870 = ~n11849 & n11869;
  assign n11871 = ~n11848 & n11870;
  assign n11872 = n2569 & n11810;
  assign n11873 = n11871 & ~n11872;
  assign n11874 = pi0110 & pi0993;
  assign n11875 = n2576 & n11874;
  assign n11876 = n2598 & n11810;
  assign n11877 = ~n11875 & ~n11876;
  assign n11878 = n11873 & n11877;
  assign n11879 = ~n11847 & n11878;
  assign n11880 = ~n11846 & n11879;
  assign n11881 = n11844 & n11880;
  assign n11882 = pi0110 & n4089;
  assign n11883 = pi0110 & n4091;
  assign n11884 = pi0110 & n3128;
  assign n11885 = ~n4094 & n11884;
  assign n11886 = ~n4097 & n11835;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = n3397 & ~n11887;
  assign n11889 = ~n11883 & ~n11888;
  assign n11890 = ~n11882 & n11889;
  assign n11891 = n4087 & ~n11890;
  assign n11892 = n3057 & n11810;
  assign n11893 = pi0110 & ~n3057;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = n4083 & ~n11894;
  assign n11896 = n2901 & n11806;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = n2881 & n11835;
  assign n11899 = n2726 & n11898;
  assign n11900 = n2854 & n11810;
  assign n11901 = ~n11899 & ~n11900;
  assign n11902 = n2858 & n11804;
  assign n11903 = pi0110 & n4124;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = n11901 & n11904;
  assign n11906 = n2681 & n11810;
  assign n11907 = ~n4077 & n11804;
  assign n11908 = ~n11906 & ~n11907;
  assign n11909 = n11905 & n11908;
  assign n11910 = n11897 & n11909;
  assign n11911 = ~n11891 & n11910;
  assign n11912 = ~n4133 & n11804;
  assign n11913 = n11911 & ~n11912;
  assign n11914 = n11881 & n11913;
  assign n11915 = n11815 & n11914;
  assign po0268 = ~n11812 | ~n11915;
  assign n11917 = pi0111 & pi0841;
  assign n11918 = n2847 & n11917;
  assign n11919 = pi0111 & ~pi0314;
  assign n11920 = pi1044 & n11919;
  assign n11921 = n2834 & n11920;
  assign n11922 = ~n11918 & ~n11921;
  assign n11923 = pi0024 & pi0111;
  assign n11924 = ~n3072 & n11923;
  assign n11925 = n11922 & ~n11924;
  assign n11926 = n2851 & n11919;
  assign n11927 = n3066 & n11923;
  assign n11928 = ~n11926 & ~n11927;
  assign n11929 = pi0111 & n2741;
  assign n11930 = pi0111 & n4708;
  assign n11931 = ~n3973 & n11930;
  assign n11932 = ~n3998 & n11917;
  assign n11933 = pi0111 & n3989;
  assign n11934 = ~n11923 & ~n11933;
  assign n11935 = n2563 & ~n11934;
  assign n11936 = n2795 & n11923;
  assign n11937 = ~n11935 & ~n11936;
  assign n11938 = ~n11932 & n11937;
  assign n11939 = ~n11931 & n11938;
  assign n11940 = ~n11929 & n11939;
  assign n11941 = n2619 & n11920;
  assign n11942 = n2644 & n11917;
  assign n11943 = ~n11941 & ~n11942;
  assign n11944 = pi0111 & n4336;
  assign n11945 = pi0111 & n4006;
  assign n11946 = pi0111 & ~n4014;
  assign n11947 = n3110 & n11923;
  assign n11948 = ~n11946 & ~n11947;
  assign n11949 = pi0111 & po0740;
  assign n11950 = n2651 & n11949;
  assign n11951 = ~n3102 & n11950;
  assign n11952 = n11948 & ~n11951;
  assign n11953 = ~n11945 & n11952;
  assign n11954 = n2591 & n11923;
  assign n11955 = n11953 & ~n11954;
  assign n11956 = ~n11944 & n11955;
  assign n11957 = n11943 & n11956;
  assign n11958 = n11940 & n11957;
  assign n11959 = n2662 & n11919;
  assign n11960 = n3033 & n11923;
  assign n11961 = ~n11959 & ~n11960;
  assign n11962 = pi0111 & n4504;
  assign n11963 = n3042 & n11923;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = pi0111 & n5491;
  assign n11966 = pi0111 & ~n3553;
  assign n11967 = n4497 & n11966;
  assign n11968 = n2917 & n11917;
  assign n11969 = n2913 & n11923;
  assign n11970 = ~n11968 & ~n11969;
  assign n11971 = n2936 & n11919;
  assign n11972 = n11970 & ~n11971;
  assign n11973 = ~n4402 & n11919;
  assign n11974 = n11972 & ~n11973;
  assign n11975 = ~n11967 & n11974;
  assign n11976 = ~n11965 & n11975;
  assign n11977 = n11964 & n11976;
  assign n11978 = n2598 & n11923;
  assign n11979 = n2656 & n11919;
  assign n11980 = ~n11978 & ~n11979;
  assign n11981 = n2910 & n11923;
  assign n11982 = pi0111 & n4067;
  assign n11983 = ~n11981 & ~n11982;
  assign n11984 = n11980 & n11983;
  assign n11985 = pi0111 & n4060;
  assign n11986 = ~n4061 & n11985;
  assign n11987 = pi0111 & pi0993;
  assign n11988 = n2576 & n11987;
  assign n11989 = pi0024 & ~pi0111;
  assign n11990 = n2569 & ~n11989;
  assign n11991 = ~n11988 & ~n11990;
  assign n11992 = ~n11986 & n11991;
  assign n11993 = n11984 & n11992;
  assign n11994 = n11977 & n11993;
  assign n11995 = n11961 & n11994;
  assign n11996 = n11958 & n11995;
  assign n11997 = pi0111 & n4089;
  assign n11998 = pi0111 & n4091;
  assign n11999 = pi0111 & n3128;
  assign n12000 = ~n4094 & n11999;
  assign n12001 = ~n4097 & n11949;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = n3397 & ~n12002;
  assign n12004 = ~n11998 & ~n12003;
  assign n12005 = ~n11997 & n12004;
  assign n12006 = n4087 & ~n12005;
  assign n12007 = n3057 & n11923;
  assign n12008 = pi0111 & ~n3057;
  assign n12009 = ~n12007 & ~n12008;
  assign n12010 = n4083 & ~n12009;
  assign n12011 = n2901 & n11919;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = n2881 & n11949;
  assign n12014 = n2726 & n12013;
  assign n12015 = n2854 & n11923;
  assign n12016 = ~n12014 & ~n12015;
  assign n12017 = n2858 & n11917;
  assign n12018 = pi0111 & n4124;
  assign n12019 = ~n12017 & ~n12018;
  assign n12020 = n12016 & n12019;
  assign n12021 = n2681 & n11923;
  assign n12022 = ~n4077 & n11917;
  assign n12023 = ~n12021 & ~n12022;
  assign n12024 = n12020 & n12023;
  assign n12025 = n12012 & n12024;
  assign n12026 = ~n12006 & n12025;
  assign n12027 = ~n4133 & n11917;
  assign n12028 = n12026 & ~n12027;
  assign n12029 = n11996 & n12028;
  assign n12030 = n11928 & n12029;
  assign po0269 = ~n11925 | ~n12030;
  assign po0270 = ~pi0124 | pi0468;
  assign n12033 = pi0113 & n4953;
  assign n12034 = ~pi0113 & ~n4953;
  assign n12035 = ~n12033 & ~n12034;
  assign n12036 = n4939 & n12035;
  assign n12037 = pi0113 & ~n4939;
  assign n12038 = ~n12036 & ~n12037;
  assign po0271 = n10873 & ~n12038;
  assign n12040 = n2753 & n4941;
  assign n12041 = pi0114 & n12040;
  assign n12042 = ~pi0114 & ~n12040;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = n4939 & n12043;
  assign n12045 = pi0114 & ~n4939;
  assign n12046 = ~n12044 & ~n12045;
  assign po0272 = n10873 & ~n12046;
  assign n12048 = pi0115 & n5837;
  assign n12049 = ~pi0115 & ~n5837;
  assign n12050 = ~n12048 & ~n12049;
  assign n12051 = n4939 & n12050;
  assign n12052 = pi0115 & ~n4939;
  assign n12053 = ~n12051 & ~n12052;
  assign po0273 = n10873 & ~n12053;
  assign n12055 = pi0116 & n4993;
  assign n12056 = ~pi0116 & ~n4993;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = n4939 & n12057;
  assign n12059 = pi0116 & ~n4939;
  assign n12060 = ~n12058 & ~n12059;
  assign po0274 = n10873 & ~n12060;
  assign n12062 = ~n2556 & n2585;
  assign n12063 = n2904 & n12062;
  assign n12064 = n2842 & n12063;
  assign n12065 = n2884 & n2943;
  assign n12066 = n2547 & n12065;
  assign n12067 = n2688 & n12066;
  assign n12068 = n12064 & n12067;
  assign po0275 = ~n2816 | ~n12068;
  assign n12070 = ~n4152 & ~n4171;
  assign n12071 = ~n3163 & n3481;
  assign n12072 = ~n4155 & ~n12071;
  assign n12073 = ~pi0185 & n2429;
  assign n12074 = ~pi0150 & ~n2429;
  assign n12075 = ~n12073 & ~n12074;
  assign n12076 = n3481 & n12075;
  assign n12077 = n4163 & ~n4182;
  assign n12078 = ~n12076 & n12077;
  assign n12079 = ~pi0143 & n2429;
  assign n12080 = ~pi0165 & ~n2429;
  assign n12081 = ~n12079 & ~n12080;
  assign n12082 = n3481 & n12081;
  assign n12083 = ~n4186 & ~n12082;
  assign n12084 = n4186 & n4198;
  assign n12085 = pi0118 & ~n8760;
  assign n12086 = ~pi0118 & n8760;
  assign n12087 = ~n12085 & ~n12086;
  assign n12088 = n4194 & ~n12087;
  assign n12089 = pi0118 & ~n4194;
  assign n12090 = ~n12088 & ~n12089;
  assign n12091 = n12084 & ~n12090;
  assign n12092 = ~n12083 & ~n12091;
  assign n12093 = n8753 & ~n12092;
  assign n12094 = n4163 & n12093;
  assign n12095 = ~n12078 & ~n12094;
  assign n12096 = n4162 & ~n12095;
  assign n12097 = ~n8748 & ~n8775;
  assign n12098 = n12076 & n12097;
  assign n12099 = ~n12076 & ~n12097;
  assign n12100 = ~n12098 & ~n12099;
  assign n12101 = n4162 & ~n12100;
  assign n12102 = ~n4163 & n12101;
  assign n12103 = ~n3481 & ~n4162;
  assign n12104 = ~n3271 & ~n4162;
  assign n12105 = ~n12103 & ~n12104;
  assign n12106 = ~n12102 & n12105;
  assign n12107 = ~n12096 & n12106;
  assign n12108 = n4155 & ~n12107;
  assign n12109 = ~n12072 & ~n12108;
  assign n12110 = n4152 & ~n12109;
  assign po0276 = n12070 | n12110;
  assign n12112 = pi0128 & pi0228;
  assign n12113 = ~n2740 & ~n3042;
  assign n12114 = ~n2656 & ~n2941;
  assign n12115 = ~n3549 & ~n10127;
  assign n12116 = ~n9440 & n12115;
  assign n12117 = n3397 & ~n12116;
  assign n12118 = n3467 & n12117;
  assign n12119 = ~n3498 & ~n12118;
  assign n12120 = ~n2619 & n12119;
  assign n12121 = ~n10024 & n12120;
  assign n12122 = ~n8472 & n12121;
  assign n12123 = n12114 & n12122;
  assign n12124 = ~n2563 & n12123;
  assign n12125 = n12113 & n12124;
  assign po0288 = n2826 | ~n12125;
  assign n12127 = ~pi0228 & po0288;
  assign po0277 = n12112 | n12127;
  assign n12129 = ~pi0031 & ~pi0080;
  assign n12130 = pi0818 & n12129;
  assign n12131 = pi0982 & n3539;
  assign n12132 = n2721 & n12131;
  assign n12133 = pi0951 & n12132;
  assign po0975 = n12130 | n12133;
  assign n12135 = pi1087 & po0975;
  assign n12136 = ~pi0120 & ~n12135;
  assign po0278 = ~po0280 & ~n12136;
  assign n12138 = ~n2656 & n2941;
  assign n12139 = pi0024 & n2656;
  assign n12140 = ~n12138 & ~n12139;
  assign n12141 = ~n8742 & ~n12140;
  assign n12142 = n11734 & n12140;
  assign n12143 = ~n3495 & n12142;
  assign n12144 = pi0087 & ~n11734;
  assign n12145 = ~n8748 & n12144;
  assign n12146 = ~pi0084 & n2476;
  assign n12147 = ~pi0068 & n12146;
  assign n12148 = ~n4272 & ~n12147;
  assign n12149 = ~pi0125 & ~pi0133;
  assign n12150 = ~pi0121 & n12149;
  assign n12151 = pi0121 & ~n12149;
  assign n12152 = ~n12150 & ~n12151;
  assign n12153 = ~pi0126 & ~pi0132;
  assign n12154 = n12150 & n12153;
  assign n12155 = ~pi0130 & n12154;
  assign n12156 = ~pi0136 & n12155;
  assign n12157 = ~pi0134 & ~pi0135;
  assign n12158 = n12156 & n12157;
  assign n12159 = ~n12152 & ~n12158;
  assign n12160 = n12147 & n12159;
  assign n12161 = ~n12148 & ~n12160;
  assign n12162 = ~pi0051 & ~pi0087;
  assign n12163 = ~n12161 & n12162;
  assign n12164 = pi0051 & ~n3481;
  assign n12165 = pi0051 & ~n2702;
  assign n12166 = ~n12164 & ~n12165;
  assign n12167 = ~pi0087 & ~n12166;
  assign n12168 = ~n12163 & ~n12167;
  assign n12169 = ~n11734 & ~n12168;
  assign n12170 = ~n12145 & ~n12169;
  assign n12171 = n12140 & ~n12170;
  assign n12172 = ~n12143 & ~n12171;
  assign n12173 = n2777 & n3402;
  assign n12174 = n2569 & ~n2777;
  assign n12175 = ~n12173 & ~n12174;
  assign n12176 = ~n3481 & ~n12140;
  assign n12177 = n12175 & ~n12176;
  assign n12178 = n12172 & n12177;
  assign n12179 = ~n12141 & n12178;
  assign n12180 = n2777 & n3398;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = ~n3486 & n12180;
  assign po0279 = n12181 | n12182;
  assign n12184 = pi0039 & pi0110;
  assign n12185 = ~pi0039 & ~pi0110;
  assign n12186 = ~n12184 & ~n12185;
  assign n12187 = ~n3967 & n12186;
  assign n12188 = ~n3469 & ~n8236;
  assign n12189 = n3397 & ~n12188;
  assign n12190 = n3466 & n12189;
  assign n12191 = n3464 & n12190;
  assign n12192 = n12187 & ~n12191;
  assign n12193 = ~pi0083 & n2868;
  assign n12194 = ~pi0067 & ~pi0085;
  assign n12195 = ~pi0069 & ~pi0071;
  assign n12196 = ~pi0087 & ~pi0109;
  assign n12197 = ~pi0077 & n12196;
  assign n12198 = ~pi0103 & n12197;
  assign n12199 = ~pi0072 & n12198;
  assign n12200 = ~pi0086 & n12199;
  assign n12201 = ~pi0036 & ~pi0110;
  assign n12202 = n2497 & n12201;
  assign n12203 = ~pi0073 & n12202;
  assign n12204 = ~pi0091 & n12203;
  assign n12205 = ~pi0090 & n2511;
  assign n12206 = ~pi0047 & n12205;
  assign n12207 = n12204 & n12206;
  assign n12208 = ~pi0111 & n12207;
  assign n12209 = n12200 & n12208;
  assign n12210 = n12195 & n12209;
  assign n12211 = n12194 & n12210;
  assign n12212 = n12193 & n12211;
  assign n12213 = ~pi0066 & n12212;
  assign n12214 = pi0081 & n12213;
  assign n12215 = n2862 & n12211;
  assign n12216 = ~pi0083 & n12215;
  assign n12217 = n2479 & n12216;
  assign n12218 = pi0067 & n12210;
  assign n12219 = ~pi0085 & n12218;
  assign n12220 = pi0071 & ~pi0085;
  assign n12221 = ~pi0069 & n12220;
  assign n12222 = pi0069 & n2971;
  assign n12223 = ~n12221 & ~n12222;
  assign n12224 = n12209 & ~n12223;
  assign n12225 = pi0085 & n12195;
  assign n12226 = n12209 & n12225;
  assign n12227 = ~n12224 & ~n12226;
  assign n12228 = pi0072 & ~n12208;
  assign n12229 = pi0111 & n12207;
  assign n12230 = n2511 & n2820;
  assign n12231 = pi0073 & n12205;
  assign n12232 = ~n12230 & ~n12231;
  assign n12233 = n3000 & ~n12232;
  assign n12234 = ~pi0111 & n2502;
  assign n12235 = n12233 & n12234;
  assign n12236 = ~n12229 & ~n12235;
  assign n12237 = ~pi0072 & n12236;
  assign n12238 = ~n12228 & ~n12237;
  assign n12239 = n2996 & n12238;
  assign n12240 = n2971 & n2995;
  assign n12241 = n12239 & n12240;
  assign n12242 = n12227 & ~n12241;
  assign n12243 = ~pi0067 & ~n12242;
  assign n12244 = ~n12219 & ~n12243;
  assign n12245 = ~pi0083 & ~n12244;
  assign n12246 = pi0083 & n12211;
  assign n12247 = ~n12245 & ~n12246;
  assign n12248 = n2481 & ~n12247;
  assign n12249 = ~n12217 & ~n12248;
  assign n12250 = pi0066 & n12212;
  assign n12251 = n12249 & ~n12250;
  assign n12252 = ~pi0081 & ~n12251;
  assign n12253 = ~n12214 & ~n12252;
  assign n12254 = ~pi0048 & ~pi0068;
  assign n12255 = ~n12253 & n12254;
  assign n12256 = pi0068 & ~pi0081;
  assign n12257 = ~pi0048 & n12256;
  assign n12258 = n12213 & n12257;
  assign n12259 = ~n12255 & ~n12258;
  assign n12260 = ~pi0059 & ~pi0062;
  assign n12261 = ~po1049 & n12260;
  assign n12262 = ~pi0065 & n2978;
  assign n12263 = n2983 & n12262;
  assign n12264 = n2962 & n12263;
  assign n12265 = ~pi0057 & n12264;
  assign n12266 = n12261 & n12265;
  assign n12267 = ~n12259 & n12266;
  assign n12268 = n2967 & n12267;
  assign n12269 = ~pi0074 & ~pi0094;
  assign n12270 = n2468 & n12269;
  assign n12271 = ~pi0096 & ~pi0097;
  assign n12272 = n12270 & n12271;
  assign n12273 = n4163 & n12272;
  assign n12274 = n12268 & n12273;
  assign n12275 = ~pi0045 & ~pi0055;
  assign n12276 = n2987 & n12275;
  assign n12277 = ~pi0038 & ~pi0053;
  assign n12278 = n2446 & n12277;
  assign n12279 = n12276 & n12278;
  assign n12280 = ~pi0056 & n12279;
  assign n12281 = n12274 & n12280;
  assign n12282 = ~n12186 & ~n12281;
  assign n12283 = pi0039 & ~pi0110;
  assign n12284 = n12187 & ~n12283;
  assign n12285 = ~pi0039 & pi0110;
  assign n12286 = ~n12191 & ~n12285;
  assign n12287 = n12186 & n12286;
  assign n12288 = ~n12284 & ~n12287;
  assign n12289 = ~n12282 & n12288;
  assign po0281 = n12192 | ~n12289;
  assign n12291 = ~n3495 & n12180;
  assign n12292 = ~n4219 & ~n12147;
  assign n12293 = pi0125 & pi0133;
  assign n12294 = ~n12149 & ~n12293;
  assign n12295 = n12147 & ~n12294;
  assign n12296 = ~n12158 & n12295;
  assign n12297 = ~n12292 & ~n12296;
  assign n12298 = n12162 & ~n12297;
  assign n12299 = pi0051 & ~n3186;
  assign n12300 = ~n12164 & ~n12299;
  assign n12301 = ~pi0087 & ~n12300;
  assign n12302 = ~n12298 & ~n12301;
  assign n12303 = ~n11734 & ~n12302;
  assign n12304 = ~n4238 & n12144;
  assign n12305 = ~n12303 & ~n12304;
  assign n12306 = n12140 & ~n12305;
  assign n12307 = ~n3482 & n12142;
  assign n12308 = ~n12306 & ~n12307;
  assign n12309 = ~n4232 & ~n12140;
  assign n12310 = n12308 & ~n12309;
  assign n12311 = ~n12176 & n12310;
  assign n12312 = n12175 & ~n12180;
  assign n12313 = ~n12311 & n12312;
  assign po0282 = n12291 | n12313;
  assign n12315 = ~n4171 & n12175;
  assign n12316 = ~n12140 & n12315;
  assign n12317 = ~n3486 & n12142;
  assign n12318 = ~n12076 & n12144;
  assign n12319 = ~n4922 & ~n12147;
  assign n12320 = pi0126 & ~n12150;
  assign n12321 = ~pi0126 & n12150;
  assign n12322 = ~n12320 & ~n12321;
  assign n12323 = ~n12158 & ~n12322;
  assign n12324 = pi0126 & n12158;
  assign n12325 = ~n12323 & ~n12324;
  assign n12326 = n12147 & ~n12325;
  assign n12327 = ~n12319 & ~n12326;
  assign n12328 = n12162 & ~n12327;
  assign n12329 = pi0051 & ~n2444;
  assign n12330 = ~n12164 & ~n12329;
  assign n12331 = ~pi0087 & ~n12330;
  assign n12332 = ~n12328 & ~n12331;
  assign n12333 = ~n11734 & ~n12332;
  assign n12334 = ~n12318 & ~n12333;
  assign n12335 = n12140 & ~n12334;
  assign n12336 = ~n12317 & ~n12335;
  assign n12337 = n12175 & ~n12336;
  assign n12338 = ~n12316 & ~n12337;
  assign n12339 = ~n12180 & ~n12338;
  assign n12340 = ~n3491 & n12180;
  assign po0283 = n12339 | n12340;
  assign n12342 = n3540 & ~n4058;
  assign n12343 = pi0250 & n12342;
  assign n12344 = ~po0740 & n12343;
  assign n12345 = pi0127 & ~n12343;
  assign n12346 = ~n12344 & ~n12345;
  assign n12347 = n2813 & ~n12346;
  assign n12348 = ~n2795 & n3998;
  assign n12349 = ~n2694 & n12348;
  assign n12350 = ~n2740 & ~n2813;
  assign n12351 = n2570 & n12350;
  assign n12352 = n3009 & n12351;
  assign n12353 = n12349 & n12352;
  assign n12354 = n2686 & n2903;
  assign n12355 = ~n2788 & ~n3066;
  assign n12356 = ~n2841 & n2883;
  assign n12357 = ~n3071 & n3418;
  assign n12358 = ~n2851 & n12357;
  assign n12359 = n2836 & n12358;
  assign n12360 = n12356 & n12359;
  assign n12361 = ~n2854 & n12360;
  assign n12362 = n12355 & n12361;
  assign n12363 = n2517 & n2534;
  assign n12364 = n2942 & n12363;
  assign n12365 = n2545 & n12364;
  assign n12366 = n3035 & n12365;
  assign n12367 = ~n2922 & ~n3042;
  assign n12368 = ~n2913 & ~n2930;
  assign n12369 = n12367 & n12368;
  assign n12370 = n12366 & n12369;
  assign n12371 = n2673 & ~n3110;
  assign n12372 = n12370 & n12371;
  assign n12373 = n5327 & n12372;
  assign n12374 = n12362 & n12373;
  assign n12375 = n12354 & n12374;
  assign n12376 = n2778 & n12375;
  assign n12377 = n12353 & n12376;
  assign n12378 = ~n2813 & ~n12377;
  assign n12379 = ~n12347 & ~n12378;
  assign po0284 = pi0129 & ~n12379;
  assign n12381 = n3540 & n4927;
  assign n12382 = pi0129 & ~n12381;
  assign n12383 = ~po0740 & n12381;
  assign n12384 = ~n12382 & ~n12383;
  assign n12385 = ~n2740 & n3042;
  assign n12386 = ~n12384 & n12385;
  assign n12387 = n2740 & n3042;
  assign n12388 = ~n12113 & ~n12387;
  assign n12389 = ~n2694 & n3998;
  assign n12390 = ~n2576 & n12389;
  assign n12391 = n12352 & n12390;
  assign n12392 = n12374 & n12391;
  assign n12393 = n2778 & n12392;
  assign n12394 = n12354 & n12393;
  assign n12395 = ~n12388 & ~n12394;
  assign n12396 = ~pi0250 & ~po0740;
  assign n12397 = pi0129 & pi0250;
  assign n12398 = ~n12396 & ~n12397;
  assign n12399 = n2740 & ~n12398;
  assign n12400 = ~n3042 & n12399;
  assign n12401 = ~n12395 & ~n12400;
  assign po0286 = n12386 | ~n12401;
  assign n12403 = ~n4238 & n12180;
  assign n12404 = ~pi0051 & ~n4208;
  assign n12405 = ~n12147 & n12404;
  assign n12406 = pi0130 & ~n12154;
  assign n12407 = ~n12155 & ~n12406;
  assign n12408 = ~n12158 & ~n12407;
  assign n12409 = n12147 & n12408;
  assign n12410 = ~pi0051 & n12409;
  assign n12411 = ~n12405 & ~n12410;
  assign n12412 = ~pi0087 & n12411;
  assign n12413 = pi0087 & n4258;
  assign n12414 = ~n12412 & ~n12413;
  assign n12415 = ~n11734 & ~n12180;
  assign n12416 = n12175 & n12415;
  assign n12417 = n12140 & n12416;
  assign n12418 = n12414 & n12417;
  assign po0287 = n12403 | n12418;
  assign n12420 = ~n4167 & n12180;
  assign n12421 = n12140 & n12312;
  assign n12422 = ~n3491 & n11734;
  assign n12423 = ~n4204 & n12144;
  assign n12424 = ~n12422 & ~n12423;
  assign n12425 = pi0051 & ~n12071;
  assign n12426 = ~n3271 & ~n12147;
  assign n12427 = ~n3481 & ~n12147;
  assign n12428 = ~n12426 & ~n12427;
  assign n12429 = ~pi0051 & ~n12428;
  assign n12430 = pi0132 & n12158;
  assign n12431 = ~pi0121 & ~pi0126;
  assign n12432 = n12149 & n12431;
  assign n12433 = pi0132 & ~n12432;
  assign n12434 = ~pi0132 & n12432;
  assign n12435 = ~n12433 & ~n12434;
  assign n12436 = ~n12158 & ~n12435;
  assign n12437 = ~n12430 & ~n12436;
  assign n12438 = ~pi0051 & n12147;
  assign n12439 = ~n12437 & n12438;
  assign n12440 = ~n12429 & ~n12439;
  assign n12441 = ~n12425 & n12440;
  assign n12442 = ~pi0087 & ~n11734;
  assign n12443 = ~n12441 & n12442;
  assign n12444 = n12424 & ~n12443;
  assign n12445 = n12421 & ~n12444;
  assign po0289 = n12420 | n12445;
  assign n12447 = ~n11734 & n12140;
  assign n12448 = pi0133 & ~n12158;
  assign n12449 = ~pi0133 & n12158;
  assign n12450 = ~n12448 & ~n12449;
  assign n12451 = n12438 & ~n12450;
  assign n12452 = ~pi0087 & ~n12451;
  assign n12453 = pi0087 & ~n4167;
  assign n12454 = ~n12452 & ~n12453;
  assign n12455 = n12447 & ~n12454;
  assign n12456 = ~n3148 & ~n12140;
  assign n12457 = ~n12455 & ~n12456;
  assign n12458 = ~n12176 & n12457;
  assign n12459 = n12312 & ~n12458;
  assign n12460 = ~n3482 & n12180;
  assign po0290 = n12459 | n12460;
  assign n12462 = ~pi0130 & ~pi0132;
  assign n12463 = ~pi0135 & ~pi0136;
  assign n12464 = n12432 & n12463;
  assign n12465 = n12462 & n12464;
  assign n12466 = pi0134 & ~n12465;
  assign n12467 = ~pi0134 & n12465;
  assign n12468 = ~n12466 & ~n12467;
  assign n12469 = ~n12158 & ~n12468;
  assign n12470 = pi0134 & n12158;
  assign n12471 = ~n12469 & ~n12470;
  assign n12472 = n12147 & ~n12471;
  assign n12473 = ~n3203 & ~n12147;
  assign n12474 = ~n12472 & ~n12473;
  assign n12475 = ~n12427 & n12474;
  assign n12476 = n12140 & ~n12475;
  assign n12477 = ~n11734 & n12162;
  assign n12478 = n12476 & n12477;
  assign n12479 = n12312 & n12478;
  assign n12480 = ~n4204 & n12180;
  assign po0291 = n12479 | n12480;
  assign n12482 = ~pi0130 & n12150;
  assign n12483 = ~pi0136 & n12153;
  assign n12484 = n12482 & n12483;
  assign n12485 = pi0135 & ~n12484;
  assign n12486 = ~pi0135 & n12484;
  assign n12487 = ~n12485 & ~n12486;
  assign n12488 = ~n12158 & ~n12487;
  assign n12489 = pi0135 & n12158;
  assign n12490 = ~n12488 & ~n12489;
  assign n12491 = n12147 & ~n12490;
  assign n12492 = ~n3220 & ~n12147;
  assign n12493 = ~n12491 & ~n12492;
  assign n12494 = ~n12427 & n12493;
  assign n12495 = n12140 & ~n12494;
  assign n12496 = n12477 & n12495;
  assign n12497 = n12312 & n12496;
  assign n12498 = ~n12076 & n12180;
  assign po0292 = n12497 | n12498;
  assign n12500 = ~n8748 & n12180;
  assign n12501 = pi0136 & n12158;
  assign n12502 = n12431 & n12462;
  assign n12503 = n12149 & n12502;
  assign n12504 = pi0136 & ~n12503;
  assign n12505 = ~pi0136 & n12503;
  assign n12506 = ~n12504 & ~n12505;
  assign n12507 = ~n12158 & ~n12506;
  assign n12508 = ~n12501 & ~n12507;
  assign n12509 = n12147 & ~n12508;
  assign n12510 = ~n4262 & ~n12147;
  assign n12511 = ~n12509 & ~n12510;
  assign n12512 = ~n12180 & ~n12511;
  assign n12513 = n12140 & n12512;
  assign n12514 = n12175 & n12513;
  assign n12515 = n12477 & n12514;
  assign po0293 = n12500 | n12515;
  assign n12517 = n3018 & n5010;
  assign n12518 = ~pi0039 & pi0137;
  assign po0294 = n12517 | n12518;
  assign n12520 = n4152 & n4155;
  assign n12521 = ~n4162 & ~n4262;
  assign n12522 = pi0138 & ~n4190;
  assign n12523 = ~n4191 & ~n12522;
  assign n12524 = n4194 & ~n12523;
  assign n12525 = pi0138 & ~n4194;
  assign n12526 = ~n12524 & ~n12525;
  assign n12527 = n4163 & n4198;
  assign n12528 = n8753 & n12527;
  assign n12529 = n4162 & n12528;
  assign n12530 = n4186 & n12529;
  assign n12531 = ~n12526 & n12530;
  assign n12532 = ~n12521 & ~n12531;
  assign po0295 = n12520 & ~n12532;
  assign n12534 = ~n4162 & ~n4208;
  assign n12535 = n4187 & n4247;
  assign n12536 = pi0139 & ~n12535;
  assign n12537 = ~pi0139 & n12535;
  assign n12538 = ~n12536 & ~n12537;
  assign n12539 = n4194 & ~n12538;
  assign n12540 = pi0139 & ~n4194;
  assign n12541 = ~n12539 & ~n12540;
  assign n12542 = n12530 & ~n12541;
  assign n12543 = ~n12534 & ~n12542;
  assign po0296 = n12520 & ~n12543;
  assign n12545 = ~n2788 & ~n2841;
  assign n12546 = pi0252 & n4009;
  assign n12547 = n2614 & n12546;
  assign n12548 = n12545 & ~n12547;
  assign n12549 = ~pi0841 & ~po0740;
  assign n12550 = n2831 & n12549;
  assign n12551 = ~n2626 & ~n12550;
  assign n12552 = pi0252 & ~n12551;
  assign n12553 = ~pi0120 & po0740;
  assign n12554 = pi0120 & n3128;
  assign n12555 = n4097 & ~n12554;
  assign n12556 = ~n12553 & ~n12555;
  assign n12557 = n3397 & n12556;
  assign n12558 = pi0120 & ~n3397;
  assign n12559 = ~n12557 & ~n12558;
  assign n12560 = ~pi0979 & n3466;
  assign n12561 = n12559 & n12560;
  assign n12562 = n3547 & ~n12561;
  assign n12563 = n2685 & n4003;
  assign n12564 = n3053 & n12563;
  assign n12565 = ~po0950 & n12564;
  assign n12566 = pi0120 & pi0287;
  assign n12567 = n2777 & n12566;
  assign n12568 = ~n2679 & ~n12567;
  assign n12569 = ~n2926 & n12568;
  assign n12570 = ~n12565 & n12569;
  assign n12571 = ~n8145 & n12570;
  assign n12572 = ~n12562 & n12571;
  assign n12573 = ~n12552 & n12572;
  assign po0387 = ~n12548 | ~n12573;
  assign n12575 = n2721 & po0387;
  assign n12576 = pi0832 & n2721;
  assign n12577 = ~n12575 & ~n12576;
  assign n12578 = pi0788 & pi1152;
  assign n12579 = pi0626 & pi0788;
  assign n12580 = n12578 & n12579;
  assign n12581 = ~pi0788 & ~n12578;
  assign n12582 = ~pi0626 & ~n12578;
  assign n12583 = ~n12581 & ~n12582;
  assign n12584 = ~n12580 & n12583;
  assign n12585 = pi0789 & pi1153;
  assign n12586 = pi0619 & n12585;
  assign n12587 = pi0789 & n12586;
  assign n12588 = ~pi0619 & ~n12585;
  assign n12589 = ~n12587 & ~n12588;
  assign n12590 = ~pi0789 & ~n12585;
  assign n12591 = n12589 & ~n12590;
  assign n12592 = ~n12584 & ~n12591;
  assign n12593 = pi0630 & pi0787;
  assign n12594 = pi0787 & pi1151;
  assign n12595 = ~n12593 & n12594;
  assign n12596 = pi0630 & ~n12594;
  assign n12597 = ~n12595 & ~n12596;
  assign n12598 = ~pi0787 & ~n12594;
  assign n12599 = ~n12597 & ~n12598;
  assign n12600 = n12592 & ~n12599;
  assign n12601 = pi0790 & pi1154;
  assign n12602 = pi0644 & pi0790;
  assign n12603 = n12601 & n12602;
  assign n12604 = ~pi0790 & ~n12601;
  assign n12605 = ~pi0644 & ~n12601;
  assign n12606 = ~n12604 & ~n12605;
  assign n12607 = ~n12603 & n12606;
  assign n12608 = pi0603 & ~n12607;
  assign n12609 = pi0629 & pi0792;
  assign n12610 = pi0792 & pi1150;
  assign n12611 = ~n12609 & n12610;
  assign n12612 = pi0629 & ~n12610;
  assign n12613 = ~n12611 & ~n12612;
  assign n12614 = ~pi0792 & ~n12610;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = n12608 & ~n12615;
  assign n12617 = pi0778 & pi1147;
  assign n12618 = pi0778 & n12617;
  assign n12619 = pi0608 & n12618;
  assign n12620 = ~pi0608 & ~n12617;
  assign n12621 = ~n12619 & ~n12620;
  assign n12622 = ~pi0778 & ~n12617;
  assign n12623 = n12621 & ~n12622;
  assign n12624 = pi0609 & pi0785;
  assign n12625 = pi0785 & pi1149;
  assign n12626 = ~n12624 & n12625;
  assign n12627 = pi0609 & ~n12625;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = ~pi0785 & ~n12625;
  assign n12630 = ~n12628 & ~n12629;
  assign n12631 = ~n12623 & ~n12630;
  assign n12632 = pi0781 & pi1148;
  assign n12633 = pi0618 & n12632;
  assign n12634 = pi0781 & n12633;
  assign n12635 = ~pi0781 & ~n12632;
  assign n12636 = ~pi0618 & ~n12632;
  assign n12637 = ~n12635 & ~n12636;
  assign n12638 = ~n12634 & n12637;
  assign n12639 = n12631 & ~n12638;
  assign n12640 = n12616 & n12639;
  assign n12641 = n12600 & n12640;
  assign n12642 = pi0621 & pi1085;
  assign n12643 = n12641 & ~n12642;
  assign n12644 = ~pi0761 & n12643;
  assign n12645 = ~n12577 & n12644;
  assign n12646 = ~pi0738 & ~n12577;
  assign n12647 = pi0647 & n12594;
  assign n12648 = pi0787 & n12647;
  assign n12649 = ~pi0647 & ~n12594;
  assign n12650 = ~n12598 & ~n12649;
  assign n12651 = ~n12648 & n12650;
  assign n12652 = pi0648 & n12585;
  assign n12653 = pi0789 & n12652;
  assign n12654 = ~pi0648 & ~n12585;
  assign n12655 = ~n12653 & ~n12654;
  assign n12656 = ~n12590 & n12655;
  assign n12657 = ~n12651 & ~n12656;
  assign n12658 = pi0641 & pi0788;
  assign n12659 = n12578 & ~n12658;
  assign n12660 = pi0641 & ~n12578;
  assign n12661 = ~n12659 & ~n12660;
  assign n12662 = ~n12581 & ~n12661;
  assign n12663 = n12657 & ~n12662;
  assign n12664 = pi0625 & n12618;
  assign n12665 = ~pi0625 & ~n12617;
  assign n12666 = ~n12664 & ~n12665;
  assign n12667 = ~n12622 & n12666;
  assign n12668 = pi0680 & ~n12667;
  assign n12669 = pi0715 & pi0790;
  assign n12670 = n12601 & ~n12669;
  assign n12671 = pi0715 & ~n12601;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = ~n12604 & ~n12672;
  assign n12674 = n12668 & ~n12673;
  assign n12675 = pi0628 & pi0792;
  assign n12676 = n12610 & ~n12675;
  assign n12677 = pi0628 & ~n12610;
  assign n12678 = ~n12676 & ~n12677;
  assign n12679 = ~n12614 & ~n12678;
  assign n12680 = pi0627 & pi0781;
  assign n12681 = n12632 & ~n12680;
  assign n12682 = pi0627 & ~n12632;
  assign n12683 = ~n12681 & ~n12682;
  assign n12684 = ~n12635 & ~n12683;
  assign n12685 = ~n12679 & ~n12684;
  assign n12686 = pi0660 & n12625;
  assign n12687 = pi0785 & n12686;
  assign n12688 = ~pi0660 & ~n12625;
  assign n12689 = ~n12629 & ~n12688;
  assign n12690 = ~n12687 & n12689;
  assign n12691 = n12685 & ~n12690;
  assign n12692 = n12674 & n12691;
  assign n12693 = n12663 & n12692;
  assign n12694 = pi0665 & pi1085;
  assign n12695 = n12693 & ~n12694;
  assign n12696 = ~n12643 & n12695;
  assign n12697 = n12646 & n12696;
  assign n12698 = ~n12645 & ~n12697;
  assign n12699 = ~pi0140 & n12577;
  assign po0297 = ~n12698 | n12699;
  assign n12701 = pi0749 & n12643;
  assign n12702 = ~n12577 & n12701;
  assign n12703 = pi0706 & ~n12577;
  assign n12704 = n12696 & n12703;
  assign n12705 = ~n12702 & ~n12704;
  assign n12706 = ~pi0141 & n12577;
  assign po0298 = ~n12705 | n12706;
  assign n12708 = pi0743 & n12643;
  assign n12709 = ~n12577 & n12708;
  assign n12710 = pi0735 & ~n12577;
  assign n12711 = n12696 & n12710;
  assign n12712 = ~n12709 & ~n12711;
  assign n12713 = pi0142 & n12577;
  assign po0299 = ~n12712 | n12713;
  assign n12715 = ~pi0774 & n12643;
  assign n12716 = ~n12577 & n12715;
  assign n12717 = pi0687 & ~n12577;
  assign n12718 = n12696 & n12717;
  assign n12719 = ~n12716 & ~n12718;
  assign n12720 = ~pi0143 & n12577;
  assign po0300 = ~n12719 | n12720;
  assign n12722 = pi0758 & n12643;
  assign n12723 = ~n12577 & n12722;
  assign n12724 = pi0736 & ~n12577;
  assign n12725 = n12696 & n12724;
  assign n12726 = ~n12723 & ~n12725;
  assign n12727 = pi0144 & n12577;
  assign po0301 = ~n12726 | n12727;
  assign n12729 = ~pi0767 & n12643;
  assign n12730 = ~n12577 & n12729;
  assign n12731 = ~pi0698 & ~n12577;
  assign n12732 = n12696 & n12731;
  assign n12733 = ~n12730 & ~n12732;
  assign n12734 = ~pi0145 & n12577;
  assign po0302 = ~n12733 | n12734;
  assign n12736 = pi0743 & pi0947;
  assign n12737 = ~n12577 & n12736;
  assign n12738 = pi0907 & ~pi0947;
  assign n12739 = n12710 & n12738;
  assign n12740 = ~n12737 & ~n12739;
  assign n12741 = pi0146 & n12577;
  assign po0303 = ~n12740 | n12741;
  assign n12743 = ~pi0770 & pi0947;
  assign n12744 = ~n12577 & n12743;
  assign n12745 = pi0726 & ~n12577;
  assign n12746 = n12738 & n12745;
  assign n12747 = ~n12744 & ~n12746;
  assign n12748 = ~pi0147 & n12577;
  assign po0304 = ~n12747 | n12748;
  assign n12750 = pi0749 & pi0947;
  assign n12751 = ~n12577 & n12750;
  assign n12752 = n12703 & n12738;
  assign n12753 = ~n12751 & ~n12752;
  assign n12754 = ~pi0148 & n12577;
  assign po0305 = ~n12753 | n12754;
  assign n12756 = ~pi0755 & pi0947;
  assign n12757 = ~n12577 & n12756;
  assign n12758 = ~pi0725 & ~n12577;
  assign n12759 = n12738 & n12758;
  assign n12760 = ~n12757 & ~n12759;
  assign n12761 = ~pi0149 & n12577;
  assign po0306 = ~n12760 | n12761;
  assign n12763 = ~pi0751 & pi0947;
  assign n12764 = ~n12577 & n12763;
  assign n12765 = ~pi0701 & ~n12577;
  assign n12766 = n12738 & n12765;
  assign n12767 = ~n12764 & ~n12766;
  assign n12768 = ~pi0150 & n12577;
  assign po0307 = ~n12767 | n12768;
  assign n12770 = ~pi0745 & pi0947;
  assign n12771 = ~n12577 & n12770;
  assign n12772 = ~pi0723 & ~n12577;
  assign n12773 = n12738 & n12772;
  assign n12774 = ~n12771 & ~n12773;
  assign n12775 = ~pi0151 & n12577;
  assign po0308 = ~n12774 | n12775;
  assign n12777 = pi0759 & pi0947;
  assign n12778 = ~n12577 & n12777;
  assign n12779 = pi0696 & ~n12577;
  assign n12780 = n12738 & n12779;
  assign n12781 = ~n12778 & ~n12780;
  assign n12782 = pi0152 & n12577;
  assign po0309 = ~n12781 | n12782;
  assign n12784 = pi0766 & pi0947;
  assign n12785 = ~n12577 & n12784;
  assign n12786 = pi0700 & ~n12577;
  assign n12787 = n12738 & n12786;
  assign n12788 = ~n12785 & ~n12787;
  assign n12789 = ~pi0153 & n12577;
  assign po0310 = ~n12788 | n12789;
  assign n12791 = ~pi0742 & pi0947;
  assign n12792 = ~n12577 & n12791;
  assign n12793 = ~pi0704 & ~n12577;
  assign n12794 = n12738 & n12793;
  assign n12795 = ~n12792 & ~n12794;
  assign n12796 = ~pi0154 & n12577;
  assign po0311 = ~n12795 | n12796;
  assign n12798 = ~pi0757 & pi0947;
  assign n12799 = ~n12577 & n12798;
  assign n12800 = ~pi0686 & ~n12577;
  assign n12801 = n12738 & n12800;
  assign n12802 = ~n12799 & ~n12801;
  assign n12803 = ~pi0155 & n12577;
  assign po0312 = ~n12802 | n12803;
  assign n12805 = ~pi0741 & pi0947;
  assign n12806 = ~n12577 & n12805;
  assign n12807 = ~pi0724 & ~n12577;
  assign n12808 = n12738 & n12807;
  assign n12809 = ~n12806 & ~n12808;
  assign n12810 = ~pi0156 & n12577;
  assign po0313 = ~n12809 | n12810;
  assign n12812 = ~pi0760 & pi0947;
  assign n12813 = ~n12577 & n12812;
  assign n12814 = ~pi0688 & ~n12577;
  assign n12815 = n12738 & n12814;
  assign n12816 = ~n12813 & ~n12815;
  assign n12817 = ~pi0157 & n12577;
  assign po0314 = ~n12816 | n12817;
  assign n12819 = ~pi0753 & pi0947;
  assign n12820 = ~n12577 & n12819;
  assign n12821 = ~pi0702 & ~n12577;
  assign n12822 = n12738 & n12821;
  assign n12823 = ~n12820 & ~n12822;
  assign n12824 = ~pi0158 & n12577;
  assign po0315 = ~n12823 | n12824;
  assign n12826 = ~pi0754 & pi0947;
  assign n12827 = ~n12577 & n12826;
  assign n12828 = ~pi0709 & ~n12577;
  assign n12829 = n12738 & n12828;
  assign n12830 = ~n12827 & ~n12829;
  assign n12831 = ~pi0159 & n12577;
  assign po0316 = ~n12830 | n12831;
  assign n12833 = ~pi0756 & pi0947;
  assign n12834 = ~n12577 & n12833;
  assign n12835 = ~pi0734 & ~n12577;
  assign n12836 = n12738 & n12835;
  assign n12837 = ~n12834 & ~n12836;
  assign n12838 = ~pi0160 & n12577;
  assign po0317 = ~n12837 | n12838;
  assign n12840 = pi0758 & pi0947;
  assign n12841 = ~n12577 & n12840;
  assign n12842 = n12724 & n12738;
  assign n12843 = ~n12841 & ~n12842;
  assign n12844 = pi0161 & n12577;
  assign po0318 = ~n12843 | n12844;
  assign n12846 = ~pi0761 & pi0947;
  assign n12847 = ~n12577 & n12846;
  assign n12848 = n12646 & n12738;
  assign n12849 = ~n12847 & ~n12848;
  assign n12850 = ~pi0162 & n12577;
  assign po0319 = ~n12849 | n12850;
  assign n12852 = ~pi0777 & pi0947;
  assign n12853 = ~n12577 & n12852;
  assign n12854 = ~pi0737 & ~n12577;
  assign n12855 = n12738 & n12854;
  assign n12856 = ~n12853 & ~n12855;
  assign n12857 = ~pi0163 & n12577;
  assign po0320 = ~n12856 | n12857;
  assign n12859 = ~pi0752 & pi0947;
  assign n12860 = ~n12577 & n12859;
  assign n12861 = pi0703 & ~n12577;
  assign n12862 = n12738 & n12861;
  assign n12863 = ~n12860 & ~n12862;
  assign n12864 = ~pi0164 & n12577;
  assign po0321 = ~n12863 | n12864;
  assign n12866 = ~pi0774 & pi0947;
  assign n12867 = ~n12577 & n12866;
  assign n12868 = n12717 & n12738;
  assign n12869 = ~n12867 & ~n12868;
  assign n12870 = ~pi0165 & n12577;
  assign po0322 = ~n12869 | n12870;
  assign n12872 = pi0772 & pi0947;
  assign n12873 = ~n12577 & n12872;
  assign n12874 = pi0727 & ~n12577;
  assign n12875 = n12738 & n12874;
  assign n12876 = ~n12873 & ~n12875;
  assign n12877 = pi0166 & n12577;
  assign po0323 = ~n12876 | n12877;
  assign n12879 = ~pi0768 & pi0947;
  assign n12880 = ~n12577 & n12879;
  assign n12881 = pi0705 & ~n12577;
  assign n12882 = n12738 & n12881;
  assign n12883 = ~n12880 & ~n12882;
  assign n12884 = ~pi0167 & n12577;
  assign po0324 = ~n12883 | n12884;
  assign n12886 = pi0763 & pi0947;
  assign n12887 = ~n12577 & n12886;
  assign n12888 = pi0699 & ~n12577;
  assign n12889 = n12738 & n12888;
  assign n12890 = ~n12887 & ~n12889;
  assign n12891 = ~pi0168 & n12577;
  assign po0325 = ~n12890 | n12891;
  assign n12893 = pi0746 & pi0947;
  assign n12894 = ~n12577 & n12893;
  assign n12895 = pi0729 & ~n12577;
  assign n12896 = n12738 & n12895;
  assign n12897 = ~n12894 & ~n12896;
  assign n12898 = ~pi0169 & n12577;
  assign po0326 = ~n12897 | n12898;
  assign n12900 = pi0748 & pi0947;
  assign n12901 = ~n12577 & n12900;
  assign n12902 = pi0730 & ~n12577;
  assign n12903 = n12738 & n12902;
  assign n12904 = ~n12901 & ~n12903;
  assign n12905 = ~pi0170 & n12577;
  assign po0327 = ~n12904 | n12905;
  assign n12907 = pi0764 & pi0947;
  assign n12908 = ~n12577 & n12907;
  assign n12909 = pi0691 & ~n12577;
  assign n12910 = n12738 & n12909;
  assign n12911 = ~n12908 & ~n12910;
  assign n12912 = ~pi0171 & n12577;
  assign po0328 = ~n12911 | n12912;
  assign n12914 = pi0739 & pi0947;
  assign n12915 = ~n12577 & n12914;
  assign n12916 = pi0690 & ~n12577;
  assign n12917 = n12738 & n12916;
  assign n12918 = ~n12915 & ~n12917;
  assign n12919 = ~pi0172 & n12577;
  assign po0329 = ~n12918 | n12919;
  assign n12921 = ~pi0745 & n12643;
  assign n12922 = ~n12577 & n12921;
  assign n12923 = n12696 & n12772;
  assign n12924 = ~n12922 & ~n12923;
  assign n12925 = ~pi0173 & n12577;
  assign po0330 = ~n12924 | n12925;
  assign n12927 = pi0759 & n12643;
  assign n12928 = ~n12577 & n12927;
  assign n12929 = n12696 & n12779;
  assign n12930 = ~n12928 & ~n12929;
  assign n12931 = pi0174 & n12577;
  assign po0331 = ~n12930 | n12931;
  assign n12933 = pi0766 & n12643;
  assign n12934 = ~n12577 & n12933;
  assign n12935 = n12696 & n12786;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = ~pi0175 & n12577;
  assign po0332 = ~n12936 | n12937;
  assign n12939 = ~pi0742 & n12643;
  assign n12940 = ~n12577 & n12939;
  assign n12941 = n12696 & n12793;
  assign n12942 = ~n12940 & ~n12941;
  assign n12943 = ~pi0176 & n12577;
  assign po0333 = ~n12942 | n12943;
  assign n12945 = ~pi0757 & n12643;
  assign n12946 = ~n12577 & n12945;
  assign n12947 = n12696 & n12800;
  assign n12948 = ~n12946 & ~n12947;
  assign n12949 = ~pi0177 & n12577;
  assign po0334 = ~n12948 | n12949;
  assign n12951 = ~pi0760 & n12643;
  assign n12952 = ~n12577 & n12951;
  assign n12953 = n12696 & n12814;
  assign n12954 = ~n12952 & ~n12953;
  assign n12955 = ~pi0178 & n12577;
  assign po0335 = ~n12954 | n12955;
  assign n12957 = ~pi0741 & n12643;
  assign n12958 = ~n12577 & n12957;
  assign n12959 = n12696 & n12807;
  assign n12960 = ~n12958 & ~n12959;
  assign n12961 = ~pi0179 & n12577;
  assign po0336 = ~n12960 | n12961;
  assign n12963 = ~pi0753 & n12643;
  assign n12964 = ~n12577 & n12963;
  assign n12965 = n12696 & n12821;
  assign n12966 = ~n12964 & ~n12965;
  assign n12967 = ~pi0180 & n12577;
  assign po0337 = ~n12966 | n12967;
  assign n12969 = ~pi0754 & n12643;
  assign n12970 = ~n12577 & n12969;
  assign n12971 = n12696 & n12828;
  assign n12972 = ~n12970 & ~n12971;
  assign n12973 = ~pi0181 & n12577;
  assign po0338 = ~n12972 | n12973;
  assign n12975 = ~pi0756 & n12643;
  assign n12976 = ~n12577 & n12975;
  assign n12977 = n12696 & n12835;
  assign n12978 = ~n12976 & ~n12977;
  assign n12979 = ~pi0182 & n12577;
  assign po0339 = ~n12978 | n12979;
  assign n12981 = ~pi0755 & n12643;
  assign n12982 = ~n12577 & n12981;
  assign n12983 = n12696 & n12758;
  assign n12984 = ~n12982 & ~n12983;
  assign n12985 = ~pi0183 & n12577;
  assign po0340 = ~n12984 | n12985;
  assign n12987 = ~pi0777 & n12643;
  assign n12988 = ~n12577 & n12987;
  assign n12989 = n12696 & n12854;
  assign n12990 = ~n12988 & ~n12989;
  assign n12991 = ~pi0184 & n12577;
  assign po0341 = ~n12990 | n12991;
  assign n12993 = ~pi0751 & n12643;
  assign n12994 = ~n12577 & n12993;
  assign n12995 = n12696 & n12765;
  assign n12996 = ~n12994 & ~n12995;
  assign n12997 = ~pi0185 & n12577;
  assign po0342 = ~n12996 | n12997;
  assign n12999 = ~pi0752 & n12643;
  assign n13000 = ~n12577 & n12999;
  assign n13001 = n12696 & n12861;
  assign n13002 = ~n13000 & ~n13001;
  assign n13003 = ~pi0186 & n12577;
  assign po0343 = ~n13002 | n13003;
  assign n13005 = ~pi0770 & n12643;
  assign n13006 = ~n12577 & n13005;
  assign n13007 = n12696 & n12745;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~pi0187 & n12577;
  assign po0344 = ~n13008 | n13009;
  assign n13011 = ~pi0768 & n12643;
  assign n13012 = ~n12577 & n13011;
  assign n13013 = n12696 & n12881;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = ~pi0188 & n12577;
  assign po0345 = ~n13014 | n13015;
  assign n13017 = pi0772 & n12643;
  assign n13018 = ~n12577 & n13017;
  assign n13019 = n12696 & n12874;
  assign n13020 = ~n13018 & ~n13019;
  assign n13021 = pi0189 & n12577;
  assign po0346 = ~n13020 | n13021;
  assign n13023 = pi0763 & n12643;
  assign n13024 = ~n12577 & n13023;
  assign n13025 = n12696 & n12888;
  assign n13026 = ~n13024 & ~n13025;
  assign n13027 = ~pi0190 & n12577;
  assign po0347 = ~n13026 | n13027;
  assign n13029 = pi0746 & n12643;
  assign n13030 = ~n12577 & n13029;
  assign n13031 = n12696 & n12895;
  assign n13032 = ~n13030 & ~n13031;
  assign n13033 = ~pi0191 & n12577;
  assign po0348 = ~n13032 | n13033;
  assign n13035 = pi0764 & n12643;
  assign n13036 = ~n12577 & n13035;
  assign n13037 = n12696 & n12909;
  assign n13038 = ~n13036 & ~n13037;
  assign n13039 = ~pi0192 & n12577;
  assign po0349 = ~n13038 | n13039;
  assign n13041 = pi0739 & n12643;
  assign n13042 = ~n12577 & n13041;
  assign n13043 = n12696 & n12916;
  assign n13044 = ~n13042 & ~n13043;
  assign n13045 = ~pi0193 & n12577;
  assign po0350 = ~n13044 | n13045;
  assign n13047 = pi0748 & n12643;
  assign n13048 = ~n12577 & n13047;
  assign n13049 = n12696 & n12902;
  assign n13050 = ~n13048 & ~n13049;
  assign n13051 = ~pi0194 & n12577;
  assign po0351 = ~n13050 | n13051;
  assign n13053 = ~pi0138 & ~pi0196;
  assign n13054 = ~pi0139 & n8760;
  assign n13055 = ~pi0118 & n13054;
  assign n13056 = n13053 & n13055;
  assign n13057 = pi0195 & n13056;
  assign n13058 = ~pi0195 & ~n13056;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = n4194 & n13059;
  assign n13061 = pi0195 & ~n4194;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = n4186 & ~n13062;
  assign n13064 = n4162 & n13063;
  assign n13065 = n4198 & n13064;
  assign n13066 = n8752 & n13065;
  assign n13067 = n4163 & n4182;
  assign n13068 = n13066 & n13067;
  assign n13069 = ~n3203 & ~n4162;
  assign n13070 = ~n13068 & ~n13069;
  assign n13071 = ~n12103 & n13070;
  assign po0352 = n12520 & ~n13071;
  assign n13073 = ~pi0139 & n4247;
  assign n13074 = ~pi0138 & n13073;
  assign n13075 = n4187 & n13074;
  assign n13076 = pi0196 & n13075;
  assign n13077 = ~pi0196 & ~n13075;
  assign n13078 = ~n13076 & ~n13077;
  assign n13079 = n4194 & n13078;
  assign n13080 = pi0196 & ~n4194;
  assign n13081 = ~n13079 & ~n13080;
  assign n13082 = n4186 & ~n13081;
  assign n13083 = n4162 & n13082;
  assign n13084 = n12528 & n13083;
  assign n13085 = ~n3220 & ~n4162;
  assign n13086 = ~n13084 & ~n13085;
  assign n13087 = ~n12103 & n13086;
  assign po0353 = n12520 & ~n13087;
  assign n13089 = ~pi0767 & pi0947;
  assign n13090 = ~n12577 & n13089;
  assign n13091 = n12731 & n12738;
  assign n13092 = ~n13090 & ~n13091;
  assign n13093 = ~pi0197 & n12577;
  assign po0354 = ~n13092 | n13093;
  assign n13095 = n12575 & n12643;
  assign n13096 = pi0633 & n13095;
  assign n13097 = pi0198 & ~n12575;
  assign n13098 = pi0634 & n12575;
  assign n13099 = n12696 & n13098;
  assign n13100 = ~n13097 & ~n13099;
  assign po0355 = n13096 | ~n13100;
  assign n13102 = pi0617 & n13095;
  assign n13103 = pi0199 & ~n12575;
  assign n13104 = pi0637 & n12575;
  assign n13105 = n12696 & n13104;
  assign n13106 = ~n13103 & ~n13105;
  assign po0356 = n13102 | ~n13106;
  assign n13108 = pi0606 & n13095;
  assign n13109 = pi0200 & ~n12575;
  assign n13110 = pi0643 & n12575;
  assign n13111 = n12696 & n13110;
  assign n13112 = ~n13109 & ~n13111;
  assign po0357 = n13108 | ~n13112;
  assign n13114 = pi0233 & pi0237;
  assign n13115 = n3375 & n10571;
  assign n13116 = n13114 & n13115;
  assign n13117 = ~pi0032 & pi0070;
  assign n13118 = ~pi0332 & n13117;
  assign n13119 = pi0032 & ~pi0070;
  assign n13120 = n3461 & n13119;
  assign n13121 = ~n13118 & ~n13120;
  assign n13122 = n3375 & ~n13121;
  assign n13123 = n13114 & n13122;
  assign n13124 = ~pi0201 & ~pi0332;
  assign n13125 = ~n13123 & n13124;
  assign n13126 = ~pi0053 & ~pi0106;
  assign n13127 = ~pi0103 & n2994;
  assign n13128 = n2992 & n13127;
  assign n13129 = ~pi0087 & n13128;
  assign n13130 = n2451 & n2454;
  assign n13131 = ~pi0063 & n13130;
  assign n13132 = n2481 & n2974;
  assign n13133 = n2971 & n2993;
  assign n13134 = ~pi0107 & n13133;
  assign n13135 = n2978 & n13134;
  assign n13136 = n13132 & n13135;
  assign n13137 = n13131 & n13136;
  assign n13138 = n13129 & n13137;
  assign n13139 = n2958 & n2998;
  assign n13140 = ~pi0088 & n13139;
  assign n13141 = n2502 & n13140;
  assign n13142 = ~pi0092 & n13141;
  assign n13143 = ~pi0047 & n13142;
  assign n13144 = n2501 & n13143;
  assign n13145 = ~pi0058 & n13144;
  assign n13146 = n2972 & n13145;
  assign n13147 = n13138 & n13146;
  assign n13148 = ~pi0060 & n13147;
  assign n13149 = n2980 & n13148;
  assign n13150 = n12260 & n13149;
  assign n13151 = ~pi0045 & pi0055;
  assign n13152 = n13150 & n13151;
  assign n13153 = n2906 & n13147;
  assign n13154 = pi0059 & n13148;
  assign n13155 = ~n13153 & ~n13154;
  assign n13156 = n2448 & ~n13155;
  assign n13157 = ~pi0045 & n13156;
  assign n13158 = n2425 & n13157;
  assign n13159 = ~n13152 & ~n13158;
  assign n13160 = ~pi0054 & ~n13159;
  assign n13161 = n12275 & n13150;
  assign n13162 = pi0054 & n13161;
  assign n13163 = ~n13160 & ~n13162;
  assign n13164 = n13126 & ~n13163;
  assign n13165 = pi0053 & n2446;
  assign n13166 = n13161 & n13165;
  assign n13167 = ~n13164 & ~n13166;
  assign n13168 = ~pi0070 & n2962;
  assign n13169 = ~pi0096 & n13168;
  assign n13170 = ~n13167 & n13169;
  assign n13171 = n2467 & n2956;
  assign n13172 = n13170 & n13171;
  assign n13173 = n2466 & n13172;
  assign n13174 = ~pi0108 & n2475;
  assign n13175 = ~pi0035 & n13174;
  assign n13176 = n13173 & n13175;
  assign n13177 = n2954 & n2955;
  assign n13178 = ~pi0070 & n13177;
  assign n13179 = n13176 & n13178;
  assign n13180 = pi0070 & pi0332;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = n3375 & ~n13181;
  assign n13183 = n13125 & ~n13182;
  assign po0358 = n13116 | n13183;
  assign n13185 = ~pi0233 & pi0237;
  assign n13186 = n13122 & n13185;
  assign n13187 = ~pi0332 & ~n13182;
  assign n13188 = ~n13186 & n13187;
  assign n13189 = ~pi0202 & n13188;
  assign n13190 = n13115 & n13185;
  assign po0359 = n13189 | n13190;
  assign n13192 = ~pi0233 & ~pi0237;
  assign n13193 = n13122 & n13192;
  assign n13194 = n13187 & ~n13193;
  assign n13195 = ~pi0203 & n13194;
  assign n13196 = n13115 & n13192;
  assign po0360 = n13195 | n13196;
  assign n13198 = ~n3384 & n10571;
  assign n13199 = n13114 & n13198;
  assign n13200 = ~n3384 & ~n13121;
  assign n13201 = n13114 & n13200;
  assign n13202 = ~pi0204 & ~pi0332;
  assign n13203 = ~n13201 & n13202;
  assign n13204 = ~n3384 & ~n13181;
  assign n13205 = n13203 & ~n13204;
  assign po0361 = n13199 | n13205;
  assign n13207 = n13185 & n13200;
  assign n13208 = ~pi0332 & ~n13204;
  assign n13209 = ~n13207 & n13208;
  assign n13210 = ~pi0205 & n13209;
  assign n13211 = n13185 & n13198;
  assign po0362 = n13210 | n13211;
  assign n13213 = pi0233 & ~pi0237;
  assign n13214 = n13200 & n13213;
  assign n13215 = n13208 & ~n13214;
  assign n13216 = ~pi0206 & n13215;
  assign n13217 = n13198 & n13213;
  assign po0363 = n13216 | n13217;
  assign n13219 = pi0623 & n12575;
  assign n13220 = n12643 & n13219;
  assign n13221 = pi0710 & n12575;
  assign n13222 = n12696 & n13221;
  assign n13223 = ~n13220 & ~n13222;
  assign n13224 = ~pi0207 & ~n12575;
  assign po0364 = ~n13223 | n13224;
  assign n13226 = pi0607 & n12575;
  assign n13227 = n12643 & n13226;
  assign n13228 = pi0638 & n12575;
  assign n13229 = n12696 & n13228;
  assign n13230 = ~n13227 & ~n13229;
  assign n13231 = ~pi0208 & ~n12575;
  assign po0365 = ~n13230 | n13231;
  assign n13233 = pi0622 & n12575;
  assign n13234 = n12643 & n13233;
  assign n13235 = pi0639 & n12575;
  assign n13236 = n12696 & n13235;
  assign n13237 = ~n13234 & ~n13236;
  assign n13238 = ~pi0209 & ~n12575;
  assign po0366 = ~n13237 | n13238;
  assign n13240 = pi0633 & n12575;
  assign n13241 = pi0947 & n13240;
  assign n13242 = pi0210 & ~n12575;
  assign n13243 = n12738 & n13098;
  assign n13244 = ~n13242 & ~n13243;
  assign po0367 = n13241 | ~n13244;
  assign n13246 = pi0606 & n12575;
  assign n13247 = pi0947 & n13246;
  assign n13248 = pi0211 & ~n12575;
  assign n13249 = n12738 & n13110;
  assign n13250 = ~n13248 & ~n13249;
  assign po0368 = n13247 | ~n13250;
  assign n13252 = pi0607 & pi0947;
  assign n13253 = n12575 & n13252;
  assign n13254 = n12738 & n13228;
  assign n13255 = ~n13253 & ~n13254;
  assign n13256 = ~pi0212 & ~n12575;
  assign po0369 = ~n13255 | n13256;
  assign n13258 = pi0622 & pi0947;
  assign n13259 = n12575 & n13258;
  assign n13260 = n12738 & n13235;
  assign n13261 = ~n13259 & ~n13260;
  assign n13262 = ~pi0213 & ~n12575;
  assign po0370 = ~n13261 | n13262;
  assign n13264 = pi0623 & pi0947;
  assign n13265 = n12575 & n13264;
  assign n13266 = n12738 & n13221;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = ~pi0214 & ~n12575;
  assign po0371 = ~n13267 | n13268;
  assign n13270 = pi0907 & n12575;
  assign n13271 = pi0681 & n13270;
  assign n13272 = ~pi0947 & n13271;
  assign n13273 = pi0215 & ~n12575;
  assign n13274 = pi0947 & n12575;
  assign n13275 = pi0642 & n13274;
  assign n13276 = ~n13273 & ~n13275;
  assign po0372 = n13272 | ~n13276;
  assign n13278 = pi0662 & n13270;
  assign n13279 = ~pi0947 & n13278;
  assign n13280 = pi0216 & ~n12575;
  assign n13281 = pi0614 & n13274;
  assign n13282 = ~n13280 & ~n13281;
  assign po0373 = n13279 | ~n13282;
  assign n13284 = pi0612 & n12643;
  assign n13285 = ~pi0695 & n12696;
  assign n13286 = ~n13284 & ~n13285;
  assign n13287 = n12575 & ~n13286;
  assign n13288 = ~pi0217 & ~n12575;
  assign po0374 = n13287 | n13288;
  assign n13290 = n13192 & n13200;
  assign n13291 = n13208 & ~n13290;
  assign n13292 = ~pi0218 & n13291;
  assign n13293 = n13192 & n13198;
  assign po0375 = n13292 | n13293;
  assign n13295 = pi0617 & n12575;
  assign n13296 = pi0947 & n13295;
  assign n13297 = pi0219 & ~n12575;
  assign n13298 = n12738 & n13104;
  assign n13299 = ~n13297 & ~n13298;
  assign po0376 = n13296 | ~n13299;
  assign n13301 = n13122 & n13213;
  assign n13302 = n13187 & ~n13301;
  assign n13303 = ~pi0220 & n13302;
  assign n13304 = n13115 & n13213;
  assign po0377 = n13303 | n13304;
  assign n13306 = pi0661 & n13270;
  assign n13307 = ~pi0947 & n13306;
  assign n13308 = pi0221 & ~n12575;
  assign n13309 = pi0616 & n13274;
  assign n13310 = ~n13308 & ~n13309;
  assign po0378 = n13307 | ~n13310;
  assign n13312 = pi0222 & ~n12575;
  assign n13313 = pi0616 & n12643;
  assign n13314 = pi0661 & n12696;
  assign n13315 = ~n13313 & ~n13314;
  assign n13316 = n12575 & ~n13315;
  assign po0379 = n13312 | n13316;
  assign n13318 = pi0223 & ~n12575;
  assign n13319 = pi0642 & n12643;
  assign n13320 = pi0681 & n12696;
  assign n13321 = ~n13319 & ~n13320;
  assign n13322 = n12575 & ~n13321;
  assign po0380 = n13318 | n13322;
  assign n13324 = pi0224 & ~n12575;
  assign n13325 = pi0614 & n12643;
  assign n13326 = pi0662 & n12696;
  assign n13327 = ~n13325 & ~n13326;
  assign n13328 = n12575 & ~n13327;
  assign po0381 = n13324 | n13328;
  assign n13330 = pi0228 & pi0231;
  assign n13331 = pi0479 & n2681;
  assign n13332 = n3349 & n12370;
  assign n13333 = n12360 & n13332;
  assign n13334 = ~n13331 & n13333;
  assign n13335 = n2672 & n13334;
  assign n13336 = n2904 & n13335;
  assign po0393 = ~n12391 | ~n13336;
  assign n13338 = ~pi0228 & po0393;
  assign po0383 = n13330 | n13338;
  assign n13340 = ~n2626 & ~n2881;
  assign n13341 = ~n3468 & ~n5312;
  assign n13342 = n2570 & ~n2777;
  assign n13343 = n13341 & n13342;
  assign n13344 = n13340 & n13343;
  assign n13345 = ~n2626 & n13342;
  assign n13346 = n2726 & ~n3468;
  assign n13347 = ~n5312 & n13346;
  assign n13348 = n13345 & n13347;
  assign n13349 = n3402 & n4160;
  assign n13350 = ~pi0287 & n3404;
  assign n13351 = n13349 & n13350;
  assign n13352 = ~n5312 & ~n13351;
  assign n13353 = ~n2569 & ~n2626;
  assign n13354 = ~n2563 & n13353;
  assign n13355 = n13346 & n13354;
  assign n13356 = n13352 & n13355;
  assign n13357 = ~n2626 & ~n13351;
  assign n13358 = ~n2569 & ~n2881;
  assign n13359 = ~n2563 & n13358;
  assign n13360 = n13357 & n13359;
  assign n13361 = n13341 & n13360;
  assign n13362 = ~n2516 & n2570;
  assign n13363 = n13346 & n13357;
  assign n13364 = n13362 & n13363;
  assign n13365 = ~n13351 & n13362;
  assign n13366 = ~n3468 & n13340;
  assign n13367 = n13365 & n13366;
  assign n13368 = ~n13364 & ~n13367;
  assign n13369 = ~n2888 & ~n13351;
  assign n13370 = n13340 & n13369;
  assign n13371 = n13362 & n13370;
  assign n13372 = ~n2626 & ~n2888;
  assign n13373 = n2726 & n13372;
  assign n13374 = n13365 & n13373;
  assign n13375 = ~n13371 & ~n13374;
  assign n13376 = n13368 & n13375;
  assign n13377 = n13352 & n13372;
  assign n13378 = n13359 & n13377;
  assign n13379 = n2726 & ~n5312;
  assign n13380 = n13369 & n13379;
  assign n13381 = n13354 & n13380;
  assign n13382 = ~n13378 & ~n13381;
  assign n13383 = n13376 & n13382;
  assign n13384 = ~n13361 & n13383;
  assign n13385 = ~n13356 & n13384;
  assign n13386 = ~n2563 & ~n2777;
  assign n13387 = ~n2516 & n13386;
  assign n13388 = n13346 & n13353;
  assign n13389 = n13387 & n13388;
  assign n13390 = ~n2626 & n13387;
  assign n13391 = ~n3468 & n13358;
  assign n13392 = n13390 & n13391;
  assign n13393 = ~n13389 & ~n13392;
  assign n13394 = n13385 & n13393;
  assign n13395 = n13342 & n13379;
  assign n13396 = n13372 & n13395;
  assign n13397 = ~n2888 & n13340;
  assign n13398 = ~n5312 & n13342;
  assign n13399 = n13397 & n13398;
  assign n13400 = ~n13396 & ~n13399;
  assign n13401 = n13358 & n13372;
  assign n13402 = n13387 & n13401;
  assign n13403 = n2726 & n13353;
  assign n13404 = ~n2888 & n13387;
  assign n13405 = n13403 & n13404;
  assign n13406 = ~n13402 & ~n13405;
  assign n13407 = n13400 & n13406;
  assign n13408 = n13394 & n13407;
  assign n13409 = ~n13348 & n13408;
  assign po0384 = n13344 | ~n13409;
  assign n13411 = ~n2651 & ~n2858;
  assign n13412 = ~po0840 & ~n3578;
  assign n13413 = ~n2651 & ~n2777;
  assign n13414 = ~n13412 & n13413;
  assign n13415 = ~n13411 & n13414;
  assign n13416 = n13411 & ~n13413;
  assign n13417 = n3397 & n4094;
  assign n13418 = ~n13412 & n13417;
  assign n13419 = n3128 & n13418;
  assign n13420 = n13416 & n13419;
  assign n13421 = ~pi0287 & ~n3405;
  assign n13422 = n13420 & n13421;
  assign n13423 = n3404 & n13422;
  assign n13424 = ~pi0039 & pi0228;
  assign n13425 = ~n13412 & ~n13413;
  assign n13426 = ~n13411 & n13425;
  assign n13427 = ~n13424 & ~n13426;
  assign n13428 = ~n13423 & n13427;
  assign po0385 = n13415 | ~n13428;
  assign n13430 = n2942 & n12367;
  assign n13431 = ~n2917 & ~n3033;
  assign n13432 = n13430 & n13431;
  assign n13433 = ~n2910 & n13432;
  assign n13434 = ~n4504 & n13433;
  assign n13435 = n2547 & n12368;
  assign n13436 = n13434 & n13435;
  assign n13437 = n2570 & n13436;
  assign n13438 = n3010 & n13437;
  assign n13439 = n12350 & n13438;
  assign n13440 = n12389 & n13439;
  assign n13441 = ~n2888 & n12371;
  assign n13442 = ~n2770 & ~n2901;
  assign n13443 = n2896 & n13442;
  assign n13444 = n2686 & n13443;
  assign n13445 = n12362 & n13444;
  assign n13446 = pi0786 & n4088;
  assign n13447 = n3404 & n13446;
  assign n13448 = n13421 & n13447;
  assign n13449 = n2777 & ~n13448;
  assign n13450 = n13445 & ~n13449;
  assign n13451 = n13441 & n13450;
  assign po0389 = ~n13440 | ~n13451;
  assign n13453 = ~pi0230 & ~pi0233;
  assign n13454 = ~n4970 & n4983;
  assign n13455 = n4973 & n13454;
  assign n13456 = pi1138 & n13455;
  assign n13457 = n4974 & n7400;
  assign n13458 = pi1136 & n13457;
  assign n13459 = ~n13456 & ~n13458;
  assign n13460 = n4964 & n4967;
  assign n13461 = n4974 & n13460;
  assign n13462 = ~n4970 & n13460;
  assign n13463 = n4973 & n13462;
  assign n13464 = n4970 & ~n4973;
  assign n13465 = n13460 & n13464;
  assign n13466 = ~n13463 & ~n13465;
  assign n13467 = ~n13461 & n13466;
  assign n13468 = pi1136 & ~n13467;
  assign n13469 = ~n4970 & n4973;
  assign n13470 = n7400 & n13469;
  assign n13471 = n4970 & n7400;
  assign n13472 = ~n4973 & n13471;
  assign n13473 = ~n13470 & ~n13472;
  assign n13474 = pi1137 & ~n13473;
  assign n13475 = ~n13468 & ~n13474;
  assign n13476 = n4970 & n4983;
  assign n13477 = ~n4973 & n13476;
  assign n13478 = pi1138 & n13477;
  assign n13479 = pi1137 & n4984;
  assign n13480 = ~n13478 & ~n13479;
  assign n13481 = n13475 & n13480;
  assign n13482 = n13459 & n13481;
  assign n13483 = ~pi0209 & n2429;
  assign n13484 = ~pi0213 & ~n2429;
  assign n13485 = ~n13483 & ~n13484;
  assign n13486 = ~n13482 & n13485;
  assign n13487 = pi1151 & n13455;
  assign n13488 = pi1147 & n13461;
  assign n13489 = pi1148 & n13465;
  assign n13490 = pi1149 & n13463;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = pi1149 & n13472;
  assign n13493 = pi1148 & n13457;
  assign n13494 = ~n13492 & ~n13493;
  assign n13495 = pi1150 & n13477;
  assign n13496 = pi1149 & n4984;
  assign n13497 = ~n13495 & ~n13496;
  assign n13498 = n13494 & n13497;
  assign n13499 = n13491 & n13498;
  assign n13500 = pi1150 & n13470;
  assign n13501 = n13499 & ~n13500;
  assign n13502 = ~n13488 & n13501;
  assign n13503 = ~n13487 & n13502;
  assign n13504 = ~n13485 & ~n13503;
  assign n13505 = ~n13486 & ~n13504;
  assign n13506 = pi0230 & ~n13505;
  assign po0390 = n13453 | n13506;
  assign n13508 = ~pi0230 & pi0234;
  assign n13509 = pi1148 & n13461;
  assign n13510 = pi1150 & n13455;
  assign n13511 = pi1149 & n13470;
  assign n13512 = ~n13510 & ~n13511;
  assign n13513 = pi1148 & n13463;
  assign n13514 = n13512 & ~n13513;
  assign n13515 = n13498 & n13514;
  assign n13516 = ~n13509 & n13515;
  assign n13517 = ~n13489 & n13516;
  assign n13518 = n13485 & ~n13517;
  assign n13519 = pi1148 & n13455;
  assign n13520 = pi1146 & n13457;
  assign n13521 = ~n13519 & ~n13520;
  assign n13522 = pi1146 & ~n13467;
  assign n13523 = pi1147 & ~n13473;
  assign n13524 = ~n13522 & ~n13523;
  assign n13525 = pi1148 & n13477;
  assign n13526 = pi1147 & n4984;
  assign n13527 = ~n13525 & ~n13526;
  assign n13528 = n13524 & n13527;
  assign n13529 = n13521 & n13528;
  assign n13530 = ~n13485 & ~n13529;
  assign n13531 = ~n13518 & ~n13530;
  assign n13532 = pi0230 & ~n13531;
  assign po0391 = n13508 | n13532;
  assign n13534 = ~pi0230 & pi0235;
  assign n13535 = pi1150 & n13472;
  assign n13536 = pi1149 & n13465;
  assign n13537 = ~n13535 & ~n13536;
  assign n13538 = pi1150 & n4984;
  assign n13539 = ~n13490 & ~n13538;
  assign n13540 = ~n13487 & n13539;
  assign n13541 = ~n13500 & n13540;
  assign n13542 = pi1151 & n13477;
  assign n13543 = pi1149 & n13457;
  assign n13544 = ~n13542 & ~n13543;
  assign n13545 = n13541 & n13544;
  assign n13546 = n13537 & n13545;
  assign n13547 = n13485 & ~n13546;
  assign n13548 = pi1149 & n13455;
  assign n13549 = pi1147 & n13457;
  assign n13550 = ~n13548 & ~n13549;
  assign n13551 = pi1149 & n13477;
  assign n13552 = pi1148 & n4984;
  assign n13553 = ~n13551 & ~n13552;
  assign n13554 = pi1148 & ~n13473;
  assign n13555 = pi1147 & ~n13466;
  assign n13556 = ~n13554 & ~n13555;
  assign n13557 = n13553 & n13556;
  assign n13558 = n13550 & n13557;
  assign n13559 = ~n13485 & ~n13558;
  assign n13560 = ~n13547 & ~n13559;
  assign n13561 = pi0230 & ~n13560;
  assign po0392 = n13534 | n13561;
  assign n13563 = ~pi0230 & ~pi0237;
  assign n13564 = pi1139 & n13455;
  assign n13565 = pi1137 & n13457;
  assign n13566 = ~n13564 & ~n13565;
  assign n13567 = pi1137 & ~n13467;
  assign n13568 = pi1138 & ~n13473;
  assign n13569 = ~n13567 & ~n13568;
  assign n13570 = pi1139 & n13477;
  assign n13571 = pi1138 & n4984;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = n13569 & n13572;
  assign n13574 = n13566 & n13573;
  assign n13575 = n13485 & ~n13574;
  assign n13576 = ~n13509 & ~n13538;
  assign n13577 = pi1152 & n13455;
  assign n13578 = pi1151 & n13470;
  assign n13579 = ~n13577 & ~n13578;
  assign n13580 = pi1150 & n13463;
  assign n13581 = n13579 & ~n13580;
  assign n13582 = n13544 & n13581;
  assign n13583 = n13537 & n13582;
  assign n13584 = n13576 & n13583;
  assign n13585 = ~n13485 & ~n13584;
  assign n13586 = ~n13575 & ~n13585;
  assign n13587 = pi0230 & ~n13586;
  assign po0394 = n13563 | n13587;
  assign n13589 = ~pi0230 & pi0238;
  assign n13590 = n13485 & ~n13488;
  assign n13591 = n13558 & n13590;
  assign n13592 = pi1147 & n13455;
  assign n13593 = pi1145 & n13457;
  assign n13594 = ~n13592 & ~n13593;
  assign n13595 = pi1145 & ~n13467;
  assign n13596 = pi1146 & ~n13473;
  assign n13597 = ~n13595 & ~n13596;
  assign n13598 = pi1147 & n13477;
  assign n13599 = pi1146 & n4984;
  assign n13600 = ~n13598 & ~n13599;
  assign n13601 = n13597 & n13600;
  assign n13602 = n13594 & n13601;
  assign n13603 = ~n13485 & n13602;
  assign n13604 = ~n13591 & ~n13603;
  assign n13605 = pi0230 & n13604;
  assign po0395 = n13589 | n13605;
  assign n13607 = ~pi0230 & pi0239;
  assign n13608 = ~n13485 & ~n13514;
  assign n13609 = n13485 & ~n13581;
  assign n13610 = ~n13608 & ~n13609;
  assign n13611 = pi0230 & ~n13610;
  assign po0396 = n13607 | n13611;
  assign n13613 = ~pi0230 & pi0240;
  assign n13614 = pi1143 & n13455;
  assign n13615 = pi1141 & n13457;
  assign n13616 = ~n13614 & ~n13615;
  assign n13617 = pi1141 & ~n13467;
  assign n13618 = pi1142 & ~n13473;
  assign n13619 = ~n13617 & ~n13618;
  assign n13620 = pi1143 & n13477;
  assign n13621 = pi1142 & n4984;
  assign n13622 = ~n13620 & ~n13621;
  assign n13623 = n13619 & n13622;
  assign n13624 = n13616 & n13623;
  assign n13625 = n13485 & ~n13624;
  assign n13626 = pi1141 & n13455;
  assign n13627 = pi1139 & n13457;
  assign n13628 = ~n13626 & ~n13627;
  assign n13629 = pi1139 & ~n13467;
  assign n13630 = pi1140 & ~n13473;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = pi1141 & n13477;
  assign n13633 = pi1140 & n4984;
  assign n13634 = ~n13632 & ~n13633;
  assign n13635 = n13631 & n13634;
  assign n13636 = n13628 & n13635;
  assign n13637 = ~n13485 & ~n13636;
  assign n13638 = ~n13625 & ~n13637;
  assign n13639 = pi0230 & ~n13638;
  assign po0397 = n13613 | n13639;
  assign n13641 = ~pi0230 & pi0241;
  assign n13642 = n13485 & ~n13602;
  assign n13643 = pi1145 & n13455;
  assign n13644 = pi1143 & n13457;
  assign n13645 = ~n13643 & ~n13644;
  assign n13646 = pi1143 & ~n13467;
  assign n13647 = pi1144 & ~n13473;
  assign n13648 = ~n13646 & ~n13647;
  assign n13649 = pi1145 & n13477;
  assign n13650 = pi1144 & n4984;
  assign n13651 = ~n13649 & ~n13650;
  assign n13652 = n13648 & n13651;
  assign n13653 = n13645 & n13652;
  assign n13654 = ~n13485 & ~n13653;
  assign n13655 = ~n13642 & ~n13654;
  assign n13656 = pi0230 & ~n13655;
  assign po0398 = n13641 | n13656;
  assign n13658 = ~pi0230 & pi0242;
  assign n13659 = pi1140 & n13455;
  assign n13660 = pi1138 & n13457;
  assign n13661 = ~n13659 & ~n13660;
  assign n13662 = pi1138 & ~n13467;
  assign n13663 = pi1139 & ~n13473;
  assign n13664 = ~n13662 & ~n13663;
  assign n13665 = pi1140 & n13477;
  assign n13666 = pi1139 & n4984;
  assign n13667 = ~n13665 & ~n13666;
  assign n13668 = n13664 & n13667;
  assign n13669 = n13661 & n13668;
  assign n13670 = n13485 & ~n13669;
  assign n13671 = ~n13482 & ~n13485;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = pi0230 & ~n13672;
  assign po0399 = n13658 | n13673;
  assign n13675 = pi0314 & ~n2477;
  assign n13676 = ~pi0081 & ~pi0085;
  assign n13677 = ~n4983 & ~n7400;
  assign n13678 = pi0314 & n2477;
  assign n13679 = ~n13677 & n13678;
  assign n13680 = ~n13676 & n13679;
  assign n13681 = ~n13675 & ~n13680;
  assign n13682 = pi0268 & pi0275;
  assign n13683 = pi0276 & pi0802;
  assign n13684 = pi0271 & n13683;
  assign n13685 = pi0273 & n13684;
  assign n13686 = pi0283 & n13685;
  assign n13687 = n13682 & n13686;
  assign n13688 = pi0272 & n13687;
  assign n13689 = pi0253 & pi0254;
  assign n13690 = n13688 & n13689;
  assign n13691 = ~pi0263 & n13690;
  assign n13692 = pi0267 & n13691;
  assign n13693 = ~pi0243 & n13692;
  assign n13694 = pi0243 & ~n13692;
  assign n13695 = ~n13693 & ~n13694;
  assign n13696 = ~n13681 & n13695;
  assign n13697 = ~pi0243 & n13681;
  assign n13698 = ~n13696 & ~n13697;
  assign n13699 = ~pi0230 & ~pi1085;
  assign n13700 = ~n13698 & n13699;
  assign n13701 = pi1149 & n4983;
  assign n13702 = pi1151 & n13460;
  assign n13703 = pi1150 & n7400;
  assign n13704 = ~n13702 & ~n13703;
  assign n13705 = ~n13701 & n13704;
  assign n13706 = ~n13699 & ~n13705;
  assign po0400 = n13700 | n13706;
  assign n13708 = ~pi0230 & pi0244;
  assign n13709 = n13485 & ~n13636;
  assign n13710 = ~n13485 & ~n13574;
  assign n13711 = ~n13709 & ~n13710;
  assign n13712 = pi0230 & ~n13711;
  assign po0401 = n13708 | n13712;
  assign n13714 = ~pi0230 & pi0245;
  assign n13715 = pi1142 & n13455;
  assign n13716 = pi1140 & n13457;
  assign n13717 = ~n13715 & ~n13716;
  assign n13718 = pi1140 & ~n13467;
  assign n13719 = pi1141 & ~n13473;
  assign n13720 = ~n13718 & ~n13719;
  assign n13721 = pi1142 & n13477;
  assign n13722 = pi1141 & n4984;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = n13720 & n13723;
  assign n13725 = n13717 & n13724;
  assign n13726 = n13485 & ~n13725;
  assign n13727 = ~n13485 & ~n13669;
  assign n13728 = ~n13726 & ~n13727;
  assign n13729 = pi0230 & ~n13728;
  assign po0402 = n13714 | n13729;
  assign n13731 = ~pi0230 & pi0246;
  assign n13732 = pi1144 & n13455;
  assign n13733 = pi1142 & n13457;
  assign n13734 = ~n13732 & ~n13733;
  assign n13735 = pi1142 & ~n13467;
  assign n13736 = pi1143 & ~n13473;
  assign n13737 = ~n13735 & ~n13736;
  assign n13738 = pi1144 & n13477;
  assign n13739 = pi1143 & n4984;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = n13737 & n13740;
  assign n13742 = n13734 & n13741;
  assign n13743 = n13485 & ~n13742;
  assign n13744 = ~n13485 & ~n13725;
  assign n13745 = ~n13743 & ~n13744;
  assign n13746 = pi0230 & ~n13745;
  assign po0403 = n13731 | n13746;
  assign n13748 = ~pi0230 & pi0247;
  assign n13749 = n13485 & ~n13653;
  assign n13750 = ~n13485 & ~n13624;
  assign n13751 = ~n13749 & ~n13750;
  assign n13752 = pi0230 & ~n13751;
  assign po0404 = n13748 | n13752;
  assign n13754 = ~pi0230 & pi0248;
  assign n13755 = pi1146 & n13455;
  assign n13756 = pi1144 & n13457;
  assign n13757 = ~n13755 & ~n13756;
  assign n13758 = pi1144 & ~n13467;
  assign n13759 = pi1145 & ~n13473;
  assign n13760 = ~n13758 & ~n13759;
  assign n13761 = pi1146 & n13477;
  assign n13762 = pi1145 & n4984;
  assign n13763 = ~n13761 & ~n13762;
  assign n13764 = n13760 & n13763;
  assign n13765 = n13757 & n13764;
  assign n13766 = n13485 & ~n13765;
  assign n13767 = ~n13485 & ~n13742;
  assign n13768 = ~n13766 & ~n13767;
  assign n13769 = pi0230 & ~n13768;
  assign po0405 = n13754 | n13769;
  assign n13771 = ~pi0230 & pi0249;
  assign n13772 = n13485 & ~n13529;
  assign n13773 = ~n13485 & ~n13765;
  assign n13774 = ~n13772 & ~n13773;
  assign n13775 = pi0230 & ~n13774;
  assign po0406 = n13771 | n13775;
  assign n13777 = ~n2813 & ~n3042;
  assign n13778 = ~pi0250 & n12350;
  assign n13779 = ~n13777 & ~n13778;
  assign n13780 = ~pi0250 & ~n12350;
  assign n13781 = n13777 & ~n13780;
  assign n13782 = ~n13779 & ~n13781;
  assign n13783 = ~n13777 & n13780;
  assign po0407 = n13782 | n13783;
  assign n13785 = ~pi0199 & ~pi0200;
  assign n13786 = pi0897 & n13785;
  assign n13787 = pi1047 & n13786;
  assign n13788 = ~pi0199 & pi0200;
  assign n13789 = ~pi0476 & n13788;
  assign n13790 = pi1033 & n13789;
  assign n13791 = pi0251 & ~n13789;
  assign n13792 = ~n13790 & ~n13791;
  assign n13793 = ~n13786 & ~n13792;
  assign po0408 = n13787 | n13793;
  assign n13795 = pi1087 & ~n3539;
  assign n13796 = pi1086 & ~n13795;
  assign n13797 = pi0252 & n13796;
  assign n13798 = n3397 & n4087;
  assign po0409 = n13797 | n13798;
  assign n13800 = pi0253 & n13688;
  assign n13801 = ~pi0253 & ~n13688;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~n13681 & n13802;
  assign n13804 = pi0253 & n13681;
  assign n13805 = ~n13803 & ~n13804;
  assign n13806 = n13699 & ~n13805;
  assign n13807 = pi1145 & n4983;
  assign n13808 = pi1147 & n13460;
  assign n13809 = pi1146 & n7400;
  assign n13810 = ~n13808 & ~n13809;
  assign n13811 = ~n13807 & n13810;
  assign n13812 = ~n13699 & ~n13811;
  assign po0410 = n13806 | n13812;
  assign n13814 = pi0272 & pi0275;
  assign n13815 = pi0253 & pi0268;
  assign n13816 = n13814 & n13815;
  assign n13817 = n13686 & n13816;
  assign n13818 = pi0254 & n13817;
  assign n13819 = ~pi0254 & ~n13817;
  assign n13820 = ~n13818 & ~n13819;
  assign n13821 = ~n13681 & n13820;
  assign n13822 = pi0254 & n13681;
  assign n13823 = ~n13821 & ~n13822;
  assign n13824 = n13699 & ~n13823;
  assign n13825 = pi1146 & n4983;
  assign n13826 = pi1148 & n13460;
  assign n13827 = pi1147 & n7400;
  assign n13828 = ~n13826 & ~n13827;
  assign n13829 = ~n13825 & n13828;
  assign n13830 = ~n13699 & ~n13829;
  assign po0411 = n13824 | n13830;
  assign n13832 = pi1043 & n13786;
  assign n13833 = pi1030 & n13789;
  assign n13834 = pi0255 & ~n13789;
  assign n13835 = ~n13833 & ~n13834;
  assign n13836 = ~n13786 & ~n13835;
  assign po0412 = n13832 | n13836;
  assign n13838 = pi1042 & n13786;
  assign n13839 = pi1064 & n13789;
  assign n13840 = pi0256 & ~n13789;
  assign n13841 = ~n13839 & ~n13840;
  assign n13842 = ~n13786 & ~n13841;
  assign po0413 = n13838 | n13842;
  assign n13844 = pi1078 & n13786;
  assign n13845 = pi1059 & n13789;
  assign n13846 = pi0257 & ~n13789;
  assign n13847 = ~n13845 & ~n13846;
  assign n13848 = ~n13786 & ~n13847;
  assign po0414 = n13844 | n13848;
  assign n13850 = pi1066 & n13786;
  assign n13851 = pi1056 & n13789;
  assign n13852 = pi0258 & ~n13789;
  assign n13853 = ~n13851 & ~n13852;
  assign n13854 = ~n13786 & ~n13853;
  assign po0415 = n13850 | n13854;
  assign n13856 = pi1053 & n13786;
  assign n13857 = pi1063 & n13789;
  assign n13858 = pi0259 & ~n13789;
  assign n13859 = ~n13857 & ~n13858;
  assign n13860 = ~n13786 & ~n13859;
  assign po0416 = n13856 | n13860;
  assign n13862 = pi1038 & n13786;
  assign n13863 = pi1061 & n13789;
  assign n13864 = pi0260 & ~n13789;
  assign n13865 = ~n13863 & ~n13864;
  assign n13866 = ~n13786 & ~n13865;
  assign po0417 = n13862 | n13866;
  assign n13868 = pi1031 & n13786;
  assign n13869 = pi1034 & n13789;
  assign n13870 = pi0261 & ~n13789;
  assign n13871 = ~n13869 & ~n13870;
  assign n13872 = ~n13786 & ~n13871;
  assign po0418 = n13868 | n13872;
  assign n13874 = ~pi0123 & pi0228;
  assign n13875 = ~pi0228 & pi1087;
  assign n13876 = ~n13874 & ~n13875;
  assign n13877 = ~pi0262 & n13876;
  assign n13878 = ~n13472 & ~n13477;
  assign n13879 = ~n4984 & n13878;
  assign n13880 = pi1136 & ~n13879;
  assign n13881 = ~n13455 & ~n13470;
  assign n13882 = pi1136 & ~n13881;
  assign n13883 = ~n13880 & ~n13882;
  assign n13884 = ~n13876 & ~n13883;
  assign po0419 = n13877 | n13884;
  assign n13886 = n13686 & n13814;
  assign n13887 = n13815 & n13886;
  assign n13888 = pi0267 & n13887;
  assign n13889 = pi0254 & n13888;
  assign n13890 = ~pi0263 & n13889;
  assign n13891 = pi0263 & ~n13889;
  assign n13892 = ~n13890 & ~n13891;
  assign n13893 = ~n13681 & n13892;
  assign n13894 = ~pi0263 & n13681;
  assign n13895 = ~n13893 & ~n13894;
  assign n13896 = n13699 & ~n13895;
  assign n13897 = pi1148 & n4983;
  assign n13898 = pi1150 & n13460;
  assign n13899 = pi1149 & n7400;
  assign n13900 = ~n13898 & ~n13899;
  assign n13901 = ~n13897 & n13900;
  assign n13902 = ~n13699 & ~n13901;
  assign po0420 = n13896 | n13902;
  assign n13904 = pi1135 & n4983;
  assign n13905 = pi1137 & n13460;
  assign n13906 = pi1136 & n7400;
  assign n13907 = ~n13905 & ~n13906;
  assign n13908 = ~n13904 & n13907;
  assign n13909 = ~n13699 & ~n13908;
  assign n13910 = pi0796 & ~n13681;
  assign n13911 = ~pi0264 & n13681;
  assign n13912 = ~n13910 & ~n13911;
  assign n13913 = n13699 & ~n13912;
  assign po0421 = n13909 | n13913;
  assign n13915 = pi1136 & n4983;
  assign n13916 = pi1138 & n13460;
  assign n13917 = pi1137 & n7400;
  assign n13918 = ~n13916 & ~n13917;
  assign n13919 = ~n13915 & n13918;
  assign n13920 = ~n13699 & ~n13919;
  assign n13921 = pi0819 & ~n13681;
  assign n13922 = ~pi0265 & n13681;
  assign n13923 = ~n13921 & ~n13922;
  assign n13924 = n13699 & ~n13923;
  assign po0422 = n13920 | n13924;
  assign n13926 = pi1128 & n4983;
  assign n13927 = pi1130 & n13460;
  assign n13928 = pi1129 & n7400;
  assign n13929 = ~n13927 & ~n13928;
  assign n13930 = ~n13926 & n13929;
  assign n13931 = ~n13699 & ~n13930;
  assign n13932 = pi0948 & ~n13681;
  assign n13933 = pi0266 & n13681;
  assign n13934 = ~n13932 & ~n13933;
  assign n13935 = n13699 & ~n13934;
  assign po0423 = n13931 | n13935;
  assign n13937 = pi1149 & n13460;
  assign n13938 = pi1148 & n7400;
  assign n13939 = ~n13937 & ~n13938;
  assign n13940 = pi1147 & n4983;
  assign n13941 = n13939 & ~n13940;
  assign n13942 = ~n13699 & ~n13941;
  assign n13943 = pi0271 & pi0273;
  assign n13944 = pi0272 & n13943;
  assign n13945 = pi0283 & n13944;
  assign n13946 = n13683 & n13945;
  assign n13947 = n13682 & n13946;
  assign n13948 = n13689 & n13947;
  assign n13949 = pi0267 & n13948;
  assign n13950 = ~pi0267 & ~n13948;
  assign n13951 = ~n13949 & ~n13950;
  assign n13952 = ~n13681 & n13951;
  assign n13953 = pi0267 & n13681;
  assign n13954 = ~n13952 & ~n13953;
  assign n13955 = n13699 & ~n13954;
  assign po0424 = n13942 | n13955;
  assign n13957 = pi1144 & n4983;
  assign n13958 = pi1146 & n13460;
  assign n13959 = pi1145 & n7400;
  assign n13960 = ~n13958 & ~n13959;
  assign n13961 = ~n13957 & n13960;
  assign n13962 = ~n13699 & ~n13961;
  assign n13963 = pi0268 & ~n13886;
  assign n13964 = ~pi0268 & n13886;
  assign n13965 = ~n13963 & ~n13964;
  assign n13966 = ~n13681 & ~n13965;
  assign n13967 = pi0268 & n13681;
  assign n13968 = ~n13966 & ~n13967;
  assign n13969 = n13699 & ~n13968;
  assign po0425 = n13962 | n13969;
  assign n13971 = pi1130 & n4983;
  assign n13972 = pi1132 & n13460;
  assign n13973 = pi1131 & n7400;
  assign n13974 = ~n13972 & ~n13973;
  assign n13975 = ~n13971 & n13974;
  assign n13976 = ~n13699 & ~n13975;
  assign n13977 = pi0817 & ~n13681;
  assign n13978 = ~pi0269 & n13681;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = n13699 & ~n13979;
  assign po0426 = n13976 | n13980;
  assign n13982 = pi1133 & n4983;
  assign n13983 = pi1135 & n13460;
  assign n13984 = pi1134 & n7400;
  assign n13985 = ~n13983 & ~n13984;
  assign n13986 = ~n13982 & n13985;
  assign n13987 = ~n13699 & ~n13986;
  assign n13988 = pi0805 & ~n13681;
  assign n13989 = ~pi0270 & n13681;
  assign n13990 = ~n13988 & ~n13989;
  assign n13991 = n13699 & ~n13990;
  assign po0427 = n13987 | n13991;
  assign n13993 = pi1139 & n4983;
  assign n13994 = pi1141 & n13460;
  assign n13995 = pi1140 & n7400;
  assign n13996 = ~n13994 & ~n13995;
  assign n13997 = ~n13993 & n13996;
  assign n13998 = ~n13699 & ~n13997;
  assign n13999 = pi0271 & ~n13683;
  assign n14000 = ~pi0271 & n13683;
  assign n14001 = ~n13999 & ~n14000;
  assign n14002 = ~n13681 & ~n14001;
  assign n14003 = pi0271 & n13681;
  assign n14004 = ~n14002 & ~n14003;
  assign n14005 = n13699 & ~n14004;
  assign po0428 = n13998 | n14005;
  assign n14007 = pi1142 & n4983;
  assign n14008 = pi1144 & n13460;
  assign n14009 = pi1143 & n7400;
  assign n14010 = ~n14008 & ~n14009;
  assign n14011 = ~n14007 & n14010;
  assign n14012 = ~n13699 & ~n14011;
  assign n14013 = pi0272 & ~n13686;
  assign n14014 = ~pi0272 & n13686;
  assign n14015 = ~n14013 & ~n14014;
  assign n14016 = ~n13681 & ~n14015;
  assign n14017 = pi0272 & n13681;
  assign n14018 = ~n14016 & ~n14017;
  assign n14019 = n13699 & ~n14018;
  assign po0429 = n14012 | n14019;
  assign n14021 = pi1140 & n4983;
  assign n14022 = pi1142 & n13460;
  assign n14023 = pi1141 & n7400;
  assign n14024 = ~n14022 & ~n14023;
  assign n14025 = ~n14021 & n14024;
  assign n14026 = ~n13699 & ~n14025;
  assign n14027 = pi0273 & ~n13684;
  assign n14028 = ~pi0273 & n13684;
  assign n14029 = ~n14027 & ~n14028;
  assign n14030 = ~n13681 & ~n14029;
  assign n14031 = pi0273 & n13681;
  assign n14032 = ~n14030 & ~n14031;
  assign n14033 = n13699 & ~n14032;
  assign po0430 = n14026 | n14033;
  assign n14035 = pi1137 & n4983;
  assign n14036 = pi1139 & n13460;
  assign n14037 = pi1138 & n7400;
  assign n14038 = ~n14036 & ~n14037;
  assign n14039 = ~n14035 & n14038;
  assign n14040 = ~n13699 & ~n14039;
  assign n14041 = pi0659 & ~n13681;
  assign n14042 = ~pi0274 & n13681;
  assign n14043 = ~n14041 & ~n14042;
  assign n14044 = n13699 & ~n14043;
  assign po0431 = n14040 | n14044;
  assign n14046 = pi1143 & n4983;
  assign n14047 = pi1145 & n13460;
  assign n14048 = pi1144 & n7400;
  assign n14049 = ~n14047 & ~n14048;
  assign n14050 = ~n14046 & n14049;
  assign n14051 = ~n13699 & ~n14050;
  assign n14052 = pi0275 & ~n13946;
  assign n14053 = ~pi0275 & n13946;
  assign n14054 = ~n14052 & ~n14053;
  assign n14055 = ~n13681 & ~n14054;
  assign n14056 = pi0275 & n13681;
  assign n14057 = ~n14055 & ~n14056;
  assign n14058 = n13699 & ~n14057;
  assign po0432 = n14051 | n14058;
  assign n14060 = pi1138 & n4983;
  assign n14061 = pi1140 & n13460;
  assign n14062 = pi1139 & n7400;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = ~n14060 & n14063;
  assign n14065 = ~n13699 & ~n14064;
  assign n14066 = ~pi0276 & pi0802;
  assign n14067 = pi0276 & ~pi0802;
  assign n14068 = ~n14066 & ~n14067;
  assign n14069 = ~n13681 & ~n14068;
  assign n14070 = pi0276 & n13681;
  assign n14071 = ~n14069 & ~n14070;
  assign n14072 = n13699 & ~n14071;
  assign po0433 = n14065 | n14072;
  assign n14074 = pi1134 & n4983;
  assign n14075 = pi1136 & n13460;
  assign n14076 = pi1135 & n7400;
  assign n14077 = ~n14075 & ~n14076;
  assign n14078 = ~n14074 & n14077;
  assign n14079 = ~n13699 & ~n14078;
  assign n14080 = pi0820 & ~n13681;
  assign n14081 = ~pi0277 & n13681;
  assign n14082 = ~n14080 & ~n14081;
  assign n14083 = n13699 & ~n14082;
  assign po0434 = n14079 | n14083;
  assign n14085 = pi1128 & n13460;
  assign n14086 = pi1126 & n4983;
  assign n14087 = pi1127 & n7400;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n14085 & n14088;
  assign n14090 = ~n13699 & ~n14089;
  assign n14091 = pi0976 & ~n13681;
  assign n14092 = pi0278 & n13681;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = n13699 & ~n14093;
  assign po0435 = n14090 | n14094;
  assign n14096 = pi1128 & n7400;
  assign n14097 = pi1127 & n4983;
  assign n14098 = pi1129 & n13460;
  assign n14099 = ~n14097 & ~n14098;
  assign n14100 = ~n14096 & n14099;
  assign n14101 = ~n13699 & ~n14100;
  assign n14102 = pi0958 & ~n13681;
  assign n14103 = pi0279 & n13681;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = n13699 & ~n14104;
  assign po0436 = n14101 | n14105;
  assign n14107 = pi1129 & n4983;
  assign n14108 = pi1131 & n13460;
  assign n14109 = pi1130 & n7400;
  assign n14110 = ~n14108 & ~n14109;
  assign n14111 = ~n14107 & n14110;
  assign n14112 = ~n13699 & ~n14111;
  assign n14113 = pi0914 & ~n13681;
  assign n14114 = ~pi0280 & n13681;
  assign n14115 = ~n14113 & ~n14114;
  assign n14116 = n13699 & ~n14115;
  assign po0437 = n14112 | n14116;
  assign n14118 = pi1131 & n4983;
  assign n14119 = pi1133 & n13460;
  assign n14120 = pi1132 & n7400;
  assign n14121 = ~n14119 & ~n14120;
  assign n14122 = ~n14118 & n14121;
  assign n14123 = ~n13699 & ~n14122;
  assign n14124 = pi0830 & ~n13681;
  assign n14125 = ~pi0281 & n13681;
  assign n14126 = ~n14124 & ~n14125;
  assign n14127 = n13699 & ~n14126;
  assign po0438 = n14123 | n14127;
  assign n14129 = pi1132 & n4983;
  assign n14130 = pi1134 & n13460;
  assign n14131 = pi1133 & n7400;
  assign n14132 = ~n14130 & ~n14131;
  assign n14133 = ~n14129 & n14132;
  assign n14134 = ~n13699 & ~n14133;
  assign n14135 = pi0836 & ~n13681;
  assign n14136 = ~pi0282 & n13681;
  assign n14137 = ~n14135 & ~n14136;
  assign n14138 = n13699 & ~n14137;
  assign po0439 = n14134 | n14138;
  assign n14140 = pi1141 & n4983;
  assign n14141 = pi1143 & n13460;
  assign n14142 = pi1142 & n7400;
  assign n14143 = ~n14141 & ~n14142;
  assign n14144 = ~n14140 & n14143;
  assign n14145 = ~n13699 & ~n14144;
  assign n14146 = pi0283 & ~n13685;
  assign n14147 = ~pi0283 & n13685;
  assign n14148 = ~n14146 & ~n14147;
  assign n14149 = ~n13681 & ~n14148;
  assign n14150 = pi0283 & n13681;
  assign n14151 = ~n14149 & ~n14150;
  assign n14152 = n13699 & ~n14151;
  assign po0440 = n14145 | n14152;
  assign n14154 = pi1137 & ~n13876;
  assign n14155 = ~n13455 & ~n13477;
  assign n14156 = n14154 & ~n14155;
  assign n14157 = ~pi0284 & n13876;
  assign po0441 = n14156 | n14157;
  assign n14159 = pi0286 & pi0288;
  assign n14160 = pi0289 & n14159;
  assign n14161 = pi0285 & n14160;
  assign n14162 = ~pi0285 & ~n14160;
  assign n14163 = ~n14161 & ~n14162;
  assign n14164 = ~n3581 & po0637;
  assign n14165 = ~n14163 & n14164;
  assign n14166 = n3581 & ~po0637;
  assign n14167 = ~pi0285 & ~n14166;
  assign n14168 = pi0285 & ~n3576;
  assign n14169 = ~n3577 & ~n14168;
  assign n14170 = n14166 & n14169;
  assign n14171 = ~n14167 & ~n14170;
  assign n14172 = ~n14164 & ~n14171;
  assign n14173 = ~n14165 & ~n14172;
  assign po0442 = ~pi0793 & n14173;
  assign n14175 = pi0286 & ~n14166;
  assign n14176 = ~n3575 & ~n14159;
  assign n14177 = n14166 & ~n14176;
  assign n14178 = ~n14175 & ~n14177;
  assign n14179 = ~n14164 & ~n14178;
  assign n14180 = pi0286 & ~pi0288;
  assign n14181 = ~pi0286 & pi0288;
  assign n14182 = ~n14180 & ~n14181;
  assign n14183 = n14164 & ~n14182;
  assign n14184 = ~n14179 & ~n14183;
  assign po0443 = ~pi0793 & ~n14184;
  assign n14186 = ~pi0287 & pi0457;
  assign po0444 = ~pi0332 & ~n14186;
  assign n14188 = ~pi0288 & n14164;
  assign n14189 = pi0288 & ~n14166;
  assign n14190 = ~pi0288 & n14166;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = ~n14164 & ~n14191;
  assign n14193 = ~n14188 & ~n14192;
  assign po0445 = ~pi0793 & ~n14193;
  assign n14195 = ~pi0289 & ~n14159;
  assign n14196 = ~n14160 & ~n14195;
  assign n14197 = n14164 & ~n14196;
  assign n14198 = ~pi0289 & ~n14166;
  assign n14199 = pi0289 & ~n3575;
  assign n14200 = ~n3576 & ~n14199;
  assign n14201 = n14166 & n14200;
  assign n14202 = ~n14198 & ~n14201;
  assign n14203 = ~n14164 & ~n14202;
  assign n14204 = ~n14197 & ~n14203;
  assign po0446 = ~pi0793 & n14204;
  assign n14206 = ~pi0476 & pi1042;
  assign n14207 = pi0290 & pi0476;
  assign po0447 = n14206 | n14207;
  assign n14209 = ~pi0476 & pi1043;
  assign n14210 = pi0291 & pi0476;
  assign po0448 = n14209 | n14210;
  assign n14212 = ~pi0476 & pi1078;
  assign n14213 = pi0292 & pi0476;
  assign po0449 = n14212 | n14213;
  assign n14215 = ~pi0476 & pi1053;
  assign n14216 = pi0293 & pi0476;
  assign po0450 = n14215 | n14216;
  assign n14218 = ~pi0476 & pi1066;
  assign n14219 = pi0294 & pi0476;
  assign po0451 = n14218 | n14219;
  assign n14221 = ~pi0476 & pi1047;
  assign n14222 = pi0295 & pi0476;
  assign po0452 = n14221 | n14222;
  assign n14224 = ~pi0476 & pi1031;
  assign n14225 = pi0296 & pi0476;
  assign po0453 = n14224 | n14225;
  assign n14227 = ~pi0476 & pi1038;
  assign n14228 = pi0297 & pi0476;
  assign po0454 = n14227 | n14228;
  assign n14230 = ~pi0478 & pi1038;
  assign n14231 = pi0298 & pi0478;
  assign po0455 = n14230 | n14231;
  assign n14233 = pi0039 & n5891;
  assign n14234 = n13169 & n13175;
  assign n14235 = n2868 & n12262;
  assign n14236 = ~pi0087 & n2992;
  assign n14237 = n13133 & n14236;
  assign n14238 = n2972 & n14237;
  assign n14239 = n13127 & n14238;
  assign n14240 = n14235 & n14239;
  assign n14241 = n2974 & n14240;
  assign n14242 = ~pi0066 & n14241;
  assign n14243 = ~po1049 & n14242;
  assign n14244 = n13145 & n14243;
  assign n14245 = n2980 & n12275;
  assign n14246 = n14244 & n14245;
  assign n14247 = n12260 & n14246;
  assign n14248 = n2983 & n14247;
  assign n14249 = n13165 & n14248;
  assign n14250 = ~n2639 & ~n3107;
  assign n14251 = n14248 & ~n14250;
  assign n14252 = ~pi0053 & n14251;
  assign n14253 = ~n14249 & ~n14252;
  assign n14254 = n14234 & ~n14253;
  assign n14255 = n2466 & n14254;
  assign n14256 = n13171 & n14255;
  assign n14257 = ~pi0039 & n14256;
  assign n14258 = n13177 & n14257;
  assign po0456 = n14233 | n14258;
  assign n14260 = ~pi0300 & ~pi0312;
  assign n14261 = pi0300 & pi0312;
  assign n14262 = ~n14260 & ~n14261;
  assign n14263 = n6892 & ~n14262;
  assign n14264 = pi0300 & ~n6892;
  assign n14265 = ~n14263 & ~n14264;
  assign po0457 = pi0055 | ~n14265;
  assign n14267 = pi0301 & n14260;
  assign n14268 = ~pi0301 & ~n14260;
  assign n14269 = ~n14267 & ~n14268;
  assign n14270 = n6892 & ~n14269;
  assign n14271 = ~pi0301 & ~n6892;
  assign n14272 = ~n14270 & ~n14271;
  assign po0458 = ~pi0055 & ~n14272;
  assign n14274 = pi0273 & n2440;
  assign n14275 = ~pi0237 & n3128;
  assign n14276 = ~n14274 & ~n14275;
  assign n14277 = pi0937 & n3132;
  assign n14278 = pi1142 & ~n3132;
  assign n14279 = ~n14277 & ~n14278;
  assign n14280 = ~n2439 & ~n14279;
  assign po0459 = ~n14276 | n14280;
  assign n14282 = ~pi0478 & pi1043;
  assign n14283 = pi0303 & pi0478;
  assign po0460 = n14282 | n14283;
  assign n14285 = ~pi0478 & pi1042;
  assign n14286 = pi0304 & pi0478;
  assign po0461 = n14285 | n14286;
  assign n14288 = ~pi0478 & pi1078;
  assign n14289 = pi0305 & pi0478;
  assign po0462 = n14288 | n14289;
  assign n14291 = ~pi0478 & pi1053;
  assign n14292 = pi0306 & pi0478;
  assign po0463 = n14291 | n14292;
  assign n14294 = ~pi0478 & pi1047;
  assign n14295 = pi0307 & pi0478;
  assign po0464 = n14294 | n14295;
  assign n14297 = ~pi0478 & pi1031;
  assign n14298 = pi0308 & pi0478;
  assign po0465 = n14297 | n14298;
  assign n14300 = ~pi0478 & pi1066;
  assign n14301 = pi0309 & pi0478;
  assign po0466 = n14300 | n14301;
  assign n14303 = pi0271 & n2440;
  assign n14304 = ~pi0233 & n3128;
  assign n14305 = ~n14303 & ~n14304;
  assign n14306 = pi0934 & n3132;
  assign n14307 = pi1141 & ~n3132;
  assign n14308 = ~n14306 & ~n14307;
  assign n14309 = ~n2439 & ~n14308;
  assign po0467 = ~n14305 | n14309;
  assign n14311 = ~pi0311 & ~n6892;
  assign n14312 = ~pi0311 & n14267;
  assign n14313 = pi0311 & ~n14267;
  assign n14314 = ~n14312 & ~n14313;
  assign n14315 = n6892 & n14314;
  assign n14316 = ~n14311 & ~n14315;
  assign po0468 = ~pi0055 & ~n14316;
  assign n14318 = pi0312 & n6892;
  assign n14319 = ~pi0312 & ~n6892;
  assign n14320 = ~n14318 & ~n14319;
  assign po0469 = ~pi0055 & n14320;
  assign n14322 = pi0314 & po0740;
  assign n14323 = ~n2604 & ~n14322;
  assign n14324 = n2662 & n14323;
  assign n14325 = ~n2662 & ~po0740;
  assign n14326 = n2604 & n14325;
  assign po0634 = ~n14324 & ~n14326;
  assign n14328 = ~pi0954 & ~po0634;
  assign n14329 = ~pi0313 & pi0954;
  assign po0470 = n14328 | n14329;
  assign n14331 = n12147 & n12158;
  assign n14332 = ~pi0051 & n14331;
  assign n14333 = n12140 & ~n12180;
  assign n14334 = n12442 & n14333;
  assign po0471 = n14332 & n14334;
  assign n14336 = ~pi0340 & po0637;
  assign n14337 = pi1074 & n14336;
  assign n14338 = pi0315 & ~n14336;
  assign po0472 = n14337 | n14338;
  assign n14340 = pi1041 & n14336;
  assign n14341 = pi0316 & ~n14336;
  assign po0473 = n14340 | n14341;
  assign n14343 = ~pi0330 & po0637;
  assign n14344 = pi1072 & n14343;
  assign n14345 = pi0317 & ~n14343;
  assign po0474 = n14344 | n14345;
  assign n14347 = ~pi0341 & po0637;
  assign n14348 = pi1068 & n14347;
  assign n14349 = pi0318 & ~n14347;
  assign po0475 = n14348 | n14349;
  assign n14351 = pi1066 & n14347;
  assign n14352 = pi0319 & ~n14347;
  assign po0476 = n14351 | n14352;
  assign n14354 = pi1042 & n14336;
  assign n14355 = pi0320 & ~n14336;
  assign po0477 = n14354 | n14355;
  assign n14357 = pi1052 & n14336;
  assign n14358 = pi0321 & ~n14336;
  assign po0478 = n14357 | n14358;
  assign n14360 = pi1045 & n14336;
  assign n14361 = pi0322 & ~n14336;
  assign po0479 = n14360 | n14361;
  assign n14363 = pi1059 & n14336;
  assign n14364 = pi0323 & ~n14336;
  assign po0480 = n14363 | n14364;
  assign n14366 = pi1080 & n14347;
  assign n14367 = pi0324 & ~n14347;
  assign po0481 = n14366 | n14367;
  assign n14369 = pi1057 & n14347;
  assign n14370 = pi0325 & ~n14347;
  assign po0482 = n14369 | n14370;
  assign n14372 = pi1051 & n14347;
  assign n14373 = pi0326 & ~n14347;
  assign po0483 = n14372 | n14373;
  assign n14375 = pi1034 & n14336;
  assign n14376 = pi0327 & ~n14336;
  assign po0484 = n14375 | n14376;
  assign n14378 = pi1052 & n14347;
  assign n14379 = pi0328 & ~n14347;
  assign po0485 = n14378 | n14379;
  assign n14381 = pi1037 & n14347;
  assign n14382 = pi0329 & ~n14347;
  assign po0486 = n14381 | n14382;
  assign n14384 = pi1086 & ~n3578;
  assign n14385 = ~pi0330 & ~po0637;
  assign n14386 = ~n14336 & ~n14385;
  assign po0487 = n14384 & ~n14386;
  assign n14388 = ~pi0331 & ~po0637;
  assign n14389 = ~n14347 & ~n14388;
  assign po0488 = n14384 & ~n14389;
  assign n14391 = ~n2780 & ~n2798;
  assign po0489 = n2784 | ~n14391;
  assign n14393 = pi1034 & n14347;
  assign n14394 = pi0333 & ~n14347;
  assign po0490 = n14393 | n14394;
  assign n14396 = pi1059 & n14347;
  assign n14397 = pi0334 & ~n14347;
  assign po0491 = n14396 | n14397;
  assign n14399 = pi1063 & n14347;
  assign n14400 = pi0335 & ~n14347;
  assign po0492 = n14399 | n14400;
  assign n14402 = pi1064 & n14343;
  assign n14403 = pi0336 & ~n14343;
  assign po0493 = n14402 | n14403;
  assign n14405 = pi1038 & n14343;
  assign n14406 = pi0337 & ~n14343;
  assign po0494 = n14405 | n14406;
  assign n14408 = pi1066 & n14343;
  assign n14409 = pi0338 & ~n14343;
  assign po0495 = n14408 | n14409;
  assign n14411 = pi1080 & n14343;
  assign n14412 = pi0339 & ~n14343;
  assign po0496 = n14411 | n14412;
  assign n14414 = ~pi0331 & po0637;
  assign n14415 = ~pi0340 & ~po0637;
  assign n14416 = n14384 & ~n14415;
  assign po0497 = n14414 | ~n14416;
  assign n14418 = ~pi0341 & ~po0637;
  assign n14419 = ~n14343 & ~n14418;
  assign po0498 = n14384 & ~n14419;
  assign n14421 = pi1043 & n14336;
  assign n14422 = pi0342 & ~n14336;
  assign po0499 = n14421 | n14422;
  assign n14424 = pi1056 & n14336;
  assign n14425 = pi0343 & ~n14336;
  assign po0500 = n14424 | n14425;
  assign n14427 = pi1063 & n14336;
  assign n14428 = pi0344 & ~n14336;
  assign po0501 = n14427 | n14428;
  assign n14430 = pi1033 & n14336;
  assign n14431 = pi0345 & ~n14336;
  assign po0502 = n14430 | n14431;
  assign n14433 = pi1061 & n14336;
  assign n14434 = pi0346 & ~n14336;
  assign po0503 = n14433 | n14434;
  assign n14436 = pi1049 & n14336;
  assign n14437 = pi0347 & ~n14336;
  assign po0504 = n14436 | n14437;
  assign n14439 = pi1081 & n14336;
  assign n14440 = pi0348 & ~n14336;
  assign po0505 = n14439 | n14440;
  assign n14442 = pi1037 & n14336;
  assign n14443 = pi0349 & ~n14336;
  assign po0506 = n14442 | n14443;
  assign n14445 = pi1029 & n14336;
  assign n14446 = pi0350 & ~n14336;
  assign po0507 = n14445 | n14446;
  assign n14448 = pi1073 & n14336;
  assign n14449 = pi0351 & ~n14336;
  assign po0508 = n14448 | n14449;
  assign n14451 = pi1072 & n14336;
  assign n14452 = pi0352 & ~n14336;
  assign po0509 = n14451 | n14452;
  assign n14454 = pi1057 & n14336;
  assign n14455 = pi0353 & ~n14336;
  assign po0510 = n14454 | n14455;
  assign n14457 = pi1039 & n14336;
  assign n14458 = pi0354 & ~n14336;
  assign po0511 = n14457 | n14458;
  assign n14460 = pi1078 & n14336;
  assign n14461 = pi0355 & ~n14336;
  assign po0512 = n14460 | n14461;
  assign n14463 = pi1075 & n14336;
  assign n14464 = pi0356 & ~n14336;
  assign po0513 = n14463 | n14464;
  assign n14466 = pi1070 & n14336;
  assign n14467 = pi0357 & ~n14336;
  assign po0514 = n14466 | n14467;
  assign n14469 = pi1065 & n14336;
  assign n14470 = pi0358 & ~n14336;
  assign po0515 = n14469 | n14470;
  assign n14472 = pi1062 & n14336;
  assign n14473 = pi0359 & ~n14336;
  assign po0516 = n14472 | n14473;
  assign n14475 = pi1036 & n14336;
  assign n14476 = pi0360 & ~n14336;
  assign po0517 = n14475 | n14476;
  assign n14478 = pi1053 & n14336;
  assign n14479 = pi0361 & ~n14336;
  assign po0518 = n14478 | n14479;
  assign n14481 = pi1064 & n14336;
  assign n14482 = pi0362 & ~n14336;
  assign po0519 = n14481 | n14482;
  assign n14484 = pi1043 & n14343;
  assign n14485 = pi0363 & ~n14343;
  assign po0520 = n14484 | n14485;
  assign n14487 = pi1056 & n14343;
  assign n14488 = pi0364 & ~n14343;
  assign po0521 = n14487 | n14488;
  assign n14490 = pi1059 & n14343;
  assign n14491 = pi0365 & ~n14343;
  assign po0522 = n14490 | n14491;
  assign n14493 = pi1063 & n14343;
  assign n14494 = pi0366 & ~n14343;
  assign po0523 = n14493 | n14494;
  assign n14496 = pi1033 & n14343;
  assign n14497 = pi0367 & ~n14343;
  assign po0524 = n14496 | n14497;
  assign n14499 = pi1061 & n14343;
  assign n14500 = pi0368 & ~n14343;
  assign po0525 = n14499 | n14500;
  assign n14502 = pi1074 & n14343;
  assign n14503 = pi0369 & ~n14343;
  assign po0526 = n14502 | n14503;
  assign n14505 = pi1049 & n14343;
  assign n14506 = pi0370 & ~n14343;
  assign po0527 = n14505 | n14506;
  assign n14508 = pi1045 & n14343;
  assign n14509 = pi0371 & ~n14343;
  assign po0528 = n14508 | n14509;
  assign n14511 = pi1042 & n14343;
  assign n14512 = pi0372 & ~n14343;
  assign po0529 = n14511 | n14512;
  assign n14514 = pi1081 & n14343;
  assign n14515 = pi0373 & ~n14343;
  assign po0530 = n14514 | n14515;
  assign n14517 = pi1029 & n14343;
  assign n14518 = pi0374 & ~n14343;
  assign po0531 = n14517 | n14518;
  assign n14520 = pi1041 & n14343;
  assign n14521 = pi0375 & ~n14343;
  assign po0532 = n14520 | n14521;
  assign n14523 = pi1073 & n14343;
  assign n14524 = pi0376 & ~n14343;
  assign po0533 = n14523 | n14524;
  assign n14526 = pi1068 & n14343;
  assign n14527 = pi0377 & ~n14343;
  assign po0534 = n14526 | n14527;
  assign n14529 = pi1057 & n14343;
  assign n14530 = pi0378 & ~n14343;
  assign po0535 = n14529 | n14530;
  assign n14532 = pi1039 & n14343;
  assign n14533 = pi0379 & ~n14343;
  assign po0536 = n14532 | n14533;
  assign n14535 = pi1078 & n14343;
  assign n14536 = pi0380 & ~n14343;
  assign po0537 = n14535 | n14536;
  assign n14538 = pi1075 & n14343;
  assign n14539 = pi0381 & ~n14343;
  assign po0538 = n14538 | n14539;
  assign n14541 = pi1070 & n14343;
  assign n14542 = pi0382 & ~n14343;
  assign po0539 = n14541 | n14542;
  assign n14544 = pi1065 & n14343;
  assign n14545 = pi0383 & ~n14343;
  assign po0540 = n14544 | n14545;
  assign n14547 = pi1062 & n14343;
  assign n14548 = pi0384 & ~n14343;
  assign po0541 = n14547 | n14548;
  assign n14550 = pi1036 & n14343;
  assign n14551 = pi0385 & ~n14343;
  assign po0542 = n14550 | n14551;
  assign n14553 = pi1053 & n14343;
  assign n14554 = pi0386 & ~n14343;
  assign po0543 = n14553 | n14554;
  assign n14556 = pi1047 & n14343;
  assign n14557 = pi0387 & ~n14343;
  assign po0544 = n14556 | n14557;
  assign n14559 = pi1031 & n14343;
  assign n14560 = pi0388 & ~n14343;
  assign po0545 = n14559 | n14560;
  assign n14562 = pi1030 & n14343;
  assign n14563 = pi0389 & ~n14343;
  assign po0546 = n14562 | n14563;
  assign n14565 = pi1043 & n14347;
  assign n14566 = pi0390 & ~n14347;
  assign po0547 = n14565 | n14566;
  assign n14568 = pi1056 & n14347;
  assign n14569 = pi0391 & ~n14347;
  assign po0548 = n14568 | n14569;
  assign n14571 = pi1033 & n14347;
  assign n14572 = pi0392 & ~n14347;
  assign po0549 = n14571 | n14572;
  assign n14574 = pi1061 & n14347;
  assign n14575 = pi0393 & ~n14347;
  assign po0550 = n14574 | n14575;
  assign n14577 = pi1074 & n14347;
  assign n14578 = pi0394 & ~n14347;
  assign po0551 = n14577 | n14578;
  assign n14580 = pi1049 & n14347;
  assign n14581 = pi0395 & ~n14347;
  assign po0552 = n14580 | n14581;
  assign n14583 = pi1045 & n14347;
  assign n14584 = pi0396 & ~n14347;
  assign po0553 = n14583 | n14584;
  assign n14586 = pi1042 & n14347;
  assign n14587 = pi0397 & ~n14347;
  assign po0554 = n14586 | n14587;
  assign n14589 = pi1081 & n14347;
  assign n14590 = pi0398 & ~n14347;
  assign po0555 = n14589 | n14590;
  assign n14592 = pi1041 & n14347;
  assign n14593 = pi0399 & ~n14347;
  assign po0556 = n14592 | n14593;
  assign n14595 = pi1029 & n14347;
  assign n14596 = pi0400 & ~n14347;
  assign po0557 = n14595 | n14596;
  assign n14598 = pi1073 & n14347;
  assign n14599 = pi0401 & ~n14347;
  assign po0558 = n14598 | n14599;
  assign n14601 = pi1072 & n14347;
  assign n14602 = pi0402 & ~n14347;
  assign po0559 = n14601 | n14602;
  assign n14604 = pi1039 & n14347;
  assign n14605 = pi0403 & ~n14347;
  assign po0560 = n14604 | n14605;
  assign n14607 = pi1078 & n14347;
  assign n14608 = pi0404 & ~n14347;
  assign po0561 = n14607 | n14608;
  assign n14610 = pi1075 & n14347;
  assign n14611 = pi0405 & ~n14347;
  assign po0562 = n14610 | n14611;
  assign n14613 = pi1070 & n14347;
  assign n14614 = pi0406 & ~n14347;
  assign po0563 = n14613 | n14614;
  assign n14616 = pi1065 & n14347;
  assign n14617 = pi0407 & ~n14347;
  assign po0564 = n14616 | n14617;
  assign n14619 = pi1062 & n14347;
  assign n14620 = pi0408 & ~n14347;
  assign po0565 = n14619 | n14620;
  assign n14622 = pi1036 & n14347;
  assign n14623 = pi0409 & ~n14347;
  assign po0566 = n14622 | n14623;
  assign n14625 = pi1053 & n14347;
  assign n14626 = pi0410 & ~n14347;
  assign po0567 = n14625 | n14626;
  assign n14628 = pi1047 & n14347;
  assign n14629 = pi0411 & ~n14347;
  assign po0568 = n14628 | n14629;
  assign n14631 = pi1031 & n14347;
  assign n14632 = pi0412 & ~n14347;
  assign po0569 = n14631 | n14632;
  assign n14634 = pi1030 & n14347;
  assign n14635 = pi0413 & ~n14347;
  assign po0570 = n14634 | n14635;
  assign n14637 = pi1043 & n14414;
  assign n14638 = pi0414 & ~n14414;
  assign po0571 = n14637 | n14638;
  assign n14640 = pi1056 & n14414;
  assign n14641 = pi0415 & ~n14414;
  assign po0572 = n14640 | n14641;
  assign n14643 = pi1063 & n14414;
  assign n14644 = pi0416 & ~n14414;
  assign po0573 = n14643 | n14644;
  assign n14646 = pi1033 & n14414;
  assign n14647 = pi0417 & ~n14414;
  assign po0574 = n14646 | n14647;
  assign n14649 = pi1061 & n14414;
  assign n14650 = pi0418 & ~n14414;
  assign po0575 = n14649 | n14650;
  assign n14652 = pi1074 & n14414;
  assign n14653 = pi0419 & ~n14414;
  assign po0576 = n14652 | n14653;
  assign n14655 = pi1049 & n14414;
  assign n14656 = pi0420 & ~n14414;
  assign po0577 = n14655 | n14656;
  assign n14658 = pi1045 & n14414;
  assign n14659 = pi0421 & ~n14414;
  assign po0578 = n14658 | n14659;
  assign n14661 = pi1042 & n14414;
  assign n14662 = pi0422 & ~n14414;
  assign po0579 = n14661 | n14662;
  assign n14664 = pi1081 & n14414;
  assign n14665 = pi0423 & ~n14414;
  assign po0580 = n14664 | n14665;
  assign n14667 = pi1041 & n14414;
  assign n14668 = pi0424 & ~n14414;
  assign po0581 = n14667 | n14668;
  assign n14670 = pi1029 & n14414;
  assign n14671 = pi0425 & ~n14414;
  assign po0582 = n14670 | n14671;
  assign n14673 = pi1073 & n14414;
  assign n14674 = pi0426 & ~n14414;
  assign po0583 = n14673 | n14674;
  assign n14676 = pi1072 & n14414;
  assign n14677 = pi0427 & ~n14414;
  assign po0584 = n14676 | n14677;
  assign n14679 = pi1039 & n14414;
  assign n14680 = pi0428 & ~n14414;
  assign po0585 = n14679 | n14680;
  assign n14682 = pi1078 & n14414;
  assign n14683 = pi0429 & ~n14414;
  assign po0586 = n14682 | n14683;
  assign n14685 = pi1070 & n14414;
  assign n14686 = pi0430 & ~n14414;
  assign po0587 = n14685 | n14686;
  assign n14688 = pi1065 & n14414;
  assign n14689 = pi0431 & ~n14414;
  assign po0588 = n14688 | n14689;
  assign n14691 = pi1062 & n14414;
  assign n14692 = pi0432 & ~n14414;
  assign po0589 = n14691 | n14692;
  assign n14694 = pi1036 & n14414;
  assign n14695 = pi0433 & ~n14414;
  assign po0590 = n14694 | n14695;
  assign n14697 = pi1053 & n14414;
  assign n14698 = pi0434 & ~n14414;
  assign po0591 = n14697 | n14698;
  assign n14700 = pi1047 & n14414;
  assign n14701 = pi0435 & ~n14414;
  assign po0592 = n14700 | n14701;
  assign n14703 = pi1031 & n14414;
  assign n14704 = pi0436 & ~n14414;
  assign po0593 = n14703 | n14704;
  assign n14706 = pi1064 & n14414;
  assign n14707 = pi0437 & ~n14414;
  assign po0594 = n14706 | n14707;
  assign n14709 = pi1030 & n14414;
  assign n14710 = pi0438 & ~n14414;
  assign po0595 = n14709 | n14710;
  assign n14712 = pi1051 & n14343;
  assign n14713 = pi0439 & ~n14343;
  assign po0596 = n14712 | n14713;
  assign n14715 = pi1037 & n14343;
  assign n14716 = pi0440 & ~n14343;
  assign po0597 = n14715 | n14716;
  assign n14718 = pi1038 & n14336;
  assign n14719 = pi0441 & ~n14336;
  assign po0598 = n14718 | n14719;
  assign n14721 = pi1052 & n14343;
  assign n14722 = pi0442 & ~n14343;
  assign po0599 = n14721 | n14722;
  assign n14724 = pi1038 & n14414;
  assign n14725 = pi0443 & ~n14414;
  assign po0600 = n14724 | n14725;
  assign n14727 = pi1066 & n14414;
  assign n14728 = pi0444 & ~n14414;
  assign po0601 = n14727 | n14728;
  assign n14730 = pi1075 & n14414;
  assign n14731 = pi0445 & ~n14414;
  assign po0602 = n14730 | n14731;
  assign n14733 = pi1080 & n14414;
  assign n14734 = pi0446 & ~n14414;
  assign po0603 = n14733 | n14734;
  assign n14736 = pi1034 & n14343;
  assign n14737 = pi0447 & ~n14343;
  assign po0604 = n14736 | n14737;
  assign n14739 = pi1068 & n14414;
  assign n14740 = pi0448 & ~n14414;
  assign po0605 = n14739 | n14740;
  assign n14742 = pi1051 & n14414;
  assign n14743 = pi0449 & ~n14414;
  assign po0606 = n14742 | n14743;
  assign n14745 = pi1030 & n14336;
  assign n14746 = pi0450 & ~n14336;
  assign po0607 = n14745 | n14746;
  assign n14748 = pi1057 & n14414;
  assign n14749 = pi0451 & ~n14414;
  assign po0608 = n14748 | n14749;
  assign n14751 = pi1047 & n14336;
  assign n14752 = pi0452 & ~n14336;
  assign po0609 = n14751 | n14752;
  assign n14754 = pi1034 & n14414;
  assign n14755 = pi0453 & ~n14414;
  assign po0610 = n14754 | n14755;
  assign n14757 = pi1037 & n14414;
  assign n14758 = pi0454 & ~n14414;
  assign po0611 = n14757 | n14758;
  assign n14760 = pi1031 & n14336;
  assign n14761 = pi0455 & ~n14336;
  assign po0612 = n14760 | n14761;
  assign n14763 = pi1038 & n14347;
  assign n14764 = pi0456 & ~n14347;
  assign po0613 = n14763 | n14764;
  assign n14766 = pi0605 & pi0821;
  assign n14767 = ~pi0804 & ~pi0810;
  assign n14768 = n14766 & n14767;
  assign n14769 = ~pi0815 & n14768;
  assign n14770 = pi0804 & ~pi0810;
  assign n14771 = pi0600 & pi0601;
  assign n14772 = pi0821 & n14771;
  assign n14773 = pi0595 & pi0597;
  assign n14774 = n14772 & n14773;
  assign n14775 = pi0594 & pi0605;
  assign n14776 = pi0596 & n14775;
  assign n14777 = n14774 & n14776;
  assign n14778 = n14770 & n14777;
  assign n14779 = pi0815 & n14778;
  assign n14780 = pi0595 & pi0596;
  assign n14781 = pi0804 & pi0810;
  assign n14782 = pi0605 & n14772;
  assign n14783 = pi0599 & n14782;
  assign n14784 = pi0594 & n14783;
  assign n14785 = pi0597 & n14784;
  assign n14786 = n14781 & n14785;
  assign n14787 = pi0815 & n14786;
  assign n14788 = n14780 & n14787;
  assign n14789 = ~pi0804 & pi0810;
  assign n14790 = n14766 & n14789;
  assign n14791 = ~pi0815 & n14790;
  assign n14792 = pi0601 & n14791;
  assign n14793 = pi0601 & pi0605;
  assign n14794 = pi0600 & n14793;
  assign n14795 = pi0594 & n14794;
  assign n14796 = pi0821 & n14781;
  assign n14797 = ~pi0815 & n14796;
  assign n14798 = n14795 & n14797;
  assign n14799 = pi0594 & pi0597;
  assign n14800 = n14766 & n14771;
  assign n14801 = n14767 & n14800;
  assign n14802 = pi0815 & n14801;
  assign n14803 = n14799 & n14802;
  assign n14804 = ~n14798 & ~n14803;
  assign n14805 = ~n14792 & n14804;
  assign n14806 = ~n14788 & n14805;
  assign n14807 = ~pi0815 & n14800;
  assign n14808 = n14770 & n14807;
  assign n14809 = n14806 & ~n14808;
  assign n14810 = pi0601 & pi0815;
  assign n14811 = pi0594 & pi0600;
  assign n14812 = n14810 & n14811;
  assign n14813 = n14789 & n14812;
  assign n14814 = n14773 & n14813;
  assign n14815 = n14766 & n14814;
  assign n14816 = n14809 & ~n14815;
  assign n14817 = ~n14779 & n14816;
  assign po0614 = n14769 | ~n14817;
  assign n14819 = pi1066 & n14336;
  assign n14820 = pi0458 & ~n14336;
  assign po0615 = n14819 | n14820;
  assign n14822 = pi1052 & n14414;
  assign n14823 = pi0459 & ~n14414;
  assign po0616 = n14822 | n14823;
  assign n14825 = pi1080 & n14336;
  assign n14826 = pi0460 & ~n14336;
  assign po0617 = n14825 | n14826;
  assign n14828 = pi1051 & n14336;
  assign n14829 = pi0461 & ~n14336;
  assign po0618 = n14828 | n14829;
  assign n14831 = pi1068 & n14336;
  assign n14832 = pi0462 & ~n14336;
  assign po0619 = n14831 | n14832;
  assign n14834 = pi1064 & n14347;
  assign n14835 = pi0463 & ~n14347;
  assign po0620 = n14834 | n14835;
  assign n14837 = pi1059 & n14414;
  assign n14838 = pi0464 & ~n14414;
  assign po0621 = n14837 | n14838;
  assign n14840 = pi0926 & n3132;
  assign n14841 = pi1151 & ~n3132;
  assign n14842 = ~n14840 & ~n14841;
  assign n14843 = ~n2439 & ~n14842;
  assign n14844 = ~pi0243 & n2440;
  assign po0622 = n14843 | n14844;
  assign n14846 = pi0943 & n3132;
  assign n14847 = pi1145 & ~n3132;
  assign n14848 = ~n14846 & ~n14847;
  assign n14849 = ~n2439 & ~n14848;
  assign n14850 = pi0275 & n2440;
  assign po0623 = n14849 | n14850;
  assign n14852 = ~pi0048 & n2967;
  assign n14853 = ~pi0040 & n2501;
  assign n14854 = n2971 & n2997;
  assign n14855 = n3000 & n14854;
  assign n14856 = n2959 & n14855;
  assign n14857 = n14853 & n14856;
  assign n14858 = n2972 & n13132;
  assign n14859 = n14857 & n14858;
  assign n14860 = n2962 & n14859;
  assign n14861 = n2502 & n14860;
  assign n14862 = n2992 & n14861;
  assign n14863 = ~pi0065 & ~pi0102;
  assign n14864 = pi0065 & pi0102;
  assign n14865 = ~n14863 & ~n14864;
  assign n14866 = n14862 & n14865;
  assign n14867 = n2980 & n2983;
  assign n14868 = n14866 & n14867;
  assign n14869 = n14852 & n14868;
  assign n14870 = n12260 & n14869;
  assign n14871 = ~pi0040 & n14870;
  assign n14872 = ~po1049 & n14871;
  assign n14873 = n12273 & n12279;
  assign n14874 = n14872 & n14873;
  assign n14875 = pi0995 & n3464;
  assign n14876 = pi0040 & po0950;
  assign n14877 = ~pi0984 & n14876;
  assign n14878 = n14875 & n14877;
  assign po0624 = n14874 | n14878;
  assign n14880 = n3465 & n6745;
  assign n14881 = ~pi0024 & n2788;
  assign n14882 = pi0468 & ~n14881;
  assign po0625 = n14880 | n14882;
  assign n14884 = pi0942 & n3132;
  assign n14885 = pi1150 & ~n3132;
  assign n14886 = ~n14884 & ~n14885;
  assign n14887 = ~n2439 & ~n14886;
  assign n14888 = ~pi0263 & n2440;
  assign po0626 = n14887 | n14888;
  assign n14890 = pi0925 & n3132;
  assign n14891 = pi1149 & ~n3132;
  assign n14892 = ~n14890 & ~n14891;
  assign n14893 = ~n2439 & ~n14892;
  assign n14894 = pi0267 & n2440;
  assign po0627 = n14893 | n14894;
  assign n14896 = pi0941 & n3132;
  assign n14897 = pi1147 & ~n3132;
  assign n14898 = ~n14896 & ~n14897;
  assign n14899 = ~n2439 & ~n14898;
  assign n14900 = pi0253 & n2440;
  assign po0628 = n14899 | n14900;
  assign n14902 = pi0923 & n3132;
  assign n14903 = pi1148 & ~n3132;
  assign n14904 = ~n14902 & ~n14903;
  assign n14905 = ~n2439 & ~n14904;
  assign n14906 = pi0254 & n2440;
  assign po0629 = n14905 | n14906;
  assign n14908 = pi0922 & n3132;
  assign n14909 = pi1146 & ~n3132;
  assign n14910 = ~n14908 & ~n14909;
  assign n14911 = ~n2439 & ~n14910;
  assign n14912 = pi0268 & n2440;
  assign po0630 = n14911 | n14912;
  assign n14914 = pi0931 & n3132;
  assign n14915 = pi1144 & ~n3132;
  assign n14916 = ~n14914 & ~n14915;
  assign n14917 = ~n2439 & ~n14916;
  assign n14918 = pi0272 & n2440;
  assign po0631 = n14917 | n14918;
  assign n14920 = pi0936 & n3132;
  assign n14921 = pi1143 & ~n3132;
  assign n14922 = ~n14920 & ~n14921;
  assign n14923 = ~n2439 & ~n14922;
  assign n14924 = pi0283 & n2440;
  assign po0632 = n14923 | n14924;
  assign n14926 = pi0071 & n7400;
  assign n14927 = ~pi0060 & ~pi0061;
  assign n14928 = n12278 & n14927;
  assign n14929 = n12260 & n14928;
  assign n14930 = n14245 & n14929;
  assign n14931 = n2987 & n4163;
  assign n14932 = n14930 & n14931;
  assign n14933 = n2959 & n12270;
  assign n14934 = n2962 & n14933;
  assign n14935 = ~pi0048 & n14934;
  assign n14936 = pi0084 & n14935;
  assign n14937 = n3003 & n14936;
  assign n14938 = n14932 & n14937;
  assign n14939 = n12271 & n14938;
  assign n14940 = n2967 & n14939;
  assign n14941 = ~pi0051 & ~pi0081;
  assign n14942 = n2973 & n12262;
  assign n14943 = n2479 & n14942;
  assign n14944 = n14941 & n14943;
  assign n14945 = ~po1049 & n14944;
  assign n14946 = ~pi0071 & n14945;
  assign n14947 = ~pi0046 & n14946;
  assign n14948 = ~pi0068 & n14947;
  assign n14949 = n14940 & n14948;
  assign po0633 = n14926 | n14949;
  assign po0635 = pi0071 & n4983;
  assign n14952 = pi0248 & n13116;
  assign n14953 = pi0481 & ~n13116;
  assign po0638 = n14952 | n14953;
  assign n14955 = pi0249 & n13196;
  assign n14956 = pi0482 & ~n13196;
  assign po0639 = n14955 | n14956;
  assign n14958 = pi0242 & n13217;
  assign n14959 = pi0483 & ~n13217;
  assign po0640 = n14958 | n14959;
  assign n14961 = pi0249 & n13217;
  assign n14962 = pi0484 & ~n13217;
  assign po0641 = n14961 | n14962;
  assign n14964 = pi0234 & n13293;
  assign n14965 = pi0485 & ~n13293;
  assign po0642 = n14964 | n14965;
  assign n14967 = pi0244 & n13293;
  assign n14968 = pi0486 & ~n13293;
  assign po0643 = n14967 | n14968;
  assign n14970 = pi0246 & n13116;
  assign n14971 = pi0487 & ~n13116;
  assign po0644 = n14970 | n14971;
  assign n14973 = pi0239 & n13116;
  assign n14974 = ~pi0488 & ~n13116;
  assign po0645 = n14973 | n14974;
  assign n14976 = pi0242 & n13293;
  assign n14977 = pi0489 & ~n13293;
  assign po0646 = n14976 | n14977;
  assign n14979 = pi0241 & n13217;
  assign n14980 = pi0490 & ~n13217;
  assign po0647 = n14979 | n14980;
  assign n14982 = pi0238 & n13217;
  assign n14983 = pi0491 & ~n13217;
  assign po0648 = n14982 | n14983;
  assign n14985 = pi0240 & n13217;
  assign n14986 = pi0492 & ~n13217;
  assign po0649 = n14985 | n14986;
  assign n14988 = pi0244 & n13217;
  assign n14989 = pi0493 & ~n13217;
  assign po0650 = n14988 | n14989;
  assign n14991 = pi0239 & n13217;
  assign n14992 = ~pi0494 & ~n13217;
  assign po0651 = n14991 | n14992;
  assign n14994 = pi0235 & n13217;
  assign n14995 = pi0495 & ~n13217;
  assign po0652 = n14994 | n14995;
  assign n14997 = pi0249 & n13211;
  assign n14998 = pi0496 & ~n13211;
  assign po0653 = n14997 | n14998;
  assign n15000 = pi0239 & n13211;
  assign n15001 = ~pi0497 & ~n13211;
  assign po0654 = n15000 | n15001;
  assign n15003 = pi0238 & n13196;
  assign n15004 = pi0498 & ~n13196;
  assign po0655 = n15003 | n15004;
  assign n15006 = pi0246 & n13211;
  assign n15007 = pi0499 & ~n13211;
  assign po0656 = n15006 | n15007;
  assign n15009 = pi0241 & n13211;
  assign n15010 = pi0500 & ~n13211;
  assign po0657 = n15009 | n15010;
  assign n15012 = pi0248 & n13211;
  assign n15013 = pi0501 & ~n13211;
  assign po0658 = n15012 | n15013;
  assign n15015 = pi0247 & n13211;
  assign n15016 = pi0502 & ~n13211;
  assign po0659 = n15015 | n15016;
  assign n15018 = pi0245 & n13211;
  assign n15019 = pi0503 & ~n13211;
  assign po0660 = n15018 | n15019;
  assign n15021 = pi0242 & n13199;
  assign n15022 = pi0504 & ~n13199;
  assign po0661 = n15021 | n15022;
  assign n15024 = pi0234 & n13211;
  assign n15025 = pi0505 & ~n13211;
  assign po0662 = n15024 | n15025;
  assign n15027 = pi0241 & n13199;
  assign n15028 = pi0506 & ~n13199;
  assign po0663 = n15027 | n15028;
  assign n15030 = pi0238 & n13199;
  assign n15031 = pi0507 & ~n13199;
  assign po0664 = n15030 | n15031;
  assign n15033 = pi0247 & n13199;
  assign n15034 = pi0508 & ~n13199;
  assign po0665 = n15033 | n15034;
  assign n15036 = pi0245 & n13199;
  assign n15037 = pi0509 & ~n13199;
  assign po0666 = n15036 | n15037;
  assign n15039 = pi0242 & n13116;
  assign n15040 = pi0510 & ~n13116;
  assign po0667 = n15039 | n15040;
  assign n15042 = pi0234 & n13116;
  assign n15043 = pi0511 & ~n13116;
  assign po0668 = n15042 | n15043;
  assign n15045 = pi0235 & n13116;
  assign n15046 = pi0512 & ~n13116;
  assign po0669 = n15045 | n15046;
  assign n15048 = pi0244 & n13116;
  assign n15049 = pi0513 & ~n13116;
  assign po0670 = n15048 | n15049;
  assign n15051 = pi0245 & n13116;
  assign n15052 = pi0514 & ~n13116;
  assign po0671 = n15051 | n15052;
  assign n15054 = pi0240 & n13116;
  assign n15055 = pi0515 & ~n13116;
  assign po0672 = n15054 | n15055;
  assign n15057 = pi0247 & n13116;
  assign n15058 = pi0516 & ~n13116;
  assign po0673 = n15057 | n15058;
  assign n15060 = pi0238 & n13116;
  assign n15061 = pi0517 & ~n13116;
  assign po0674 = n15060 | n15061;
  assign n15063 = pi0234 & n13190;
  assign n15064 = pi0518 & ~n13190;
  assign po0675 = n15063 | n15064;
  assign n15066 = pi0239 & n13190;
  assign n15067 = ~pi0519 & ~n13190;
  assign po0676 = n15066 | n15067;
  assign n15069 = pi0246 & n13190;
  assign n15070 = pi0520 & ~n13190;
  assign po0677 = n15069 | n15070;
  assign n15072 = pi0248 & n13190;
  assign n15073 = pi0521 & ~n13190;
  assign po0678 = n15072 | n15073;
  assign n15075 = pi0238 & n13190;
  assign n15076 = pi0522 & ~n13190;
  assign po0679 = n15075 | n15076;
  assign n15078 = pi0234 & n13304;
  assign n15079 = pi0523 & ~n13304;
  assign po0680 = n15078 | n15079;
  assign n15081 = pi0239 & n13304;
  assign n15082 = ~pi0524 & ~n13304;
  assign po0681 = n15081 | n15082;
  assign n15084 = pi0245 & n13304;
  assign n15085 = pi0525 & ~n13304;
  assign po0682 = n15084 | n15085;
  assign n15087 = pi0246 & n13304;
  assign n15088 = pi0526 & ~n13304;
  assign po0683 = n15087 | n15088;
  assign n15090 = pi0247 & n13304;
  assign n15091 = pi0527 & ~n13304;
  assign po0684 = n15090 | n15091;
  assign n15093 = pi0249 & n13304;
  assign n15094 = pi0528 & ~n13304;
  assign po0685 = n15093 | n15094;
  assign n15096 = pi0238 & n13304;
  assign n15097 = pi0529 & ~n13304;
  assign po0686 = n15096 | n15097;
  assign n15099 = pi0240 & n13304;
  assign n15100 = pi0530 & ~n13304;
  assign po0687 = n15099 | n15100;
  assign n15102 = pi0235 & n13196;
  assign n15103 = pi0531 & ~n13196;
  assign po0688 = n15102 | n15103;
  assign n15105 = pi0247 & n13196;
  assign n15106 = pi0532 & ~n13196;
  assign po0689 = n15105 | n15106;
  assign n15108 = pi0235 & n13199;
  assign n15109 = pi0533 & ~n13199;
  assign po0690 = n15108 | n15109;
  assign n15111 = pi0239 & n13199;
  assign n15112 = ~pi0534 & ~n13199;
  assign po0691 = n15111 | n15112;
  assign n15114 = pi0240 & n13199;
  assign n15115 = pi0535 & ~n13199;
  assign po0692 = n15114 | n15115;
  assign n15117 = pi0246 & n13199;
  assign n15118 = pi0536 & ~n13199;
  assign po0693 = n15117 | n15118;
  assign n15120 = pi0248 & n13199;
  assign n15121 = pi0537 & ~n13199;
  assign po0694 = n15120 | n15121;
  assign n15123 = pi0249 & n13199;
  assign n15124 = pi0538 & ~n13199;
  assign po0695 = n15123 | n15124;
  assign n15126 = pi0242 & n13211;
  assign n15127 = pi0539 & ~n13211;
  assign po0696 = n15126 | n15127;
  assign n15129 = pi0235 & n13211;
  assign n15130 = pi0540 & ~n13211;
  assign po0697 = n15129 | n15130;
  assign n15132 = pi0244 & n13211;
  assign n15133 = pi0541 & ~n13211;
  assign po0698 = n15132 | n15133;
  assign n15135 = pi0240 & n13211;
  assign n15136 = pi0542 & ~n13211;
  assign po0699 = n15135 | n15136;
  assign n15138 = pi0238 & n13211;
  assign n15139 = pi0543 & ~n13211;
  assign po0700 = n15138 | n15139;
  assign n15141 = pi0234 & n13217;
  assign n15142 = pi0544 & ~n13217;
  assign po0701 = n15141 | n15142;
  assign n15144 = pi0245 & n13217;
  assign n15145 = pi0545 & ~n13217;
  assign po0702 = n15144 | n15145;
  assign n15147 = pi0246 & n13217;
  assign n15148 = pi0546 & ~n13217;
  assign po0703 = n15147 | n15148;
  assign n15150 = pi0247 & n13217;
  assign n15151 = pi0547 & ~n13217;
  assign po0704 = n15150 | n15151;
  assign n15153 = pi0248 & n13217;
  assign n15154 = pi0548 & ~n13217;
  assign po0705 = n15153 | n15154;
  assign n15156 = pi0235 & n13293;
  assign n15157 = pi0549 & ~n13293;
  assign po0706 = n15156 | n15157;
  assign n15159 = pi0239 & n13293;
  assign n15160 = ~pi0550 & ~n13293;
  assign po0707 = n15159 | n15160;
  assign n15162 = pi0240 & n13293;
  assign n15163 = pi0551 & ~n13293;
  assign po0708 = n15162 | n15163;
  assign n15165 = pi0247 & n13293;
  assign n15166 = pi0552 & ~n13293;
  assign po0709 = n15165 | n15166;
  assign n15168 = pi0241 & n13293;
  assign n15169 = pi0553 & ~n13293;
  assign po0710 = n15168 | n15169;
  assign n15171 = pi0248 & n13293;
  assign n15172 = pi0554 & ~n13293;
  assign po0711 = n15171 | n15172;
  assign n15174 = pi0249 & n13293;
  assign n15175 = pi0555 & ~n13293;
  assign po0712 = n15174 | n15175;
  assign n15177 = pi0242 & n13196;
  assign n15178 = pi0556 & ~n13196;
  assign po0713 = n15177 | n15178;
  assign n15180 = pi0234 & n13199;
  assign n15181 = pi0557 & ~n13199;
  assign po0714 = n15180 | n15181;
  assign n15183 = pi0244 & n13199;
  assign n15184 = pi0558 & ~n13199;
  assign po0715 = n15183 | n15184;
  assign n15186 = pi0241 & n13116;
  assign n15187 = pi0559 & ~n13116;
  assign po0716 = n15186 | n15187;
  assign n15189 = pi0240 & n13196;
  assign n15190 = pi0560 & ~n13196;
  assign po0717 = n15189 | n15190;
  assign n15192 = pi0247 & n13190;
  assign n15193 = pi0561 & ~n13190;
  assign po0718 = n15192 | n15193;
  assign n15195 = pi0241 & n13196;
  assign n15196 = pi0562 & ~n13196;
  assign po0719 = n15195 | n15196;
  assign n15198 = pi0246 & n13293;
  assign n15199 = pi0563 & ~n13293;
  assign po0720 = n15198 | n15199;
  assign n15201 = pi0246 & n13196;
  assign n15202 = pi0564 & ~n13196;
  assign po0721 = n15201 | n15202;
  assign n15204 = pi0248 & n13196;
  assign n15205 = pi0565 & ~n13196;
  assign po0722 = n15204 | n15205;
  assign n15207 = pi0244 & n13196;
  assign n15208 = pi0566 & ~n13196;
  assign po0723 = n15207 | n15208;
  assign po1102 = pi0230 & n2721;
  assign n15211 = ~pi0567 & ~po1102;
  assign n15212 = pi1086 & n15211;
  assign n15213 = pi0665 & n12693;
  assign n15214 = pi0621 & n12641;
  assign n15215 = ~n15213 & ~n15214;
  assign n15216 = po1102 & ~n15215;
  assign n15217 = pi1085 & n15216;
  assign po0724 = n15212 | n15217;
  assign n15219 = pi0245 & n13196;
  assign n15220 = pi0568 & ~n13196;
  assign po0725 = n15219 | n15220;
  assign n15222 = pi0239 & n13196;
  assign n15223 = ~pi0569 & ~n13196;
  assign po0726 = n15222 | n15223;
  assign n15225 = pi0234 & n13196;
  assign n15226 = pi0570 & ~n13196;
  assign po0727 = n15225 | n15226;
  assign n15228 = pi0241 & n13304;
  assign n15229 = pi0571 & ~n13304;
  assign po0728 = n15228 | n15229;
  assign n15231 = pi0244 & n13304;
  assign n15232 = pi0572 & ~n13304;
  assign po0729 = n15231 | n15232;
  assign n15234 = pi0242 & n13304;
  assign n15235 = pi0573 & ~n13304;
  assign po0730 = n15234 | n15235;
  assign n15237 = pi0241 & n13190;
  assign n15238 = pi0574 & ~n13190;
  assign po0731 = n15237 | n15238;
  assign n15240 = pi0235 & n13304;
  assign n15241 = pi0575 & ~n13304;
  assign po0732 = n15240 | n15241;
  assign n15243 = pi0248 & n13304;
  assign n15244 = pi0576 & ~n13304;
  assign po0733 = n15243 | n15244;
  assign n15246 = pi0238 & n13293;
  assign n15247 = pi0577 & ~n13293;
  assign po0734 = n15246 | n15247;
  assign n15249 = pi0249 & n13190;
  assign n15250 = pi0578 & ~n13190;
  assign po0735 = n15249 | n15250;
  assign n15252 = pi0249 & n13116;
  assign n15253 = pi0579 & ~n13116;
  assign po0736 = n15252 | n15253;
  assign n15255 = pi0245 & n13293;
  assign n15256 = pi0580 & ~n13293;
  assign po0737 = n15255 | n15256;
  assign n15258 = pi0235 & n13190;
  assign n15259 = pi0581 & ~n13190;
  assign po0738 = n15258 | n15259;
  assign n15261 = pi0240 & n13190;
  assign n15262 = pi0582 & ~n13190;
  assign po0739 = n15261 | n15262;
  assign n15264 = pi0245 & n13190;
  assign n15265 = pi0584 & ~n13190;
  assign po0741 = n15264 | n15265;
  assign n15267 = pi0244 & n13190;
  assign n15268 = pi0585 & ~n13190;
  assign po0742 = n15267 | n15268;
  assign n15270 = pi0242 & n13190;
  assign n15271 = pi0586 & ~n13190;
  assign po0743 = n15270 | n15271;
  assign n15273 = ~pi0230 & pi0587;
  assign n15274 = pi0230 & n12643;
  assign po0744 = n15273 | n15274;
  assign n15276 = ~pi0123 & n2726;
  assign n15277 = pi0588 & ~n15276;
  assign n15278 = pi0591 & n15276;
  assign n15279 = ~n15277 & ~n15278;
  assign po0745 = n14384 & ~n15279;
  assign n15281 = ~pi0201 & n13114;
  assign n15282 = ~pi0202 & n13185;
  assign n15283 = ~n15281 & ~n15282;
  assign n15284 = ~pi0220 & n13213;
  assign n15285 = ~pi0203 & n13192;
  assign n15286 = ~n15284 & ~n15285;
  assign n15287 = n15283 & n15286;
  assign n15288 = n3375 & ~n15287;
  assign n15289 = ~pi0204 & n13114;
  assign n15290 = ~pi0205 & n13185;
  assign n15291 = ~n15289 & ~n15290;
  assign n15292 = ~pi0218 & n13192;
  assign n15293 = n15291 & ~n15292;
  assign n15294 = ~pi0206 & n13213;
  assign n15295 = n15293 & ~n15294;
  assign n15296 = ~n3384 & ~n15295;
  assign po0746 = n15288 | n15296;
  assign n15298 = pi0588 & n15276;
  assign n15299 = pi0590 & ~n15276;
  assign n15300 = ~n15298 & ~n15299;
  assign po0747 = ~n14384 | ~n15300;
  assign n15302 = pi0591 & ~n15276;
  assign n15303 = pi0592 & n15276;
  assign n15304 = ~n15302 & ~n15303;
  assign po0748 = n14384 & ~n15304;
  assign n15306 = pi0592 & ~n15276;
  assign n15307 = pi0590 & n15276;
  assign n15308 = ~n15306 & ~n15307;
  assign po0749 = n14384 & ~n15308;
  assign n15310 = ~pi0234 & pi0557;
  assign n15311 = pi0234 & ~pi0557;
  assign n15312 = ~n15310 & ~n15311;
  assign n15313 = ~pi0235 & pi0533;
  assign n15314 = pi0235 & ~pi0533;
  assign n15315 = ~n15313 & ~n15314;
  assign n15316 = n15312 & n15315;
  assign n15317 = ~pi0238 & pi0507;
  assign n15318 = pi0238 & ~pi0507;
  assign n15319 = ~n15317 & ~n15318;
  assign n15320 = ~pi0249 & pi0538;
  assign n15321 = pi0249 & ~pi0538;
  assign n15322 = ~n15320 & ~n15321;
  assign n15323 = n15319 & n15322;
  assign n15324 = pi0246 & pi0536;
  assign n15325 = ~pi0246 & ~pi0536;
  assign n15326 = ~n15324 & ~n15325;
  assign n15327 = n13114 & ~n15326;
  assign n15328 = ~pi0247 & pi0508;
  assign n15329 = pi0247 & ~pi0508;
  assign n15330 = ~n15328 & ~n15329;
  assign n15331 = n15327 & n15330;
  assign n15332 = ~pi0241 & pi0506;
  assign n15333 = pi0241 & ~pi0506;
  assign n15334 = ~n15332 & ~n15333;
  assign n15335 = ~pi0248 & pi0537;
  assign n15336 = pi0248 & ~pi0537;
  assign n15337 = ~n15335 & ~n15336;
  assign n15338 = n15334 & n15337;
  assign n15339 = n15331 & n15338;
  assign n15340 = n15323 & n15339;
  assign n15341 = n15316 & n15340;
  assign n15342 = ~pi0244 & pi0558;
  assign n15343 = pi0244 & ~pi0558;
  assign n15344 = ~n15342 & ~n15343;
  assign n15345 = ~pi0242 & pi0504;
  assign n15346 = pi0242 & ~pi0504;
  assign n15347 = ~n15345 & ~n15346;
  assign n15348 = ~pi0240 & pi0535;
  assign n15349 = pi0240 & ~pi0535;
  assign n15350 = ~n15348 & ~n15349;
  assign n15351 = ~pi0245 & pi0509;
  assign n15352 = pi0245 & ~pi0509;
  assign n15353 = ~n15351 & ~n15352;
  assign n15354 = n15350 & n15353;
  assign n15355 = n15347 & n15354;
  assign n15356 = n15344 & n15355;
  assign n15357 = ~pi0239 & ~pi0534;
  assign n15358 = pi0239 & pi0534;
  assign n15359 = ~n15357 & ~n15358;
  assign n15360 = n15356 & n15359;
  assign n15361 = n15341 & n15360;
  assign n15362 = ~pi0239 & ~pi0497;
  assign n15363 = pi0239 & pi0497;
  assign n15364 = ~n15362 & ~n15363;
  assign n15365 = ~pi0249 & pi0496;
  assign n15366 = pi0249 & ~pi0496;
  assign n15367 = ~n15365 & ~n15366;
  assign n15368 = ~pi0234 & pi0505;
  assign n15369 = pi0234 & ~pi0505;
  assign n15370 = ~n15368 & ~n15369;
  assign n15371 = n15367 & n15370;
  assign n15372 = ~pi0235 & pi0540;
  assign n15373 = pi0235 & ~pi0540;
  assign n15374 = ~n15372 & ~n15373;
  assign n15375 = ~pi0238 & pi0543;
  assign n15376 = pi0238 & ~pi0543;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = n15374 & n15377;
  assign n15379 = pi0246 & pi0499;
  assign n15380 = ~pi0246 & ~pi0499;
  assign n15381 = ~n15379 & ~n15380;
  assign n15382 = n13185 & ~n15381;
  assign n15383 = ~pi0248 & pi0501;
  assign n15384 = pi0248 & ~pi0501;
  assign n15385 = ~n15383 & ~n15384;
  assign n15386 = n15382 & n15385;
  assign n15387 = ~pi0247 & pi0502;
  assign n15388 = pi0247 & ~pi0502;
  assign n15389 = ~n15387 & ~n15388;
  assign n15390 = ~pi0241 & pi0500;
  assign n15391 = pi0241 & ~pi0500;
  assign n15392 = ~n15390 & ~n15391;
  assign n15393 = n15389 & n15392;
  assign n15394 = n15386 & n15393;
  assign n15395 = n15378 & n15394;
  assign n15396 = n15371 & n15395;
  assign n15397 = ~pi0245 & pi0503;
  assign n15398 = pi0245 & ~pi0503;
  assign n15399 = ~n15397 & ~n15398;
  assign n15400 = ~pi0242 & pi0539;
  assign n15401 = pi0242 & ~pi0539;
  assign n15402 = ~n15400 & ~n15401;
  assign n15403 = ~pi0240 & pi0542;
  assign n15404 = pi0240 & ~pi0542;
  assign n15405 = ~n15403 & ~n15404;
  assign n15406 = ~pi0244 & pi0541;
  assign n15407 = pi0244 & ~pi0541;
  assign n15408 = ~n15406 & ~n15407;
  assign n15409 = n15405 & n15408;
  assign n15410 = n15402 & n15409;
  assign n15411 = n15399 & n15410;
  assign n15412 = n15396 & n15411;
  assign n15413 = n15364 & n15412;
  assign n15414 = ~n15361 & ~n15413;
  assign n15415 = ~pi0249 & pi0484;
  assign n15416 = pi0249 & ~pi0484;
  assign n15417 = ~n15415 & ~n15416;
  assign n15418 = ~pi0235 & pi0495;
  assign n15419 = pi0235 & ~pi0495;
  assign n15420 = ~n15418 & ~n15419;
  assign n15421 = n15417 & n15420;
  assign n15422 = ~pi0238 & pi0491;
  assign n15423 = pi0238 & ~pi0491;
  assign n15424 = ~n15422 & ~n15423;
  assign n15425 = ~pi0234 & pi0544;
  assign n15426 = pi0234 & ~pi0544;
  assign n15427 = ~n15425 & ~n15426;
  assign n15428 = n15424 & n15427;
  assign n15429 = pi0248 & pi0548;
  assign n15430 = ~pi0248 & ~pi0548;
  assign n15431 = ~n15429 & ~n15430;
  assign n15432 = n13213 & ~n15431;
  assign n15433 = ~pi0241 & pi0490;
  assign n15434 = pi0241 & ~pi0490;
  assign n15435 = ~n15433 & ~n15434;
  assign n15436 = n15432 & n15435;
  assign n15437 = ~pi0247 & pi0547;
  assign n15438 = pi0247 & ~pi0547;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = ~pi0246 & pi0546;
  assign n15441 = pi0246 & ~pi0546;
  assign n15442 = ~n15440 & ~n15441;
  assign n15443 = n15439 & n15442;
  assign n15444 = n15436 & n15443;
  assign n15445 = n15428 & n15444;
  assign n15446 = n15421 & n15445;
  assign n15447 = ~pi0245 & pi0545;
  assign n15448 = pi0245 & ~pi0545;
  assign n15449 = ~n15447 & ~n15448;
  assign n15450 = ~pi0244 & pi0493;
  assign n15451 = pi0244 & ~pi0493;
  assign n15452 = ~n15450 & ~n15451;
  assign n15453 = ~pi0242 & pi0483;
  assign n15454 = pi0242 & ~pi0483;
  assign n15455 = ~n15453 & ~n15454;
  assign n15456 = ~pi0240 & pi0492;
  assign n15457 = pi0240 & ~pi0492;
  assign n15458 = ~n15456 & ~n15457;
  assign n15459 = n15455 & n15458;
  assign n15460 = n15452 & n15459;
  assign n15461 = n15449 & n15460;
  assign n15462 = ~pi0239 & ~pi0494;
  assign n15463 = pi0239 & pi0494;
  assign n15464 = ~n15462 & ~n15463;
  assign n15465 = n15461 & n15464;
  assign n15466 = n15446 & n15465;
  assign n15467 = ~pi0239 & ~pi0550;
  assign n15468 = pi0239 & pi0550;
  assign n15469 = ~n15467 & ~n15468;
  assign n15470 = ~pi0235 & pi0549;
  assign n15471 = pi0235 & ~pi0549;
  assign n15472 = ~n15470 & ~n15471;
  assign n15473 = ~pi0234 & pi0485;
  assign n15474 = pi0234 & ~pi0485;
  assign n15475 = ~n15473 & ~n15474;
  assign n15476 = n15472 & n15475;
  assign n15477 = ~pi0238 & pi0577;
  assign n15478 = pi0238 & ~pi0577;
  assign n15479 = ~n15477 & ~n15478;
  assign n15480 = ~pi0249 & pi0555;
  assign n15481 = pi0249 & ~pi0555;
  assign n15482 = ~n15480 & ~n15481;
  assign n15483 = n15479 & n15482;
  assign n15484 = pi0246 & pi0563;
  assign n15485 = ~pi0246 & ~pi0563;
  assign n15486 = ~n15484 & ~n15485;
  assign n15487 = n13192 & ~n15486;
  assign n15488 = ~pi0247 & pi0552;
  assign n15489 = pi0247 & ~pi0552;
  assign n15490 = ~n15488 & ~n15489;
  assign n15491 = n15487 & n15490;
  assign n15492 = ~pi0241 & pi0553;
  assign n15493 = pi0241 & ~pi0553;
  assign n15494 = ~n15492 & ~n15493;
  assign n15495 = ~pi0248 & pi0554;
  assign n15496 = pi0248 & ~pi0554;
  assign n15497 = ~n15495 & ~n15496;
  assign n15498 = n15494 & n15497;
  assign n15499 = n15491 & n15498;
  assign n15500 = n15483 & n15499;
  assign n15501 = n15476 & n15500;
  assign n15502 = ~pi0244 & pi0486;
  assign n15503 = pi0244 & ~pi0486;
  assign n15504 = ~n15502 & ~n15503;
  assign n15505 = ~pi0242 & pi0489;
  assign n15506 = pi0242 & ~pi0489;
  assign n15507 = ~n15505 & ~n15506;
  assign n15508 = ~pi0240 & pi0551;
  assign n15509 = pi0240 & ~pi0551;
  assign n15510 = ~n15508 & ~n15509;
  assign n15511 = ~pi0245 & pi0580;
  assign n15512 = pi0245 & ~pi0580;
  assign n15513 = ~n15511 & ~n15512;
  assign n15514 = n15510 & n15513;
  assign n15515 = n15507 & n15514;
  assign n15516 = n15504 & n15515;
  assign n15517 = n15501 & n15516;
  assign n15518 = n15469 & n15517;
  assign n15519 = ~n15466 & ~n15518;
  assign n15520 = n15414 & n15519;
  assign n15521 = ~n3384 & ~n15520;
  assign n15522 = ~pi0235 & pi0575;
  assign n15523 = pi0235 & ~pi0575;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = ~pi0238 & pi0529;
  assign n15526 = pi0238 & ~pi0529;
  assign n15527 = ~n15525 & ~n15526;
  assign n15528 = n15524 & n15527;
  assign n15529 = ~pi0249 & pi0528;
  assign n15530 = pi0249 & ~pi0528;
  assign n15531 = ~n15529 & ~n15530;
  assign n15532 = ~pi0234 & pi0523;
  assign n15533 = pi0234 & ~pi0523;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = n15531 & n15534;
  assign n15536 = pi0247 & pi0527;
  assign n15537 = ~pi0247 & ~pi0527;
  assign n15538 = ~n15536 & ~n15537;
  assign n15539 = n13213 & ~n15538;
  assign n15540 = ~pi0248 & pi0576;
  assign n15541 = pi0248 & ~pi0576;
  assign n15542 = ~n15540 & ~n15541;
  assign n15543 = n15539 & n15542;
  assign n15544 = ~pi0246 & pi0526;
  assign n15545 = pi0246 & ~pi0526;
  assign n15546 = ~n15544 & ~n15545;
  assign n15547 = ~pi0241 & pi0571;
  assign n15548 = pi0241 & ~pi0571;
  assign n15549 = ~n15547 & ~n15548;
  assign n15550 = n15546 & n15549;
  assign n15551 = n15543 & n15550;
  assign n15552 = n15535 & n15551;
  assign n15553 = n15528 & n15552;
  assign n15554 = ~pi0244 & pi0572;
  assign n15555 = pi0244 & ~pi0572;
  assign n15556 = ~n15554 & ~n15555;
  assign n15557 = ~pi0242 & pi0573;
  assign n15558 = pi0242 & ~pi0573;
  assign n15559 = ~n15557 & ~n15558;
  assign n15560 = ~pi0240 & pi0530;
  assign n15561 = pi0240 & ~pi0530;
  assign n15562 = ~n15560 & ~n15561;
  assign n15563 = ~pi0245 & pi0525;
  assign n15564 = pi0245 & ~pi0525;
  assign n15565 = ~n15563 & ~n15564;
  assign n15566 = n15562 & n15565;
  assign n15567 = n15559 & n15566;
  assign n15568 = n15556 & n15567;
  assign n15569 = ~pi0239 & ~pi0524;
  assign n15570 = pi0239 & pi0524;
  assign n15571 = ~n15569 & ~n15570;
  assign n15572 = n15568 & n15571;
  assign n15573 = n15553 & n15572;
  assign n15574 = ~pi0239 & ~pi0569;
  assign n15575 = pi0239 & pi0569;
  assign n15576 = ~n15574 & ~n15575;
  assign n15577 = ~pi0234 & pi0570;
  assign n15578 = pi0234 & ~pi0570;
  assign n15579 = ~n15577 & ~n15578;
  assign n15580 = ~pi0235 & pi0531;
  assign n15581 = pi0235 & ~pi0531;
  assign n15582 = ~n15580 & ~n15581;
  assign n15583 = n15579 & n15582;
  assign n15584 = ~pi0238 & pi0498;
  assign n15585 = pi0238 & ~pi0498;
  assign n15586 = ~n15584 & ~n15585;
  assign n15587 = ~pi0249 & pi0482;
  assign n15588 = pi0249 & ~pi0482;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = n15586 & n15589;
  assign n15591 = pi0246 & pi0564;
  assign n15592 = ~pi0246 & ~pi0564;
  assign n15593 = ~n15591 & ~n15592;
  assign n15594 = n13192 & ~n15593;
  assign n15595 = ~pi0247 & pi0532;
  assign n15596 = pi0247 & ~pi0532;
  assign n15597 = ~n15595 & ~n15596;
  assign n15598 = n15594 & n15597;
  assign n15599 = ~pi0248 & pi0565;
  assign n15600 = pi0248 & ~pi0565;
  assign n15601 = ~n15599 & ~n15600;
  assign n15602 = ~pi0241 & pi0562;
  assign n15603 = pi0241 & ~pi0562;
  assign n15604 = ~n15602 & ~n15603;
  assign n15605 = n15601 & n15604;
  assign n15606 = n15598 & n15605;
  assign n15607 = n15590 & n15606;
  assign n15608 = n15583 & n15607;
  assign n15609 = ~pi0244 & pi0566;
  assign n15610 = pi0244 & ~pi0566;
  assign n15611 = ~n15609 & ~n15610;
  assign n15612 = ~pi0242 & pi0556;
  assign n15613 = pi0242 & ~pi0556;
  assign n15614 = ~n15612 & ~n15613;
  assign n15615 = ~pi0240 & pi0560;
  assign n15616 = pi0240 & ~pi0560;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = ~pi0245 & pi0568;
  assign n15619 = pi0245 & ~pi0568;
  assign n15620 = ~n15618 & ~n15619;
  assign n15621 = n15617 & n15620;
  assign n15622 = n15614 & n15621;
  assign n15623 = n15611 & n15622;
  assign n15624 = n15608 & n15623;
  assign n15625 = n15576 & n15624;
  assign n15626 = ~n15573 & ~n15625;
  assign n15627 = ~pi0249 & pi0578;
  assign n15628 = pi0249 & ~pi0578;
  assign n15629 = ~n15627 & ~n15628;
  assign n15630 = ~pi0235 & pi0581;
  assign n15631 = pi0235 & ~pi0581;
  assign n15632 = ~n15630 & ~n15631;
  assign n15633 = n15629 & n15632;
  assign n15634 = ~pi0234 & pi0518;
  assign n15635 = pi0234 & ~pi0518;
  assign n15636 = ~n15634 & ~n15635;
  assign n15637 = ~pi0238 & pi0522;
  assign n15638 = pi0238 & ~pi0522;
  assign n15639 = ~n15637 & ~n15638;
  assign n15640 = n15636 & n15639;
  assign n15641 = pi0246 & pi0520;
  assign n15642 = ~pi0246 & ~pi0520;
  assign n15643 = ~n15641 & ~n15642;
  assign n15644 = n13185 & ~n15643;
  assign n15645 = ~pi0247 & pi0561;
  assign n15646 = pi0247 & ~pi0561;
  assign n15647 = ~n15645 & ~n15646;
  assign n15648 = n15644 & n15647;
  assign n15649 = ~pi0241 & pi0574;
  assign n15650 = pi0241 & ~pi0574;
  assign n15651 = ~n15649 & ~n15650;
  assign n15652 = ~pi0248 & pi0521;
  assign n15653 = pi0248 & ~pi0521;
  assign n15654 = ~n15652 & ~n15653;
  assign n15655 = n15651 & n15654;
  assign n15656 = n15648 & n15655;
  assign n15657 = n15640 & n15656;
  assign n15658 = n15633 & n15657;
  assign n15659 = ~pi0242 & pi0586;
  assign n15660 = pi0242 & ~pi0586;
  assign n15661 = ~n15659 & ~n15660;
  assign n15662 = ~pi0244 & pi0585;
  assign n15663 = pi0244 & ~pi0585;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = ~pi0245 & pi0584;
  assign n15666 = pi0245 & ~pi0584;
  assign n15667 = ~n15665 & ~n15666;
  assign n15668 = ~pi0240 & pi0582;
  assign n15669 = pi0240 & ~pi0582;
  assign n15670 = ~n15668 & ~n15669;
  assign n15671 = n15667 & n15670;
  assign n15672 = n15664 & n15671;
  assign n15673 = n15661 & n15672;
  assign n15674 = n15658 & n15673;
  assign n15675 = pi0239 & ~pi0519;
  assign n15676 = ~pi0239 & pi0519;
  assign n15677 = ~n15675 & ~n15676;
  assign n15678 = n15674 & ~n15677;
  assign n15679 = n15626 & ~n15678;
  assign n15680 = ~pi0240 & pi0515;
  assign n15681 = pi0240 & ~pi0515;
  assign n15682 = ~n15680 & ~n15681;
  assign n15683 = ~pi0244 & pi0513;
  assign n15684 = pi0244 & ~pi0513;
  assign n15685 = ~n15683 & ~n15684;
  assign n15686 = n15682 & n15685;
  assign n15687 = ~pi0245 & pi0514;
  assign n15688 = pi0245 & ~pi0514;
  assign n15689 = ~n15687 & ~n15688;
  assign n15690 = ~pi0242 & pi0510;
  assign n15691 = pi0242 & ~pi0510;
  assign n15692 = ~n15690 & ~n15691;
  assign n15693 = n15689 & n15692;
  assign n15694 = ~pi0234 & pi0511;
  assign n15695 = pi0234 & ~pi0511;
  assign n15696 = ~n15694 & ~n15695;
  assign n15697 = ~pi0249 & pi0579;
  assign n15698 = pi0249 & ~pi0579;
  assign n15699 = ~n15697 & ~n15698;
  assign n15700 = n15696 & n15699;
  assign n15701 = ~pi0247 & pi0516;
  assign n15702 = pi0247 & ~pi0516;
  assign n15703 = ~n15701 & ~n15702;
  assign n15704 = ~pi0248 & pi0481;
  assign n15705 = pi0248 & ~pi0481;
  assign n15706 = ~n15704 & ~n15705;
  assign n15707 = n15703 & n15706;
  assign n15708 = ~pi0235 & pi0512;
  assign n15709 = pi0235 & ~pi0512;
  assign n15710 = ~n15708 & ~n15709;
  assign n15711 = ~pi0238 & pi0517;
  assign n15712 = pi0238 & ~pi0517;
  assign n15713 = ~n15711 & ~n15712;
  assign n15714 = n15710 & n15713;
  assign n15715 = n15707 & n15714;
  assign n15716 = n15700 & n15715;
  assign n15717 = pi0241 & pi0559;
  assign n15718 = ~pi0241 & ~pi0559;
  assign n15719 = ~n15717 & ~n15718;
  assign n15720 = pi0246 & pi0487;
  assign n15721 = ~pi0246 & ~pi0487;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = ~n15719 & ~n15722;
  assign n15724 = n13114 & n15723;
  assign n15725 = n15716 & n15724;
  assign n15726 = pi0239 & ~pi0488;
  assign n15727 = ~pi0239 & pi0488;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = n15725 & ~n15728;
  assign n15730 = n15693 & n15729;
  assign n15731 = n15686 & n15730;
  assign n15732 = n15679 & ~n15731;
  assign n15733 = n3375 & ~n15732;
  assign po0750 = n15521 | n15733;
  assign n15735 = ~pi0594 & ~n14794;
  assign n15736 = ~n14795 & ~n15735;
  assign n15737 = ~pi0806 & n15736;
  assign n15738 = pi0594 & pi0806;
  assign n15739 = ~n15737 & ~n15738;
  assign po0751 = ~pi0332 & ~n15739;
  assign n15741 = pi0605 & n14771;
  assign n15742 = n14799 & n15741;
  assign n15743 = pi0595 & n15742;
  assign n15744 = ~pi0595 & ~n15742;
  assign n15745 = ~n15743 & ~n15744;
  assign n15746 = ~pi0806 & n15745;
  assign n15747 = pi0595 & pi0806;
  assign n15748 = ~n15746 & ~n15747;
  assign po0752 = ~pi0332 & ~n15748;
  assign n15750 = n14773 & n14811;
  assign n15751 = n14793 & n15750;
  assign n15752 = pi0596 & n15751;
  assign n15753 = ~pi0596 & ~n15751;
  assign n15754 = ~n15752 & ~n15753;
  assign n15755 = ~pi0806 & n15754;
  assign n15756 = pi0596 & pi0806;
  assign n15757 = ~n15755 & ~n15756;
  assign po0753 = ~pi0332 & ~n15757;
  assign n15759 = ~pi0597 & ~n14795;
  assign n15760 = pi0597 & n14795;
  assign n15761 = ~n15759 & ~n15760;
  assign n15762 = ~pi0806 & n15761;
  assign n15763 = pi0597 & pi0806;
  assign n15764 = ~n15762 & ~n15763;
  assign po0754 = ~pi0332 & ~n15764;
  assign po1038 = ~n2587 | ~n2981;
  assign n15767 = ~pi0882 & ~po1038;
  assign n15768 = pi0947 & n15767;
  assign n15769 = pi0598 & ~n15768;
  assign n15770 = pi0740 & pi0780;
  assign n15771 = pi0603 & n15770;
  assign n15772 = n3368 & n15771;
  assign po0755 = n15769 | n15772;
  assign n15774 = n14794 & n14799;
  assign n15775 = n14780 & n15774;
  assign n15776 = pi0599 & n15775;
  assign n15777 = ~pi0599 & ~n15775;
  assign n15778 = ~n15776 & ~n15777;
  assign n15779 = ~pi0806 & n15778;
  assign n15780 = pi0599 & pi0806;
  assign n15781 = ~n15779 & ~n15780;
  assign po0756 = ~pi0332 & ~n15781;
  assign n15783 = ~pi0600 & ~n14793;
  assign n15784 = ~n14794 & ~n15783;
  assign n15785 = ~pi0806 & n15784;
  assign n15786 = pi0600 & pi0806;
  assign n15787 = ~n15785 & ~n15786;
  assign po0757 = ~pi0332 & ~n15787;
  assign n15789 = pi0601 & pi0806;
  assign n15790 = ~pi0601 & pi0605;
  assign n15791 = pi0601 & ~pi0605;
  assign n15792 = ~n15790 & ~n15791;
  assign n15793 = ~pi0806 & ~n15792;
  assign n15794 = ~n15789 & ~n15793;
  assign po0758 = ~pi0332 & ~n15794;
  assign n15796 = ~pi0230 & pi0602;
  assign n15797 = pi0230 & n12695;
  assign po0759 = n15796 | n15797;
  assign n15799 = pi0872 & pi0966;
  assign n15800 = pi0871 & pi0966;
  assign n15801 = ~pi0980 & ~pi1055;
  assign n15802 = pi1032 & n15801;
  assign n15803 = pi0832 & n15802;
  assign n15804 = pi1054 & n15803;
  assign po0897 = pi0952 & n15804;
  assign n15806 = pi1094 & po0897;
  assign n15807 = pi0603 & ~po0897;
  assign n15808 = ~n15806 & ~n15807;
  assign n15809 = ~pi0966 & ~n15808;
  assign n15810 = ~n15800 & ~n15809;
  assign po0760 = n15799 | ~n15810;
  assign n15812 = ~pi0661 & n3377;
  assign n15813 = pi0823 & n15812;
  assign n15814 = ~pi0779 & n15813;
  assign n15815 = ~pi0299 & pi0983;
  assign n15816 = pi0907 & n15815;
  assign n15817 = ~n15813 & ~n15816;
  assign n15818 = pi0604 & n15817;
  assign po0761 = n15814 | n15818;
  assign n15820 = pi0605 & ~pi0806;
  assign n15821 = ~pi0605 & pi0806;
  assign n15822 = ~n15820 & ~n15821;
  assign po0762 = ~pi0332 & n15822;
  assign n15824 = pi1098 & po0897;
  assign n15825 = pi0606 & ~po0897;
  assign n15826 = ~n15824 & ~n15825;
  assign n15827 = ~pi0966 & ~n15826;
  assign n15828 = pi0837 & pi0966;
  assign po0763 = n15827 | n15828;
  assign n15830 = pi0607 & ~po0897;
  assign n15831 = pi1101 & po0897;
  assign n15832 = ~n15830 & ~n15831;
  assign po0764 = ~pi0966 & ~n15832;
  assign n15834 = pi0608 & ~po0897;
  assign n15835 = pi1110 & po0897;
  assign n15836 = ~n15834 & ~n15835;
  assign po0765 = ~pi0966 & ~n15836;
  assign n15838 = pi0609 & ~po0897;
  assign n15839 = pi1112 & po0897;
  assign n15840 = ~n15838 & ~n15839;
  assign po0766 = ~pi0966 & ~n15840;
  assign n15842 = pi0610 & ~po0897;
  assign n15843 = pi1107 & po0897;
  assign n15844 = ~n15842 & ~n15843;
  assign po0767 = ~pi0966 & ~n15844;
  assign n15846 = pi0611 & ~po0897;
  assign n15847 = pi1108 & po0897;
  assign n15848 = ~n15846 & ~n15847;
  assign po0768 = ~pi0966 & ~n15848;
  assign n15850 = pi0612 & ~po0897;
  assign n15851 = pi1105 & po0897;
  assign n15852 = ~n15850 & ~n15851;
  assign po0769 = ~pi0966 & ~n15852;
  assign n15854 = pi0613 & ~po0897;
  assign n15855 = pi1109 & po0897;
  assign n15856 = ~n15854 & ~n15855;
  assign po0770 = ~pi0966 & ~n15856;
  assign n15858 = pi1096 & po0897;
  assign n15859 = pi0614 & ~po0897;
  assign n15860 = ~n15858 & ~n15859;
  assign n15861 = ~pi0966 & ~n15860;
  assign po0771 = n15800 | n15861;
  assign n15863 = pi0779 & pi0797;
  assign n15864 = pi0680 & n15863;
  assign n15865 = n15812 & n15864;
  assign n15866 = pi0907 & n15767;
  assign n15867 = ~pi0615 & ~n15866;
  assign po0772 = n15865 | n15867;
  assign n15869 = pi1095 & po0897;
  assign n15870 = pi0616 & ~po0897;
  assign n15871 = ~n15869 & ~n15870;
  assign n15872 = ~pi0966 & ~n15871;
  assign po0773 = n15799 | n15872;
  assign n15874 = pi1099 & po0897;
  assign n15875 = pi0617 & ~po0897;
  assign n15876 = ~n15874 & ~n15875;
  assign n15877 = ~pi0966 & ~n15876;
  assign n15878 = pi0850 & pi0966;
  assign po0774 = n15877 | n15878;
  assign n15880 = pi0618 & ~po0897;
  assign n15881 = pi1111 & po0897;
  assign n15882 = ~n15880 & ~n15881;
  assign po0775 = ~pi0966 & ~n15882;
  assign n15884 = pi0619 & ~po0897;
  assign n15885 = pi1116 & po0897;
  assign n15886 = ~n15884 & ~n15885;
  assign po0776 = ~pi0966 & ~n15886;
  assign n15888 = pi0620 & ~po0897;
  assign n15889 = pi1106 & po0897;
  assign n15890 = ~n15888 & ~n15889;
  assign po0777 = ~pi0966 & ~n15890;
  assign n15892 = pi0621 & ~po0897;
  assign n15893 = pi1102 & po0897;
  assign n15894 = ~n15892 & ~n15893;
  assign po0778 = ~pi0966 & ~n15894;
  assign n15896 = pi0622 & ~po0897;
  assign n15897 = pi1103 & po0897;
  assign n15898 = ~n15896 & ~n15897;
  assign po0779 = ~pi0966 & ~n15898;
  assign n15900 = pi0623 & ~po0897;
  assign n15901 = pi1100 & po0897;
  assign n15902 = ~n15900 & ~n15901;
  assign po0780 = ~pi0966 & ~n15902;
  assign n15904 = pi0831 & n3368;
  assign n15905 = ~pi0780 & n15904;
  assign n15906 = pi0947 & n15815;
  assign n15907 = ~n15904 & ~n15906;
  assign n15908 = pi0624 & n15907;
  assign po0781 = n15905 | n15908;
  assign n15910 = ~pi0973 & ~pi1048;
  assign n15911 = pi1082 & n15910;
  assign n15912 = pi0832 & n15911;
  assign n15913 = pi1060 & n15912;
  assign po0954 = ~pi0953 & n15913;
  assign n15915 = pi0625 & ~po0954;
  assign n15916 = pi1110 & po0954;
  assign n15917 = ~n15915 & ~n15916;
  assign po0782 = ~pi0962 & ~n15917;
  assign n15919 = pi0626 & ~po0897;
  assign n15920 = pi1115 & po0897;
  assign n15921 = ~n15919 & ~n15920;
  assign po0783 = ~pi0966 & ~n15921;
  assign n15923 = pi0627 & ~po0954;
  assign n15924 = pi1111 & po0954;
  assign n15925 = ~n15923 & ~n15924;
  assign po0784 = ~pi0962 & ~n15925;
  assign n15927 = pi0628 & ~po0954;
  assign n15928 = pi1113 & po0954;
  assign n15929 = ~n15927 & ~n15928;
  assign po0785 = ~pi0962 & ~n15929;
  assign n15931 = pi0629 & ~po0897;
  assign n15932 = pi1113 & po0897;
  assign n15933 = ~n15931 & ~n15932;
  assign po0786 = ~pi0966 & ~n15933;
  assign n15935 = pi0630 & ~po0897;
  assign n15936 = pi1114 & po0897;
  assign n15937 = ~n15935 & ~n15936;
  assign po0787 = ~pi0966 & ~n15937;
  assign n15939 = ~pi0631 & ~po0954;
  assign n15940 = pi1107 & po0954;
  assign n15941 = ~n15939 & ~n15940;
  assign po0788 = ~pi0962 & ~n15941;
  assign n15943 = ~pi0632 & ~po0954;
  assign n15944 = pi1109 & po0954;
  assign n15945 = ~n15943 & ~n15944;
  assign po0789 = ~pi0962 & ~n15945;
  assign n15947 = pi0633 & ~po0897;
  assign n15948 = pi1104 & po0897;
  assign n15949 = ~n15947 & ~n15948;
  assign po0790 = ~pi0966 & ~n15949;
  assign n15951 = pi0634 & ~po0954;
  assign n15952 = pi1104 & po0954;
  assign n15953 = ~n15951 & ~n15952;
  assign po0791 = ~pi0962 & ~n15953;
  assign n15955 = ~pi0635 & ~po0954;
  assign n15956 = pi1106 & po0954;
  assign n15957 = ~n15955 & ~n15956;
  assign po0792 = ~pi0962 & ~n15957;
  assign n15959 = pi0636 & ~po0897;
  assign n15960 = pi1121 & po0897;
  assign n15961 = ~n15959 & ~n15960;
  assign po0793 = ~pi0966 & ~n15961;
  assign n15963 = pi0637 & ~po0954;
  assign n15964 = pi1099 & po0954;
  assign n15965 = ~n15963 & ~n15964;
  assign po0794 = ~pi0962 & ~n15965;
  assign n15967 = pi0638 & ~po0954;
  assign n15968 = pi1101 & po0954;
  assign n15969 = ~n15967 & ~n15968;
  assign po0795 = ~pi0962 & ~n15969;
  assign n15971 = pi0639 & ~po0954;
  assign n15972 = pi1103 & po0954;
  assign n15973 = ~n15971 & ~n15972;
  assign po0796 = ~pi0962 & ~n15973;
  assign n15975 = pi0640 & ~po0897;
  assign n15976 = pi1122 & po0897;
  assign n15977 = ~n15975 & ~n15976;
  assign po0797 = ~pi0966 & ~n15977;
  assign n15979 = pi0641 & ~po0954;
  assign n15980 = pi1115 & po0954;
  assign n15981 = ~n15979 & ~n15980;
  assign po0798 = ~pi0962 & ~n15981;
  assign n15983 = pi0642 & ~po0897;
  assign n15984 = pi1097 & po0897;
  assign n15985 = ~n15983 & ~n15984;
  assign po0799 = ~pi0966 & ~n15985;
  assign n15987 = pi0643 & ~po0954;
  assign n15988 = pi1098 & po0954;
  assign n15989 = ~n15987 & ~n15988;
  assign po0800 = ~pi0962 & ~n15989;
  assign n15991 = pi0644 & ~po0897;
  assign n15992 = pi1117 & po0897;
  assign n15993 = ~n15991 & ~n15992;
  assign po0801 = ~pi0966 & ~n15993;
  assign n15995 = pi0645 & ~po0897;
  assign n15996 = pi1119 & po0897;
  assign n15997 = ~n15995 & ~n15996;
  assign po0802 = ~pi0966 & ~n15997;
  assign n15999 = ~pi0646 & ~po0954;
  assign n16000 = pi1108 & po0954;
  assign n16001 = ~n15999 & ~n16000;
  assign po0803 = ~pi0962 & ~n16001;
  assign n16003 = pi0647 & ~po0954;
  assign n16004 = pi1114 & po0954;
  assign n16005 = ~n16003 & ~n16004;
  assign po0804 = ~pi0962 & ~n16005;
  assign n16007 = pi0648 & ~po0954;
  assign n16008 = pi1116 & po0954;
  assign n16009 = ~n16007 & ~n16008;
  assign po0805 = ~pi0962 & ~n16009;
  assign n16011 = ~pi0649 & ~po0954;
  assign n16012 = pi1120 & po0954;
  assign n16013 = ~n16011 & ~n16012;
  assign po0806 = ~pi0962 & ~n16013;
  assign n16015 = ~pi0650 & ~po0954;
  assign n16016 = pi1121 & po0954;
  assign n16017 = ~n16015 & ~n16016;
  assign po0807 = ~pi0962 & ~n16017;
  assign n16019 = pi0651 & ~po0897;
  assign n16020 = pi1124 & po0897;
  assign n16021 = ~n16019 & ~n16020;
  assign po0808 = ~pi0966 & ~n16021;
  assign n16023 = pi0652 & ~po0897;
  assign n16024 = pi1125 & po0897;
  assign n16025 = ~n16023 & ~n16024;
  assign po0809 = ~pi0966 & ~n16025;
  assign n16027 = pi0653 & ~po0897;
  assign n16028 = pi1123 & po0897;
  assign n16029 = ~n16027 & ~n16028;
  assign po0810 = ~pi0966 & ~n16029;
  assign n16031 = ~pi0654 & ~po0954;
  assign n16032 = pi1124 & po0954;
  assign n16033 = ~n16031 & ~n16032;
  assign po0811 = ~pi0962 & ~n16033;
  assign n16035 = ~pi0655 & ~po0954;
  assign n16036 = pi1118 & po0954;
  assign n16037 = ~n16035 & ~n16036;
  assign po0812 = ~pi0962 & ~n16037;
  assign n16039 = pi0656 & ~po0897;
  assign n16040 = pi1120 & po0897;
  assign n16041 = ~n16039 & ~n16040;
  assign po0813 = ~pi0966 & ~n16041;
  assign n16043 = ~pi0657 & ~po0954;
  assign n16044 = pi1125 & po0954;
  assign n16045 = ~n16043 & ~n16044;
  assign po0814 = ~pi0962 & ~n16045;
  assign n16047 = pi0658 & ~po0897;
  assign n16048 = pi1118 & po0897;
  assign n16049 = ~n16047 & ~n16048;
  assign po0815 = ~pi0966 & ~n16049;
  assign n16051 = pi0278 & pi0279;
  assign n16052 = pi0266 & n16051;
  assign n16053 = ~pi0280 & n16052;
  assign n16054 = ~pi0269 & n16053;
  assign n16055 = ~pi0282 & n16054;
  assign n16056 = ~pi0281 & n16055;
  assign n16057 = ~pi0264 & ~pi0277;
  assign n16058 = n16056 & n16057;
  assign n16059 = ~pi0265 & n16058;
  assign n16060 = ~pi0270 & n16059;
  assign n16061 = ~pi0274 & ~n16060;
  assign n16062 = pi0274 & n16060;
  assign po0816 = n16061 | n16062;
  assign n16064 = pi0660 & ~po0954;
  assign n16065 = pi1112 & po0954;
  assign n16066 = ~n16064 & ~n16065;
  assign po0817 = ~pi0962 & ~n16066;
  assign n16068 = pi0661 & ~po0954;
  assign n16069 = pi1095 & po0954;
  assign n16070 = ~n16068 & ~n16069;
  assign po0818 = ~pi0962 & ~n16070;
  assign n16072 = pi0662 & ~po0954;
  assign n16073 = pi1096 & po0954;
  assign n16074 = ~n16072 & ~n16073;
  assign po0819 = ~pi0962 & ~n16074;
  assign n16076 = ~pi1131 & ~pi1132;
  assign n16077 = ~pi1128 & n16076;
  assign n16078 = pi1129 & ~pi1130;
  assign n16079 = n16077 & n16078;
  assign n16080 = pi0784 & n16079;
  assign n16081 = ~pi1129 & ~pi1130;
  assign n16082 = n16076 & n16081;
  assign n16083 = ~pi1128 & n16082;
  assign n16084 = pi0815 & n16083;
  assign n16085 = ~n16080 & ~n16084;
  assign n16086 = pi1128 & n16082;
  assign n16087 = pi0855 & n16086;
  assign n16088 = ~pi1129 & n16076;
  assign n16089 = pi1130 & n16088;
  assign n16090 = pi1128 & n16089;
  assign n16091 = pi0766 & n16090;
  assign n16092 = ~pi1128 & n16089;
  assign n16093 = pi0633 & n16092;
  assign n16094 = ~n16091 & ~n16093;
  assign n16095 = pi1129 & n16076;
  assign n16096 = pi1130 & n16095;
  assign n16097 = pi1128 & n16096;
  assign n16098 = pi0700 & n16097;
  assign n16099 = ~pi1128 & n16096;
  assign n16100 = pi0634 & n16099;
  assign n16101 = ~n16098 & ~n16100;
  assign n16102 = n16094 & n16101;
  assign n16103 = ~n16087 & n16102;
  assign n16104 = n16085 & n16103;
  assign n16105 = ~n3539 & ~n16104;
  assign n16106 = ~pi0223 & ~pi0224;
  assign n16107 = pi0222 & n16106;
  assign n16108 = ~pi0222 & ~pi0223;
  assign n16109 = ~pi0224 & n16108;
  assign n16110 = ~n16107 & ~n16109;
  assign n16111 = ~n3667 & ~n16110;
  assign n16112 = ~n13785 & ~n13788;
  assign n16113 = pi0257 & ~n16112;
  assign n16114 = pi0199 & pi1059;
  assign n16115 = ~n16113 & ~n16114;
  assign n16116 = n16110 & ~n16115;
  assign n16117 = ~n16111 & ~n16116;
  assign n16118 = n3539 & ~n16117;
  assign po0820 = n16105 | n16118;
  assign n16120 = pi0785 & n16079;
  assign n16121 = pi0872 & n16086;
  assign n16122 = ~n16120 & ~n16121;
  assign n16123 = pi0811 & n16083;
  assign n16124 = pi0772 & n16090;
  assign n16125 = pi0614 & n16092;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = pi0727 & n16097;
  assign n16128 = pi0662 & n16099;
  assign n16129 = ~n16127 & ~n16128;
  assign n16130 = n16126 & n16129;
  assign n16131 = ~n16123 & n16130;
  assign n16132 = n16122 & n16131;
  assign n16133 = ~n3539 & ~n16132;
  assign n16134 = ~n3806 & ~n16110;
  assign n16135 = pi0292 & ~n16112;
  assign n16136 = pi0199 & pi1078;
  assign n16137 = ~n16135 & ~n16136;
  assign n16138 = n16110 & ~n16137;
  assign n16139 = ~n16134 & ~n16138;
  assign n16140 = n3539 & ~n16139;
  assign po0821 = n16133 | n16140;
  assign n16142 = pi0665 & ~po0954;
  assign n16143 = pi1102 & po0954;
  assign n16144 = ~n16142 & ~n16143;
  assign po0822 = ~pi0962 & ~n16144;
  assign n16146 = pi0790 & n16079;
  assign n16147 = ~pi0799 & n16083;
  assign n16148 = ~n16146 & ~n16147;
  assign n16149 = pi0873 & n16086;
  assign n16150 = pi0764 & n16090;
  assign n16151 = pi0607 & n16092;
  assign n16152 = ~n16150 & ~n16151;
  assign n16153 = pi0691 & n16097;
  assign n16154 = pi0638 & n16099;
  assign n16155 = ~n16153 & ~n16154;
  assign n16156 = n16152 & n16155;
  assign n16157 = ~n16149 & n16156;
  assign n16158 = n16148 & n16157;
  assign n16159 = ~n3539 & ~n16158;
  assign n16160 = ~n3789 & ~n16110;
  assign n16161 = pi0297 & ~n16112;
  assign n16162 = pi0199 & pi1038;
  assign n16163 = ~n16161 & ~n16162;
  assign n16164 = n16110 & ~n16163;
  assign n16165 = ~n16160 & ~n16164;
  assign n16166 = n3539 & ~n16165;
  assign po0823 = n16159 | n16166;
  assign n16168 = pi0763 & n16090;
  assign n16169 = pi0642 & n16092;
  assign n16170 = ~n16168 & ~n16169;
  assign n16171 = pi0699 & n16097;
  assign n16172 = pi0681 & n16099;
  assign n16173 = ~n16171 & ~n16172;
  assign n16174 = pi0792 & n16079;
  assign n16175 = pi0871 & n16086;
  assign n16176 = ~n16174 & ~n16175;
  assign n16177 = ~pi0809 & n16083;
  assign n16178 = n16176 & ~n16177;
  assign n16179 = n16173 & n16178;
  assign n16180 = n16170 & n16179;
  assign n16181 = ~n3539 & ~n16180;
  assign n16182 = ~n3826 & ~n16110;
  assign n16183 = pi0294 & ~n16112;
  assign n16184 = pi0199 & pi1066;
  assign n16185 = ~n16183 & ~n16184;
  assign n16186 = n16110 & ~n16185;
  assign n16187 = ~n16182 & ~n16186;
  assign n16188 = n3539 & ~n16187;
  assign po0824 = n16181 | n16188;
  assign n16190 = pi0778 & n16079;
  assign n16191 = pi0981 & n16083;
  assign n16192 = ~n16190 & ~n16191;
  assign n16193 = pi0837 & n16086;
  assign n16194 = pi0759 & n16090;
  assign n16195 = pi0603 & n16092;
  assign n16196 = ~n16194 & ~n16195;
  assign n16197 = pi0696 & n16097;
  assign n16198 = pi0680 & n16099;
  assign n16199 = ~n16197 & ~n16198;
  assign n16200 = n16196 & n16199;
  assign n16201 = ~n16193 & n16200;
  assign n16202 = n16192 & n16201;
  assign n16203 = ~n3539 & ~n16202;
  assign n16204 = ~n3796 & ~n16110;
  assign n16205 = pi0291 & ~n16112;
  assign n16206 = pi0199 & pi1043;
  assign n16207 = ~n16205 & ~n16206;
  assign n16208 = n16110 & ~n16207;
  assign n16209 = ~n16204 & ~n16208;
  assign n16210 = n3539 & ~n16209;
  assign po0825 = n16203 | n16210;
  assign n16212 = ~pi0669 & ~po0954;
  assign n16213 = pi1119 & po0954;
  assign n16214 = ~n16212 & ~n16213;
  assign po0826 = ~pi0962 & ~n16214;
  assign n16216 = pi0612 & n16092;
  assign n16217 = pi0852 & n16086;
  assign n16218 = ~n16216 & ~n16217;
  assign n16219 = ~pi0723 & n16097;
  assign n16220 = ~pi0695 & n16099;
  assign n16221 = ~n16219 & ~n16220;
  assign n16222 = ~pi0745 & n16090;
  assign n16223 = n16221 & ~n16222;
  assign n16224 = n16218 & n16223;
  assign n16225 = ~n3539 & ~n16224;
  assign n16226 = ~n3613 & ~n16110;
  assign n16227 = pi0258 & ~n16112;
  assign n16228 = pi0199 & pi1056;
  assign n16229 = ~n16227 & ~n16228;
  assign n16230 = n16110 & ~n16229;
  assign n16231 = ~n16226 & ~n16230;
  assign n16232 = n3539 & ~n16231;
  assign po0827 = n16225 | n16232;
  assign n16234 = pi0611 & n16092;
  assign n16235 = pi0865 & n16086;
  assign n16236 = ~n16234 & ~n16235;
  assign n16237 = ~pi0724 & n16097;
  assign n16238 = ~pi0646 & n16099;
  assign n16239 = ~n16237 & ~n16238;
  assign n16240 = ~pi0741 & n16090;
  assign n16241 = n16239 & ~n16240;
  assign n16242 = n16236 & n16241;
  assign n16243 = ~n3539 & ~n16242;
  assign n16244 = ~n3637 & ~n16110;
  assign n16245 = pi0261 & ~n16112;
  assign n16246 = pi0199 & pi1034;
  assign n16247 = ~n16245 & ~n16246;
  assign n16248 = n16110 & ~n16247;
  assign n16249 = ~n16244 & ~n16248;
  assign n16250 = n3539 & ~n16249;
  assign po0828 = n16243 | n16250;
  assign n16252 = pi0736 & n16097;
  assign n16253 = pi0661 & n16099;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = pi0758 & n16090;
  assign n16256 = pi0616 & n16092;
  assign n16257 = ~n16255 & ~n16256;
  assign n16258 = pi0781 & n16079;
  assign n16259 = pi0850 & n16086;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = pi0808 & n16083;
  assign n16262 = n16260 & ~n16261;
  assign n16263 = n16257 & n16262;
  assign n16264 = n16254 & n16263;
  assign n16265 = ~n3539 & ~n16264;
  assign n16266 = ~n3843 & ~n16110;
  assign n16267 = pi0290 & ~n16112;
  assign n16268 = pi0199 & pi1042;
  assign n16269 = ~n16267 & ~n16268;
  assign n16270 = n16110 & ~n16269;
  assign n16271 = ~n16266 & ~n16270;
  assign n16272 = n3539 & ~n16271;
  assign po0829 = n16265 | n16272;
  assign n16274 = pi0749 & n16090;
  assign n16275 = pi0617 & n16092;
  assign n16276 = ~n16274 & ~n16275;
  assign n16277 = pi0706 & n16097;
  assign n16278 = pi0637 & n16099;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = pi0788 & n16079;
  assign n16281 = pi0866 & n16086;
  assign n16282 = ~n16280 & ~n16281;
  assign n16283 = ~pi0814 & n16083;
  assign n16284 = n16282 & ~n16283;
  assign n16285 = n16279 & n16284;
  assign n16286 = n16276 & n16285;
  assign n16287 = ~n3539 & ~n16286;
  assign n16288 = ~n3833 & ~n16110;
  assign n16289 = pi0295 & ~n16112;
  assign n16290 = pi0199 & pi1047;
  assign n16291 = ~n16289 & ~n16290;
  assign n16292 = n16110 & ~n16291;
  assign n16293 = ~n16288 & ~n16292;
  assign n16294 = n3539 & ~n16293;
  assign po0830 = n16287 | n16294;
  assign n16296 = pi0735 & n16097;
  assign n16297 = pi0639 & n16099;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = pi0743 & n16090;
  assign n16300 = pi0622 & n16092;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = pi0783 & n16079;
  assign n16303 = pi0859 & n16086;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = pi0804 & n16083;
  assign n16306 = n16304 & ~n16305;
  assign n16307 = n16301 & n16306;
  assign n16308 = n16298 & n16307;
  assign n16309 = ~n3539 & ~n16308;
  assign n16310 = ~n3630 & ~n16110;
  assign n16311 = pi0256 & ~n16112;
  assign n16312 = pi0199 & pi1064;
  assign n16313 = ~n16311 & ~n16312;
  assign n16314 = n16110 & ~n16313;
  assign n16315 = ~n16310 & ~n16314;
  assign n16316 = n3539 & ~n16315;
  assign po0831 = n16309 | n16316;
  assign n16318 = pi0730 & n16097;
  assign n16319 = pi0710 & n16099;
  assign n16320 = ~n16318 & ~n16319;
  assign n16321 = pi0748 & n16090;
  assign n16322 = pi0623 & n16092;
  assign n16323 = ~n16321 & ~n16322;
  assign n16324 = pi0789 & n16079;
  assign n16325 = pi0876 & n16086;
  assign n16326 = ~n16324 & ~n16325;
  assign n16327 = ~pi0803 & n16083;
  assign n16328 = n16326 & ~n16327;
  assign n16329 = n16323 & n16328;
  assign n16330 = n16320 & n16329;
  assign n16331 = ~n3539 & ~n16330;
  assign n16332 = ~n3850 & ~n16110;
  assign n16333 = pi0296 & ~n16112;
  assign n16334 = pi0199 & pi1031;
  assign n16335 = ~n16333 & ~n16334;
  assign n16336 = n16110 & ~n16335;
  assign n16337 = ~n16332 & ~n16336;
  assign n16338 = n3539 & ~n16337;
  assign po0832 = n16331 | n16338;
  assign n16340 = pi0729 & n16097;
  assign n16341 = pi0643 & n16099;
  assign n16342 = ~n16340 & ~n16341;
  assign n16343 = pi0746 & n16090;
  assign n16344 = pi0606 & n16092;
  assign n16345 = ~n16343 & ~n16344;
  assign n16346 = pi0787 & n16079;
  assign n16347 = pi0881 & n16086;
  assign n16348 = ~n16346 & ~n16347;
  assign n16349 = ~pi0812 & n16083;
  assign n16350 = n16348 & ~n16349;
  assign n16351 = n16345 & n16350;
  assign n16352 = n16342 & n16351;
  assign n16353 = ~n3539 & ~n16352;
  assign n16354 = ~n3813 & ~n16110;
  assign n16355 = pi0293 & ~n16112;
  assign n16356 = pi0199 & pi1053;
  assign n16357 = ~n16355 & ~n16356;
  assign n16358 = n16110 & ~n16357;
  assign n16359 = ~n16354 & ~n16358;
  assign n16360 = n3539 & ~n16359;
  assign po0833 = n16353 | n16360;
  assign n16362 = pi0620 & n16092;
  assign n16363 = pi0870 & n16086;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = ~pi0704 & n16097;
  assign n16366 = ~pi0635 & n16099;
  assign n16367 = ~n16365 & ~n16366;
  assign n16368 = ~pi0742 & n16090;
  assign n16369 = n16367 & ~n16368;
  assign n16370 = n16364 & n16369;
  assign n16371 = ~n3539 & ~n16370;
  assign n16372 = ~n3674 & ~n16110;
  assign n16373 = pi0259 & ~n16112;
  assign n16374 = pi0199 & pi1063;
  assign n16375 = ~n16373 & ~n16374;
  assign n16376 = n16110 & ~n16375;
  assign n16377 = ~n16372 & ~n16376;
  assign n16378 = n3539 & ~n16377;
  assign po0834 = n16371 | n16378;
  assign n16380 = pi0613 & n16092;
  assign n16381 = pi0856 & n16086;
  assign n16382 = ~n16380 & ~n16381;
  assign n16383 = ~pi0688 & n16097;
  assign n16384 = ~pi0632 & n16099;
  assign n16385 = ~n16383 & ~n16384;
  assign n16386 = ~pi0760 & n16090;
  assign n16387 = n16385 & ~n16386;
  assign n16388 = n16382 & n16387;
  assign n16389 = ~n3539 & ~n16388;
  assign n16390 = ~n3650 & ~n16110;
  assign n16391 = pi0260 & ~n16112;
  assign n16392 = pi0199 & pi1061;
  assign n16393 = ~n16391 & ~n16392;
  assign n16394 = n16110 & ~n16393;
  assign n16395 = ~n16390 & ~n16394;
  assign n16396 = n3539 & ~n16395;
  assign po0835 = n16389 | n16396;
  assign n16398 = pi0791 & n16079;
  assign n16399 = pi0810 & n16083;
  assign n16400 = ~n16398 & ~n16399;
  assign n16401 = pi0874 & n16086;
  assign n16402 = pi0739 & n16090;
  assign n16403 = pi0621 & n16092;
  assign n16404 = ~n16402 & ~n16403;
  assign n16405 = pi0690 & n16097;
  assign n16406 = pi0665 & n16099;
  assign n16407 = ~n16405 & ~n16406;
  assign n16408 = n16404 & n16407;
  assign n16409 = ~n16401 & n16408;
  assign n16410 = n16400 & n16409;
  assign n16411 = ~n3539 & ~n16410;
  assign n16412 = ~n3657 & ~n16110;
  assign n16413 = pi0255 & ~n16112;
  assign n16414 = pi0199 & pi1030;
  assign n16415 = ~n16413 & ~n16414;
  assign n16416 = n16110 & ~n16415;
  assign n16417 = ~n16412 & ~n16416;
  assign n16418 = n3539 & ~n16417;
  assign po0836 = n16411 | n16418;
  assign n16420 = pi0680 & ~po0954;
  assign n16421 = pi1094 & po0954;
  assign n16422 = ~n16420 & ~n16421;
  assign po0837 = ~pi0962 & ~n16422;
  assign n16424 = pi0681 & ~po0954;
  assign n16425 = pi1097 & po0954;
  assign n16426 = ~n16424 & ~n16425;
  assign po0838 = ~pi0962 & ~n16426;
  assign n16428 = pi0610 & n16092;
  assign n16429 = pi0848 & n16086;
  assign n16430 = ~n16428 & ~n16429;
  assign n16431 = ~pi0686 & n16097;
  assign n16432 = ~pi0631 & n16099;
  assign n16433 = ~n16431 & ~n16432;
  assign n16434 = ~pi0757 & n16090;
  assign n16435 = n16433 & ~n16434;
  assign n16436 = n16430 & n16435;
  assign n16437 = ~n3539 & ~n16436;
  assign n16438 = ~n3620 & ~n16110;
  assign n16439 = pi0251 & ~n16112;
  assign n16440 = pi0199 & pi1033;
  assign n16441 = ~n16439 & ~n16440;
  assign n16442 = n16110 & ~n16441;
  assign n16443 = ~n16438 & ~n16442;
  assign n16444 = n3539 & ~n16443;
  assign po0839 = n16437 | n16444;
  assign po0980 = pi0953 & n15913;
  assign n16447 = ~pi0684 & ~po0980;
  assign n16448 = pi1124 & po0980;
  assign n16449 = ~n16447 & ~n16448;
  assign po0841 = ~pi0962 & ~n16449;
  assign n16451 = ~pi0728 & n16097;
  assign n16452 = ~pi0657 & n16099;
  assign n16453 = ~n16451 & ~n16452;
  assign n16454 = ~pi0744 & n16090;
  assign n16455 = pi0652 & n16092;
  assign n16456 = pi0860 & n16086;
  assign n16457 = ~n16455 & ~n16456;
  assign n16458 = pi0813 & n16083;
  assign n16459 = n16457 & ~n16458;
  assign n16460 = ~n16454 & n16459;
  assign n16461 = n16453 & n16460;
  assign n16462 = ~n3539 & ~n16461;
  assign n16463 = pi1038 & n13785;
  assign n16464 = pi1061 & n13788;
  assign n16465 = pi0199 & pi1070;
  assign n16466 = ~n16464 & ~n16465;
  assign n16467 = ~n16463 & n16466;
  assign n16468 = n16110 & ~n16467;
  assign n16469 = ~n3738 & ~n16110;
  assign n16470 = ~n16468 & ~n16469;
  assign n16471 = n3539 & ~n16470;
  assign po0842 = n16462 | n16471;
  assign n16473 = ~pi0686 & ~po0980;
  assign n16474 = pi1107 & po0980;
  assign n16475 = ~n16473 & ~n16474;
  assign po0843 = ~pi0962 & ~n16475;
  assign n16477 = pi0687 & ~po0980;
  assign n16478 = pi1121 & po0980;
  assign n16479 = ~n16477 & ~n16478;
  assign po0844 = ~pi0962 & ~n16479;
  assign n16481 = ~pi0688 & ~po0980;
  assign n16482 = pi1109 & po0980;
  assign n16483 = ~n16481 & ~n16482;
  assign po0845 = ~pi0962 & ~n16483;
  assign n16485 = pi0658 & n16092;
  assign n16486 = pi0798 & n16083;
  assign n16487 = ~n16485 & ~n16486;
  assign n16488 = pi0843 & n16086;
  assign n16489 = pi0703 & n16097;
  assign n16490 = ~pi0655 & n16099;
  assign n16491 = ~n16489 & ~n16490;
  assign n16492 = ~pi0752 & n16090;
  assign n16493 = n16491 & ~n16492;
  assign n16494 = ~n16488 & n16493;
  assign n16495 = n16487 & n16494;
  assign n16496 = ~n3539 & ~n16495;
  assign n16497 = pi1030 & n13788;
  assign n16498 = pi1043 & n13785;
  assign n16499 = pi0199 & pi1073;
  assign n16500 = ~n16498 & ~n16499;
  assign n16501 = ~n16497 & n16500;
  assign n16502 = n16110 & ~n16501;
  assign n16503 = ~n3745 & ~n16110;
  assign n16504 = ~n16502 & ~n16503;
  assign n16505 = n3539 & ~n16504;
  assign po0846 = n16496 | n16505;
  assign n16507 = pi0690 & ~po0980;
  assign n16508 = pi1102 & po0980;
  assign n16509 = ~n16507 & ~n16508;
  assign po0847 = ~pi0962 & ~n16509;
  assign n16511 = pi0691 & ~po0980;
  assign n16512 = pi1101 & po0980;
  assign n16513 = ~n16511 & ~n16512;
  assign po0848 = ~pi0962 & ~n16513;
  assign n16515 = pi0656 & n16092;
  assign n16516 = pi0801 & n16083;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = pi0844 & n16086;
  assign n16519 = pi0726 & n16097;
  assign n16520 = ~pi0649 & n16099;
  assign n16521 = ~n16519 & ~n16520;
  assign n16522 = ~pi0770 & n16090;
  assign n16523 = n16521 & ~n16522;
  assign n16524 = ~n16518 & n16523;
  assign n16525 = n16517 & n16524;
  assign n16526 = ~n3539 & ~n16525;
  assign n16527 = pi1078 & n13785;
  assign n16528 = pi1059 & n13788;
  assign n16529 = pi0199 & pi1072;
  assign n16530 = ~n16528 & ~n16529;
  assign n16531 = ~n16527 & n16530;
  assign n16532 = n16110 & ~n16531;
  assign n16533 = ~n3755 & ~n16110;
  assign n16534 = ~n16532 & ~n16533;
  assign n16535 = n3539 & ~n16534;
  assign po0849 = n16526 | n16535;
  assign n16537 = ~pi0693 & ~po0954;
  assign n16538 = pi1123 & po0954;
  assign n16539 = ~n16537 & ~n16538;
  assign po0850 = ~pi0962 & ~n16539;
  assign n16541 = ~pi0694 & ~po0980;
  assign n16542 = pi1122 & po0980;
  assign n16543 = ~n16541 & ~n16542;
  assign po0851 = ~pi0962 & ~n16543;
  assign n16545 = ~pi0695 & ~po0954;
  assign n16546 = pi1105 & po0954;
  assign n16547 = ~n16545 & ~n16546;
  assign po0852 = ~pi0962 & ~n16547;
  assign n16549 = pi0696 & ~po0980;
  assign n16550 = pi1094 & po0980;
  assign n16551 = ~n16549 & ~n16550;
  assign po0853 = ~pi0962 & ~n16551;
  assign n16553 = ~pi0697 & ~po0980;
  assign n16554 = pi1123 & po0980;
  assign n16555 = ~n16553 & ~n16554;
  assign po0854 = ~pi0962 & ~n16555;
  assign n16557 = ~pi0698 & ~po0980;
  assign n16558 = pi1110 & po0980;
  assign n16559 = ~n16557 & ~n16558;
  assign po0855 = ~pi0962 & ~n16559;
  assign n16561 = pi0699 & ~po0980;
  assign n16562 = pi1097 & po0980;
  assign n16563 = ~n16561 & ~n16562;
  assign po0856 = ~pi0962 & ~n16563;
  assign n16565 = pi0700 & ~po0980;
  assign n16566 = pi1104 & po0980;
  assign n16567 = ~n16565 & ~n16566;
  assign po0857 = ~pi0962 & ~n16567;
  assign n16569 = ~pi0701 & ~po0980;
  assign n16570 = pi1117 & po0980;
  assign n16571 = ~n16569 & ~n16570;
  assign po0858 = ~pi0962 & ~n16571;
  assign n16573 = ~pi0702 & ~po0980;
  assign n16574 = pi1111 & po0980;
  assign n16575 = ~n16573 & ~n16574;
  assign po0859 = ~pi0962 & ~n16575;
  assign n16577 = pi0703 & ~po0980;
  assign n16578 = pi1118 & po0980;
  assign n16579 = ~n16577 & ~n16578;
  assign po0860 = ~pi0962 & ~n16579;
  assign n16581 = ~pi0704 & ~po0980;
  assign n16582 = pi1106 & po0980;
  assign n16583 = ~n16581 & ~n16582;
  assign po0861 = ~pi0962 & ~n16583;
  assign n16585 = pi0705 & ~po0980;
  assign n16586 = pi1119 & po0980;
  assign n16587 = ~n16585 & ~n16586;
  assign po0862 = ~pi0962 & ~n16587;
  assign n16589 = pi0706 & ~po0980;
  assign n16590 = pi1099 & po0980;
  assign n16591 = ~n16589 & ~n16590;
  assign po0863 = ~pi0962 & ~n16591;
  assign n16593 = pi0618 & n16092;
  assign n16594 = pi0847 & n16086;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = ~pi0702 & n16097;
  assign n16597 = pi0627 & n16099;
  assign n16598 = ~n16596 & ~n16597;
  assign n16599 = ~pi0753 & n16090;
  assign n16600 = n16598 & ~n16599;
  assign n16601 = n16595 & n16600;
  assign n16602 = ~n3539 & ~n16601;
  assign n16603 = pi1042 & n13788;
  assign n16604 = pi0304 & n13785;
  assign n16605 = pi0199 & pi1049;
  assign n16606 = ~n16604 & ~n16605;
  assign n16607 = ~n16603 & n16606;
  assign n16608 = n16110 & ~n16607;
  assign n16609 = ~n3894 & ~n16110;
  assign n16610 = ~n16608 & ~n16609;
  assign n16611 = n3539 & ~n16610;
  assign po0864 = n16602 | n16611;
  assign n16613 = pi0609 & n16092;
  assign n16614 = pi0857 & n16086;
  assign n16615 = ~n16613 & ~n16614;
  assign n16616 = ~pi0709 & n16097;
  assign n16617 = pi0660 & n16099;
  assign n16618 = ~n16616 & ~n16617;
  assign n16619 = ~pi0754 & n16090;
  assign n16620 = n16618 & ~n16619;
  assign n16621 = n16615 & n16620;
  assign n16622 = ~n3539 & ~n16621;
  assign n16623 = pi1078 & n13788;
  assign n16624 = pi0305 & n13785;
  assign n16625 = pi0199 & pi1052;
  assign n16626 = ~n16624 & ~n16625;
  assign n16627 = ~n16623 & n16626;
  assign n16628 = n16110 & ~n16627;
  assign n16629 = ~n3931 & ~n16110;
  assign n16630 = ~n16628 & ~n16629;
  assign n16631 = n3539 & ~n16630;
  assign po0865 = n16622 | n16631;
  assign n16633 = ~pi0709 & ~po0980;
  assign n16634 = pi1112 & po0980;
  assign n16635 = ~n16633 & ~n16634;
  assign po0866 = ~pi0962 & ~n16635;
  assign n16637 = pi0710 & ~po0954;
  assign n16638 = pi1100 & po0954;
  assign n16639 = ~n16637 & ~n16638;
  assign po0867 = ~pi0962 & ~n16639;
  assign n16641 = pi0630 & n16092;
  assign n16642 = pi0858 & n16086;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = ~pi0725 & n16097;
  assign n16645 = pi0647 & n16099;
  assign n16646 = ~n16644 & ~n16645;
  assign n16647 = ~pi0755 & n16090;
  assign n16648 = n16646 & ~n16647;
  assign n16649 = n16643 & n16648;
  assign n16650 = ~n3539 & ~n16649;
  assign n16651 = pi1053 & n13788;
  assign n16652 = pi0306 & n13785;
  assign n16653 = pi0199 & pi1081;
  assign n16654 = ~n16652 & ~n16653;
  assign n16655 = ~n16651 & n16654;
  assign n16656 = n16110 & ~n16655;
  assign n16657 = ~n3938 & ~n16110;
  assign n16658 = ~n16656 & ~n16657;
  assign n16659 = n3539 & ~n16658;
  assign po0868 = n16650 | n16659;
  assign n16661 = pi0644 & n16092;
  assign n16662 = pi0842 & n16086;
  assign n16663 = ~n16661 & ~n16662;
  assign n16664 = ~pi0701 & n16097;
  assign n16665 = pi0715 & n16099;
  assign n16666 = ~n16664 & ~n16665;
  assign n16667 = ~pi0751 & n16090;
  assign n16668 = n16666 & ~n16667;
  assign n16669 = n16663 & n16668;
  assign n16670 = ~n3539 & ~n16669;
  assign n16671 = pi1038 & n13788;
  assign n16672 = pi0298 & n13785;
  assign n16673 = pi0199 & pi1029;
  assign n16674 = ~n16672 & ~n16673;
  assign n16675 = ~n16671 & n16674;
  assign n16676 = n16110 & ~n16675;
  assign n16677 = ~n3914 & ~n16110;
  assign n16678 = ~n16676 & ~n16677;
  assign n16679 = n3539 & ~n16678;
  assign po0869 = n16670 | n16679;
  assign n16681 = pi0629 & n16092;
  assign n16682 = pi0854 & n16086;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = ~pi0734 & n16097;
  assign n16685 = pi0628 & n16099;
  assign n16686 = ~n16684 & ~n16685;
  assign n16687 = ~pi0756 & n16090;
  assign n16688 = n16686 & ~n16687;
  assign n16689 = n16683 & n16688;
  assign n16690 = ~n3539 & ~n16689;
  assign n16691 = pi1066 & n13788;
  assign n16692 = pi0309 & n13785;
  assign n16693 = pi0199 & pi1045;
  assign n16694 = ~n16692 & ~n16693;
  assign n16695 = ~n16691 & n16694;
  assign n16696 = n16110 & ~n16695;
  assign n16697 = ~n3877 & ~n16110;
  assign n16698 = ~n16696 & ~n16697;
  assign n16699 = n3539 & ~n16698;
  assign po0870 = n16690 | n16699;
  assign n16701 = pi0653 & n16092;
  assign n16702 = pi0816 & n16083;
  assign n16703 = ~n16701 & ~n16702;
  assign n16704 = pi0867 & n16086;
  assign n16705 = ~pi0697 & n16097;
  assign n16706 = ~pi0693 & n16099;
  assign n16707 = ~n16705 & ~n16706;
  assign n16708 = ~pi0762 & n16090;
  assign n16709 = n16707 & ~n16708;
  assign n16710 = ~n16704 & n16709;
  assign n16711 = n16703 & n16710;
  assign n16712 = ~n3539 & ~n16711;
  assign n16713 = pi1047 & n13785;
  assign n16714 = pi1033 & n13788;
  assign n16715 = pi0199 & pi1051;
  assign n16716 = ~n16714 & ~n16715;
  assign n16717 = ~n16713 & n16716;
  assign n16718 = n16110 & ~n16717;
  assign n16719 = ~n3718 & ~n16110;
  assign n16720 = ~n16718 & ~n16719;
  assign n16721 = n3539 & ~n16720;
  assign po0871 = n16712 | n16721;
  assign n16723 = pi0715 & ~po0954;
  assign n16724 = pi1117 & po0954;
  assign n16725 = ~n16723 & ~n16724;
  assign po0872 = ~pi0962 & ~n16725;
  assign n16727 = pi0626 & n16092;
  assign n16728 = pi0845 & n16086;
  assign n16729 = ~n16727 & ~n16728;
  assign n16730 = ~pi0738 & n16097;
  assign n16731 = pi0641 & n16099;
  assign n16732 = ~n16730 & ~n16731;
  assign n16733 = ~pi0761 & n16090;
  assign n16734 = n16732 & ~n16733;
  assign n16735 = n16729 & n16734;
  assign n16736 = ~n3539 & ~n16735;
  assign n16737 = pi1047 & n13788;
  assign n16738 = pi0307 & n13785;
  assign n16739 = pi0199 & pi1037;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = ~n16737 & n16740;
  assign n16742 = n16110 & ~n16741;
  assign n16743 = ~n3884 & ~n16110;
  assign n16744 = ~n16742 & ~n16743;
  assign n16745 = n3539 & ~n16744;
  assign po0873 = n16736 | n16745;
  assign n16747 = pi0645 & n16092;
  assign n16748 = pi0800 & n16083;
  assign n16749 = ~n16747 & ~n16748;
  assign n16750 = pi0839 & n16086;
  assign n16751 = pi0705 & n16097;
  assign n16752 = ~pi0669 & n16099;
  assign n16753 = ~n16751 & ~n16752;
  assign n16754 = ~pi0768 & n16090;
  assign n16755 = n16753 & ~n16754;
  assign n16756 = ~n16750 & n16755;
  assign n16757 = n16749 & n16756;
  assign n16758 = ~n3539 & ~n16757;
  assign n16759 = pi1064 & n13788;
  assign n16760 = pi1042 & n13785;
  assign n16761 = pi0199 & pi1068;
  assign n16762 = ~n16760 & ~n16761;
  assign n16763 = ~n16759 & n16762;
  assign n16764 = n16110 & ~n16763;
  assign n16765 = ~n3701 & ~n16110;
  assign n16766 = ~n16764 & ~n16765;
  assign n16767 = n3539 & ~n16766;
  assign po0874 = n16758 | n16767;
  assign n16769 = pi0608 & n16092;
  assign n16770 = pi0853 & n16086;
  assign n16771 = ~n16769 & ~n16770;
  assign n16772 = ~pi0698 & n16097;
  assign n16773 = pi0625 & n16099;
  assign n16774 = ~n16772 & ~n16773;
  assign n16775 = ~pi0767 & n16090;
  assign n16776 = n16774 & ~n16775;
  assign n16777 = n16771 & n16776;
  assign n16778 = ~n3539 & ~n16777;
  assign n16779 = pi1043 & n13788;
  assign n16780 = pi0303 & n13785;
  assign n16781 = pi0199 & pi1074;
  assign n16782 = ~n16780 & ~n16781;
  assign n16783 = ~n16779 & n16782;
  assign n16784 = n16110 & ~n16783;
  assign n16785 = ~n3921 & ~n16110;
  assign n16786 = ~n16784 & ~n16785;
  assign n16787 = n3539 & ~n16786;
  assign po0875 = n16778 | n16787;
  assign n16789 = pi0636 & n16092;
  assign n16790 = pi0807 & n16083;
  assign n16791 = ~n16789 & ~n16790;
  assign n16792 = pi0868 & n16086;
  assign n16793 = pi0687 & n16097;
  assign n16794 = ~pi0650 & n16099;
  assign n16795 = ~n16793 & ~n16794;
  assign n16796 = ~pi0774 & n16090;
  assign n16797 = n16795 & ~n16796;
  assign n16798 = ~n16792 & n16797;
  assign n16799 = n16791 & n16798;
  assign n16800 = ~n3539 & ~n16799;
  assign n16801 = pi1066 & n13785;
  assign n16802 = pi1056 & n13788;
  assign n16803 = pi0199 & pi1057;
  assign n16804 = ~n16802 & ~n16803;
  assign n16805 = ~n16801 & n16804;
  assign n16806 = n16110 & ~n16805;
  assign n16807 = ~n3725 & ~n16110;
  assign n16808 = ~n16806 & ~n16807;
  assign n16809 = n3539 & ~n16808;
  assign po0876 = n16800 | n16809;
  assign n16811 = pi0651 & n16092;
  assign n16812 = pi0794 & n16083;
  assign n16813 = ~n16811 & ~n16812;
  assign n16814 = pi0880 & n16086;
  assign n16815 = ~pi0684 & n16097;
  assign n16816 = ~pi0654 & n16099;
  assign n16817 = ~n16815 & ~n16816;
  assign n16818 = ~pi0750 & n16090;
  assign n16819 = n16817 & ~n16818;
  assign n16820 = ~n16814 & n16819;
  assign n16821 = n16813 & n16820;
  assign n16822 = ~n3539 & ~n16821;
  assign n16823 = pi1031 & n13785;
  assign n16824 = pi1034 & n13788;
  assign n16825 = pi0199 & pi1075;
  assign n16826 = ~n16824 & ~n16825;
  assign n16827 = ~n16823 & n16826;
  assign n16828 = n16110 & ~n16827;
  assign n16829 = ~n3708 & ~n16110;
  assign n16830 = ~n16828 & ~n16829;
  assign n16831 = n3539 & ~n16830;
  assign po0877 = n16822 | n16831;
  assign n16833 = pi0765 & pi0771;
  assign n16834 = pi0773 & n16833;
  assign n16835 = pi0731 & pi0775;
  assign n16836 = n16834 & n16835;
  assign n16837 = pi0769 & n16836;
  assign n16838 = pi0747 & n16837;
  assign n16839 = pi0721 & n16838;
  assign n16840 = ~pi0721 & ~n16838;
  assign n16841 = ~n16839 & ~n16840;
  assign n16842 = ~pi0945 & n16841;
  assign n16843 = pi0721 & pi0945;
  assign n16844 = ~n16842 & ~n16843;
  assign n16845 = ~pi0773 & pi0801;
  assign n16846 = pi0773 & ~pi0801;
  assign n16847 = ~n16845 & ~n16846;
  assign n16848 = ~pi0771 & pi0800;
  assign n16849 = pi0771 & ~pi0800;
  assign n16850 = ~n16848 & ~n16849;
  assign n16851 = n16847 & n16850;
  assign n16852 = pi0721 & pi0813;
  assign n16853 = ~pi0721 & ~pi0813;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = ~pi0747 & pi0807;
  assign n16856 = pi0747 & ~pi0807;
  assign n16857 = ~n16855 & ~n16856;
  assign n16858 = pi0765 & ~pi0798;
  assign n16859 = ~pi0765 & pi0798;
  assign n16860 = ~n16858 & ~n16859;
  assign n16861 = n16857 & n16860;
  assign n16862 = ~n16854 & n16861;
  assign n16863 = n16851 & n16862;
  assign n16864 = ~pi0769 & pi0794;
  assign n16865 = pi0769 & ~pi0794;
  assign n16866 = ~n16864 & ~n16865;
  assign n16867 = ~pi0775 & pi0816;
  assign n16868 = pi0775 & ~pi0816;
  assign n16869 = ~n16867 & ~n16868;
  assign n16870 = ~pi0731 & pi0795;
  assign n16871 = pi0731 & ~pi0795;
  assign n16872 = ~n16870 & ~n16871;
  assign n16873 = n16869 & n16872;
  assign n16874 = n16866 & n16873;
  assign po0978 = n16863 & n16874;
  assign n16876 = ~pi0795 & ~pi0816;
  assign n16877 = ~pi0794 & ~pi0813;
  assign n16878 = n16876 & n16877;
  assign n16879 = ~pi0798 & ~pi0800;
  assign n16880 = ~pi0801 & ~pi0807;
  assign n16881 = n16879 & n16880;
  assign n16882 = n16878 & n16881;
  assign po0963 = po0978 & ~n16882;
  assign po0878 = ~n16844 & ~po0963;
  assign n16885 = pi0640 & n16092;
  assign n16886 = pi0795 & n16083;
  assign n16887 = ~n16885 & ~n16886;
  assign n16888 = pi0851 & n16086;
  assign n16889 = ~pi0694 & n16097;
  assign n16890 = ~pi0732 & n16099;
  assign n16891 = ~n16889 & ~n16890;
  assign n16892 = ~pi0776 & n16090;
  assign n16893 = n16891 & ~n16892;
  assign n16894 = ~n16888 & n16893;
  assign n16895 = n16887 & n16894;
  assign n16896 = ~n3539 & ~n16895;
  assign n16897 = pi1053 & n13785;
  assign n16898 = pi1063 & n13788;
  assign n16899 = pi0199 & pi1039;
  assign n16900 = ~n16898 & ~n16899;
  assign n16901 = ~n16897 & n16900;
  assign n16902 = n16110 & ~n16901;
  assign n16903 = ~n3762 & ~n16110;
  assign n16904 = ~n16902 & ~n16903;
  assign n16905 = n3539 & ~n16904;
  assign po0879 = n16896 | n16905;
  assign n16907 = ~pi0723 & ~po0980;
  assign n16908 = pi1105 & po0980;
  assign n16909 = ~n16907 & ~n16908;
  assign po0880 = ~pi0962 & ~n16909;
  assign n16911 = ~pi0724 & ~po0980;
  assign n16912 = pi1108 & po0980;
  assign n16913 = ~n16911 & ~n16912;
  assign po0881 = ~pi0962 & ~n16913;
  assign n16915 = ~pi0725 & ~po0980;
  assign n16916 = pi1114 & po0980;
  assign n16917 = ~n16915 & ~n16916;
  assign po0882 = ~pi0962 & ~n16917;
  assign n16919 = pi0726 & ~po0980;
  assign n16920 = pi1120 & po0980;
  assign n16921 = ~n16919 & ~n16920;
  assign po0883 = ~pi0962 & ~n16921;
  assign n16923 = pi0727 & ~po0980;
  assign n16924 = pi1096 & po0980;
  assign n16925 = ~n16923 & ~n16924;
  assign po0884 = ~pi0962 & ~n16925;
  assign n16927 = ~pi0728 & ~po0980;
  assign n16928 = pi1125 & po0980;
  assign n16929 = ~n16927 & ~n16928;
  assign po0885 = ~pi0962 & ~n16929;
  assign n16931 = pi0729 & ~po0980;
  assign n16932 = pi1098 & po0980;
  assign n16933 = ~n16931 & ~n16932;
  assign po0886 = ~pi0962 & ~n16933;
  assign n16935 = pi0730 & ~po0980;
  assign n16936 = pi1100 & po0980;
  assign n16937 = ~n16935 & ~n16936;
  assign po0887 = ~pi0962 & ~n16937;
  assign n16939 = pi0747 & n16834;
  assign n16940 = pi0731 & n16939;
  assign n16941 = ~pi0731 & ~n16939;
  assign n16942 = ~n16940 & ~n16941;
  assign n16943 = ~pi0945 & n16942;
  assign n16944 = pi0731 & pi0945;
  assign n16945 = ~n16943 & ~n16944;
  assign po0888 = ~po0963 & ~n16945;
  assign n16947 = ~pi0732 & ~po0954;
  assign n16948 = pi1122 & po0954;
  assign n16949 = ~n16947 & ~n16948;
  assign po0889 = ~pi0962 & ~n16949;
  assign n16951 = pi0619 & n16092;
  assign n16952 = pi0838 & n16086;
  assign n16953 = ~n16951 & ~n16952;
  assign n16954 = ~pi0737 & n16097;
  assign n16955 = pi0648 & n16099;
  assign n16956 = ~n16954 & ~n16955;
  assign n16957 = ~pi0777 & n16090;
  assign n16958 = n16956 & ~n16957;
  assign n16959 = n16953 & n16958;
  assign n16960 = ~n3539 & ~n16959;
  assign n16961 = pi1031 & n13788;
  assign n16962 = pi0308 & n13785;
  assign n16963 = pi0199 & pi1041;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = ~n16961 & n16964;
  assign n16966 = n16110 & ~n16965;
  assign n16967 = ~n3901 & ~n16110;
  assign n16968 = ~n16966 & ~n16967;
  assign n16969 = n3539 & ~n16968;
  assign po0890 = n16960 | n16969;
  assign n16971 = ~pi0734 & ~po0980;
  assign n16972 = pi1113 & po0980;
  assign n16973 = ~n16971 & ~n16972;
  assign po0891 = ~pi0962 & ~n16973;
  assign n16975 = pi0735 & ~po0980;
  assign n16976 = pi1103 & po0980;
  assign n16977 = ~n16975 & ~n16976;
  assign po0892 = ~pi0962 & ~n16977;
  assign n16979 = pi0736 & ~po0980;
  assign n16980 = pi1095 & po0980;
  assign n16981 = ~n16979 & ~n16980;
  assign po0893 = ~pi0962 & ~n16981;
  assign n16983 = ~pi0737 & ~po0980;
  assign n16984 = pi1116 & po0980;
  assign n16985 = ~n16983 & ~n16984;
  assign po0894 = ~pi0962 & ~n16985;
  assign n16987 = ~pi0738 & ~po0980;
  assign n16988 = pi1115 & po0980;
  assign n16989 = ~n16987 & ~n16988;
  assign po0895 = ~pi0962 & ~n16989;
  assign po0988 = ~pi0952 & n15804;
  assign n16992 = pi0739 & ~po0988;
  assign n16993 = pi1102 & po0988;
  assign n16994 = ~n16992 & ~n16993;
  assign po0896 = pi0966 | ~n16994;
  assign n16996 = ~pi0741 & ~po0988;
  assign n16997 = pi1108 & po0988;
  assign n16998 = ~n16996 & ~n16997;
  assign po0898 = pi0966 | ~n16998;
  assign n17000 = ~pi0742 & ~po0988;
  assign n17001 = pi1106 & po0988;
  assign n17002 = ~n17000 & ~n17001;
  assign po0899 = pi0966 | ~n17002;
  assign n17004 = pi0743 & ~po0988;
  assign n17005 = pi1103 & po0988;
  assign n17006 = ~n17004 & ~n17005;
  assign po0900 = pi0966 | ~n17006;
  assign n17008 = ~pi0744 & ~po0988;
  assign n17009 = pi1125 & po0988;
  assign n17010 = ~n17008 & ~n17009;
  assign po0901 = pi0966 | ~n17010;
  assign n17012 = ~pi0745 & ~po0988;
  assign n17013 = pi1105 & po0988;
  assign n17014 = ~n17012 & ~n17013;
  assign po0902 = pi0966 | ~n17014;
  assign n17016 = pi0746 & ~po0988;
  assign n17017 = pi1098 & po0988;
  assign n17018 = ~n17016 & ~n17017;
  assign po0903 = pi0966 | ~n17018;
  assign n17020 = ~pi0747 & ~n16834;
  assign n17021 = ~n16939 & ~n17020;
  assign n17022 = ~pi0945 & n17021;
  assign n17023 = pi0747 & pi0945;
  assign n17024 = ~n17022 & ~n17023;
  assign po0904 = ~po0963 & ~n17024;
  assign n17026 = pi0748 & ~po0988;
  assign n17027 = pi1100 & po0988;
  assign n17028 = ~n17026 & ~n17027;
  assign po0905 = pi0966 | ~n17028;
  assign n17030 = pi0749 & ~po0988;
  assign n17031 = pi1099 & po0988;
  assign n17032 = ~n17030 & ~n17031;
  assign po0906 = pi0966 | ~n17032;
  assign n17034 = ~pi0750 & ~po0988;
  assign n17035 = pi1124 & po0988;
  assign n17036 = ~n17034 & ~n17035;
  assign po0907 = pi0966 | ~n17036;
  assign n17038 = ~pi0751 & ~po0988;
  assign n17039 = pi1117 & po0988;
  assign n17040 = ~n17038 & ~n17039;
  assign po0908 = pi0966 | ~n17040;
  assign n17042 = ~pi0752 & ~po0988;
  assign n17043 = pi1118 & po0988;
  assign n17044 = ~n17042 & ~n17043;
  assign po0909 = pi0966 | ~n17044;
  assign n17046 = ~pi0753 & ~po0988;
  assign n17047 = pi1111 & po0988;
  assign n17048 = ~n17046 & ~n17047;
  assign po0910 = pi0966 | ~n17048;
  assign n17050 = ~pi0754 & ~po0988;
  assign n17051 = pi1112 & po0988;
  assign n17052 = ~n17050 & ~n17051;
  assign po0911 = pi0966 | ~n17052;
  assign n17054 = ~pi0755 & ~po0988;
  assign n17055 = pi1114 & po0988;
  assign n17056 = ~n17054 & ~n17055;
  assign po0912 = pi0966 | ~n17056;
  assign n17058 = ~pi0756 & ~po0988;
  assign n17059 = pi1113 & po0988;
  assign n17060 = ~n17058 & ~n17059;
  assign po0913 = pi0966 | ~n17060;
  assign n17062 = ~pi0757 & ~po0988;
  assign n17063 = pi1107 & po0988;
  assign n17064 = ~n17062 & ~n17063;
  assign po0914 = pi0966 | ~n17064;
  assign n17066 = pi0758 & ~po0988;
  assign n17067 = pi1095 & po0988;
  assign n17068 = ~n17066 & ~n17067;
  assign po0915 = pi0966 | ~n17068;
  assign n17070 = pi0759 & ~po0988;
  assign n17071 = pi1094 & po0988;
  assign n17072 = ~n17070 & ~n17071;
  assign po0916 = pi0966 | ~n17072;
  assign n17074 = ~pi0760 & ~po0988;
  assign n17075 = pi1109 & po0988;
  assign n17076 = ~n17074 & ~n17075;
  assign po0917 = pi0966 | ~n17076;
  assign n17078 = ~pi0761 & ~po0988;
  assign n17079 = pi1115 & po0988;
  assign n17080 = ~n17078 & ~n17079;
  assign po0918 = pi0966 | ~n17080;
  assign n17082 = ~pi0762 & ~po0988;
  assign n17083 = pi1123 & po0988;
  assign n17084 = ~n17082 & ~n17083;
  assign po0919 = pi0966 | ~n17084;
  assign n17086 = pi0763 & ~po0988;
  assign n17087 = pi1097 & po0988;
  assign n17088 = ~n17086 & ~n17087;
  assign po0920 = pi0966 | ~n17088;
  assign n17090 = pi0764 & ~po0988;
  assign n17091 = pi1101 & po0988;
  assign n17092 = ~n17090 & ~n17091;
  assign po0921 = pi0966 | ~n17092;
  assign n17094 = pi0765 & ~pi0945;
  assign n17095 = ~pi0765 & pi0945;
  assign n17096 = ~n17094 & ~n17095;
  assign po0922 = ~po0963 & n17096;
  assign n17098 = pi0766 & ~po0988;
  assign n17099 = pi1104 & po0988;
  assign n17100 = ~n17098 & ~n17099;
  assign po0923 = pi0966 | ~n17100;
  assign n17102 = ~pi0767 & ~po0988;
  assign n17103 = pi1110 & po0988;
  assign n17104 = ~n17102 & ~n17103;
  assign po0924 = pi0966 | ~n17104;
  assign n17106 = ~pi0768 & ~po0988;
  assign n17107 = pi1119 & po0988;
  assign n17108 = ~n17106 & ~n17107;
  assign po0925 = pi0966 | ~n17108;
  assign n17110 = pi0747 & pi0773;
  assign n17111 = n16833 & n17110;
  assign n17112 = n16835 & n17111;
  assign n17113 = pi0769 & n17112;
  assign n17114 = ~pi0769 & ~n17112;
  assign n17115 = ~n17113 & ~n17114;
  assign n17116 = ~pi0945 & n17115;
  assign n17117 = pi0769 & pi0945;
  assign n17118 = ~n17116 & ~n17117;
  assign po0926 = ~po0963 & ~n17118;
  assign n17120 = ~pi0770 & ~po0988;
  assign n17121 = pi1120 & po0988;
  assign n17122 = ~n17120 & ~n17121;
  assign po0927 = pi0966 | ~n17122;
  assign n17124 = pi0771 & pi0945;
  assign n17125 = ~pi0765 & pi0771;
  assign n17126 = pi0765 & ~pi0771;
  assign n17127 = ~n17125 & ~n17126;
  assign n17128 = ~pi0945 & ~n17127;
  assign n17129 = ~n17124 & ~n17128;
  assign po0928 = ~po0963 & ~n17129;
  assign n17131 = pi0772 & ~po0988;
  assign n17132 = pi1096 & po0988;
  assign n17133 = ~n17131 & ~n17132;
  assign po0929 = pi0966 | ~n17133;
  assign n17135 = ~pi0773 & ~n16833;
  assign n17136 = ~n16834 & ~n17135;
  assign n17137 = ~pi0945 & n17136;
  assign n17138 = pi0773 & pi0945;
  assign n17139 = ~n17137 & ~n17138;
  assign po0930 = ~po0963 & ~n17139;
  assign n17141 = ~pi0774 & ~po0988;
  assign n17142 = pi1121 & po0988;
  assign n17143 = ~n17141 & ~n17142;
  assign po0931 = pi0966 | ~n17143;
  assign n17145 = pi0771 & n17110;
  assign n17146 = pi0731 & n17145;
  assign n17147 = pi0765 & n17146;
  assign n17148 = pi0775 & n17147;
  assign n17149 = ~pi0775 & ~n17147;
  assign n17150 = ~n17148 & ~n17149;
  assign n17151 = ~pi0945 & n17150;
  assign n17152 = pi0775 & pi0945;
  assign n17153 = ~n17151 & ~n17152;
  assign po0932 = ~po0963 & ~n17153;
  assign n17155 = ~pi0776 & ~po0988;
  assign n17156 = pi1122 & po0988;
  assign n17157 = ~n17155 & ~n17156;
  assign po0933 = pi0966 | ~n17157;
  assign n17159 = ~pi0777 & ~po0988;
  assign n17160 = pi1116 & po0988;
  assign n17161 = ~n17159 & ~n17160;
  assign po0934 = pi0966 | ~n17161;
  assign n17163 = pi0956 & pi1079;
  assign n17164 = pi0832 & n17163;
  assign n17165 = ~pi1040 & ~pi1077;
  assign n17166 = n17164 & n17165;
  assign n17167 = ~pi0968 & n17166;
  assign n17168 = pi1094 & n17167;
  assign n17169 = pi0778 & ~n17167;
  assign po0935 = n17168 | n17169;
  assign po0936 = ~pi0779 | n15866;
  assign po0937 = ~pi0780 | n15768;
  assign n17173 = pi1095 & n17167;
  assign n17174 = pi0781 & ~n17167;
  assign po0938 = n17173 | n17174;
  assign n17176 = ~pi0979 & ~pi0984;
  assign n17177 = ~n15815 & ~n17176;
  assign po0939 = n15767 | ~n17177;
  assign n17179 = pi1103 & n17167;
  assign n17180 = pi0783 & ~n17167;
  assign po0940 = n17179 | n17180;
  assign n17182 = pi1104 & n17167;
  assign n17183 = pi0784 & ~n17167;
  assign po0941 = n17182 | n17183;
  assign n17185 = pi1096 & n17167;
  assign n17186 = pi0785 & ~n17167;
  assign po0942 = n17185 | n17186;
  assign n17188 = ~pi0786 & pi0954;
  assign n17189 = ~pi0024 & ~pi0954;
  assign po0943 = n17188 | n17189;
  assign n17191 = pi1098 & n17167;
  assign n17192 = pi0787 & ~n17167;
  assign po0944 = n17191 | n17192;
  assign n17194 = pi1099 & n17167;
  assign n17195 = pi0788 & ~n17167;
  assign po0945 = n17194 | n17195;
  assign n17197 = pi1100 & n17167;
  assign n17198 = pi0789 & ~n17167;
  assign po0946 = n17197 | n17198;
  assign n17200 = pi1101 & n17167;
  assign n17201 = pi0790 & ~n17167;
  assign po0947 = n17200 | n17201;
  assign n17203 = pi1102 & n17167;
  assign n17204 = pi0791 & ~n17167;
  assign po0948 = n17203 | n17204;
  assign n17206 = pi1097 & n17167;
  assign n17207 = pi0792 & ~n17167;
  assign po0949 = n17206 | n17207;
  assign n17209 = pi0968 & n17165;
  assign n17210 = n17164 & n17209;
  assign n17211 = pi0794 & ~n17210;
  assign n17212 = pi1124 & n17210;
  assign po0951 = n17211 | n17212;
  assign n17214 = pi0795 & ~n17210;
  assign n17215 = pi1122 & n17210;
  assign po0952 = n17214 | n17215;
  assign n17217 = pi0278 & ~pi0281;
  assign n17218 = pi0266 & pi0279;
  assign n17219 = ~pi0269 & n17218;
  assign n17220 = ~pi0280 & n17219;
  assign n17221 = n17217 & n17220;
  assign n17222 = ~pi0282 & n17221;
  assign n17223 = ~pi0277 & n17222;
  assign n17224 = ~pi0270 & n17223;
  assign n17225 = ~pi0264 & ~n17224;
  assign n17226 = pi0264 & n17224;
  assign po0953 = n17225 | n17226;
  assign n17228 = pi0798 & ~n17210;
  assign n17229 = pi1118 & n17210;
  assign po0955 = n17228 | n17229;
  assign n17231 = ~pi0799 & ~n17210;
  assign n17232 = pi1101 & n17210;
  assign po0956 = n17231 | n17232;
  assign n17234 = pi0800 & ~n17210;
  assign n17235 = pi1119 & n17210;
  assign po0957 = n17234 | n17235;
  assign n17237 = pi0801 & ~n17210;
  assign n17238 = pi1120 & n17210;
  assign po0958 = n17237 | n17238;
  assign n17240 = n16053 & n16057;
  assign n17241 = ~pi0269 & ~pi0281;
  assign n17242 = ~pi0270 & ~pi0282;
  assign n17243 = n17241 & n17242;
  assign n17244 = n17240 & n17243;
  assign n17245 = ~pi0274 & n17244;
  assign po0959 = ~pi0265 & n17245;
  assign n17247 = ~pi0803 & ~n17210;
  assign n17248 = pi1100 & n17210;
  assign po0960 = n17247 | n17248;
  assign n17250 = pi0804 & ~n17210;
  assign n17251 = pi1103 & n17210;
  assign po0961 = n17250 | n17251;
  assign n17253 = ~pi0270 & ~n16056;
  assign n17254 = pi0270 & n16056;
  assign po0962 = n17253 | n17254;
  assign n17256 = pi0807 & ~n17210;
  assign n17257 = pi1121 & n17210;
  assign po0964 = n17256 | n17257;
  assign n17259 = pi0808 & ~n17210;
  assign n17260 = pi1095 & n17210;
  assign po0965 = n17259 | n17260;
  assign n17262 = ~pi0809 & ~n17210;
  assign n17263 = pi1097 & n17210;
  assign po0966 = n17262 | n17263;
  assign n17265 = pi0810 & ~n17210;
  assign n17266 = pi1102 & n17210;
  assign po0967 = n17265 | n17266;
  assign n17268 = pi0811 & ~n17210;
  assign n17269 = pi1096 & n17210;
  assign po0968 = n17268 | n17269;
  assign n17271 = ~pi0812 & ~n17210;
  assign n17272 = pi1098 & n17210;
  assign po0969 = n17271 | n17272;
  assign n17274 = pi0813 & ~n17210;
  assign n17275 = pi1125 & n17210;
  assign po0970 = n17274 | n17275;
  assign n17277 = ~pi0814 & ~n17210;
  assign n17278 = pi1099 & n17210;
  assign po0971 = n17277 | n17278;
  assign n17280 = pi0815 & ~n17210;
  assign n17281 = pi1104 & n17210;
  assign po0972 = n17280 | n17281;
  assign n17283 = pi0816 & ~n17210;
  assign n17284 = pi1123 & n17210;
  assign po0973 = n17283 | n17284;
  assign n17286 = ~pi0269 & ~n16053;
  assign n17287 = pi0269 & n16053;
  assign po0974 = n17286 | n17287;
  assign n17289 = n16057 & n17242;
  assign n17290 = ~pi0280 & n17241;
  assign n17291 = n16052 & n17290;
  assign n17292 = n17289 & n17291;
  assign n17293 = ~pi0265 & ~n17292;
  assign n17294 = pi0265 & n17292;
  assign po0976 = n17293 | n17294;
  assign n17296 = n16053 & n17243;
  assign n17297 = ~pi0277 & ~n17296;
  assign n17298 = pi0277 & n17296;
  assign po0977 = n17297 | n17298;
  assign po0979 = ~pi0811 & ~pi0893;
  assign n17301 = pi1086 & n2725;
  assign n17302 = n2727 & n3539;
  assign n17303 = pi0982 & ~n17302;
  assign po0981 = n17301 & ~n17303;
  assign n17305 = ~pi1121 & pi1123;
  assign n17306 = pi1121 & ~pi1123;
  assign n17307 = ~n17305 & ~n17306;
  assign n17308 = ~pi1119 & pi1124;
  assign n17309 = pi1119 & ~pi1124;
  assign n17310 = ~n17308 & ~n17309;
  assign n17311 = ~n17307 & n17310;
  assign n17312 = n17307 & ~n17310;
  assign n17313 = ~n17311 & ~n17312;
  assign n17314 = ~pi1120 & pi1122;
  assign n17315 = pi1120 & ~pi1122;
  assign n17316 = ~n17314 & ~n17315;
  assign n17317 = ~pi1118 & pi1125;
  assign n17318 = pi1118 & ~pi1125;
  assign n17319 = ~n17317 & ~n17318;
  assign n17320 = ~n17316 & n17319;
  assign n17321 = n17316 & ~n17319;
  assign n17322 = ~n17320 & ~n17321;
  assign n17323 = ~n17313 & n17322;
  assign n17324 = n17313 & ~n17322;
  assign n17325 = ~n17323 & ~n17324;
  assign n17326 = pi0123 & n16109;
  assign n17327 = ~n17325 & ~n17326;
  assign n17328 = ~pi0825 & n17326;
  assign po0982 = n17327 | n17328;
  assign n17330 = ~pi1111 & pi1116;
  assign n17331 = pi1111 & ~pi1116;
  assign n17332 = ~n17330 & ~n17331;
  assign n17333 = ~pi1113 & pi1115;
  assign n17334 = pi1113 & ~pi1115;
  assign n17335 = ~n17333 & ~n17334;
  assign n17336 = ~n17332 & n17335;
  assign n17337 = n17332 & ~n17335;
  assign n17338 = ~n17336 & ~n17337;
  assign n17339 = ~pi1112 & pi1114;
  assign n17340 = pi1112 & ~pi1114;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = ~pi1110 & pi1117;
  assign n17343 = pi1110 & ~pi1117;
  assign n17344 = ~n17342 & ~n17343;
  assign n17345 = ~n17341 & n17344;
  assign n17346 = n17341 & ~n17344;
  assign n17347 = ~n17345 & ~n17346;
  assign n17348 = ~n17338 & n17347;
  assign n17349 = n17338 & ~n17347;
  assign n17350 = ~n17348 & ~n17349;
  assign n17351 = ~n17326 & ~n17350;
  assign n17352 = ~pi0826 & n17326;
  assign po0983 = n17351 | n17352;
  assign n17354 = ~pi1095 & pi1100;
  assign n17355 = pi1095 & ~pi1100;
  assign n17356 = ~n17354 & ~n17355;
  assign n17357 = ~pi1097 & pi1099;
  assign n17358 = pi1097 & ~pi1099;
  assign n17359 = ~n17357 & ~n17358;
  assign n17360 = ~n17356 & n17359;
  assign n17361 = n17356 & ~n17359;
  assign n17362 = ~n17360 & ~n17361;
  assign n17363 = ~pi1094 & pi1101;
  assign n17364 = pi1094 & ~pi1101;
  assign n17365 = ~n17363 & ~n17364;
  assign n17366 = ~pi1096 & pi1098;
  assign n17367 = pi1096 & ~pi1098;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = ~n17365 & n17368;
  assign n17370 = n17365 & ~n17368;
  assign n17371 = ~n17369 & ~n17370;
  assign n17372 = ~n17362 & n17371;
  assign n17373 = n17362 & ~n17371;
  assign n17374 = ~n17372 & ~n17373;
  assign n17375 = ~n17326 & ~n17374;
  assign n17376 = ~pi0827 & n17326;
  assign po0984 = n17375 | n17376;
  assign n17378 = ~pi1105 & pi1107;
  assign n17379 = pi1105 & ~pi1107;
  assign n17380 = ~n17378 & ~n17379;
  assign n17381 = ~pi1103 & pi1108;
  assign n17382 = pi1103 & ~pi1108;
  assign n17383 = ~n17381 & ~n17382;
  assign n17384 = ~n17380 & n17383;
  assign n17385 = n17380 & ~n17383;
  assign n17386 = ~n17384 & ~n17385;
  assign n17387 = ~pi1104 & pi1106;
  assign n17388 = pi1104 & ~pi1106;
  assign n17389 = ~n17387 & ~n17388;
  assign n17390 = ~pi1102 & pi1109;
  assign n17391 = pi1102 & ~pi1109;
  assign n17392 = ~n17390 & ~n17391;
  assign n17393 = ~n17389 & n17392;
  assign n17394 = n17389 & ~n17392;
  assign n17395 = ~n17393 & ~n17394;
  assign n17396 = ~n17386 & n17395;
  assign n17397 = n17386 & ~n17395;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = ~n17326 & ~n17398;
  assign n17400 = ~pi0828 & n17326;
  assign po0985 = n17399 | n17400;
  assign n17402 = n3539 & n3578;
  assign n17403 = pi0951 & ~n17402;
  assign po0986 = pi1086 & ~n17403;
  assign n17405 = pi0278 & n17220;
  assign n17406 = ~pi0281 & ~n17405;
  assign n17407 = pi0281 & n17405;
  assign po0987 = n17406 | n17407;
  assign n17409 = pi1085 & n2721;
  assign n17410 = ~pi0832 & n17409;
  assign po0989 = n3962 & n17410;
  assign n17412 = pi0833 & ~n2721;
  assign po0990 = n17409 | n17412;
  assign po0991 = pi0946 & n2721;
  assign n17415 = ~pi0282 & ~n17291;
  assign n17416 = pi0282 & n17291;
  assign po0992 = n17415 | n17416;
  assign n17418 = ~pi0955 & pi1043;
  assign n17419 = pi0837 & pi0955;
  assign po0993 = n17418 | n17419;
  assign n17421 = ~pi0955 & pi1041;
  assign n17422 = pi0838 & pi0955;
  assign po0994 = n17421 | n17422;
  assign n17424 = ~pi0955 & pi1068;
  assign n17425 = pi0839 & pi0955;
  assign po0995 = n17424 | n17425;
  assign n17427 = pi0840 & ~n2721;
  assign n17428 = pi1190 & n2721;
  assign po0996 = n17427 | n17428;
  assign n17430 = ~pi0955 & pi1029;
  assign n17431 = pi0842 & pi0955;
  assign po0998 = n17430 | n17431;
  assign n17433 = ~pi0955 & pi1073;
  assign n17434 = pi0843 & pi0955;
  assign po0999 = n17433 | n17434;
  assign n17436 = ~pi0955 & pi1072;
  assign n17437 = pi0844 & pi0955;
  assign po1000 = n17436 | n17437;
  assign n17439 = ~pi0955 & pi1037;
  assign n17440 = pi0845 & pi0955;
  assign po1001 = n17439 | n17440;
  assign n17442 = pi1128 & ~n13876;
  assign n17443 = pi0846 & n13876;
  assign po1002 = n17442 | n17443;
  assign n17445 = ~pi0955 & pi1049;
  assign n17446 = pi0847 & pi0955;
  assign po1003 = n17445 | n17446;
  assign n17448 = ~pi0955 & pi1033;
  assign n17449 = pi0848 & pi0955;
  assign po1004 = n17448 | n17449;
  assign n17451 = pi0849 & ~n2721;
  assign n17452 = pi1192 & n2721;
  assign po1005 = n17451 | n17452;
  assign n17454 = ~pi0955 & pi1042;
  assign n17455 = pi0850 & pi0955;
  assign po1006 = n17454 | n17455;
  assign n17457 = ~pi0955 & pi1039;
  assign n17458 = pi0851 & pi0955;
  assign po1007 = n17457 | n17458;
  assign n17460 = ~pi0955 & pi1056;
  assign n17461 = pi0852 & pi0955;
  assign po1008 = n17460 | n17461;
  assign n17463 = ~pi0955 & pi1074;
  assign n17464 = pi0853 & pi0955;
  assign po1009 = n17463 | n17464;
  assign n17466 = ~pi0955 & pi1045;
  assign n17467 = pi0854 & pi0955;
  assign po1010 = n17466 | n17467;
  assign n17469 = ~pi0955 & pi1059;
  assign n17470 = pi0855 & pi0955;
  assign po1011 = n17469 | n17470;
  assign n17472 = ~pi0955 & pi1061;
  assign n17473 = pi0856 & pi0955;
  assign po1012 = n17472 | n17473;
  assign n17475 = ~pi0955 & pi1052;
  assign n17476 = pi0857 & pi0955;
  assign po1013 = n17475 | n17476;
  assign n17478 = ~pi0955 & pi1081;
  assign n17479 = pi0858 & pi0955;
  assign po1014 = n17478 | n17479;
  assign n17481 = ~pi0955 & pi1064;
  assign n17482 = pi0859 & pi0955;
  assign po1015 = n17481 | n17482;
  assign n17484 = ~pi0955 & pi1070;
  assign n17485 = pi0860 & pi0955;
  assign po1016 = n17484 | n17485;
  assign n17487 = pi1135 & ~n13876;
  assign n17488 = pi0861 & n13876;
  assign po1017 = n17487 | n17488;
  assign n17490 = pi1133 & ~n13876;
  assign n17491 = pi0862 & n13876;
  assign po1018 = n17490 | n17491;
  assign n17493 = pi0863 & ~n2721;
  assign n17494 = pi1193 & n2721;
  assign po1019 = n17493 | n17494;
  assign n17496 = pi0864 & ~n2721;
  assign n17497 = pi1191 & n2721;
  assign po1020 = n17496 | n17497;
  assign n17499 = ~pi0955 & pi1034;
  assign n17500 = pi0865 & pi0955;
  assign po1021 = n17499 | n17500;
  assign n17502 = ~pi0955 & pi1047;
  assign n17503 = pi0866 & pi0955;
  assign po1022 = n17502 | n17503;
  assign n17505 = ~pi0955 & pi1051;
  assign n17506 = pi0867 & pi0955;
  assign po1023 = n17505 | n17506;
  assign n17508 = ~pi0955 & pi1057;
  assign n17509 = pi0868 & pi0955;
  assign po1024 = n17508 | n17509;
  assign n17511 = pi1134 & ~n13876;
  assign n17512 = pi0869 & n13876;
  assign po1025 = n17511 | n17512;
  assign n17514 = ~pi0955 & pi1063;
  assign n17515 = pi0870 & pi0955;
  assign po1026 = n17514 | n17515;
  assign n17517 = ~pi0955 & pi1066;
  assign n17518 = pi0871 & pi0955;
  assign po1027 = n17517 | n17518;
  assign n17520 = ~pi0955 & pi1078;
  assign n17521 = pi0872 & pi0955;
  assign po1028 = n17520 | n17521;
  assign n17523 = ~pi0955 & pi1038;
  assign n17524 = pi0873 & pi0955;
  assign po1029 = n17523 | n17524;
  assign n17526 = ~pi0955 & pi1030;
  assign n17527 = pi0874 & pi0955;
  assign po1030 = n17526 | n17527;
  assign n17529 = pi1130 & ~n13876;
  assign n17530 = pi0875 & n13876;
  assign po1031 = n17529 | n17530;
  assign n17532 = ~pi0955 & pi1031;
  assign n17533 = pi0876 & pi0955;
  assign po1032 = n17532 | n17533;
  assign n17535 = pi1132 & ~n13876;
  assign n17536 = pi0877 & n13876;
  assign po1033 = n17535 | n17536;
  assign n17538 = pi1131 & ~n13876;
  assign n17539 = pi0878 & n13876;
  assign po1034 = n17538 | n17539;
  assign n17541 = pi1129 & ~n13876;
  assign n17542 = pi0879 & n13876;
  assign po1035 = n17541 | n17542;
  assign n17544 = ~pi0955 & pi1075;
  assign n17545 = pi0880 & pi0955;
  assign po1036 = n17544 | n17545;
  assign n17547 = ~pi0955 & pi1053;
  assign n17548 = pi0881 & pi0955;
  assign po1037 = n17547 | n17548;
  assign n17550 = pi1101 & ~n17326;
  assign n17551 = ~pi0883 & n17326;
  assign po1039 = n17550 | n17551;
  assign n17553 = pi1118 & ~n17326;
  assign n17554 = ~pi0884 & n17326;
  assign po1040 = n17553 | n17554;
  assign n17556 = pi1119 & ~n17326;
  assign n17557 = ~pi0885 & n17326;
  assign po1041 = n17556 | n17557;
  assign n17559 = pi1103 & ~n17326;
  assign n17560 = ~pi0886 & n17326;
  assign po1042 = n17559 | n17560;
  assign n17562 = pi1094 & ~n17326;
  assign n17563 = ~pi0887 & n17326;
  assign po1043 = n17562 | n17563;
  assign n17565 = pi1114 & ~n17326;
  assign n17566 = ~pi0888 & n17326;
  assign po1044 = n17565 | n17566;
  assign n17568 = pi1097 & ~n17326;
  assign n17569 = ~pi0889 & n17326;
  assign po1045 = n17568 | n17569;
  assign n17571 = pi1120 & ~n17326;
  assign n17572 = ~pi0890 & n17326;
  assign po1046 = n17571 | n17572;
  assign n17574 = pi1110 & ~n17326;
  assign n17575 = ~pi0891 & n17326;
  assign po1047 = n17574 | n17575;
  assign n17577 = pi1095 & ~n17326;
  assign n17578 = ~pi0892 & n17326;
  assign po1048 = n17577 | n17578;
  assign n17580 = pi1113 & ~n17326;
  assign n17581 = ~pi0894 & n17326;
  assign po1050 = n17580 | n17581;
  assign n17583 = pi1107 & ~n17326;
  assign n17584 = ~pi0895 & n17326;
  assign po1051 = n17583 | n17584;
  assign n17586 = pi1112 & ~n17326;
  assign n17587 = ~pi0896 & n17326;
  assign po1052 = n17586 | n17587;
  assign n17589 = pi1123 & ~n17326;
  assign n17590 = ~pi0898 & n17326;
  assign po1054 = n17589 | n17590;
  assign n17592 = pi1109 & ~n17326;
  assign n17593 = ~pi0899 & n17326;
  assign po1055 = n17592 | n17593;
  assign n17595 = pi1104 & ~n17326;
  assign n17596 = ~pi0900 & n17326;
  assign po1056 = n17595 | n17596;
  assign n17598 = pi1105 & ~n17326;
  assign n17599 = ~pi0902 & n17326;
  assign po1058 = n17598 | n17599;
  assign n17601 = pi1115 & ~n17326;
  assign n17602 = ~pi0903 & n17326;
  assign po1059 = n17601 | n17602;
  assign n17604 = pi1121 & ~n17326;
  assign n17605 = ~pi0904 & n17326;
  assign po1060 = n17604 | n17605;
  assign n17607 = pi1125 & ~n17326;
  assign n17608 = ~pi0905 & n17326;
  assign po1061 = n17607 | n17608;
  assign n17610 = pi1122 & ~n17326;
  assign n17611 = ~pi0906 & n17326;
  assign po1062 = n17610 | n17611;
  assign n17613 = ~pi0604 & ~pi0979;
  assign n17614 = pi0615 & pi0979;
  assign n17615 = ~n17613 & ~n17614;
  assign n17616 = pi0624 & ~pi0979;
  assign n17617 = pi0598 & pi0979;
  assign n17618 = ~n17616 & ~n17617;
  assign n17619 = n17615 & n17618;
  assign n17620 = pi0782 & n17619;
  assign n17621 = ~pi0782 & pi0907;
  assign po1063 = n17620 | n17621;
  assign n17623 = pi1116 & ~n17326;
  assign n17624 = ~pi0908 & n17326;
  assign po1064 = n17623 | n17624;
  assign n17626 = pi1099 & ~n17326;
  assign n17627 = ~pi0909 & n17326;
  assign po1065 = n17626 | n17627;
  assign n17629 = pi1111 & ~n17326;
  assign n17630 = ~pi0910 & n17326;
  assign po1066 = n17629 | n17630;
  assign n17632 = pi1124 & ~n17326;
  assign n17633 = ~pi0911 & n17326;
  assign po1067 = n17632 | n17633;
  assign n17635 = pi1108 & ~n17326;
  assign n17636 = ~pi0912 & n17326;
  assign po1068 = n17635 | n17636;
  assign n17638 = pi1100 & ~n17326;
  assign n17639 = ~pi0913 & n17326;
  assign po1069 = n17638 | n17639;
  assign n17641 = ~pi0280 & ~n16052;
  assign n17642 = pi0280 & n16052;
  assign po1070 = n17641 | n17642;
  assign n17644 = pi1102 & ~n17326;
  assign n17645 = ~pi0915 & n17326;
  assign po1071 = n17644 | n17645;
  assign n17647 = pi1117 & ~n17326;
  assign n17648 = ~pi0916 & n17326;
  assign po1072 = n17647 | n17648;
  assign n17650 = pi1106 & ~n17326;
  assign n17651 = ~pi0917 & n17326;
  assign po1073 = n17650 | n17651;
  assign n17653 = pi1098 & ~n17326;
  assign n17654 = ~pi0918 & n17326;
  assign po1074 = n17653 | n17654;
  assign n17656 = pi1096 & ~n17326;
  assign n17657 = ~pi0919 & n17326;
  assign po1075 = n17656 | n17657;
  assign n17659 = pi0920 & ~pi1087;
  assign n17660 = pi1087 & pi1133;
  assign po1076 = n17659 | n17660;
  assign n17662 = pi0921 & ~pi1087;
  assign n17663 = pi1087 & pi1134;
  assign po1077 = n17662 | n17663;
  assign n17665 = pi0922 & ~pi1087;
  assign n17666 = pi1087 & pi1146;
  assign po1078 = n17665 | n17666;
  assign n17668 = pi0923 & ~pi1087;
  assign n17669 = pi1087 & pi1148;
  assign po1079 = n17668 | n17669;
  assign n17671 = pi0311 & n14260;
  assign po1080 = pi0301 & n17671;
  assign n17673 = pi0925 & ~pi1087;
  assign n17674 = pi1087 & pi1149;
  assign po1081 = n17673 | n17674;
  assign n17676 = pi0926 & ~pi1087;
  assign n17677 = pi1087 & pi1151;
  assign po1082 = n17676 | n17677;
  assign n17679 = pi0927 & ~pi1087;
  assign n17680 = pi1087 & pi1139;
  assign po1083 = n17679 | n17680;
  assign n17682 = pi0928 & ~pi1087;
  assign n17683 = pi1087 & pi1130;
  assign po1084 = n17682 | n17683;
  assign n17685 = pi0929 & ~pi1087;
  assign n17686 = pi1087 & pi1138;
  assign po1085 = n17685 | n17686;
  assign n17688 = pi0930 & ~pi1087;
  assign n17689 = pi1087 & pi1128;
  assign po1086 = n17688 | n17689;
  assign n17691 = pi0931 & ~pi1087;
  assign n17692 = pi1087 & pi1144;
  assign po1087 = n17691 | n17692;
  assign n17694 = pi0932 & ~pi1087;
  assign n17695 = pi1087 & pi1136;
  assign po1088 = n17694 | n17695;
  assign n17697 = pi0933 & ~pi1087;
  assign n17698 = pi1087 & pi1131;
  assign po1089 = n17697 | n17698;
  assign n17700 = pi0934 & ~pi1087;
  assign n17701 = pi1087 & pi1141;
  assign po1090 = n17700 | n17701;
  assign n17703 = pi0935 & ~pi1087;
  assign n17704 = pi1087 & pi1135;
  assign po1091 = n17703 | n17704;
  assign n17706 = pi0936 & ~pi1087;
  assign n17707 = pi1087 & pi1143;
  assign po1092 = n17706 | n17707;
  assign n17709 = pi0937 & ~pi1087;
  assign n17710 = pi1087 & pi1142;
  assign po1093 = n17709 | n17710;
  assign n17712 = pi0938 & ~pi1087;
  assign n17713 = pi1087 & pi1129;
  assign po1094 = n17712 | n17713;
  assign n17715 = pi0939 & ~pi1087;
  assign n17716 = pi1087 & pi1140;
  assign po1095 = n17715 | n17716;
  assign n17718 = pi0940 & ~pi1087;
  assign n17719 = pi1087 & pi1132;
  assign po1096 = n17718 | n17719;
  assign n17721 = pi0941 & ~pi1087;
  assign n17722 = pi1087 & pi1147;
  assign po1097 = n17721 | n17722;
  assign n17724 = pi0942 & ~pi1087;
  assign n17725 = pi1087 & pi1150;
  assign po1098 = n17724 | n17725;
  assign n17727 = pi0943 & ~pi1087;
  assign n17728 = pi1087 & pi1145;
  assign po1099 = n17727 | n17728;
  assign n17730 = pi0944 & ~pi1087;
  assign n17731 = pi1087 & pi1137;
  assign po1100 = n17730 | n17731;
  assign po1101 = n3369 | n3378;
  assign n17734 = pi0782 & ~n17618;
  assign n17735 = ~pi0782 & pi0947;
  assign po1103 = n17734 | n17735;
  assign n17737 = pi0266 & ~n16051;
  assign n17738 = ~pi0266 & n16051;
  assign po1104 = n17737 | n17738;
  assign n17740 = pi0949 & pi0954;
  assign n17741 = ~pi0313 & ~pi0954;
  assign po1105 = n17740 | n17741;
  assign n17743 = pi0957 & pi1086;
  assign po1112 = pi0031 | n17743;
  assign n17745 = pi0278 & ~pi0279;
  assign n17746 = ~pi0278 & pi0279;
  assign po1113 = n17745 | n17746;
  assign po1115 = ~pi0782 & pi0960;
  assign po1116 = ~pi0230 & pi0961;
  assign po1118 = ~pi0782 & pi0963;
  assign po1122 = ~pi0230 & pi0967;
  assign po1124 = ~pi0230 & pi0969;
  assign po1125 = ~pi0782 & pi0970;
  assign po1126 = ~pi0230 & pi0971;
  assign po1127 = ~pi0782 & pi0972;
  assign po1128 = ~pi0230 & pi0974;
  assign po1129 = ~pi0782 & pi0975;
  assign po1131 = ~pi0230 & pi0977;
  assign po1132 = ~pi0782 & pi0978;
  assign po1133 = pi0598 | ~pi0615;
  assign po1137 = pi0604 | pi0624;
  assign po0166 = 1'b1;
  assign po0170 = ~pi1084;
  assign po1110 = ~pi0954;
  assign po1130 = ~pi0278;
  assign po1140 = ~pi0915;
  assign po1141 = ~pi0825;
  assign po1142 = ~pi0826;
  assign po1143 = ~pi0913;
  assign po1144 = ~pi0894;
  assign po1145 = ~pi0905;
  assign po1147 = ~pi0890;
  assign po1149 = ~pi0906;
  assign po1150 = ~pi0896;
  assign po1151 = ~pi0909;
  assign po1152 = ~pi0911;
  assign po1153 = ~pi0908;
  assign po1154 = ~pi0891;
  assign po1155 = ~pi0902;
  assign po1156 = ~pi0903;
  assign po1157 = ~pi0883;
  assign po1158 = ~pi0888;
  assign po1159 = ~pi0919;
  assign po1160 = ~pi0886;
  assign po1161 = ~pi0912;
  assign po1162 = ~pi0895;
  assign po1163 = ~pi0916;
  assign po1164 = ~pi0889;
  assign po1165 = ~pi0900;
  assign po1166 = ~pi0885;
  assign po1167 = ~pi0904;
  assign po1168 = ~pi0899;
  assign po1169 = ~pi0918;
  assign po1170 = ~pi0898;
  assign po1171 = ~pi0917;
  assign po1172 = ~pi0827;
  assign po1173 = ~pi0887;
  assign po1174 = ~pi0884;
  assign po1175 = ~pi0910;
  assign po1176 = ~pi0828;
  assign po1177 = ~pi0892;
  assign po0000 = pi0668;
  assign po0001 = pi0672;
  assign po0002 = pi0664;
  assign po0003 = pi0667;
  assign po0004 = pi0676;
  assign po0005 = pi0673;
  assign po0006 = pi0675;
  assign po0007 = pi0666;
  assign po0008 = pi0679;
  assign po0009 = pi0674;
  assign po0010 = pi0663;
  assign po0011 = pi0670;
  assign po0012 = pi0677;
  assign po0013 = pi0682;
  assign po0014 = pi0671;
  assign po0015 = pi0678;
  assign po0016 = pi0718;
  assign po0017 = pi0707;
  assign po0018 = pi0708;
  assign po0019 = pi0713;
  assign po0020 = pi0711;
  assign po0021 = pi0716;
  assign po0022 = pi0733;
  assign po0023 = pi0712;
  assign po0024 = pi0689;
  assign po0025 = pi0717;
  assign po0026 = pi0692;
  assign po0027 = pi0719;
  assign po0028 = pi0722;
  assign po0029 = pi0714;
  assign po0030 = pi0720;
  assign po0031 = pi0685;
  assign po0032 = pi0837;
  assign po0033 = pi0850;
  assign po0034 = pi0872;
  assign po0035 = pi0871;
  assign po0036 = pi0881;
  assign po0037 = pi0866;
  assign po0038 = pi0876;
  assign po0039 = pi0873;
  assign po0040 = pi0874;
  assign po0041 = pi0859;
  assign po0042 = pi0855;
  assign po0043 = pi0852;
  assign po0044 = pi0870;
  assign po0045 = pi0848;
  assign po0046 = pi0865;
  assign po0047 = pi0856;
  assign po0048 = pi0853;
  assign po0049 = pi0847;
  assign po0050 = pi0857;
  assign po0051 = pi0854;
  assign po0052 = pi0858;
  assign po0053 = pi0845;
  assign po0054 = pi0838;
  assign po0055 = pi0842;
  assign po0056 = pi0843;
  assign po0057 = pi0839;
  assign po0058 = pi0844;
  assign po0059 = pi0868;
  assign po0060 = pi0851;
  assign po0061 = pi0867;
  assign po0062 = pi0880;
  assign po0063 = pi0860;
  assign po0064 = pi1024;
  assign po0065 = pi1028;
  assign po0066 = pi1009;
  assign po0067 = pi1014;
  assign po0068 = pi1019;
  assign po0069 = pi0999;
  assign po0070 = pi0990;
  assign po0071 = pi1006;
  assign po0072 = pi0987;
  assign po0073 = pi1010;
  assign po0074 = pi1015;
  assign po0075 = pi1004;
  assign po0076 = pi1021;
  assign po0077 = pi1012;
  assign po0078 = pi1011;
  assign po0079 = pi1018;
  assign po0080 = pi1003;
  assign po0081 = pi1026;
  assign po0082 = pi0997;
  assign po0083 = pi0991;
  assign po0084 = pi1007;
  assign po0085 = pi1005;
  assign po0086 = pi1002;
  assign po0087 = pi1013;
  assign po0088 = pi1025;
  assign po0089 = pi1016;
  assign po0090 = pi0994;
  assign po0091 = pi1017;
  assign po0092 = pi0996;
  assign po0093 = pi1020;
  assign po0094 = pi1000;
  assign po0095 = pi0992;
  assign po0096 = pi0031;
  assign po0097 = pi0080;
  assign po0098 = pi0893;
  assign po0099 = pi0467;
  assign po0100 = pi0078;
  assign po0101 = pi0112;
  assign po0102 = pi0013;
  assign po0103 = pi0025;
  assign po0104 = pi0226;
  assign po0105 = pi0127;
  assign po0106 = pi0822;
  assign po0107 = pi0808;
  assign po0108 = pi0227;
  assign po0109 = pi0477;
  assign po0110 = pi0834;
  assign po0111 = pi0229;
  assign po0112 = pi0012;
  assign po0113 = pi0011;
  assign po0114 = pi0010;
  assign po0115 = pi0009;
  assign po0116 = pi0008;
  assign po0117 = pi0007;
  assign po0118 = pi0006;
  assign po0119 = pi0005;
  assign po0120 = pi0004;
  assign po0121 = pi0003;
  assign po0122 = pi0000;
  assign po0123 = pi0002;
  assign po0124 = pi0001;
  assign po0125 = pi0310;
  assign po0126 = pi0302;
  assign po0127 = pi0475;
  assign po0128 = pi0474;
  assign po0129 = pi0466;
  assign po0130 = pi0473;
  assign po0131 = pi0471;
  assign po0132 = pi0472;
  assign po0133 = pi0470;
  assign po0134 = pi0469;
  assign po0135 = pi0465;
  assign po0136 = pi1022;
  assign po0137 = pi1027;
  assign po0138 = pi0989;
  assign po0139 = pi0988;
  assign po0140 = pi0028;
  assign po0141 = pi0027;
  assign po0142 = pi0026;
  assign po0143 = pi0029;
  assign po0144 = pi0015;
  assign po0145 = pi0014;
  assign po0146 = pi0021;
  assign po0147 = pi0020;
  assign po0148 = pi0019;
  assign po0149 = pi0018;
  assign po0150 = pi0017;
  assign po0151 = pi0016;
  assign po0152 = pi1090;
  assign po0168 = pi0228;
  assign po0169 = pi0022;
  assign po0179 = pi1083;
  assign po0180 = pi0023;
  assign po0181 = po0167;
  assign po0188 = pi0037;
  assign po0263 = pi0117;
  assign po0285 = pi0131;
  assign po0386 = pi0232;
  assign po0388 = pi0236;
  assign po0636 = pi0583;
  assign po1053 = pi0067;
  assign po1108 = pi1128;
  assign po1109 = pi0964;
  assign po1111 = pi0965;
  assign po1114 = pi0985;
  assign po1117 = pi1008;
  assign po1119 = pi1023;
  assign po1120 = pi0998;
  assign po1121 = pi1001;
  assign po1123 = pi1129;
  assign po1134 = pi1058;
  assign po1136 = pi0299;
  assign po1138 = pi1069;
  assign po1139 = pi1046;
  assign po1146 = pi1089;
  assign po1148 = pi1088;
  assign po1178 = pi1181;
  assign po1179 = pi1166;
  assign po1180 = pi1164;
  assign po1181 = pi1132;
  assign po1182 = pi1171;
  assign po1183 = pi1172;
  assign po1184 = pi0863;
  assign po1185 = pi1197;
  assign po1186 = pi1179;
  assign po1187 = pi1165;
  assign po1188 = pi1186;
  assign po1189 = pi1131;
  assign po1190 = pi1180;
  assign po1191 = pi1159;
  assign po1192 = pi1158;
  assign po1193 = pi1092;
  assign po1194 = pi1177;
  assign po1195 = pi0230;
  assign po1196 = pi1163;
  assign po1197 = pi1130;
  assign po1198 = pi1175;
  assign po1199 = pi0849;
  assign po1200 = pi1187;
  assign po1201 = pi1176;
  assign po1202 = pi1162;
  assign po1203 = pi1169;
  assign po1204 = pi1185;
  assign po1205 = pi1093;
  assign po1206 = pi1168;
  assign po1207 = pi1173;
  assign po1208 = pi1196;
  assign po1209 = pi1170;
  assign po1210 = pi1167;
  assign po1211 = pi1195;
  assign po1212 = pi1161;
  assign po1213 = pi0840;
  assign po1214 = pi1183;
  assign po1215 = pi1189;
  assign po1216 = pi0864;
  assign po1217 = pi1184;
  assign po1218 = pi1182;
  assign po1219 = pi1174;
  assign po1220 = pi1188;
  assign po1221 = pi1091;
  assign po1222 = pi1160;
  assign po1223 = pi1194;
  assign po1224 = pi1178;
endmodule


