module spi ( 
    pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008, pi009,
    pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018, pi019,
    pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028, pi029,
    pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038, pi039,
    pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048, pi049,
    pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058, pi059,
    pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068, pi069,
    pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078, pi079,
    pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088, pi089,
    pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098, pi099,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148, pi149,
    pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159,
    pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188, pi189,
    pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198, pi199,
    pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208, pi209,
    pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218, pi219,
    pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228, pi229,
    pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238, pi239,
    pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249,
    pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273,
    po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275  );
  input  pi000, pi001, pi002, pi003, pi004, pi005, pi006, pi007, pi008,
    pi009, pi010, pi011, pi012, pi013, pi014, pi015, pi016, pi017, pi018,
    pi019, pi020, pi021, pi022, pi023, pi024, pi025, pi026, pi027, pi028,
    pi029, pi030, pi031, pi032, pi033, pi034, pi035, pi036, pi037, pi038,
    pi039, pi040, pi041, pi042, pi043, pi044, pi045, pi046, pi047, pi048,
    pi049, pi050, pi051, pi052, pi053, pi054, pi055, pi056, pi057, pi058,
    pi059, pi060, pi061, pi062, pi063, pi064, pi065, pi066, pi067, pi068,
    pi069, pi070, pi071, pi072, pi073, pi074, pi075, pi076, pi077, pi078,
    pi079, pi080, pi081, pi082, pi083, pi084, pi085, pi086, pi087, pi088,
    pi089, pi090, pi091, pi092, pi093, pi094, pi095, pi096, pi097, pi098,
    pi099, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146, pi147, pi148,
    pi149, pi150, pi151, pi152, pi153, pi154, pi155, pi156, pi157, pi158,
    pi159, pi160, pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168,
    pi169, pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197, pi198,
    pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206, pi207, pi208,
    pi209, pi210, pi211, pi212, pi213, pi214, pi215, pi216, pi217, pi218,
    pi219, pi220, pi221, pi222, pi223, pi224, pi225, pi226, pi227, pi228,
    pi229, pi230, pi231, pi232, pi233, pi234, pi235, pi236, pi237, pi238,
    pi239, pi240, pi241, pi242, pi243, pi244, pi245, pi246, pi247, pi248,
    pi249, pi250, pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258,
    pi259, pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273;
  output po000, po001, po002, po003, po004, po005, po006, po007, po008, po009,
    po010, po011, po012, po013, po014, po015, po016, po017, po018, po019,
    po020, po021, po022, po023, po024, po025, po026, po027, po028, po029,
    po030, po031, po032, po033, po034, po035, po036, po037, po038, po039,
    po040, po041, po042, po043, po044, po045, po046, po047, po048, po049,
    po050, po051, po052, po053, po054, po055, po056, po057, po058, po059,
    po060, po061, po062, po063, po064, po065, po066, po067, po068, po069,
    po070, po071, po072, po073, po074, po075, po076, po077, po078, po079,
    po080, po081, po082, po083, po084, po085, po086, po087, po088, po089,
    po090, po091, po092, po093, po094, po095, po096, po097, po098, po099,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141, po142, po143, po144, po145, po146, po147, po148, po149,
    po150, po151, po152, po153, po154, po155, po156, po157, po158, po159,
    po160, po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188, po189,
    po190, po191, po192, po193, po194, po195, po196, po197, po198, po199,
    po200, po201, po202, po203, po204, po205, po206, po207, po208, po209,
    po210, po211, po212, po213, po214, po215, po216, po217, po218, po219,
    po220, po221, po222, po223, po224, po225, po226, po227, po228, po229,
    po230, po231, po232, po233, po234, po235, po236, po237, po238, po239,
    po240, po241, po242, po243, po244, po245, po246, po247, po248, po249,
    po250, po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275;
  wire n552, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
    n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
    n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
    n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
    n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
    n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
    n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
    n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
    n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1211, n1212, n1213,
    n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1293, n1294, n1295, n1296, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
    n1382, n1383, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
    n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
    n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
    n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
    n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
    n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
    n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
    n1742, n1743, n1744, n1745, n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
    n1763, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
    n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1856, n1857, n1858,
    n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
    n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
    n1922, n1923, n1924, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
    n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
    n1986, n1987, n1988, n1990, n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
    n2082, n2083, n2084, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
    n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
    n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
    n2306, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
    n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
    n2381, n2382, n2383, n2384, n2385, n2386, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
    n2402, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2433, n2434,
    n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2527, n2528, n2529, n2530,
    n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2600, n2601, n2602, n2603, n2604, n2605,
    n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
    n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2731, n2732, n2733, n2734, n2735,
    n2736, n2737, n2738, n2739, n2740, n2741, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
    n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2870, n2871, n2872, n2873, n2874, n2875,
    n2876, n2877, n2878, n2879, n2880, n2881, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
    n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3099, n3100, n3101,
    n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3135, n3136, n3137, n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3165, n3166,
    n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
    n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
    n3188, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
    n3702, n3703, n3704, n3705, n3706, n3707, n3709, n3710, n3711, n3712,
    n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
    n3734, n3735, n3736, n3737, n3738, n3739, n3741, n3742, n3743, n3744,
    n3745, n3746, n3748, n3749, n3750, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3773, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784, n3786, n3787, n3788, n3790,
    n3791, n3792, n3793, n3794, n3795, n3797, n3798, n3799, n3800, n3801,
    n3802, n3804, n3805, n3806, n3807, n3809, n3810, n3811, n3812, n3813,
    n3814, n3816, n3817, n3819, n3820, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3846, n3847,
    n3848, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3862, n3863, n3864, n3865, n3866, n3867, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
    n3881, n3882, n3884, n3885, n3886, n3887, n3888, n3890, n3891, n3893,
    n3894, n3896, n3897, n3898, n3899, n3900, n3901, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3911, n3912, n3913, n3915, n3916, n3918,
    n3919, n3921, n3922, n3924, n3925, n3926, n3927, n3928, n3930, n3931,
    n3933, n3934, n3936, n3937, n3938, n3939, n3941, n3942, n3944, n3945,
    n3946, n3947, n3948, n3950, n3951, n3953, n3954, n3955, n3956, n3958,
    n3959, n3960, n3961, n3963, n3964, n3965, n3966, n3967, n3969, n3970,
    n3971, n3972, n3973, n3975, n3976, n3977, n3978, n3980, n3981, n3983,
    n3984, n3986, n3987, n3989, n3990, n3992, n3993, n3995, n3996, n3998,
    n3999, n4001, n4002, n4004, n4005, n4007, n4008, n4010, n4011, n4013,
    n4014, n4016, n4017, n4019, n4020, n4022, n4023, n4025, n4026, n4027,
    n4028, n4029, n4031, n4032, n4033, n4034, n4035, n4036, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4065, n4066, n4067, n4068, n4069, n4070, n4072,
    n4073, n4074, n4075, n4076, n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4086, n4087, n4089, n4090, n4092, n4093, n4095, n4096, n4098,
    n4099, n4101, n4102, n4104, n4105, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4133,
    n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4227, n4228, n4229, n4230, n4231,
    n4232, n4233, n4234, n4235, n4236, n4238, n4239, n4240, n4241, n4242,
    n4243, n4244, n4245, n4247, n4248, n4249, n4250, n4251, n4252, n4254,
    n4255, n4256, n4257, n4258, n4259, n4261, n4262, n4263, n4264, n4265,
    n4266, n4268, n4269, n4270, n4271, n4272, n4273, n4275, n4276, n4277,
    n4278, n4279, n4280, n4282, n4283, n4284, n4285, n4286, n4287, n4289,
    n4290, n4291, n4292, n4293, n4294, n4296, n4297, n4298, n4299, n4300,
    n4301, n4303, n4304, n4305, n4306, n4307, n4308, n4310, n4311, n4312,
    n4313, n4314, n4315, n4317, n4318, n4319, n4320, n4321, n4322, n4324,
    n4325, n4326, n4327, n4328, n4329, n4331, n4332, n4333, n4334, n4335,
    n4336, n4338, n4339, n4340, n4341, n4342, n4343, n4345, n4346, n4347,
    n4348, n4349, n4350, n4352, n4353, n4354, n4355, n4356, n4357;
  assign n552 = ~pi136 & ~pi152;
  assign po036 = pi196 | n552;
  assign po037 = pi194 | n552;
  assign po038 = pi197 | n552;
  assign po039 = pi193 | n552;
  assign po040 = pi198 | n552;
  assign po041 = pi192 | n552;
  assign po042 = pi199 | n552;
  assign po043 = pi195 | n552;
  assign n561 = pi232 & pi233;
  assign n562 = ~pi236 & ~pi237;
  assign n563 = n561 & n562;
  assign n564 = pi231 & n563;
  assign n565 = ~pi136 & ~pi235;
  assign n566 = n564 & n565;
  assign n567 = ~pi136 & n564;
  assign n568 = pi235 & n567;
  assign n569 = ~n566 & n568;
  assign n570 = pi000 & ~pi270;
  assign n571 = pi245 & pi270;
  assign n572 = ~n570 & ~n571;
  assign n573 = n569 & ~n572;
  assign n574 = pi232 & ~pi235;
  assign n575 = pi231 & n574;
  assign n576 = ~pi136 & pi236;
  assign n577 = pi233 & ~pi237;
  assign n578 = n576 & n577;
  assign n579 = n575 & n578;
  assign n580 = pi000 & n579;
  assign n581 = pi232 & pi235;
  assign n582 = n576 & n581;
  assign n583 = n577 & n582;
  assign n584 = pi231 & n583;
  assign n585 = pi000 & n584;
  assign n586 = pi138 & pi146;
  assign n587 = ~pi187 & ~pi190;
  assign n588 = ~pi142 & ~pi148;
  assign n589 = n587 & n588;
  assign n590 = ~pi139 & n589;
  assign n591 = ~pi130 & ~pi133;
  assign n592 = n590 & n591;
  assign n593 = ~pi140 & n592;
  assign n594 = ~pi129 & n593;
  assign n595 = ~pi138 & ~pi145;
  assign n596 = ~n594 & ~n595;
  assign n597 = ~n586 & n596;
  assign n598 = pi234 & n597;
  assign n599 = ~pi138 & pi139;
  assign n600 = pi187 & pi190;
  assign n601 = pi142 & pi148;
  assign n602 = n600 & n601;
  assign n603 = ~pi139 & n602;
  assign n604 = pi139 & ~n602;
  assign n605 = ~n603 & ~n604;
  assign n606 = pi138 & ~n605;
  assign n607 = ~n599 & ~n606;
  assign n608 = pi177 & n607;
  assign n609 = ~pi138 & pi148;
  assign n610 = pi148 & ~n600;
  assign n611 = ~pi148 & n600;
  assign n612 = ~n610 & ~n611;
  assign n613 = pi138 & ~n612;
  assign n614 = ~n609 & ~n613;
  assign n615 = ~pi156 & ~n614;
  assign n616 = pi138 & ~pi190;
  assign n617 = ~pi138 & pi190;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~pi150 & ~n618;
  assign n620 = ~pi187 & pi190;
  assign n621 = pi187 & ~pi190;
  assign n622 = ~n620 & ~n621;
  assign n623 = pi138 & ~n622;
  assign n624 = ~pi138 & pi187;
  assign n625 = ~n623 & ~n624;
  assign n626 = ~pi171 & ~n625;
  assign n627 = ~n619 & ~n626;
  assign n628 = ~n615 & n627;
  assign n629 = ~pi138 & pi142;
  assign n630 = pi148 & n600;
  assign n631 = ~pi142 & n630;
  assign n632 = pi142 & ~n630;
  assign n633 = ~n631 & ~n632;
  assign n634 = pi138 & ~n633;
  assign n635 = ~n629 & ~n634;
  assign n636 = ~pi176 & ~n635;
  assign n637 = ~pi177 & ~n607;
  assign n638 = ~n636 & ~n637;
  assign n639 = n628 & n638;
  assign n640 = ~n608 & ~n639;
  assign n641 = pi156 & ~n609;
  assign n642 = ~n613 & n641;
  assign n643 = pi171 & n625;
  assign n644 = ~n615 & n643;
  assign n645 = ~n642 & ~n644;
  assign n646 = n638 & ~n645;
  assign n647 = pi176 & n635;
  assign n648 = ~n637 & n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = n640 & n649;
  assign n651 = ~pi138 & pi140;
  assign n652 = pi139 & n602;
  assign n653 = ~pi140 & n652;
  assign n654 = pi140 & ~n652;
  assign n655 = ~n653 & ~n654;
  assign n656 = pi138 & ~n655;
  assign n657 = ~n651 & ~n656;
  assign n658 = pi161 & n657;
  assign n659 = ~pi161 & ~n657;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n650 & n660;
  assign n662 = n650 & ~n660;
  assign n663 = ~n661 & ~n662;
  assign n664 = pi143 & n663;
  assign n665 = pi138 & pi140;
  assign n666 = ~pi139 & ~pi142;
  assign n667 = ~pi190 & n666;
  assign n668 = ~pi148 & n667;
  assign n669 = ~pi187 & n668;
  assign n670 = ~pi140 & n669;
  assign n671 = pi140 & ~n669;
  assign n672 = ~n670 & ~n671;
  assign n673 = ~pi138 & ~n672;
  assign n674 = ~n665 & ~n673;
  assign n675 = ~pi143 & ~n674;
  assign n676 = ~n664 & ~n675;
  assign n677 = ~pi148 & ~pi190;
  assign n678 = ~pi187 & n677;
  assign n679 = ~pi142 & n678;
  assign n680 = pi139 & n679;
  assign n681 = ~pi139 & ~n679;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~pi138 & n682;
  assign n684 = pi138 & pi139;
  assign n685 = ~pi143 & ~n684;
  assign n686 = ~n683 & n685;
  assign n687 = ~n627 & ~n643;
  assign n688 = ~n615 & ~n687;
  assign n689 = ~n636 & n688;
  assign n690 = ~n636 & n642;
  assign n691 = ~n647 & ~n690;
  assign n692 = ~n689 & n691;
  assign n693 = ~n608 & ~n637;
  assign n694 = ~n692 & n693;
  assign n695 = pi143 & n694;
  assign n696 = pi143 & ~n693;
  assign n697 = n692 & n696;
  assign n698 = ~n695 & ~n697;
  assign n699 = ~n686 & n698;
  assign n700 = pi138 & pi142;
  assign n701 = pi142 & ~n678;
  assign n702 = ~n679 & ~n701;
  assign n703 = ~pi138 & ~n702;
  assign n704 = ~n700 & ~n703;
  assign n705 = ~pi143 & ~n704;
  assign n706 = ~n628 & n645;
  assign n707 = ~n636 & ~n647;
  assign n708 = pi143 & n707;
  assign n709 = n706 & n708;
  assign n710 = ~n706 & ~n707;
  assign n711 = pi143 & n710;
  assign n712 = ~n709 & ~n711;
  assign n713 = ~n705 & n712;
  assign n714 = ~n615 & ~n642;
  assign n715 = ~n687 & ~n714;
  assign n716 = n687 & n714;
  assign n717 = ~n715 & ~n716;
  assign n718 = pi143 & ~n717;
  assign n719 = pi138 & pi148;
  assign n720 = pi148 & ~n587;
  assign n721 = ~n678 & ~n720;
  assign n722 = ~pi138 & ~n721;
  assign n723 = ~n719 & ~n722;
  assign n724 = ~pi143 & ~n723;
  assign n725 = ~n718 & ~n724;
  assign n726 = ~n626 & ~n643;
  assign n727 = n619 & n726;
  assign n728 = ~n619 & ~n726;
  assign n729 = ~n727 & ~n728;
  assign n730 = pi143 & ~n729;
  assign n731 = pi138 & pi187;
  assign n732 = ~n587 & ~n600;
  assign n733 = ~pi138 & ~n732;
  assign n734 = ~n731 & ~n733;
  assign n735 = ~pi143 & ~n734;
  assign n736 = ~n730 & ~n735;
  assign n737 = pi150 & n618;
  assign n738 = pi143 & ~n737;
  assign n739 = ~n619 & n738;
  assign n740 = ~pi138 & ~pi190;
  assign n741 = pi138 & pi190;
  assign n742 = ~pi143 & ~n741;
  assign n743 = ~n740 & n742;
  assign n744 = ~n739 & ~n743;
  assign n745 = pi045 & ~n744;
  assign n746 = pi041 & n744;
  assign n747 = ~n745 & ~n746;
  assign n748 = ~n736 & ~n747;
  assign n749 = ~n619 & ~n737;
  assign n750 = pi143 & ~n749;
  assign n751 = ~n740 & ~n741;
  assign n752 = ~pi143 & ~n751;
  assign n753 = ~n750 & ~n752;
  assign n754 = pi043 & ~n753;
  assign n755 = pi040 & ~n744;
  assign n756 = ~n754 & ~n755;
  assign n757 = n736 & ~n756;
  assign n758 = ~n748 & ~n757;
  assign n759 = n725 & ~n758;
  assign n760 = pi011 & n744;
  assign n761 = pi042 & ~n744;
  assign n762 = ~n760 & ~n761;
  assign n763 = n736 & ~n762;
  assign n764 = pi013 & n744;
  assign n765 = pi012 & ~n744;
  assign n766 = ~n764 & ~n765;
  assign n767 = ~n736 & ~n766;
  assign n768 = ~n763 & ~n767;
  assign n769 = ~n725 & ~n768;
  assign n770 = ~n759 & ~n769;
  assign n771 = n713 & ~n770;
  assign n772 = pi017 & ~n753;
  assign n773 = pi016 & ~n744;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~n736 & ~n774;
  assign n776 = pi015 & n744;
  assign n777 = pi031 & ~n744;
  assign n778 = ~n776 & ~n777;
  assign n779 = n736 & ~n778;
  assign n780 = ~n775 & ~n779;
  assign n781 = ~n725 & ~n780;
  assign n782 = pi046 & ~n744;
  assign n783 = pi014 & n744;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~n736 & ~n784;
  assign n786 = pi044 & ~n744;
  assign n787 = pi032 & n744;
  assign n788 = ~n786 & ~n787;
  assign n789 = n736 & ~n788;
  assign n790 = ~n785 & ~n789;
  assign n791 = n725 & ~n790;
  assign n792 = ~n781 & ~n791;
  assign n793 = ~n713 & ~n792;
  assign n794 = ~n771 & ~n793;
  assign n795 = n699 & n794;
  assign n796 = ~n705 & ~n711;
  assign n797 = ~n709 & n796;
  assign n798 = pi047 & n744;
  assign n799 = pi048 & ~n744;
  assign n800 = ~n798 & ~n799;
  assign n801 = ~n736 & ~n800;
  assign n802 = pi039 & n744;
  assign n803 = pi010 & ~n744;
  assign n804 = ~n802 & ~n803;
  assign n805 = n736 & ~n804;
  assign n806 = ~n801 & ~n805;
  assign n807 = ~n725 & ~n806;
  assign n808 = pi038 & n744;
  assign n809 = pi037 & ~n744;
  assign n810 = ~n808 & ~n809;
  assign n811 = n736 & ~n810;
  assign n812 = pi009 & n744;
  assign n813 = pi008 & ~n744;
  assign n814 = ~n812 & ~n813;
  assign n815 = ~n736 & ~n814;
  assign n816 = ~n811 & ~n815;
  assign n817 = n725 & ~n816;
  assign n818 = ~n807 & ~n817;
  assign n819 = ~n797 & ~n818;
  assign n820 = pi036 & ~n744;
  assign n821 = pi007 & n744;
  assign n822 = ~n820 & ~n821;
  assign n823 = ~n736 & ~n822;
  assign n824 = pi035 & ~n753;
  assign n825 = pi006 & ~n744;
  assign n826 = ~n824 & ~n825;
  assign n827 = n736 & ~n826;
  assign n828 = ~n823 & ~n827;
  assign n829 = ~n725 & ~n828;
  assign n830 = pi034 & ~n753;
  assign n831 = pi005 & ~n744;
  assign n832 = ~n830 & ~n831;
  assign n833 = ~n736 & ~n832;
  assign n834 = pi004 & n744;
  assign n835 = pi033 & ~n744;
  assign n836 = ~n834 & ~n835;
  assign n837 = n736 & ~n836;
  assign n838 = ~n833 & ~n837;
  assign n839 = n725 & ~n838;
  assign n840 = ~n829 & ~n839;
  assign n841 = n713 & ~n840;
  assign n842 = ~n819 & ~n841;
  assign n843 = ~n699 & n842;
  assign n844 = ~n795 & ~n843;
  assign n845 = n676 & n844;
  assign n846 = pi087 & n744;
  assign n847 = pi120 & ~n744;
  assign n848 = ~n846 & ~n847;
  assign n849 = ~n736 & ~n848;
  assign n850 = pi127 & n744;
  assign n851 = pi108 & ~n744;
  assign n852 = ~n850 & ~n851;
  assign n853 = n736 & ~n852;
  assign n854 = ~n849 & ~n853;
  assign n855 = ~n725 & ~n854;
  assign n856 = pi097 & ~n744;
  assign n857 = pi121 & n744;
  assign n858 = ~n856 & ~n857;
  assign n859 = ~n736 & ~n858;
  assign n860 = pi104 & n744;
  assign n861 = pi086 & ~n744;
  assign n862 = ~n860 & ~n861;
  assign n863 = n736 & ~n862;
  assign n864 = ~n859 & ~n863;
  assign n865 = n725 & ~n864;
  assign n866 = ~n855 & ~n865;
  assign n867 = n713 & ~n866;
  assign n868 = pi090 & n744;
  assign n869 = pi093 & ~n744;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n736 & ~n870;
  assign n872 = pi088 & n744;
  assign n873 = pi102 & ~n744;
  assign n874 = ~n872 & ~n873;
  assign n875 = n736 & ~n874;
  assign n876 = ~n871 & ~n875;
  assign n877 = n725 & ~n876;
  assign n878 = pi094 & n744;
  assign n879 = pi092 & ~n744;
  assign n880 = ~n878 & ~n879;
  assign n881 = ~n736 & ~n880;
  assign n882 = pi095 & ~n744;
  assign n883 = pi091 & n744;
  assign n884 = ~n882 & ~n883;
  assign n885 = n736 & ~n884;
  assign n886 = ~n881 & ~n885;
  assign n887 = ~n725 & ~n886;
  assign n888 = ~n877 & ~n887;
  assign n889 = ~n713 & ~n888;
  assign n890 = ~n867 & ~n889;
  assign n891 = n699 & n890;
  assign n892 = pi096 & ~n744;
  assign n893 = pi119 & n744;
  assign n894 = ~n892 & ~n893;
  assign n895 = ~n736 & ~n894;
  assign n896 = pi089 & n744;
  assign n897 = pi118 & ~n744;
  assign n898 = ~n896 & ~n897;
  assign n899 = n736 & ~n898;
  assign n900 = ~n895 & ~n899;
  assign n901 = n725 & ~n900;
  assign n902 = pi115 & ~n753;
  assign n903 = pi123 & ~n744;
  assign n904 = ~n902 & ~n903;
  assign n905 = ~n736 & ~n904;
  assign n906 = pi122 & n744;
  assign n907 = pi116 & ~n744;
  assign n908 = ~n906 & ~n907;
  assign n909 = n736 & ~n908;
  assign n910 = ~n905 & ~n909;
  assign n911 = ~n725 & ~n910;
  assign n912 = ~n901 & ~n911;
  assign n913 = n713 & ~n912;
  assign n914 = pi126 & ~n744;
  assign n915 = pi085 & ~n753;
  assign n916 = ~n914 & ~n915;
  assign n917 = ~n736 & ~n916;
  assign n918 = pi105 & ~n744;
  assign n919 = pi125 & n744;
  assign n920 = ~n918 & ~n919;
  assign n921 = n736 & ~n920;
  assign n922 = ~n917 & ~n921;
  assign n923 = ~n725 & ~n922;
  assign n924 = pi124 & ~n753;
  assign n925 = pi117 & ~n744;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n736 & ~n926;
  assign n928 = pi103 & ~n753;
  assign n929 = pi084 & ~n744;
  assign n930 = ~n928 & ~n929;
  assign n931 = n736 & ~n930;
  assign n932 = ~n927 & ~n931;
  assign n933 = n725 & ~n932;
  assign n934 = ~n923 & ~n933;
  assign n935 = ~n797 & ~n934;
  assign n936 = ~n913 & ~n935;
  assign n937 = ~n699 & n936;
  assign n938 = ~n891 & ~n937;
  assign n939 = ~n676 & n938;
  assign n940 = ~n845 & ~n939;
  assign n941 = ~pi139 & n587;
  assign n942 = ~pi140 & n588;
  assign n943 = n941 & n942;
  assign n944 = pi133 & ~n943;
  assign n945 = ~pi133 & n943;
  assign n946 = ~n944 & ~n945;
  assign n947 = ~pi138 & ~n946;
  assign n948 = pi133 & pi138;
  assign n949 = ~n947 & ~n948;
  assign n950 = ~pi143 & ~n949;
  assign n951 = ~pi133 & ~pi138;
  assign n952 = pi140 & pi142;
  assign n953 = n630 & n952;
  assign n954 = pi139 & n953;
  assign n955 = pi133 & ~n954;
  assign n956 = ~pi133 & n954;
  assign n957 = ~n955 & ~n956;
  assign n958 = pi138 & n957;
  assign n959 = ~n951 & ~n958;
  assign n960 = ~pi178 & n959;
  assign n961 = pi178 & ~n959;
  assign n962 = ~n960 & ~n961;
  assign n963 = ~n637 & ~n691;
  assign n964 = ~n608 & ~n963;
  assign n965 = ~n659 & ~n964;
  assign n966 = n638 & n688;
  assign n967 = ~n659 & n966;
  assign n968 = ~n965 & ~n967;
  assign n969 = ~n658 & n968;
  assign n970 = ~n962 & n969;
  assign n971 = n962 & ~n969;
  assign n972 = ~n970 & ~n971;
  assign n973 = pi143 & n972;
  assign n974 = ~n950 & ~n973;
  assign n975 = ~n597 & ~n974;
  assign n976 = ~n940 & n975;
  assign n977 = ~n598 & ~n976;
  assign n978 = pi063 & n744;
  assign n979 = pi056 & ~n744;
  assign n980 = ~n978 & ~n979;
  assign n981 = ~n736 & ~n980;
  assign n982 = pi064 & n744;
  assign n983 = pi022 & ~n744;
  assign n984 = ~n982 & ~n983;
  assign n985 = n736 & ~n984;
  assign n986 = ~n981 & ~n985;
  assign n987 = n725 & ~n986;
  assign n988 = pi024 & n744;
  assign n989 = pi023 & ~n744;
  assign n990 = ~n988 & ~n989;
  assign n991 = ~n736 & ~n990;
  assign n992 = pi062 & n744;
  assign n993 = pi061 & n753;
  assign n994 = ~n992 & ~n993;
  assign n995 = n736 & ~n994;
  assign n996 = ~n991 & ~n995;
  assign n997 = ~n725 & ~n996;
  assign n998 = ~n987 & ~n997;
  assign n999 = ~n713 & ~n998;
  assign n1000 = pi021 & n744;
  assign n1001 = pi060 & n753;
  assign n1002 = ~n1000 & ~n1001;
  assign n1003 = ~n736 & ~n1002;
  assign n1004 = pi058 & n744;
  assign n1005 = pi020 & n753;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = n736 & ~n1006;
  assign n1008 = ~n1003 & ~n1007;
  assign n1009 = ~n725 & ~n1008;
  assign n1010 = pi057 & n744;
  assign n1011 = pi019 & ~n744;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~n736 & ~n1012;
  assign n1014 = pi028 & n744;
  assign n1015 = pi018 & ~n744;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = n736 & ~n1016;
  assign n1018 = ~n1013 & ~n1017;
  assign n1019 = n725 & ~n1018;
  assign n1020 = ~n1009 & ~n1019;
  assign n1021 = n797 & ~n1020;
  assign n1022 = ~n999 & ~n1021;
  assign n1023 = ~n699 & ~n1022;
  assign n1024 = pi065 & n744;
  assign n1025 = pi027 & ~n744;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n736 & ~n1026;
  assign n1028 = pi026 & n744;
  assign n1029 = pi025 & ~n744;
  assign n1030 = ~n1028 & ~n1029;
  assign n1031 = n736 & ~n1030;
  assign n1032 = ~n1027 & ~n1031;
  assign n1033 = n725 & ~n1032;
  assign n1034 = pi029 & ~n744;
  assign n1035 = pi066 & n744;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = n736 & ~n1036;
  assign n1038 = pi067 & ~n744;
  assign n1039 = pi030 & ~n753;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = ~n736 & ~n1040;
  assign n1042 = ~n1037 & ~n1041;
  assign n1043 = ~n725 & ~n1042;
  assign n1044 = ~n1033 & ~n1043;
  assign n1045 = n713 & ~n1044;
  assign n1046 = pi055 & n744;
  assign n1047 = pi054 & ~n744;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n736 & ~n1048;
  assign n1050 = pi052 & n744;
  assign n1051 = pi053 & ~n744;
  assign n1052 = ~n1050 & ~n1051;
  assign n1053 = n736 & ~n1052;
  assign n1054 = ~n1049 & ~n1053;
  assign n1055 = ~n725 & ~n1054;
  assign n1056 = pi059 & ~n753;
  assign n1057 = pi051 & ~n744;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = n736 & ~n1058;
  assign n1060 = pi049 & ~n744;
  assign n1061 = pi050 & n744;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~n736 & ~n1062;
  assign n1064 = ~n1059 & ~n1063;
  assign n1065 = n725 & ~n1064;
  assign n1066 = ~n1055 & ~n1065;
  assign n1067 = ~n713 & ~n1066;
  assign n1068 = ~n1045 & ~n1067;
  assign n1069 = n699 & ~n1068;
  assign n1070 = ~n1023 & ~n1069;
  assign n1071 = n676 & ~n1070;
  assign n1072 = pi068 & n744;
  assign n1073 = pi113 & n753;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = n736 & ~n1074;
  assign n1076 = pi114 & n744;
  assign n1077 = pi069 & ~n744;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~n736 & ~n1078;
  assign n1080 = ~n1075 & ~n1079;
  assign n1081 = ~n725 & ~n1080;
  assign n1082 = pi110 & n744;
  assign n1083 = pi099 & ~n744;
  assign n1084 = ~n1082 & ~n1083;
  assign n1085 = n736 & ~n1084;
  assign n1086 = pi070 & n744;
  assign n1087 = pi111 & ~n744;
  assign n1088 = ~n1086 & ~n1087;
  assign n1089 = ~n736 & ~n1088;
  assign n1090 = ~n1085 & ~n1089;
  assign n1091 = n725 & ~n1090;
  assign n1092 = ~n1081 & ~n1091;
  assign n1093 = n797 & ~n1092;
  assign n1094 = pi081 & n744;
  assign n1095 = pi080 & ~n744;
  assign n1096 = ~n1094 & ~n1095;
  assign n1097 = ~n736 & ~n1096;
  assign n1098 = pi079 & n744;
  assign n1099 = pi001 & ~n744;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = n736 & ~n1100;
  assign n1102 = ~n1097 & ~n1101;
  assign n1103 = n725 & ~n1102;
  assign n1104 = pi083 & ~n744;
  assign n1105 = pi002 & n744;
  assign n1106 = ~n1104 & ~n1105;
  assign n1107 = ~n736 & ~n1106;
  assign n1108 = pi098 & ~n744;
  assign n1109 = pi082 & ~n753;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = n736 & ~n1110;
  assign n1112 = ~n1107 & ~n1111;
  assign n1113 = ~n725 & ~n1112;
  assign n1114 = ~n1103 & ~n1113;
  assign n1115 = ~n713 & ~n1114;
  assign n1116 = ~n1093 & ~n1115;
  assign n1117 = n699 & ~n1116;
  assign n1118 = pi078 & n744;
  assign n1119 = pi077 & ~n744;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~n736 & ~n1120;
  assign n1122 = pi076 & n744;
  assign n1123 = pi112 & ~n744;
  assign n1124 = ~n1122 & ~n1123;
  assign n1125 = n736 & ~n1124;
  assign n1126 = ~n1121 & ~n1125;
  assign n1127 = ~n725 & ~n1126;
  assign n1128 = pi109 & ~n744;
  assign n1129 = pi075 & n744;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n736 & ~n1130;
  assign n1132 = pi100 & ~n753;
  assign n1133 = pi101 & ~n744;
  assign n1134 = ~n1132 & ~n1133;
  assign n1135 = n736 & ~n1134;
  assign n1136 = ~n1131 & ~n1135;
  assign n1137 = n725 & ~n1136;
  assign n1138 = ~n1127 & ~n1137;
  assign n1139 = ~n713 & ~n1138;
  assign n1140 = pi072 & ~n744;
  assign n1141 = pi073 & n744;
  assign n1142 = ~n1140 & ~n1141;
  assign n1143 = ~n736 & ~n1142;
  assign n1144 = pi003 & ~n744;
  assign n1145 = pi071 & n744;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = n736 & ~n1146;
  assign n1148 = ~n1143 & ~n1147;
  assign n1149 = n725 & ~n1148;
  assign n1150 = pi106 & n744;
  assign n1151 = pi074 & ~n744;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = n736 & ~n1152;
  assign n1154 = pi000 & n744;
  assign n1155 = pi107 & ~n744;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = ~n736 & ~n1156;
  assign n1158 = ~n1153 & ~n1157;
  assign n1159 = ~n725 & ~n1158;
  assign n1160 = ~n1149 & ~n1159;
  assign n1161 = n713 & ~n1160;
  assign n1162 = ~n1139 & ~n1161;
  assign n1163 = ~n699 & ~n1162;
  assign n1164 = ~n1117 & ~n1163;
  assign n1165 = ~n676 & ~n1164;
  assign n1166 = ~n1071 & ~n1165;
  assign n1167 = n974 & ~n1166;
  assign n1168 = ~n597 & n1167;
  assign n1169 = n977 & ~n1168;
  assign n1170 = ~n699 & n797;
  assign n1171 = n974 & n1170;
  assign n1172 = ~n676 & ~n725;
  assign n1173 = ~n736 & ~n753;
  assign n1174 = n1172 & n1173;
  assign n1175 = n1171 & n1174;
  assign n1176 = ~n1169 & n1175;
  assign n1177 = pi000 & ~n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n584 & ~n1178;
  assign n1180 = ~n585 & ~n1179;
  assign n1181 = ~n579 & ~n1180;
  assign n1182 = ~n580 & ~n1181;
  assign n1183 = ~n566 & ~n568;
  assign n1184 = ~n1182 & n1183;
  assign n1185 = ~n573 & ~n1184;
  assign n1186 = pi000 & n566;
  assign po047 = ~n1185 | n1186;
  assign n1188 = pi001 & ~pi273;
  assign n1189 = pi262 & pi273;
  assign n1190 = ~n1188 & ~n1189;
  assign n1191 = n569 & ~n1190;
  assign n1192 = pi001 & n579;
  assign n1193 = pi001 & n584;
  assign n1194 = n736 & n753;
  assign n1195 = ~n676 & ~n797;
  assign n1196 = n699 & n1195;
  assign n1197 = n725 & n974;
  assign n1198 = n1196 & n1197;
  assign n1199 = n1194 & n1198;
  assign n1200 = ~n1169 & n1199;
  assign n1201 = pi001 & ~n1199;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n584 & ~n1202;
  assign n1204 = ~n1193 & ~n1203;
  assign n1205 = ~n579 & ~n1204;
  assign n1206 = ~n1192 & ~n1205;
  assign n1207 = n1183 & ~n1206;
  assign n1208 = ~n1191 & ~n1207;
  assign n1209 = pi001 & n566;
  assign po048 = ~n1208 | n1209;
  assign n1211 = pi002 & n566;
  assign n1212 = pi002 & ~pi273;
  assign n1213 = pi269 & pi273;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = n569 & ~n1214;
  assign n1216 = pi002 & n579;
  assign n1217 = pi002 & n584;
  assign n1218 = ~n725 & n974;
  assign n1219 = n1196 & n1218;
  assign n1220 = n1173 & n1219;
  assign n1221 = pi002 & ~n1220;
  assign n1222 = ~n584 & n1221;
  assign n1223 = ~n1217 & ~n1222;
  assign n1224 = ~n1169 & n1220;
  assign n1225 = ~n584 & n1224;
  assign n1226 = n1223 & ~n1225;
  assign n1227 = ~n579 & ~n1226;
  assign n1228 = ~n1216 & ~n1227;
  assign n1229 = n1183 & ~n1228;
  assign n1230 = ~n1215 & ~n1229;
  assign po049 = n1211 | ~n1230;
  assign n1232 = pi003 & ~pi270;
  assign n1233 = pi238 & pi270;
  assign n1234 = ~n1232 & ~n1233;
  assign n1235 = n569 & ~n1234;
  assign n1236 = pi003 & n579;
  assign n1237 = pi003 & n584;
  assign n1238 = ~n676 & n725;
  assign n1239 = n1171 & n1238;
  assign n1240 = n1194 & n1239;
  assign n1241 = ~n1169 & n1240;
  assign n1242 = pi003 & ~n1240;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n584 & ~n1243;
  assign n1245 = ~n1237 & ~n1244;
  assign n1246 = ~n579 & ~n1245;
  assign n1247 = ~n1236 & ~n1246;
  assign n1248 = n1183 & ~n1247;
  assign n1249 = ~n1235 & ~n1248;
  assign n1250 = pi003 & n566;
  assign po050 = ~n1249 | n1250;
  assign n1252 = pi239 & pi270;
  assign n1253 = pi004 & ~pi270;
  assign n1254 = ~n1252 & ~n1253;
  assign n1255 = ~n568 & n579;
  assign n1256 = ~n1254 & n1255;
  assign n1257 = pi004 & n584;
  assign n1258 = n725 & n736;
  assign n1259 = ~n753 & n1170;
  assign n1260 = n1258 & n1259;
  assign n1261 = n676 & ~n974;
  assign n1262 = n1260 & n1261;
  assign n1263 = pi004 & ~n1262;
  assign n1264 = ~n1169 & n1262;
  assign n1265 = ~n1263 & ~n1264;
  assign n1266 = ~n584 & ~n1265;
  assign n1267 = ~n1257 & ~n1266;
  assign n1268 = ~n568 & ~n579;
  assign n1269 = ~n1267 & n1268;
  assign n1270 = ~n1256 & ~n1269;
  assign n1271 = ~n566 & ~n1270;
  assign n1272 = pi004 & ~n1183;
  assign po051 = n1271 | n1272;
  assign n1274 = pi240 & pi270;
  assign n1275 = pi005 & ~pi270;
  assign n1276 = ~n1274 & ~n1275;
  assign n1277 = n1255 & ~n1276;
  assign n1278 = pi005 & n584;
  assign n1279 = n725 & n753;
  assign n1280 = ~n736 & n1170;
  assign n1281 = n1279 & n1280;
  assign n1282 = n1261 & n1281;
  assign n1283 = ~n1169 & n1282;
  assign n1284 = pi005 & ~n1282;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~n584 & ~n1285;
  assign n1287 = ~n1278 & ~n1286;
  assign n1288 = n1268 & ~n1287;
  assign n1289 = ~n1277 & ~n1288;
  assign n1290 = ~n566 & ~n1289;
  assign n1291 = pi005 & ~n1183;
  assign po052 = n1290 | n1291;
  assign n1293 = pi242 & pi270;
  assign n1294 = pi006 & ~pi270;
  assign n1295 = ~n1293 & ~n1294;
  assign n1296 = n1255 & ~n1295;
  assign n1297 = pi006 & n584;
  assign n1298 = ~n725 & n1194;
  assign n1299 = n1170 & n1298;
  assign n1300 = n1261 & n1299;
  assign n1301 = ~n1169 & n1300;
  assign n1302 = pi006 & ~n1300;
  assign n1303 = ~n1301 & ~n1302;
  assign n1304 = ~n584 & ~n1303;
  assign n1305 = ~n1297 & ~n1304;
  assign n1306 = n1268 & ~n1305;
  assign n1307 = ~n1296 & ~n1306;
  assign n1308 = ~n566 & ~n1307;
  assign n1309 = pi006 & ~n1183;
  assign po053 = n1308 | n1309;
  assign n1311 = pi007 & ~pi270;
  assign n1312 = ~n571 & ~n1311;
  assign n1313 = n1255 & ~n1312;
  assign n1314 = pi007 & n584;
  assign n1315 = n676 & n1170;
  assign n1316 = ~n725 & ~n974;
  assign n1317 = n1315 & n1316;
  assign n1318 = n1173 & n1317;
  assign n1319 = ~n1169 & n1318;
  assign n1320 = pi007 & ~n1318;
  assign n1321 = ~n1319 & ~n1320;
  assign n1322 = ~n584 & ~n1321;
  assign n1323 = ~n1314 & ~n1322;
  assign n1324 = n1268 & ~n1323;
  assign n1325 = ~n1313 & ~n1324;
  assign n1326 = ~n566 & ~n1325;
  assign n1327 = pi007 & ~n1183;
  assign po054 = n1326 | n1327;
  assign n1329 = pi248 & pi271;
  assign n1330 = pi008 & ~pi271;
  assign n1331 = ~n1329 & ~n1330;
  assign n1332 = n1255 & ~n1331;
  assign n1333 = pi008 & n584;
  assign n1334 = n676 & ~n699;
  assign n1335 = n1279 & n1334;
  assign n1336 = ~n736 & n1335;
  assign n1337 = ~n797 & ~n974;
  assign n1338 = n1336 & n1337;
  assign n1339 = pi008 & ~n1338;
  assign n1340 = ~n1169 & n1338;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = ~n584 & ~n1341;
  assign n1343 = ~n1333 & ~n1342;
  assign n1344 = n1268 & ~n1343;
  assign n1345 = ~n1332 & ~n1344;
  assign n1346 = ~n566 & ~n1345;
  assign n1347 = pi008 & ~n1183;
  assign po055 = n1346 | n1347;
  assign n1349 = pi249 & pi271;
  assign n1350 = pi009 & ~pi271;
  assign n1351 = ~n1349 & ~n1350;
  assign n1352 = n1255 & ~n1351;
  assign n1353 = pi009 & n584;
  assign n1354 = n725 & n1337;
  assign n1355 = n1173 & n1354;
  assign n1356 = n1334 & n1355;
  assign n1357 = pi009 & ~n1356;
  assign n1358 = ~n1169 & n1356;
  assign n1359 = ~n1357 & ~n1358;
  assign n1360 = ~n584 & ~n1359;
  assign n1361 = ~n1353 & ~n1360;
  assign n1362 = n1268 & ~n1361;
  assign n1363 = ~n1352 & ~n1362;
  assign n1364 = ~n566 & ~n1363;
  assign n1365 = pi009 & ~n1183;
  assign po056 = n1364 | n1365;
  assign n1367 = pi250 & pi271;
  assign n1368 = pi010 & ~pi271;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = n1255 & ~n1369;
  assign n1371 = pi010 & n584;
  assign n1372 = n1194 & n1334;
  assign n1373 = ~n725 & n1372;
  assign n1374 = n1337 & n1373;
  assign n1375 = ~n1169 & n1374;
  assign n1376 = pi010 & ~n1374;
  assign n1377 = ~n1375 & ~n1376;
  assign n1378 = ~n584 & ~n1377;
  assign n1379 = ~n1371 & ~n1378;
  assign n1380 = n1268 & ~n1379;
  assign n1381 = ~n1370 & ~n1380;
  assign n1382 = ~n566 & ~n1381;
  assign n1383 = pi010 & ~n1183;
  assign po057 = n1382 | n1383;
  assign n1385 = pi259 & pi272;
  assign n1386 = pi011 & ~pi272;
  assign n1387 = ~n1385 & ~n1386;
  assign n1388 = n1255 & ~n1387;
  assign n1389 = pi011 & n584;
  assign n1390 = n676 & n797;
  assign n1391 = ~n725 & ~n753;
  assign n1392 = n699 & ~n974;
  assign n1393 = n736 & n1392;
  assign n1394 = n1391 & n1393;
  assign n1395 = n1390 & n1394;
  assign n1396 = ~n1169 & n1395;
  assign n1397 = pi011 & ~n1395;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n584 & ~n1398;
  assign n1400 = ~n1389 & ~n1399;
  assign n1401 = n1268 & ~n1400;
  assign n1402 = ~n1388 & ~n1401;
  assign n1403 = ~n566 & ~n1402;
  assign n1404 = pi011 & ~n1183;
  assign po058 = n1403 | n1404;
  assign n1406 = pi260 & pi272;
  assign n1407 = pi012 & ~pi272;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = n1255 & ~n1408;
  assign n1410 = pi012 & n584;
  assign n1411 = ~n725 & ~n736;
  assign n1412 = n753 & n1392;
  assign n1413 = n1411 & n1412;
  assign n1414 = n1390 & n1413;
  assign n1415 = pi012 & ~n1414;
  assign n1416 = ~n1169 & n1414;
  assign n1417 = ~n1415 & ~n1416;
  assign n1418 = ~n584 & ~n1417;
  assign n1419 = ~n1410 & ~n1418;
  assign n1420 = n1268 & ~n1419;
  assign n1421 = ~n1409 & ~n1420;
  assign n1422 = ~n566 & ~n1421;
  assign n1423 = pi012 & ~n1183;
  assign po059 = n1422 | n1423;
  assign n1425 = pi261 & pi272;
  assign n1426 = pi013 & ~pi272;
  assign n1427 = ~n1425 & ~n1426;
  assign n1428 = n1255 & ~n1427;
  assign n1429 = pi013 & n584;
  assign n1430 = n699 & ~n725;
  assign n1431 = n1173 & n1430;
  assign n1432 = ~n974 & n1390;
  assign n1433 = n1431 & n1432;
  assign n1434 = ~n1169 & n1433;
  assign n1435 = pi013 & ~n1433;
  assign n1436 = ~n1434 & ~n1435;
  assign n1437 = ~n584 & ~n1436;
  assign n1438 = ~n1429 & ~n1437;
  assign n1439 = n1268 & ~n1438;
  assign n1440 = ~n1428 & ~n1439;
  assign n1441 = ~n566 & ~n1440;
  assign n1442 = pi013 & ~n1183;
  assign po060 = n1441 | n1442;
  assign n1444 = pi265 & pi273;
  assign n1445 = pi014 & ~pi273;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = n1255 & ~n1446;
  assign n1448 = pi014 & n584;
  assign n1449 = n699 & ~n797;
  assign n1450 = n725 & n1449;
  assign n1451 = n1173 & n1450;
  assign n1452 = n1261 & n1451;
  assign n1453 = ~n1169 & n1452;
  assign n1454 = pi014 & ~n1452;
  assign n1455 = ~n1453 & ~n1454;
  assign n1456 = ~n584 & ~n1455;
  assign n1457 = ~n1448 & ~n1456;
  assign n1458 = n1268 & ~n1457;
  assign n1459 = ~n1447 & ~n1458;
  assign n1460 = ~n566 & ~n1459;
  assign n1461 = pi014 & ~n1183;
  assign po061 = n1460 | n1461;
  assign n1463 = pi267 & pi273;
  assign n1464 = pi015 & ~pi273;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = n1255 & ~n1465;
  assign n1467 = pi015 & n584;
  assign n1468 = n736 & n1391;
  assign n1469 = n1449 & n1468;
  assign n1470 = n1261 & n1469;
  assign n1471 = ~n1169 & n1470;
  assign n1472 = pi015 & ~n1470;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = ~n584 & ~n1473;
  assign n1475 = ~n1467 & ~n1474;
  assign n1476 = n1268 & ~n1475;
  assign n1477 = ~n1466 & ~n1476;
  assign n1478 = ~n566 & ~n1477;
  assign n1479 = pi015 & ~n1183;
  assign po062 = n1478 | n1479;
  assign n1481 = pi268 & pi273;
  assign n1482 = pi016 & ~pi273;
  assign n1483 = ~n1481 & ~n1482;
  assign n1484 = n1255 & ~n1483;
  assign n1485 = pi016 & n584;
  assign n1486 = n753 & n1449;
  assign n1487 = n1411 & n1486;
  assign n1488 = n1261 & n1487;
  assign n1489 = pi016 & ~n1488;
  assign n1490 = ~n1169 & n1488;
  assign n1491 = ~n1489 & ~n1490;
  assign n1492 = ~n584 & ~n1491;
  assign n1493 = ~n1485 & ~n1492;
  assign n1494 = n1268 & ~n1493;
  assign n1495 = ~n1484 & ~n1494;
  assign n1496 = ~n566 & ~n1495;
  assign n1497 = pi016 & ~n1183;
  assign po063 = n1496 | n1497;
  assign n1499 = pi017 & ~pi273;
  assign n1500 = ~n1213 & ~n1499;
  assign n1501 = n1255 & ~n1500;
  assign n1502 = pi017 & n584;
  assign n1503 = n699 & n1337;
  assign n1504 = n676 & ~n725;
  assign n1505 = n1503 & n1504;
  assign n1506 = n1173 & n1505;
  assign n1507 = pi017 & ~n1506;
  assign n1508 = ~n1169 & n1506;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n584 & ~n1509;
  assign n1511 = ~n1502 & ~n1510;
  assign n1512 = n1268 & ~n1511;
  assign n1513 = ~n1501 & ~n1512;
  assign n1514 = ~n566 & ~n1513;
  assign n1515 = pi017 & ~n1183;
  assign po064 = n1514 | n1515;
  assign n1517 = n974 & n1334;
  assign n1518 = n725 & n797;
  assign n1519 = n1194 & n1518;
  assign n1520 = n1517 & n1519;
  assign n1521 = ~n1169 & n1520;
  assign n1522 = pi018 & ~n1520;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n584 & n1523;
  assign n1525 = ~pi018 & n584;
  assign n1526 = ~n1524 & ~n1525;
  assign n1527 = n1268 & n1526;
  assign n1528 = pi018 & ~n1268;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n566 & ~n1529;
  assign n1531 = pi018 & ~pi270;
  assign n1532 = ~n1233 & ~n1531;
  assign n1533 = n566 & ~n1532;
  assign po065 = n1530 | n1533;
  assign n1535 = ~n736 & n753;
  assign n1536 = n1518 & n1535;
  assign n1537 = n1517 & n1536;
  assign n1538 = ~n1169 & n1537;
  assign n1539 = pi019 & ~n1537;
  assign n1540 = ~n1538 & ~n1539;
  assign n1541 = ~n584 & n1540;
  assign n1542 = ~pi019 & n584;
  assign n1543 = ~n1541 & ~n1542;
  assign n1544 = n1268 & n1543;
  assign n1545 = pi019 & ~n1268;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~n566 & ~n1546;
  assign n1548 = pi019 & ~pi270;
  assign n1549 = ~n1274 & ~n1548;
  assign n1550 = n566 & ~n1549;
  assign po066 = n1547 | n1550;
  assign n1552 = ~n725 & n797;
  assign n1553 = n1194 & n1552;
  assign n1554 = n1517 & n1553;
  assign n1555 = ~n1169 & n1554;
  assign n1556 = pi020 & ~n1554;
  assign n1557 = ~n1555 & ~n1556;
  assign n1558 = ~n584 & n1557;
  assign n1559 = ~pi020 & n584;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = n1268 & n1560;
  assign n1562 = pi020 & ~n1268;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = ~n566 & ~n1563;
  assign n1565 = pi020 & ~pi270;
  assign n1566 = ~n1293 & ~n1565;
  assign n1567 = n566 & ~n1566;
  assign po067 = n1564 | n1567;
  assign n1569 = pi021 & ~pi270;
  assign n1570 = ~n571 & ~n1569;
  assign n1571 = n566 & ~n1570;
  assign n1572 = pi021 & n568;
  assign n1573 = ~n579 & ~n584;
  assign n1574 = pi021 & ~n1573;
  assign n1575 = ~n736 & n1517;
  assign n1576 = n1552 & n1575;
  assign n1577 = ~n753 & n1576;
  assign n1578 = n1169 & n1577;
  assign n1579 = ~pi021 & ~n1577;
  assign n1580 = n1573 & ~n1579;
  assign n1581 = ~n1578 & n1580;
  assign n1582 = ~n1574 & ~n1581;
  assign n1583 = ~n568 & ~n1582;
  assign n1584 = ~n1572 & ~n1583;
  assign n1585 = ~n566 & ~n1584;
  assign po068 = n1571 | n1585;
  assign n1587 = n725 & ~n797;
  assign n1588 = n1194 & n1587;
  assign n1589 = n1517 & n1588;
  assign n1590 = ~n1169 & n1589;
  assign n1591 = pi022 & ~n1589;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~n584 & n1592;
  assign n1594 = ~pi022 & n584;
  assign n1595 = ~n1593 & ~n1594;
  assign n1596 = n1268 & n1595;
  assign n1597 = pi022 & ~n1268;
  assign n1598 = ~n1596 & ~n1597;
  assign n1599 = ~n566 & ~n1598;
  assign n1600 = pi246 & pi271;
  assign n1601 = pi022 & ~pi271;
  assign n1602 = ~n1600 & ~n1601;
  assign n1603 = n566 & ~n1602;
  assign po069 = n1599 | n1603;
  assign n1605 = pi252 & pi271;
  assign n1606 = pi023 & ~pi271;
  assign n1607 = ~n1605 & ~n1606;
  assign n1608 = n566 & ~n1607;
  assign n1609 = pi023 & n568;
  assign n1610 = pi023 & ~n1573;
  assign n1611 = ~n725 & ~n797;
  assign n1612 = n753 & n1611;
  assign n1613 = n1575 & n1612;
  assign n1614 = n1169 & n1613;
  assign n1615 = ~pi023 & ~n1613;
  assign n1616 = n1573 & ~n1615;
  assign n1617 = ~n1614 & n1616;
  assign n1618 = ~n1610 & ~n1617;
  assign n1619 = ~n568 & ~n1618;
  assign n1620 = ~n1609 & ~n1619;
  assign n1621 = ~n566 & ~n1620;
  assign po070 = n1608 | n1621;
  assign n1623 = n1173 & n1611;
  assign n1624 = n1517 & n1623;
  assign n1625 = ~n1169 & n1624;
  assign n1626 = pi024 & ~n1624;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n584 & n1627;
  assign n1629 = ~pi024 & n584;
  assign n1630 = ~n1628 & ~n1629;
  assign n1631 = n1268 & n1630;
  assign n1632 = pi024 & ~n1268;
  assign n1633 = ~n1631 & ~n1632;
  assign n1634 = ~n566 & ~n1633;
  assign n1635 = pi253 & pi271;
  assign n1636 = pi024 & ~pi271;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = n566 & ~n1637;
  assign po071 = n1634 | n1638;
  assign n1640 = n699 & n725;
  assign n1641 = n676 & n974;
  assign n1642 = n797 & n1641;
  assign n1643 = n1640 & n1642;
  assign n1644 = n1194 & n1643;
  assign n1645 = ~n1169 & n1644;
  assign n1646 = pi025 & ~n1644;
  assign n1647 = ~n1645 & ~n1646;
  assign n1648 = ~n584 & n1647;
  assign n1649 = ~pi025 & n584;
  assign n1650 = ~n1648 & ~n1649;
  assign n1651 = n1268 & n1650;
  assign n1652 = pi025 & ~n1268;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~n566 & ~n1653;
  assign n1655 = pi254 & pi272;
  assign n1656 = pi025 & ~pi272;
  assign n1657 = ~n1655 & ~n1656;
  assign n1658 = n566 & ~n1657;
  assign po072 = n1654 | n1658;
  assign n1660 = pi255 & pi272;
  assign n1661 = pi026 & ~pi272;
  assign n1662 = ~n1660 & ~n1661;
  assign n1663 = n566 & ~n1662;
  assign n1664 = pi026 & n568;
  assign n1665 = pi026 & ~n1573;
  assign n1666 = n1258 & n1390;
  assign n1667 = ~n753 & n1666;
  assign n1668 = n699 & n974;
  assign n1669 = n1667 & n1668;
  assign n1670 = n1169 & n1669;
  assign n1671 = ~pi026 & ~n1669;
  assign n1672 = n1573 & ~n1671;
  assign n1673 = ~n1670 & n1672;
  assign n1674 = ~n1665 & ~n1673;
  assign n1675 = ~n568 & ~n1674;
  assign n1676 = ~n1664 & ~n1675;
  assign n1677 = ~n566 & ~n1676;
  assign po073 = n1663 | n1677;
  assign n1679 = pi256 & pi272;
  assign n1680 = pi027 & ~pi272;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = n566 & ~n1681;
  assign n1683 = pi027 & n568;
  assign n1684 = pi027 & ~n1573;
  assign n1685 = n1279 & n1390;
  assign n1686 = ~n736 & n1685;
  assign n1687 = n1668 & n1686;
  assign n1688 = n1169 & n1687;
  assign n1689 = ~pi027 & ~n1687;
  assign n1690 = n1573 & ~n1689;
  assign n1691 = ~n1688 & n1690;
  assign n1692 = ~n1684 & ~n1691;
  assign n1693 = ~n568 & ~n1692;
  assign n1694 = ~n1683 & ~n1693;
  assign n1695 = ~n566 & ~n1694;
  assign po074 = n1682 | n1695;
  assign n1697 = n736 & ~n753;
  assign n1698 = n1518 & n1697;
  assign n1699 = n1517 & n1698;
  assign n1700 = ~n1169 & n1699;
  assign n1701 = pi028 & ~n1699;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n584 & n1702;
  assign n1704 = ~pi028 & n584;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = n1268 & n1705;
  assign n1707 = pi028 & ~n1268;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = ~n566 & ~n1708;
  assign n1710 = pi028 & ~pi270;
  assign n1711 = ~n1252 & ~n1710;
  assign n1712 = n566 & ~n1711;
  assign po075 = n1709 | n1712;
  assign n1714 = pi258 & pi272;
  assign n1715 = pi029 & ~pi272;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = n566 & ~n1716;
  assign n1718 = pi029 & n568;
  assign n1719 = pi029 & ~n1573;
  assign n1720 = n1194 & n1390;
  assign n1721 = ~n725 & n1720;
  assign n1722 = n1668 & n1721;
  assign n1723 = n1169 & n1722;
  assign n1724 = ~pi029 & ~n1722;
  assign n1725 = n1573 & ~n1724;
  assign n1726 = ~n1723 & n1725;
  assign n1727 = ~n1719 & ~n1726;
  assign n1728 = ~n568 & ~n1727;
  assign n1729 = ~n1718 & ~n1728;
  assign n1730 = ~n566 & ~n1729;
  assign po076 = n1717 | n1730;
  assign n1732 = n1431 & n1642;
  assign n1733 = ~n1169 & n1732;
  assign n1734 = pi030 & ~n1732;
  assign n1735 = ~n1733 & ~n1734;
  assign n1736 = ~n584 & n1735;
  assign n1737 = ~pi030 & n584;
  assign n1738 = ~n1736 & ~n1737;
  assign n1739 = n1268 & n1738;
  assign n1740 = pi030 & ~n1268;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n566 & ~n1741;
  assign n1743 = pi030 & ~pi272;
  assign n1744 = ~n1425 & ~n1743;
  assign n1745 = n566 & ~n1744;
  assign po077 = n1742 | n1745;
  assign n1747 = pi266 & pi273;
  assign n1748 = pi031 & ~pi273;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = n1255 & ~n1749;
  assign n1751 = pi031 & n584;
  assign n1752 = n736 & n1503;
  assign n1753 = n753 & n1752;
  assign n1754 = n1504 & n1753;
  assign n1755 = ~n1169 & n1754;
  assign n1756 = pi031 & ~n1754;
  assign n1757 = ~n1755 & ~n1756;
  assign n1758 = ~n584 & ~n1757;
  assign n1759 = ~n1751 & ~n1758;
  assign n1760 = n1268 & ~n1759;
  assign n1761 = ~n1750 & ~n1760;
  assign n1762 = ~n566 & ~n1761;
  assign n1763 = pi031 & ~n1183;
  assign po078 = n1762 | n1763;
  assign n1765 = pi032 & ~n1183;
  assign n1766 = pi263 & pi273;
  assign n1767 = pi032 & ~pi273;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = n1255 & ~n1768;
  assign n1770 = pi032 & n584;
  assign n1771 = n676 & n725;
  assign n1772 = n1752 & n1771;
  assign n1773 = ~n753 & n1772;
  assign n1774 = pi032 & ~n1773;
  assign n1775 = ~n1169 & n1773;
  assign n1776 = ~n1774 & ~n1775;
  assign n1777 = ~n584 & ~n1776;
  assign n1778 = ~n1770 & ~n1777;
  assign n1779 = n1268 & ~n1778;
  assign n1780 = ~n1769 & ~n1779;
  assign n1781 = ~n566 & ~n1780;
  assign po079 = n1765 | n1781;
  assign n1783 = pi033 & ~pi270;
  assign n1784 = ~n1233 & ~n1783;
  assign n1785 = n1255 & ~n1784;
  assign n1786 = pi033 & n584;
  assign n1787 = n725 & ~n974;
  assign n1788 = n1315 & n1787;
  assign n1789 = n1194 & n1788;
  assign n1790 = ~n1169 & n1789;
  assign n1791 = pi033 & ~n1789;
  assign n1792 = ~n1790 & ~n1791;
  assign n1793 = ~n584 & ~n1792;
  assign n1794 = ~n1786 & ~n1793;
  assign n1795 = n1268 & ~n1794;
  assign n1796 = ~n1785 & ~n1795;
  assign n1797 = ~n566 & ~n1796;
  assign n1798 = pi033 & ~n1183;
  assign po080 = n1797 | n1798;
  assign n1800 = pi241 & pi270;
  assign n1801 = pi034 & ~pi270;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = n1255 & ~n1802;
  assign n1804 = pi034 & n584;
  assign n1805 = ~n736 & n1315;
  assign n1806 = n725 & n1805;
  assign n1807 = ~n974 & n1806;
  assign n1808 = ~n753 & n1807;
  assign n1809 = ~n1169 & n1808;
  assign n1810 = pi034 & ~n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = ~n584 & ~n1811;
  assign n1813 = ~n1804 & ~n1812;
  assign n1814 = n1268 & ~n1813;
  assign n1815 = ~n1803 & ~n1814;
  assign n1816 = ~n566 & ~n1815;
  assign n1817 = pi034 & ~n1183;
  assign po081 = n1816 | n1817;
  assign n1819 = pi243 & pi270;
  assign n1820 = pi035 & ~pi270;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = n1255 & ~n1821;
  assign n1823 = pi035 & n584;
  assign n1824 = n736 & n1315;
  assign n1825 = ~n753 & n1824;
  assign n1826 = n1316 & n1825;
  assign n1827 = ~n1169 & n1826;
  assign n1828 = pi035 & ~n1826;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~n584 & ~n1829;
  assign n1831 = ~n1823 & ~n1830;
  assign n1832 = n1268 & ~n1831;
  assign n1833 = ~n1822 & ~n1832;
  assign n1834 = ~n566 & ~n1833;
  assign n1835 = pi035 & ~n1183;
  assign po082 = n1834 | n1835;
  assign n1837 = pi036 & ~n1183;
  assign n1838 = pi244 & pi270;
  assign n1839 = pi036 & ~pi270;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = n1255 & ~n1840;
  assign n1842 = pi036 & n584;
  assign n1843 = n753 & n1805;
  assign n1844 = ~n1169 & n1316;
  assign n1845 = n1843 & n1844;
  assign n1846 = ~n584 & n1845;
  assign n1847 = n1316 & n1843;
  assign n1848 = ~n584 & ~n1847;
  assign n1849 = pi036 & n1848;
  assign n1850 = ~n1846 & ~n1849;
  assign n1851 = ~n1842 & n1850;
  assign n1852 = n1268 & ~n1851;
  assign n1853 = ~n1841 & ~n1852;
  assign n1854 = ~n566 & ~n1853;
  assign po083 = n1837 | n1854;
  assign n1856 = pi037 & ~pi271;
  assign n1857 = ~n1600 & ~n1856;
  assign n1858 = n1255 & ~n1857;
  assign n1859 = pi037 & n584;
  assign n1860 = ~n699 & n725;
  assign n1861 = n1194 & n1860;
  assign n1862 = ~n797 & n1261;
  assign n1863 = n1861 & n1862;
  assign n1864 = ~n1169 & n1863;
  assign n1865 = pi037 & ~n1863;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = ~n584 & ~n1866;
  assign n1868 = ~n1859 & ~n1867;
  assign n1869 = n1268 & ~n1868;
  assign n1870 = ~n1858 & ~n1869;
  assign n1871 = ~n566 & ~n1870;
  assign n1872 = pi037 & ~n1183;
  assign po084 = n1871 | n1872;
  assign n1874 = pi247 & pi271;
  assign n1875 = pi038 & ~pi271;
  assign n1876 = ~n1874 & ~n1875;
  assign n1877 = n1255 & ~n1876;
  assign n1878 = pi038 & n584;
  assign n1879 = n1258 & n1334;
  assign n1880 = ~n753 & n1879;
  assign n1881 = n1337 & n1880;
  assign n1882 = ~n1169 & n1881;
  assign n1883 = pi038 & ~n1881;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = ~n584 & ~n1884;
  assign n1886 = ~n1878 & ~n1885;
  assign n1887 = n1268 & ~n1886;
  assign n1888 = ~n1877 & ~n1887;
  assign n1889 = ~n566 & ~n1888;
  assign n1890 = pi038 & ~n1183;
  assign po085 = n1889 | n1890;
  assign n1892 = pi251 & pi271;
  assign n1893 = pi039 & ~pi271;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = n1255 & ~n1894;
  assign n1896 = pi039 & n584;
  assign n1897 = n1334 & n1337;
  assign n1898 = n1468 & n1897;
  assign n1899 = ~n1169 & n1898;
  assign n1900 = pi039 & ~n1898;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = ~n584 & ~n1901;
  assign n1903 = ~n1896 & ~n1902;
  assign n1904 = n1268 & ~n1903;
  assign n1905 = ~n1895 & ~n1904;
  assign n1906 = ~n566 & ~n1905;
  assign n1907 = pi039 & ~n1183;
  assign po086 = n1906 | n1907;
  assign n1909 = pi040 & ~pi272;
  assign n1910 = ~n1655 & ~n1909;
  assign n1911 = n1255 & ~n1910;
  assign n1912 = pi040 & n584;
  assign n1913 = n676 & n699;
  assign n1914 = ~n974 & n1519;
  assign n1915 = n1913 & n1914;
  assign n1916 = ~n1169 & n1915;
  assign n1917 = pi040 & ~n1915;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = ~n584 & ~n1918;
  assign n1920 = ~n1912 & ~n1919;
  assign n1921 = n1268 & ~n1920;
  assign n1922 = ~n1911 & ~n1921;
  assign n1923 = ~n566 & ~n1922;
  assign n1924 = pi040 & ~n1183;
  assign po087 = n1923 | n1924;
  assign n1926 = pi257 & pi272;
  assign n1927 = pi041 & ~pi272;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = n1255 & ~n1928;
  assign n1930 = pi041 & n584;
  assign n1931 = n725 & n1392;
  assign n1932 = n1173 & n1931;
  assign n1933 = n1390 & n1932;
  assign n1934 = ~n1169 & n1933;
  assign n1935 = pi041 & ~n1933;
  assign n1936 = ~n1934 & ~n1935;
  assign n1937 = ~n584 & ~n1936;
  assign n1938 = ~n1930 & ~n1937;
  assign n1939 = n1268 & ~n1938;
  assign n1940 = ~n1929 & ~n1939;
  assign n1941 = ~n566 & ~n1940;
  assign n1942 = pi041 & ~n1183;
  assign po088 = n1941 | n1942;
  assign n1944 = pi042 & ~pi272;
  assign n1945 = ~n1714 & ~n1944;
  assign n1946 = n1255 & ~n1945;
  assign n1947 = pi042 & n584;
  assign n1948 = n1392 & n1721;
  assign n1949 = ~n1169 & n1948;
  assign n1950 = pi042 & ~n1948;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = ~n584 & ~n1951;
  assign n1953 = ~n1947 & ~n1952;
  assign n1954 = n1268 & ~n1953;
  assign n1955 = ~n1946 & ~n1954;
  assign n1956 = ~n566 & ~n1955;
  assign n1957 = pi042 & ~n1183;
  assign po089 = n1956 | n1957;
  assign n1959 = pi043 & ~pi272;
  assign n1960 = ~n1660 & ~n1959;
  assign n1961 = n1255 & ~n1960;
  assign n1962 = pi043 & n584;
  assign n1963 = n1392 & n1667;
  assign n1964 = ~n1169 & n1963;
  assign n1965 = pi043 & ~n1963;
  assign n1966 = ~n1964 & ~n1965;
  assign n1967 = ~n584 & ~n1966;
  assign n1968 = ~n1962 & ~n1967;
  assign n1969 = n1268 & ~n1968;
  assign n1970 = ~n1961 & ~n1969;
  assign n1971 = ~n566 & ~n1970;
  assign n1972 = pi043 & ~n1183;
  assign po090 = n1971 | n1972;
  assign n1974 = pi044 & ~pi273;
  assign n1975 = ~n1189 & ~n1974;
  assign n1976 = n1255 & ~n1975;
  assign n1977 = pi044 & n584;
  assign n1978 = n1194 & n1771;
  assign n1979 = n1503 & n1978;
  assign n1980 = ~n1169 & n1979;
  assign n1981 = pi044 & ~n1979;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = ~n584 & ~n1982;
  assign n1984 = ~n1977 & ~n1983;
  assign n1985 = n1268 & ~n1984;
  assign n1986 = ~n1976 & ~n1985;
  assign n1987 = ~n566 & ~n1986;
  assign n1988 = pi044 & ~n1183;
  assign po091 = n1987 | n1988;
  assign n1990 = pi045 & ~n1183;
  assign n1991 = pi045 & ~pi272;
  assign n1992 = ~n1679 & ~n1991;
  assign n1993 = n1255 & ~n1992;
  assign n1994 = pi045 & n584;
  assign n1995 = n1392 & n1686;
  assign n1996 = pi045 & ~n1995;
  assign n1997 = ~n1169 & n1995;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = ~n584 & ~n1998;
  assign n2000 = ~n1994 & ~n1999;
  assign n2001 = n1268 & ~n2000;
  assign n2002 = ~n1993 & ~n2001;
  assign n2003 = ~n566 & ~n2002;
  assign po092 = n1990 | n2003;
  assign n2005 = pi264 & pi273;
  assign n2006 = pi046 & ~pi273;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = n1255 & ~n2007;
  assign n2009 = pi046 & n584;
  assign n2010 = n1535 & n1771;
  assign n2011 = n1503 & n2010;
  assign n2012 = ~n1169 & n2011;
  assign n2013 = pi046 & ~n2011;
  assign n2014 = ~n2012 & ~n2013;
  assign n2015 = ~n584 & ~n2014;
  assign n2016 = ~n2009 & ~n2015;
  assign n2017 = n1268 & ~n2016;
  assign n2018 = ~n2008 & ~n2017;
  assign n2019 = ~n566 & ~n2018;
  assign n2020 = pi046 & ~n1183;
  assign po093 = n2019 | n2020;
  assign n2022 = pi047 & ~pi271;
  assign n2023 = ~n1635 & ~n2022;
  assign n2024 = n1255 & ~n2023;
  assign n2025 = pi047 & n584;
  assign n2026 = ~n974 & n1334;
  assign n2027 = n1623 & n2026;
  assign n2028 = ~n1169 & n2027;
  assign n2029 = pi047 & ~n2027;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = ~n584 & ~n2030;
  assign n2032 = ~n2025 & ~n2031;
  assign n2033 = n1268 & ~n2032;
  assign n2034 = ~n2024 & ~n2033;
  assign n2035 = ~n566 & ~n2034;
  assign n2036 = pi047 & ~n1183;
  assign po094 = n2035 | n2036;
  assign n2038 = pi048 & ~pi271;
  assign n2039 = ~n1605 & ~n2038;
  assign n2040 = n1255 & ~n2039;
  assign n2041 = pi048 & n584;
  assign n2042 = n753 & n1411;
  assign n2043 = n1897 & n2042;
  assign n2044 = ~n1169 & n2043;
  assign n2045 = pi048 & ~n2043;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~n584 & ~n2046;
  assign n2048 = ~n2041 & ~n2047;
  assign n2049 = n1268 & ~n2048;
  assign n2050 = ~n2040 & ~n2049;
  assign n2051 = ~n566 & ~n2050;
  assign n2052 = pi048 & ~n1183;
  assign po095 = n2051 | n2052;
  assign n2054 = pi049 & ~pi273;
  assign n2055 = ~n2005 & ~n2054;
  assign n2056 = n566 & ~n2055;
  assign n2057 = pi049 & n568;
  assign n2058 = pi049 & ~n1573;
  assign n2059 = ~n736 & n1641;
  assign n2060 = n1279 & n2059;
  assign n2061 = n1449 & n2060;
  assign n2062 = n1169 & n2061;
  assign n2063 = ~pi049 & ~n2061;
  assign n2064 = n1573 & ~n2063;
  assign n2065 = ~n2062 & n2064;
  assign n2066 = ~n2058 & ~n2065;
  assign n2067 = ~n568 & ~n2066;
  assign n2068 = ~n2057 & ~n2067;
  assign n2069 = ~n566 & ~n2068;
  assign po096 = n2056 | n2069;
  assign n2071 = pi050 & ~pi273;
  assign n2072 = ~n1444 & ~n2071;
  assign n2073 = n566 & ~n2072;
  assign n2074 = pi050 & ~n1573;
  assign n2075 = n1451 & n1641;
  assign n2076 = n1169 & n2075;
  assign n2077 = ~pi050 & ~n2075;
  assign n2078 = n1573 & ~n2077;
  assign n2079 = ~n2076 & n2078;
  assign n2080 = ~n2074 & ~n2079;
  assign n2081 = ~n568 & ~n2080;
  assign n2082 = pi050 & n568;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n566 & ~n2083;
  assign po097 = n2073 | n2084;
  assign n2086 = pi051 & ~pi273;
  assign n2087 = ~n1189 & ~n2086;
  assign n2088 = n566 & ~n2087;
  assign n2089 = pi051 & ~n1573;
  assign n2090 = n974 & n1978;
  assign n2091 = n1449 & n2090;
  assign n2092 = n1169 & n2091;
  assign n2093 = ~pi051 & ~n2091;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = n1573 & n2094;
  assign n2096 = ~n2089 & ~n2095;
  assign n2097 = ~n568 & ~n2096;
  assign n2098 = pi051 & n568;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = ~n566 & ~n2099;
  assign po098 = n2088 | n2100;
  assign n2102 = pi052 & ~pi273;
  assign n2103 = ~n1463 & ~n2102;
  assign n2104 = n566 & ~n2103;
  assign n2105 = pi052 & n568;
  assign n2106 = pi052 & ~n1573;
  assign n2107 = n1469 & n1641;
  assign n2108 = n1169 & n2107;
  assign n2109 = ~pi052 & ~n2107;
  assign n2110 = n1573 & ~n2109;
  assign n2111 = ~n2108 & n2110;
  assign n2112 = ~n2106 & ~n2111;
  assign n2113 = ~n568 & ~n2112;
  assign n2114 = ~n2105 & ~n2113;
  assign n2115 = ~n566 & ~n2114;
  assign po099 = n2104 | n2115;
  assign n2117 = pi053 & ~pi273;
  assign n2118 = ~n1747 & ~n2117;
  assign n2119 = n566 & ~n2118;
  assign n2120 = pi053 & n568;
  assign n2121 = pi053 & ~n1573;
  assign n2122 = ~n725 & n1641;
  assign n2123 = n1194 & n1449;
  assign n2124 = n2122 & n2123;
  assign n2125 = n1169 & n2124;
  assign n2126 = ~pi053 & ~n2124;
  assign n2127 = n1573 & ~n2126;
  assign n2128 = ~n2125 & n2127;
  assign n2129 = ~n2121 & ~n2128;
  assign n2130 = ~n568 & ~n2129;
  assign n2131 = ~n2120 & ~n2130;
  assign n2132 = ~n566 & ~n2131;
  assign po100 = n2119 | n2132;
  assign n2134 = pi054 & ~pi273;
  assign n2135 = ~n1481 & ~n2134;
  assign n2136 = n566 & ~n2135;
  assign n2137 = pi054 & ~n1573;
  assign n2138 = n1487 & n1641;
  assign n2139 = n1169 & n2138;
  assign n2140 = ~pi054 & ~n2138;
  assign n2141 = n1573 & ~n2140;
  assign n2142 = ~n2139 & n2141;
  assign n2143 = ~n2137 & ~n2142;
  assign n2144 = ~n568 & ~n2143;
  assign n2145 = pi054 & n568;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = ~n566 & ~n2146;
  assign po101 = n2136 | n2147;
  assign n2149 = pi055 & ~pi273;
  assign n2150 = ~n1213 & ~n2149;
  assign n2151 = n566 & ~n2150;
  assign n2152 = pi055 & ~n1573;
  assign n2153 = n974 & n1623;
  assign n2154 = n1913 & n2153;
  assign n2155 = n1169 & n2154;
  assign n2156 = ~pi055 & ~n2154;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = n1573 & n2157;
  assign n2159 = ~n2152 & ~n2158;
  assign n2160 = ~n568 & ~n2159;
  assign n2161 = pi055 & n568;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = ~n566 & ~n2162;
  assign po102 = n2151 | n2163;
  assign n2165 = pi056 & ~pi271;
  assign n2166 = ~n1329 & ~n2165;
  assign n2167 = n566 & ~n2166;
  assign n2168 = pi056 & n568;
  assign n2169 = n568 & ~n2168;
  assign n2170 = ~n566 & ~n2169;
  assign n2171 = ~n797 & n974;
  assign n2172 = n1336 & n2171;
  assign n2173 = ~pi056 & ~n2172;
  assign n2174 = n1169 & n2172;
  assign n2175 = ~n2173 & ~n2174;
  assign n2176 = n1573 & n2175;
  assign n2177 = ~n568 & n1573;
  assign n2178 = pi056 & ~n2177;
  assign n2179 = ~n2176 & ~n2178;
  assign n2180 = n2170 & ~n2179;
  assign po103 = n2167 | n2180;
  assign n2182 = pi057 & ~pi270;
  assign n2183 = ~n1800 & ~n2182;
  assign n2184 = n566 & ~n2183;
  assign n2185 = pi057 & ~n1573;
  assign n2186 = n974 & n1806;
  assign n2187 = ~n753 & n2186;
  assign n2188 = n1169 & n2187;
  assign n2189 = ~pi057 & ~n2187;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = n1573 & n2190;
  assign n2192 = ~n2185 & ~n2191;
  assign n2193 = ~n568 & ~n2192;
  assign n2194 = pi057 & n568;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~n566 & ~n2195;
  assign po104 = n2184 | n2196;
  assign n2198 = pi058 & ~pi270;
  assign n2199 = ~n1819 & ~n2198;
  assign n2200 = n566 & ~n2199;
  assign n2201 = pi058 & n568;
  assign n2202 = pi058 & ~n1573;
  assign n2203 = n1218 & n1825;
  assign n2204 = n1169 & n2203;
  assign n2205 = ~pi058 & ~n2203;
  assign n2206 = n1573 & ~n2205;
  assign n2207 = ~n2204 & n2206;
  assign n2208 = ~n2202 & ~n2207;
  assign n2209 = ~n568 & ~n2208;
  assign n2210 = ~n2201 & ~n2209;
  assign n2211 = ~n566 & ~n2210;
  assign po105 = n2200 | n2211;
  assign n2213 = pi059 & ~pi273;
  assign n2214 = ~n1766 & ~n2213;
  assign n2215 = n566 & ~n2214;
  assign n2216 = pi059 & n568;
  assign n2217 = pi059 & ~n1573;
  assign n2218 = ~n753 & n1641;
  assign n2219 = n1258 & n1449;
  assign n2220 = n2218 & n2219;
  assign n2221 = n1169 & n2220;
  assign n2222 = ~pi059 & ~n2220;
  assign n2223 = n1573 & ~n2222;
  assign n2224 = ~n2221 & n2223;
  assign n2225 = ~n2217 & ~n2224;
  assign n2226 = ~n568 & ~n2225;
  assign n2227 = ~n2216 & ~n2226;
  assign n2228 = ~n566 & ~n2227;
  assign po106 = n2215 | n2228;
  assign n2230 = pi060 & ~pi270;
  assign n2231 = ~n1838 & ~n2230;
  assign n2232 = n566 & ~n2231;
  assign n2233 = pi060 & ~n1573;
  assign n2234 = n1218 & n1843;
  assign n2235 = n1169 & n2234;
  assign n2236 = ~pi060 & ~n2234;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = n1573 & n2237;
  assign n2239 = ~n2233 & ~n2238;
  assign n2240 = ~n568 & ~n2239;
  assign n2241 = pi060 & n568;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~n566 & ~n2242;
  assign po107 = n2232 | n2243;
  assign n2245 = pi061 & ~pi271;
  assign n2246 = ~n1367 & ~n2245;
  assign n2247 = n566 & ~n2246;
  assign n2248 = pi061 & n568;
  assign n2249 = n568 & ~n2248;
  assign n2250 = ~n566 & ~n2249;
  assign n2251 = n1373 & n2171;
  assign n2252 = ~pi061 & ~n2251;
  assign n2253 = n1169 & n2251;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = n1573 & n2254;
  assign n2256 = pi061 & ~n2177;
  assign n2257 = ~n2255 & ~n2256;
  assign n2258 = n2250 & ~n2257;
  assign po108 = n2247 | n2258;
  assign n2260 = pi062 & ~pi271;
  assign n2261 = ~n1892 & ~n2260;
  assign n2262 = n566 & ~n2261;
  assign n2263 = pi062 & n568;
  assign n2264 = pi062 & ~n1573;
  assign n2265 = ~n753 & n1517;
  assign n2266 = n736 & n1611;
  assign n2267 = n2265 & n2266;
  assign n2268 = n1169 & n2267;
  assign n2269 = ~pi062 & ~n2267;
  assign n2270 = n1573 & ~n2269;
  assign n2271 = ~n2268 & n2270;
  assign n2272 = ~n2264 & ~n2271;
  assign n2273 = ~n568 & ~n2272;
  assign n2274 = ~n2263 & ~n2273;
  assign n2275 = ~n566 & ~n2274;
  assign po109 = n2262 | n2275;
  assign n2277 = pi063 & ~pi271;
  assign n2278 = ~n1349 & ~n2277;
  assign n2279 = n566 & ~n2278;
  assign n2280 = pi063 & ~n1573;
  assign n2281 = n1575 & n1587;
  assign n2282 = ~n753 & n2281;
  assign n2283 = n1169 & n2282;
  assign n2284 = ~pi063 & ~n2282;
  assign n2285 = ~n2283 & ~n2284;
  assign n2286 = n1573 & n2285;
  assign n2287 = ~n2280 & ~n2286;
  assign n2288 = ~n568 & ~n2287;
  assign n2289 = pi063 & n568;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = ~n566 & ~n2290;
  assign po110 = n2279 | n2291;
  assign n2293 = pi064 & ~pi271;
  assign n2294 = ~n1874 & ~n2293;
  assign n2295 = n566 & ~n2294;
  assign n2296 = pi064 & ~n1573;
  assign n2297 = n1880 & n2171;
  assign n2298 = n1169 & n2297;
  assign n2299 = ~pi064 & ~n2297;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = n1573 & n2300;
  assign n2302 = ~n2296 & ~n2301;
  assign n2303 = ~n568 & ~n2302;
  assign n2304 = pi064 & n568;
  assign n2305 = ~n2303 & ~n2304;
  assign n2306 = ~n566 & ~n2305;
  assign po111 = n2295 | n2306;
  assign n2308 = pi065 & ~pi272;
  assign n2309 = ~n1926 & ~n2308;
  assign n2310 = n566 & ~n2309;
  assign n2311 = pi065 & n568;
  assign n2312 = pi065 & ~n1573;
  assign n2313 = n1173 & n1643;
  assign n2314 = n1169 & n2313;
  assign n2315 = ~pi065 & ~n2313;
  assign n2316 = n1573 & ~n2315;
  assign n2317 = ~n2314 & n2316;
  assign n2318 = ~n2312 & ~n2317;
  assign n2319 = ~n568 & ~n2318;
  assign n2320 = ~n2311 & ~n2319;
  assign n2321 = ~n566 & ~n2320;
  assign po112 = n2310 | n2321;
  assign n2323 = pi066 & ~pi272;
  assign n2324 = ~n1385 & ~n2323;
  assign n2325 = n566 & ~n2324;
  assign n2326 = pi066 & ~n1573;
  assign n2327 = n1430 & n1642;
  assign n2328 = n1697 & n2327;
  assign n2329 = n1169 & n2328;
  assign n2330 = ~pi066 & ~n2328;
  assign n2331 = n1573 & ~n2330;
  assign n2332 = ~n2329 & n2331;
  assign n2333 = ~n2326 & ~n2332;
  assign n2334 = ~n568 & ~n2333;
  assign n2335 = pi066 & n568;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = ~n566 & ~n2336;
  assign po113 = n2325 | n2337;
  assign n2339 = pi067 & ~pi272;
  assign n2340 = ~n1406 & ~n2339;
  assign n2341 = n566 & ~n2340;
  assign n2342 = pi067 & ~n1573;
  assign n2343 = n1535 & n2327;
  assign n2344 = n1169 & n2343;
  assign n2345 = ~pi067 & ~n2343;
  assign n2346 = ~n2344 & ~n2345;
  assign n2347 = n1573 & n2346;
  assign n2348 = ~n2342 & ~n2347;
  assign n2349 = ~n568 & ~n2348;
  assign n2350 = pi067 & n568;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n566 & ~n2351;
  assign po114 = n2341 | n2352;
  assign n2354 = pi068 & ~n1573;
  assign n2355 = ~n676 & n699;
  assign n2356 = n1391 & n2355;
  assign n2357 = n736 & n2356;
  assign n2358 = n797 & n974;
  assign n2359 = n2357 & n2358;
  assign n2360 = n1169 & n2359;
  assign n2361 = ~pi068 & ~n2359;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = n1573 & n2362;
  assign n2364 = ~n2354 & ~n2363;
  assign n2365 = n1183 & ~n2364;
  assign n2366 = pi068 & n566;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = pi068 & ~pi272;
  assign n2369 = ~n1385 & ~n2368;
  assign n2370 = n569 & ~n2369;
  assign po115 = ~n2367 | n2370;
  assign n2372 = pi069 & ~n1573;
  assign n2373 = n1411 & n2355;
  assign n2374 = n753 & n2373;
  assign n2375 = n2358 & n2374;
  assign n2376 = n1169 & n2375;
  assign n2377 = ~pi069 & ~n2375;
  assign n2378 = ~n2376 & ~n2377;
  assign n2379 = n1573 & n2378;
  assign n2380 = ~n2372 & ~n2379;
  assign n2381 = n1183 & ~n2380;
  assign n2382 = pi069 & n566;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = pi069 & ~pi272;
  assign n2385 = ~n1406 & ~n2384;
  assign n2386 = n569 & ~n2385;
  assign po116 = ~n2383 | n2386;
  assign n2388 = pi070 & ~n1573;
  assign n2389 = n725 & n2355;
  assign n2390 = n1173 & n2389;
  assign n2391 = n2358 & n2390;
  assign n2392 = n1169 & n2391;
  assign n2393 = ~pi070 & ~n2391;
  assign n2394 = ~n2392 & ~n2393;
  assign n2395 = n1573 & n2394;
  assign n2396 = ~n2388 & ~n2395;
  assign n2397 = n1183 & ~n2396;
  assign n2398 = pi070 & n566;
  assign n2399 = ~n2397 & ~n2398;
  assign n2400 = pi070 & ~pi272;
  assign n2401 = ~n1926 & ~n2400;
  assign n2402 = n569 & ~n2401;
  assign po117 = ~n2399 | n2402;
  assign n2404 = ~n676 & n974;
  assign n2405 = n1260 & n2404;
  assign n2406 = ~pi071 & ~n2405;
  assign n2407 = n1169 & n2405;
  assign n2408 = ~n2406 & ~n2407;
  assign n2409 = n1573 & n2408;
  assign n2410 = pi071 & ~n1573;
  assign n2411 = ~n2409 & ~n2410;
  assign n2412 = n1183 & ~n2411;
  assign n2413 = pi071 & n566;
  assign n2414 = ~n2412 & ~n2413;
  assign n2415 = pi071 & ~pi270;
  assign n2416 = ~n1252 & ~n2415;
  assign n2417 = n569 & ~n2416;
  assign po118 = ~n2414 | n2417;
  assign n2419 = n1281 & n2404;
  assign n2420 = ~pi072 & ~n2419;
  assign n2421 = n1169 & n2419;
  assign n2422 = ~n2420 & ~n2421;
  assign n2423 = n1573 & n2422;
  assign n2424 = pi072 & ~n1573;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = n1183 & ~n2425;
  assign n2427 = pi072 & n566;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = pi072 & ~pi270;
  assign n2430 = ~n1274 & ~n2429;
  assign n2431 = n569 & ~n2430;
  assign po119 = ~n2428 | n2431;
  assign n2433 = ~n736 & n1171;
  assign n2434 = n1238 & n2433;
  assign n2435 = ~n753 & n2434;
  assign n2436 = ~pi073 & ~n2435;
  assign n2437 = n1169 & n2435;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = n1573 & n2438;
  assign n2440 = pi073 & ~n1573;
  assign n2441 = ~n2439 & ~n2440;
  assign n2442 = n1183 & ~n2441;
  assign n2443 = pi073 & n566;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = pi073 & ~pi270;
  assign n2446 = ~n1800 & ~n2445;
  assign n2447 = n569 & ~n2446;
  assign po120 = ~n2444 | n2447;
  assign n2449 = n1299 & n2404;
  assign n2450 = ~pi074 & ~n2449;
  assign n2451 = n1169 & n2449;
  assign n2452 = ~n2450 & ~n2451;
  assign n2453 = n1573 & n2452;
  assign n2454 = pi074 & ~n1573;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = n1183 & ~n2455;
  assign n2457 = pi074 & n566;
  assign n2458 = ~n2456 & ~n2457;
  assign n2459 = pi074 & ~pi270;
  assign n2460 = ~n1293 & ~n2459;
  assign n2461 = n569 & ~n2460;
  assign po121 = ~n2458 | n2461;
  assign n2463 = n725 & n1195;
  assign n2464 = n1173 & n2463;
  assign n2465 = ~n699 & n974;
  assign n2466 = n2464 & n2465;
  assign n2467 = ~pi075 & ~n2466;
  assign n2468 = n1169 & n2466;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = n1573 & n2469;
  assign n2471 = pi075 & ~n1573;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = n1183 & ~n2472;
  assign n2474 = pi075 & n566;
  assign n2475 = ~n2473 & ~n2474;
  assign n2476 = pi075 & ~pi271;
  assign n2477 = ~n1349 & ~n2476;
  assign n2478 = n569 & ~n2477;
  assign po122 = ~n2475 | n2478;
  assign n2480 = n736 & n1195;
  assign n2481 = n1391 & n2480;
  assign n2482 = n2465 & n2481;
  assign n2483 = ~pi076 & ~n2482;
  assign n2484 = n1169 & n2482;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = n1573 & n2485;
  assign n2487 = pi076 & ~n1573;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n1183 & ~n2488;
  assign n2490 = pi076 & n566;
  assign n2491 = ~n2489 & ~n2490;
  assign n2492 = pi076 & ~pi271;
  assign n2493 = ~n1892 & ~n2492;
  assign n2494 = n569 & ~n2493;
  assign po123 = ~n2491 | n2494;
  assign n2496 = n753 & n1195;
  assign n2497 = n1411 & n2496;
  assign n2498 = n2465 & n2497;
  assign n2499 = ~pi077 & ~n2498;
  assign n2500 = n1169 & n2498;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = n1573 & n2501;
  assign n2503 = pi077 & ~n1573;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = n1183 & ~n2504;
  assign n2506 = pi077 & n566;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = pi077 & ~pi271;
  assign n2509 = ~n1605 & ~n2508;
  assign n2510 = n569 & ~n2509;
  assign po124 = ~n2507 | n2510;
  assign n2512 = ~n676 & ~n699;
  assign n2513 = n2153 & n2512;
  assign n2514 = ~pi078 & ~n2513;
  assign n2515 = n1169 & n2513;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = n1573 & n2516;
  assign n2518 = pi078 & ~n1573;
  assign n2519 = ~n2517 & ~n2518;
  assign n2520 = n1183 & ~n2519;
  assign n2521 = pi078 & n566;
  assign n2522 = ~n2520 & ~n2521;
  assign n2523 = pi078 & ~pi271;
  assign n2524 = ~n1635 & ~n2523;
  assign n2525 = n569 & ~n2524;
  assign po125 = ~n2522 | n2525;
  assign n2527 = n736 & n1196;
  assign n2528 = ~n753 & n2527;
  assign n2529 = n1197 & n2528;
  assign n2530 = ~pi079 & ~n2529;
  assign n2531 = n1169 & n2529;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = n1573 & n2532;
  assign n2534 = pi079 & ~n1573;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = n1183 & ~n2535;
  assign n2537 = pi079 & n566;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = pi079 & ~pi273;
  assign n2540 = ~n1766 & ~n2539;
  assign n2541 = n569 & ~n2540;
  assign po126 = ~n2538 | n2541;
  assign n2543 = n1196 & n1535;
  assign n2544 = n1197 & n2543;
  assign n2545 = ~pi080 & ~n2544;
  assign n2546 = n1169 & n2544;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n1573 & n2547;
  assign n2549 = pi080 & ~n1573;
  assign n2550 = ~n2548 & ~n2549;
  assign n2551 = n1183 & ~n2550;
  assign n2552 = pi080 & n566;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = pi080 & ~pi273;
  assign n2555 = ~n2005 & ~n2554;
  assign n2556 = n569 & ~n2555;
  assign po127 = ~n2553 | n2556;
  assign n2558 = n1451 & n2404;
  assign n2559 = ~pi081 & ~n2558;
  assign n2560 = n1169 & n2558;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = n1573 & n2561;
  assign n2563 = pi081 & ~n1573;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = n1183 & ~n2564;
  assign n2566 = pi081 & n566;
  assign n2567 = ~n2565 & ~n2566;
  assign n2568 = pi081 & ~pi273;
  assign n2569 = ~n1444 & ~n2568;
  assign n2570 = n569 & ~n2569;
  assign po128 = ~n2567 | n2570;
  assign n2572 = n1469 & n2404;
  assign n2573 = ~pi082 & ~n2572;
  assign n2574 = n1169 & n2572;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = n1573 & n2575;
  assign n2577 = pi082 & ~n1573;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = n1183 & ~n2578;
  assign n2580 = pi082 & n566;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = pi082 & ~pi273;
  assign n2583 = ~n1463 & ~n2582;
  assign n2584 = n569 & ~n2583;
  assign po129 = ~n2581 | n2584;
  assign n2586 = n1487 & n2404;
  assign n2587 = ~pi083 & ~n2586;
  assign n2588 = n1169 & n2586;
  assign n2589 = ~n2587 & ~n2588;
  assign n2590 = n1573 & n2589;
  assign n2591 = pi083 & ~n1573;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = n1183 & ~n2592;
  assign n2594 = pi083 & n566;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = pi083 & ~pi273;
  assign n2597 = ~n1481 & ~n2596;
  assign n2598 = n569 & ~n2597;
  assign po130 = ~n2595 | n2598;
  assign n2600 = ~n676 & ~n974;
  assign n2601 = ~n797 & n2600;
  assign n2602 = n1861 & n2601;
  assign n2603 = ~n1169 & n2602;
  assign n2604 = pi084 & ~n2602;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = n1573 & ~n2605;
  assign n2607 = ~n579 & n584;
  assign n2608 = pi084 & ~pi271;
  assign n2609 = ~n1600 & ~n2608;
  assign n2610 = n2607 & ~n2609;
  assign n2611 = ~n2606 & ~n2610;
  assign n2612 = n1183 & ~n2611;
  assign n2613 = ~n579 & n1183;
  assign n2614 = pi084 & ~n2613;
  assign po131 = n2612 | n2614;
  assign n2616 = ~n699 & ~n725;
  assign n2617 = n2601 & n2616;
  assign n2618 = n1173 & n2617;
  assign n2619 = ~n1169 & n2618;
  assign n2620 = pi085 & ~n2618;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = n1573 & ~n2621;
  assign n2623 = pi085 & ~pi271;
  assign n2624 = ~n1635 & ~n2623;
  assign n2625 = n2607 & ~n2624;
  assign n2626 = ~n2622 & ~n2625;
  assign n2627 = n1183 & ~n2626;
  assign n2628 = pi085 & ~n2613;
  assign po132 = n2627 | n2628;
  assign n2630 = n699 & n2600;
  assign n2631 = n1519 & n2630;
  assign n2632 = ~n1169 & n2631;
  assign n2633 = pi086 & ~n2631;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = n1573 & ~n2634;
  assign n2636 = pi086 & ~pi272;
  assign n2637 = ~n1655 & ~n2636;
  assign n2638 = n2607 & ~n2637;
  assign n2639 = ~n2635 & ~n2638;
  assign n2640 = n1183 & ~n2639;
  assign n2641 = pi086 & ~n2613;
  assign po133 = n2640 | n2641;
  assign n2643 = n1552 & n2630;
  assign n2644 = n1173 & n2643;
  assign n2645 = ~n1169 & n2644;
  assign n2646 = pi087 & ~n2644;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = n1573 & ~n2647;
  assign n2649 = pi087 & ~pi272;
  assign n2650 = ~n1425 & ~n2649;
  assign n2651 = n2607 & ~n2650;
  assign n2652 = ~n2648 & ~n2651;
  assign n2653 = n1183 & ~n2652;
  assign n2654 = pi087 & ~n2613;
  assign po134 = n2653 | n2654;
  assign n2656 = n1787 & n2528;
  assign n2657 = ~n1169 & n2656;
  assign n2658 = pi088 & ~n2656;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = n1573 & ~n2659;
  assign n2661 = pi088 & ~pi273;
  assign n2662 = ~n1766 & ~n2661;
  assign n2663 = n2607 & ~n2662;
  assign n2664 = ~n2660 & ~n2663;
  assign n2665 = n1183 & ~n2664;
  assign n2666 = pi088 & ~n2613;
  assign po135 = n2665 | n2666;
  assign n2668 = n1260 & n2600;
  assign n2669 = ~n1169 & n2668;
  assign n2670 = pi089 & ~n2668;
  assign n2671 = ~n2669 & ~n2670;
  assign n2672 = n1573 & ~n2671;
  assign n2673 = pi089 & ~pi270;
  assign n2674 = ~n1252 & ~n2673;
  assign n2675 = n2607 & ~n2674;
  assign n2676 = ~n2672 & ~n2675;
  assign n2677 = n1183 & ~n2676;
  assign n2678 = pi089 & ~n2613;
  assign po136 = n2677 | n2678;
  assign n2680 = n1587 & n2630;
  assign n2681 = n1173 & n2680;
  assign n2682 = ~n1169 & n2681;
  assign n2683 = pi090 & ~n2681;
  assign n2684 = ~n2682 & ~n2683;
  assign n2685 = n1573 & ~n2684;
  assign n2686 = pi090 & ~pi273;
  assign n2687 = ~n1444 & ~n2686;
  assign n2688 = n2607 & ~n2687;
  assign n2689 = ~n2685 & ~n2688;
  assign n2690 = n1183 & ~n2689;
  assign n2691 = pi090 & ~n2613;
  assign po137 = n2690 | n2691;
  assign n2693 = n1697 & n2630;
  assign n2694 = n1611 & n2693;
  assign n2695 = ~n1169 & n2694;
  assign n2696 = pi091 & ~n2694;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = n1573 & ~n2697;
  assign n2699 = pi091 & ~pi273;
  assign n2700 = ~n1463 & ~n2699;
  assign n2701 = n2607 & ~n2700;
  assign n2702 = ~n2698 & ~n2701;
  assign n2703 = n1183 & ~n2702;
  assign n2704 = pi091 & ~n2613;
  assign po138 = n2703 | n2704;
  assign n2706 = n1535 & n2630;
  assign n2707 = n1611 & n2706;
  assign n2708 = ~n1169 & n2707;
  assign n2709 = pi092 & ~n2707;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n1573 & ~n2710;
  assign n2712 = pi092 & ~pi273;
  assign n2713 = ~n1481 & ~n2712;
  assign n2714 = n2607 & ~n2713;
  assign n2715 = ~n2711 & ~n2714;
  assign n2716 = n1183 & ~n2715;
  assign n2717 = pi092 & ~n2613;
  assign po139 = n2716 | n2717;
  assign n2719 = n1787 & n2543;
  assign n2720 = ~n1169 & n2719;
  assign n2721 = pi093 & ~n2719;
  assign n2722 = ~n2720 & ~n2721;
  assign n2723 = n1573 & ~n2722;
  assign n2724 = pi093 & ~pi273;
  assign n2725 = ~n2005 & ~n2724;
  assign n2726 = n2607 & ~n2725;
  assign n2727 = ~n2723 & ~n2726;
  assign n2728 = n1183 & ~n2727;
  assign n2729 = pi093 & ~n2613;
  assign po140 = n2728 | n2729;
  assign n2731 = n1623 & n2630;
  assign n2732 = ~n1169 & n2731;
  assign n2733 = pi094 & ~n2731;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n1573 & ~n2734;
  assign n2736 = pi094 & ~pi273;
  assign n2737 = ~n1213 & ~n2736;
  assign n2738 = n2607 & ~n2737;
  assign n2739 = ~n2735 & ~n2738;
  assign n2740 = n1183 & ~n2739;
  assign n2741 = pi094 & ~n2613;
  assign po141 = n2740 | n2741;
  assign n2743 = ~n725 & n2527;
  assign n2744 = n753 & n2743;
  assign n2745 = ~n974 & n2744;
  assign n2746 = ~n1169 & n2745;
  assign n2747 = pi095 & ~n2745;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = n1573 & ~n2748;
  assign n2750 = pi095 & ~pi273;
  assign n2751 = ~n1747 & ~n2750;
  assign n2752 = n2607 & ~n2751;
  assign n2753 = ~n2749 & ~n2752;
  assign n2754 = n1183 & ~n2753;
  assign n2755 = pi095 & ~n2613;
  assign po142 = n2754 | n2755;
  assign n2757 = n1281 & n2600;
  assign n2758 = ~n1169 & n2757;
  assign n2759 = pi096 & ~n2757;
  assign n2760 = ~n2758 & ~n2759;
  assign n2761 = n1573 & ~n2760;
  assign n2762 = pi096 & ~pi270;
  assign n2763 = ~n1274 & ~n2762;
  assign n2764 = n2607 & ~n2763;
  assign n2765 = ~n2761 & ~n2764;
  assign n2766 = n1183 & ~n2765;
  assign n2767 = pi096 & ~n2613;
  assign po143 = n2766 | n2767;
  assign n2769 = n1518 & n2706;
  assign n2770 = ~n1169 & n2769;
  assign n2771 = pi097 & ~n2769;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = n1573 & ~n2772;
  assign n2774 = pi097 & ~pi272;
  assign n2775 = ~n1679 & ~n2774;
  assign n2776 = n2607 & ~n2775;
  assign n2777 = ~n2773 & ~n2776;
  assign n2778 = n1183 & ~n2777;
  assign n2779 = pi097 & ~n2613;
  assign po144 = n2778 | n2779;
  assign n2781 = n974 & n2744;
  assign n2782 = n1169 & n2781;
  assign n2783 = ~pi098 & ~n2781;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = n1573 & n2784;
  assign n2786 = pi098 & ~n1573;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = n1183 & ~n2787;
  assign n2789 = pi098 & n566;
  assign n2790 = ~n2788 & ~n2789;
  assign n2791 = pi098 & ~pi273;
  assign n2792 = ~n1747 & ~n2791;
  assign n2793 = n569 & ~n2792;
  assign po145 = ~n2790 | n2793;
  assign n2795 = n974 & n2355;
  assign n2796 = n1519 & n2795;
  assign n2797 = n1169 & n2796;
  assign n2798 = ~pi099 & ~n2796;
  assign n2799 = ~n2797 & ~n2798;
  assign n2800 = n1573 & n2799;
  assign n2801 = pi099 & ~n1573;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = n1183 & ~n2802;
  assign n2804 = pi099 & n566;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = pi099 & ~pi272;
  assign n2807 = ~n1655 & ~n2806;
  assign n2808 = n569 & ~n2807;
  assign po146 = ~n2805 | n2808;
  assign n2810 = ~n753 & n2465;
  assign n2811 = n1258 & n2810;
  assign n2812 = n1195 & n2811;
  assign n2813 = n1169 & n2812;
  assign n2814 = ~pi100 & ~n2812;
  assign n2815 = ~n2813 & ~n2814;
  assign n2816 = n1573 & n2815;
  assign n2817 = pi100 & ~n1573;
  assign n2818 = ~n2816 & ~n2817;
  assign n2819 = n1183 & ~n2818;
  assign n2820 = pi100 & n566;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = pi100 & ~pi271;
  assign n2823 = ~n1874 & ~n2822;
  assign n2824 = n569 & ~n2823;
  assign po147 = ~n2821 | n2824;
  assign n2826 = n974 & n1195;
  assign n2827 = n1861 & n2826;
  assign n2828 = n1169 & n2827;
  assign n2829 = ~pi101 & ~n2827;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = n1573 & n2830;
  assign n2832 = pi101 & ~n1573;
  assign n2833 = ~n2831 & ~n2832;
  assign n2834 = n1183 & ~n2833;
  assign n2835 = pi101 & n566;
  assign n2836 = ~n2834 & ~n2835;
  assign n2837 = pi101 & ~pi271;
  assign n2838 = ~n1600 & ~n2837;
  assign n2839 = n569 & ~n2838;
  assign po148 = ~n2836 | n2839;
  assign n2841 = n736 & n2630;
  assign n2842 = n753 & n1587;
  assign n2843 = n2841 & n2842;
  assign n2844 = n1573 & ~n2843;
  assign n2845 = pi102 & n2844;
  assign n2846 = n1573 & n2843;
  assign n2847 = ~n1169 & n2846;
  assign n2848 = ~n2845 & ~n2847;
  assign n2849 = pi102 & ~pi273;
  assign n2850 = ~n1189 & ~n2849;
  assign n2851 = n2607 & ~n2850;
  assign n2852 = n2848 & ~n2851;
  assign n2853 = n1183 & ~n2852;
  assign n2854 = pi102 & ~n2613;
  assign po149 = n2853 | n2854;
  assign n2856 = n736 & n2601;
  assign n2857 = ~n753 & n2856;
  assign n2858 = n1860 & n2857;
  assign n2859 = ~n1169 & n2858;
  assign n2860 = pi103 & ~n2858;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = n1573 & ~n2861;
  assign n2863 = pi103 & ~pi271;
  assign n2864 = ~n1874 & ~n2863;
  assign n2865 = n2607 & ~n2864;
  assign n2866 = ~n2862 & ~n2865;
  assign n2867 = n1183 & ~n2866;
  assign n2868 = pi103 & ~n2613;
  assign po150 = n2867 | n2868;
  assign n2870 = ~n753 & n2841;
  assign n2871 = n1518 & n2870;
  assign n2872 = ~n1169 & n2871;
  assign n2873 = pi104 & ~n2871;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = n1573 & ~n2874;
  assign n2876 = pi104 & ~pi272;
  assign n2877 = ~n1660 & ~n2876;
  assign n2878 = n2607 & ~n2877;
  assign n2879 = ~n2875 & ~n2878;
  assign n2880 = n1183 & ~n2879;
  assign n2881 = pi104 & ~n2613;
  assign po151 = n2880 | n2881;
  assign n2883 = n753 & n2856;
  assign n2884 = n2616 & n2883;
  assign n2885 = ~n1169 & n2884;
  assign n2886 = pi105 & ~n2884;
  assign n2887 = ~n2885 & ~n2886;
  assign n2888 = n1573 & ~n2887;
  assign n2889 = pi105 & ~pi271;
  assign n2890 = ~n1367 & ~n2889;
  assign n2891 = n2607 & ~n2890;
  assign n2892 = ~n2888 & ~n2891;
  assign n2893 = n1183 & ~n2892;
  assign n2894 = pi105 & ~n2613;
  assign po152 = n2893 | n2894;
  assign n2896 = n1171 & n1697;
  assign n2897 = n1172 & n2896;
  assign n2898 = n1169 & n2897;
  assign n2899 = ~pi106 & ~n2897;
  assign n2900 = ~n2898 & ~n2899;
  assign n2901 = n1573 & n2900;
  assign n2902 = pi106 & ~n1573;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = n1183 & ~n2903;
  assign n2905 = pi106 & n566;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = pi106 & ~pi270;
  assign n2908 = ~n1819 & ~n2907;
  assign n2909 = n569 & ~n2908;
  assign po153 = ~n2906 | n2909;
  assign n2911 = n753 & n2433;
  assign n2912 = n1172 & n2911;
  assign n2913 = n1169 & n2912;
  assign n2914 = ~pi107 & ~n2912;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = n1573 & n2915;
  assign n2917 = pi107 & ~n1573;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = n1183 & ~n2918;
  assign n2920 = pi107 & n566;
  assign n2921 = ~n2919 & ~n2920;
  assign n2922 = pi107 & ~pi270;
  assign n2923 = ~n1838 & ~n2922;
  assign n2924 = n569 & ~n2923;
  assign po154 = ~n2921 | n2924;
  assign n2926 = n753 & n2841;
  assign n2927 = n1552 & n2926;
  assign n2928 = ~n1169 & n2927;
  assign n2929 = pi108 & ~n2927;
  assign n2930 = ~n2928 & ~n2929;
  assign n2931 = n1573 & ~n2930;
  assign n2932 = pi108 & ~pi272;
  assign n2933 = ~n1714 & ~n2932;
  assign n2934 = n2607 & ~n2933;
  assign n2935 = ~n2931 & ~n2934;
  assign n2936 = n1183 & ~n2935;
  assign n2937 = pi108 & ~n2613;
  assign po155 = n2936 | n2937;
  assign n2939 = ~n736 & n2465;
  assign n2940 = n1279 & n2939;
  assign n2941 = n1195 & n2940;
  assign n2942 = n1169 & n2941;
  assign n2943 = ~pi109 & ~n2941;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = n1573 & n2944;
  assign n2946 = pi109 & ~n1573;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = n1183 & ~n2947;
  assign n2949 = pi109 & n566;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = pi109 & ~pi271;
  assign n2952 = ~n1329 & ~n2951;
  assign n2953 = n569 & ~n2952;
  assign po156 = ~n2950 | n2953;
  assign n2955 = ~n753 & n2358;
  assign n2956 = n1258 & n2955;
  assign n2957 = n2355 & n2956;
  assign n2958 = n1169 & n2957;
  assign n2959 = ~pi110 & ~n2957;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = n1573 & n2960;
  assign n2962 = pi110 & ~n1573;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = n1183 & ~n2963;
  assign n2965 = pi110 & n566;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = pi110 & ~pi272;
  assign n2968 = ~n1660 & ~n2967;
  assign n2969 = n569 & ~n2968;
  assign po157 = ~n2966 | n2969;
  assign n2971 = ~n736 & n2358;
  assign n2972 = n1279 & n2971;
  assign n2973 = n2355 & n2972;
  assign n2974 = n1169 & n2973;
  assign n2975 = ~pi111 & ~n2973;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = n1573 & n2976;
  assign n2978 = pi111 & ~n1573;
  assign n2979 = ~n2977 & ~n2978;
  assign n2980 = n1183 & ~n2979;
  assign n2981 = pi111 & n566;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = pi111 & ~pi272;
  assign n2984 = ~n1679 & ~n2983;
  assign n2985 = n569 & ~n2984;
  assign po158 = ~n2982 | n2985;
  assign n2987 = ~n725 & n2465;
  assign n2988 = n1194 & n2987;
  assign n2989 = n1195 & n2988;
  assign n2990 = n1169 & n2989;
  assign n2991 = ~pi112 & ~n2989;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = n1573 & n2992;
  assign n2994 = pi112 & ~n1573;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = n1183 & ~n2995;
  assign n2997 = pi112 & n566;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = pi112 & ~pi271;
  assign n3000 = ~n1367 & ~n2999;
  assign n3001 = n569 & ~n3000;
  assign po159 = ~n2998 | n3001;
  assign n3003 = ~n725 & n2358;
  assign n3004 = n1194 & n3003;
  assign n3005 = n2355 & n3004;
  assign n3006 = n1169 & n3005;
  assign n3007 = ~pi113 & ~n3005;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = n1573 & n3008;
  assign n3010 = pi113 & ~n1573;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = n1183 & ~n3011;
  assign n3013 = pi113 & n566;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = pi113 & ~pi272;
  assign n3016 = ~n1714 & ~n3015;
  assign n3017 = n569 & ~n3016;
  assign po160 = ~n3014 | n3017;
  assign n3019 = ~pi114 & ~n1573;
  assign n3020 = n1183 & ~n3019;
  assign n3021 = n797 & n1431;
  assign n3022 = n2404 & n3021;
  assign n3023 = n1169 & n3022;
  assign n3024 = ~pi114 & ~n3022;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = n1573 & ~n3025;
  assign n3027 = n3020 & ~n3026;
  assign n3028 = pi114 & ~pi272;
  assign n3029 = ~n1425 & ~n3028;
  assign n3030 = n569 & ~n3029;
  assign n3031 = pi114 & n566;
  assign n3032 = ~n3030 & ~n3031;
  assign po161 = n3027 | ~n3032;
  assign n3034 = ~n974 & n1174;
  assign n3035 = n1170 & n3034;
  assign n3036 = ~n1169 & n3035;
  assign n3037 = pi115 & ~pi270;
  assign n3038 = ~n571 & ~n3037;
  assign n3039 = n2607 & ~n3038;
  assign n3040 = pi115 & ~n3035;
  assign n3041 = ~n3039 & ~n3040;
  assign n3042 = ~n3036 & n3041;
  assign n3043 = ~n1573 & ~n3039;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = n1183 & n3044;
  assign n3046 = pi115 & ~n2613;
  assign po162 = n3045 | n3046;
  assign n3048 = n1299 & n2600;
  assign n3049 = ~n1169 & n3048;
  assign n3050 = pi116 & ~n3048;
  assign n3051 = ~n3049 & ~n3050;
  assign n3052 = n1573 & ~n3051;
  assign n3053 = pi116 & ~pi270;
  assign n3054 = ~n1293 & ~n3053;
  assign n3055 = n2607 & ~n3054;
  assign n3056 = ~n3052 & ~n3055;
  assign n3057 = n1183 & ~n3056;
  assign n3058 = pi116 & ~n2613;
  assign po163 = n3057 | n3058;
  assign n3060 = n1535 & n2601;
  assign n3061 = n1860 & n3060;
  assign n3062 = ~n1169 & n3061;
  assign n3063 = pi117 & ~n3061;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = n1573 & ~n3064;
  assign n3066 = pi117 & ~pi271;
  assign n3067 = ~n1329 & ~n3066;
  assign n3068 = n2607 & ~n3067;
  assign n3069 = ~n3065 & ~n3068;
  assign n3070 = n1183 & ~n3069;
  assign n3071 = pi117 & ~n2613;
  assign po164 = n3070 | n3071;
  assign n3073 = n1914 & n2512;
  assign n3074 = ~n1169 & n3073;
  assign n3075 = pi118 & ~n3073;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = n1573 & ~n3076;
  assign n3078 = pi118 & ~pi270;
  assign n3079 = ~n1233 & ~n3078;
  assign n3080 = n2607 & ~n3079;
  assign n3081 = ~n3077 & ~n3080;
  assign n3082 = n1183 & ~n3081;
  assign n3083 = pi118 & ~n2613;
  assign po165 = n3082 | n3083;
  assign n3085 = n725 & n1170;
  assign n3086 = n2600 & n3085;
  assign n3087 = n1173 & n3086;
  assign n3088 = ~n1169 & n3087;
  assign n3089 = pi119 & ~n3087;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = n1573 & ~n3090;
  assign n3092 = pi119 & ~pi270;
  assign n3093 = ~n1800 & ~n3092;
  assign n3094 = n2607 & ~n3093;
  assign n3095 = ~n3091 & ~n3094;
  assign n3096 = n1183 & ~n3095;
  assign n3097 = pi119 & ~n2613;
  assign po166 = n3096 | n3097;
  assign n3099 = n797 & ~n974;
  assign n3100 = n2374 & n3099;
  assign n3101 = ~n1169 & n3100;
  assign n3102 = pi120 & ~n3100;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = n1573 & ~n3103;
  assign n3105 = pi120 & ~pi272;
  assign n3106 = ~n1406 & ~n3105;
  assign n3107 = n2607 & ~n3106;
  assign n3108 = ~n3104 & ~n3107;
  assign n3109 = n1183 & ~n3108;
  assign n3110 = pi120 & ~n2613;
  assign po167 = n3109 | n3110;
  assign n3112 = n2390 & n3099;
  assign n3113 = ~n1169 & n3112;
  assign n3114 = pi121 & ~pi272;
  assign n3115 = ~n1926 & ~n3114;
  assign n3116 = n2607 & ~n3115;
  assign n3117 = pi121 & ~n3112;
  assign n3118 = ~n3116 & ~n3117;
  assign n3119 = ~n3113 & n3118;
  assign n3120 = ~n1573 & ~n3116;
  assign n3121 = ~n3119 & ~n3120;
  assign n3122 = n1183 & n3121;
  assign n3123 = pi121 & ~n2613;
  assign po168 = n3122 | n3123;
  assign n3125 = pi122 & ~pi270;
  assign n3126 = ~n1819 & ~n3125;
  assign n3127 = n2607 & ~n3126;
  assign n3128 = ~n1573 & ~n3127;
  assign n3129 = n1183 & ~n3128;
  assign n3130 = n1170 & n2600;
  assign n3131 = n1468 & n3130;
  assign n3132 = ~n1169 & n3131;
  assign n3133 = pi122 & ~n3131;
  assign n3134 = ~n3127 & ~n3133;
  assign n3135 = ~n3132 & n3134;
  assign n3136 = n3129 & ~n3135;
  assign n3137 = pi122 & ~n2613;
  assign po169 = n3136 | n3137;
  assign n3139 = n2042 & n3130;
  assign n3140 = ~n1169 & n3139;
  assign n3141 = pi123 & ~pi270;
  assign n3142 = ~n1838 & ~n3141;
  assign n3143 = n2607 & ~n3142;
  assign n3144 = pi123 & ~n3139;
  assign n3145 = ~n3143 & ~n3144;
  assign n3146 = ~n3140 & n3145;
  assign n3147 = ~n1573 & ~n3143;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = n1183 & n3148;
  assign n3150 = pi123 & ~n2613;
  assign po170 = n3149 | n3150;
  assign n3152 = ~n699 & ~n974;
  assign n3153 = n2464 & n3152;
  assign n3154 = ~n1169 & n3153;
  assign n3155 = pi124 & ~n3153;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = n1573 & ~n3156;
  assign n3158 = pi124 & ~pi271;
  assign n3159 = ~n1349 & ~n3158;
  assign n3160 = n2607 & ~n3159;
  assign n3161 = ~n3157 & ~n3160;
  assign n3162 = n1183 & ~n3161;
  assign n3163 = pi124 & ~n2613;
  assign po171 = n3162 | n3163;
  assign n3165 = pi125 & ~pi271;
  assign n3166 = ~n1892 & ~n3165;
  assign n3167 = n1183 & ~n3166;
  assign n3168 = n2607 & n3167;
  assign n3169 = pi125 & ~n2613;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = n1183 & n1573;
  assign n3172 = n2481 & n3152;
  assign n3173 = ~n1169 & n3172;
  assign n3174 = pi125 & ~n3172;
  assign n3175 = ~n3173 & ~n3174;
  assign n3176 = n3171 & ~n3175;
  assign po172 = ~n3170 | n3176;
  assign n3178 = pi126 & ~pi271;
  assign n3179 = ~n1605 & ~n3178;
  assign n3180 = n1183 & ~n3179;
  assign n3181 = n2607 & n3180;
  assign n3182 = pi126 & ~n2613;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = n2497 & n3152;
  assign n3185 = ~n1169 & n3184;
  assign n3186 = pi126 & ~n3184;
  assign n3187 = ~n3185 & ~n3186;
  assign n3188 = n3171 & ~n3187;
  assign po173 = ~n3183 | n3188;
  assign n3190 = n2357 & n3099;
  assign n3191 = ~n1169 & n3190;
  assign n3192 = pi127 & ~n3190;
  assign n3193 = ~n3191 & ~n3192;
  assign n3194 = n1573 & ~n3193;
  assign n3195 = pi127 & ~pi272;
  assign n3196 = ~n1385 & ~n3195;
  assign n3197 = n2607 & ~n3196;
  assign n3198 = ~n3194 & ~n3197;
  assign n3199 = n1183 & ~n3198;
  assign n3200 = pi127 & ~n2613;
  assign po174 = n3199 | n3200;
  assign n3202 = ~pi144 & pi145;
  assign n3203 = pi144 & ~pi146;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = ~n593 & ~n3204;
  assign n3206 = pi136 & ~n3205;
  assign n3207 = pi128 & n3206;
  assign n3208 = ~pi143 & n732;
  assign n3209 = pi171 & ~pi187;
  assign n3210 = ~pi171 & pi187;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = ~pi150 & pi190;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = n3211 & n3212;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = pi143 & n3215;
  assign n3217 = ~n3208 & ~n3216;
  assign n3218 = pi143 & ~pi150;
  assign n3219 = ~pi190 & ~n3218;
  assign n3220 = pi143 & n3212;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = pi097 & n3221;
  assign n3223 = pi121 & ~n3221;
  assign n3224 = ~n3222 & ~n3223;
  assign n3225 = n3217 & ~n3224;
  assign n3226 = pi086 & n3221;
  assign n3227 = pi104 & ~n3221;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = ~n3217 & ~n3228;
  assign n3230 = ~n3225 & ~n3229;
  assign n3231 = ~pi143 & ~n702;
  assign n3232 = pi142 & ~pi176;
  assign n3233 = ~pi142 & pi176;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = pi148 & ~pi156;
  assign n3236 = ~n3210 & ~n3212;
  assign n3237 = ~n3235 & n3236;
  assign n3238 = n3209 & ~n3235;
  assign n3239 = ~pi148 & pi156;
  assign n3240 = ~n3238 & ~n3239;
  assign n3241 = ~n3237 & n3240;
  assign n3242 = n3234 & n3241;
  assign n3243 = ~n3234 & ~n3241;
  assign n3244 = ~n3242 & ~n3243;
  assign n3245 = pi143 & ~n3244;
  assign n3246 = ~n3231 & ~n3245;
  assign n3247 = ~pi143 & ~n721;
  assign n3248 = ~n3235 & ~n3239;
  assign n3249 = ~n3209 & ~n3236;
  assign n3250 = ~n3248 & ~n3249;
  assign n3251 = n3248 & n3249;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = pi143 & ~n3252;
  assign n3254 = ~n3247 & ~n3253;
  assign n3255 = n3246 & n3254;
  assign n3256 = ~n3230 & n3255;
  assign n3257 = pi087 & ~n3221;
  assign n3258 = pi120 & n3221;
  assign n3259 = ~n3257 & ~n3258;
  assign n3260 = n3217 & ~n3259;
  assign n3261 = pi108 & n3221;
  assign n3262 = pi127 & ~n3221;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = ~n3217 & ~n3263;
  assign n3265 = ~n3260 & ~n3264;
  assign n3266 = n3246 & ~n3254;
  assign n3267 = ~n3265 & n3266;
  assign n3268 = pi092 & n3221;
  assign n3269 = pi094 & ~n3221;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = n3217 & ~n3270;
  assign n3272 = pi095 & n3221;
  assign n3273 = pi091 & ~n3221;
  assign n3274 = ~n3272 & ~n3273;
  assign n3275 = ~n3217 & ~n3274;
  assign n3276 = ~n3271 & ~n3275;
  assign n3277 = ~n3254 & ~n3276;
  assign n3278 = pi093 & n3221;
  assign n3279 = pi090 & ~n3221;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = n3217 & ~n3280;
  assign n3282 = pi088 & ~n3221;
  assign n3283 = pi102 & n3221;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = ~n3217 & ~n3284;
  assign n3286 = ~n3281 & ~n3285;
  assign n3287 = n3254 & ~n3286;
  assign n3288 = ~n3277 & ~n3287;
  assign n3289 = ~n3246 & ~n3288;
  assign n3290 = ~n3267 & ~n3289;
  assign n3291 = ~n3256 & n3290;
  assign n3292 = pi139 & ~pi177;
  assign n3293 = ~pi139 & pi177;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = ~n3232 & n3239;
  assign n3296 = ~n3233 & ~n3295;
  assign n3297 = ~n3232 & ~n3235;
  assign n3298 = ~n3249 & n3297;
  assign n3299 = n3296 & ~n3298;
  assign n3300 = ~n3294 & ~n3299;
  assign n3301 = pi143 & n3300;
  assign n3302 = ~pi143 & n682;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = pi143 & n3294;
  assign n3305 = n3299 & n3304;
  assign n3306 = n3303 & ~n3305;
  assign n3307 = n3291 & ~n3306;
  assign n3308 = pi085 & ~n3221;
  assign n3309 = pi126 & n3221;
  assign n3310 = ~n3308 & ~n3309;
  assign n3311 = n3217 & ~n3310;
  assign n3312 = pi105 & n3221;
  assign n3313 = pi125 & ~n3221;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n3217 & ~n3314;
  assign n3316 = ~n3311 & ~n3315;
  assign n3317 = ~n3254 & ~n3316;
  assign n3318 = pi124 & ~n3221;
  assign n3319 = pi117 & n3221;
  assign n3320 = ~n3318 & ~n3319;
  assign n3321 = n3217 & ~n3320;
  assign n3322 = pi084 & n3221;
  assign n3323 = pi103 & ~n3221;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3217 & ~n3324;
  assign n3326 = ~n3321 & ~n3325;
  assign n3327 = n3254 & ~n3326;
  assign n3328 = ~n3317 & ~n3327;
  assign n3329 = ~n3246 & ~n3328;
  assign n3330 = pi096 & n3221;
  assign n3331 = pi119 & ~n3221;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = n3217 & ~n3332;
  assign n3334 = pi118 & n3221;
  assign n3335 = pi089 & ~n3221;
  assign n3336 = ~n3334 & ~n3335;
  assign n3337 = ~n3217 & ~n3336;
  assign n3338 = ~n3333 & ~n3337;
  assign n3339 = n3255 & ~n3338;
  assign n3340 = ~n3329 & ~n3339;
  assign n3341 = pi123 & n3221;
  assign n3342 = pi115 & ~n3221;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = n3217 & ~n3343;
  assign n3345 = pi122 & ~n3221;
  assign n3346 = pi116 & n3221;
  assign n3347 = ~n3345 & ~n3346;
  assign n3348 = ~n3217 & ~n3347;
  assign n3349 = ~n3344 & ~n3348;
  assign n3350 = n3266 & ~n3349;
  assign n3351 = n3340 & ~n3350;
  assign n3352 = n3306 & n3351;
  assign n3353 = ~n3307 & ~n3352;
  assign n3354 = pi140 & ~pi161;
  assign n3355 = ~pi140 & pi161;
  assign n3356 = ~n3354 & ~n3355;
  assign n3357 = n3233 & ~n3292;
  assign n3358 = ~n3232 & ~n3292;
  assign n3359 = ~n3240 & n3358;
  assign n3360 = ~n3357 & ~n3359;
  assign n3361 = n3237 & n3358;
  assign n3362 = ~n3293 & ~n3361;
  assign n3363 = n3360 & n3362;
  assign n3364 = n3356 & n3363;
  assign n3365 = ~n3356 & ~n3363;
  assign n3366 = ~n3364 & ~n3365;
  assign n3367 = pi143 & ~n3366;
  assign n3368 = ~pi143 & ~n672;
  assign n3369 = ~n3367 & ~n3368;
  assign n3370 = ~n3353 & ~n3369;
  assign n3371 = pi045 & n3221;
  assign n3372 = pi041 & ~n3221;
  assign n3373 = ~n3371 & ~n3372;
  assign n3374 = n3217 & ~n3373;
  assign n3375 = pi040 & n3221;
  assign n3376 = pi043 & ~n3221;
  assign n3377 = ~n3375 & ~n3376;
  assign n3378 = ~n3217 & ~n3377;
  assign n3379 = ~n3374 & ~n3378;
  assign n3380 = n3255 & ~n3379;
  assign n3381 = pi014 & ~n3221;
  assign n3382 = pi046 & n3221;
  assign n3383 = ~n3381 & ~n3382;
  assign n3384 = n3217 & ~n3383;
  assign n3385 = pi044 & n3221;
  assign n3386 = pi032 & ~n3221;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = ~n3217 & ~n3387;
  assign n3389 = ~n3384 & ~n3388;
  assign n3390 = n3254 & ~n3389;
  assign n3391 = pi017 & ~n3221;
  assign n3392 = pi016 & n3221;
  assign n3393 = ~n3391 & ~n3392;
  assign n3394 = n3217 & ~n3393;
  assign n3395 = pi031 & n3221;
  assign n3396 = pi015 & ~n3221;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = ~n3217 & ~n3397;
  assign n3399 = ~n3394 & ~n3398;
  assign n3400 = ~n3254 & ~n3399;
  assign n3401 = ~n3390 & ~n3400;
  assign n3402 = ~n3246 & ~n3401;
  assign n3403 = pi013 & ~n3221;
  assign n3404 = pi012 & n3221;
  assign n3405 = ~n3403 & ~n3404;
  assign n3406 = n3217 & ~n3405;
  assign n3407 = pi011 & ~n3221;
  assign n3408 = pi042 & n3221;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = ~n3217 & ~n3409;
  assign n3411 = ~n3406 & ~n3410;
  assign n3412 = n3266 & ~n3411;
  assign n3413 = ~n3402 & ~n3412;
  assign n3414 = ~n3380 & n3413;
  assign n3415 = ~n3306 & ~n3414;
  assign n3416 = pi048 & n3221;
  assign n3417 = pi047 & ~n3221;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = n3217 & ~n3418;
  assign n3420 = pi010 & n3221;
  assign n3421 = pi039 & ~n3221;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = ~n3217 & ~n3422;
  assign n3424 = ~n3419 & ~n3423;
  assign n3425 = ~n3254 & ~n3424;
  assign n3426 = pi009 & ~n3221;
  assign n3427 = pi008 & n3221;
  assign n3428 = ~n3426 & ~n3427;
  assign n3429 = n3217 & ~n3428;
  assign n3430 = pi037 & n3221;
  assign n3431 = pi038 & ~n3221;
  assign n3432 = ~n3430 & ~n3431;
  assign n3433 = ~n3217 & ~n3432;
  assign n3434 = ~n3429 & ~n3433;
  assign n3435 = n3254 & ~n3434;
  assign n3436 = ~n3425 & ~n3435;
  assign n3437 = ~n3246 & ~n3436;
  assign n3438 = pi007 & ~n3221;
  assign n3439 = pi036 & n3221;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = n3217 & ~n3440;
  assign n3442 = pi006 & n3221;
  assign n3443 = pi035 & ~n3221;
  assign n3444 = ~n3442 & ~n3443;
  assign n3445 = ~n3217 & ~n3444;
  assign n3446 = ~n3441 & ~n3445;
  assign n3447 = n3266 & ~n3446;
  assign n3448 = ~n3437 & ~n3447;
  assign n3449 = pi005 & n3221;
  assign n3450 = pi034 & ~n3221;
  assign n3451 = ~n3449 & ~n3450;
  assign n3452 = n3217 & ~n3451;
  assign n3453 = pi033 & n3221;
  assign n3454 = pi004 & ~n3221;
  assign n3455 = ~n3453 & ~n3454;
  assign n3456 = ~n3217 & ~n3455;
  assign n3457 = ~n3452 & ~n3456;
  assign n3458 = n3255 & ~n3457;
  assign n3459 = n3448 & ~n3458;
  assign n3460 = n3306 & ~n3459;
  assign n3461 = ~n3415 & ~n3460;
  assign n3462 = n3369 & n3461;
  assign n3463 = ~n3370 & ~n3462;
  assign n3464 = ~pi133 & pi178;
  assign n3465 = pi133 & ~pi178;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = n3297 & ~n3354;
  assign n3468 = ~n3249 & n3467;
  assign n3469 = ~n3292 & n3468;
  assign n3470 = ~n3292 & ~n3296;
  assign n3471 = ~n3293 & ~n3470;
  assign n3472 = ~n3354 & ~n3471;
  assign n3473 = ~n3469 & ~n3472;
  assign n3474 = ~n3355 & n3473;
  assign n3475 = ~n3466 & ~n3474;
  assign n3476 = n3466 & n3474;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = pi143 & ~n3477;
  assign n3479 = ~pi143 & ~n946;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = ~n3463 & ~n3480;
  assign n3482 = pi002 & ~n3221;
  assign n3483 = pi083 & n3221;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = n3217 & ~n3484;
  assign n3486 = pi082 & ~n3221;
  assign n3487 = pi098 & n3221;
  assign n3488 = ~n3486 & ~n3487;
  assign n3489 = ~n3217 & ~n3488;
  assign n3490 = ~n3485 & ~n3489;
  assign n3491 = ~n3254 & ~n3490;
  assign n3492 = pi081 & ~n3221;
  assign n3493 = pi080 & n3221;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = n3217 & ~n3494;
  assign n3496 = pi079 & ~n3221;
  assign n3497 = pi001 & n3221;
  assign n3498 = ~n3496 & ~n3497;
  assign n3499 = ~n3217 & ~n3498;
  assign n3500 = ~n3495 & ~n3499;
  assign n3501 = n3254 & ~n3500;
  assign n3502 = ~n3491 & ~n3501;
  assign n3503 = ~n3246 & ~n3502;
  assign n3504 = pi111 & n3221;
  assign n3505 = pi070 & ~n3221;
  assign n3506 = ~n3504 & ~n3505;
  assign n3507 = n3217 & ~n3506;
  assign n3508 = pi110 & ~n3221;
  assign n3509 = pi099 & n3221;
  assign n3510 = ~n3508 & ~n3509;
  assign n3511 = ~n3217 & ~n3510;
  assign n3512 = ~n3507 & ~n3511;
  assign n3513 = n3255 & ~n3512;
  assign n3514 = ~n3503 & ~n3513;
  assign n3515 = pi114 & ~n3221;
  assign n3516 = pi069 & n3221;
  assign n3517 = ~n3515 & ~n3516;
  assign n3518 = n3217 & ~n3517;
  assign n3519 = pi068 & ~n3221;
  assign n3520 = pi113 & n3221;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = ~n3217 & ~n3521;
  assign n3523 = ~n3518 & ~n3522;
  assign n3524 = n3266 & ~n3523;
  assign n3525 = n3514 & ~n3524;
  assign n3526 = ~n3306 & ~n3525;
  assign n3527 = pi075 & ~n3221;
  assign n3528 = pi109 & n3221;
  assign n3529 = ~n3527 & ~n3528;
  assign n3530 = n3217 & ~n3529;
  assign n3531 = pi100 & ~n3221;
  assign n3532 = pi101 & n3221;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = ~n3217 & ~n3533;
  assign n3535 = ~n3530 & ~n3534;
  assign n3536 = n3254 & ~n3535;
  assign n3537 = pi077 & n3221;
  assign n3538 = pi078 & ~n3221;
  assign n3539 = ~n3537 & ~n3538;
  assign n3540 = n3217 & ~n3539;
  assign n3541 = pi112 & n3221;
  assign n3542 = pi076 & ~n3221;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = ~n3217 & ~n3543;
  assign n3545 = ~n3540 & ~n3544;
  assign n3546 = ~n3254 & ~n3545;
  assign n3547 = ~n3536 & ~n3546;
  assign n3548 = ~n3246 & ~n3547;
  assign n3549 = pi000 & ~n3221;
  assign n3550 = pi107 & n3221;
  assign n3551 = ~n3549 & ~n3550;
  assign n3552 = n3217 & ~n3551;
  assign n3553 = pi106 & ~n3221;
  assign n3554 = pi074 & n3221;
  assign n3555 = ~n3553 & ~n3554;
  assign n3556 = ~n3217 & ~n3555;
  assign n3557 = ~n3552 & ~n3556;
  assign n3558 = n3266 & ~n3557;
  assign n3559 = ~n3548 & ~n3558;
  assign n3560 = pi072 & n3221;
  assign n3561 = pi073 & ~n3221;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = n3217 & ~n3562;
  assign n3564 = pi003 & n3221;
  assign n3565 = pi071 & ~n3221;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = ~n3217 & ~n3566;
  assign n3568 = ~n3563 & ~n3567;
  assign n3569 = n3255 & ~n3568;
  assign n3570 = n3559 & ~n3569;
  assign n3571 = n3306 & ~n3570;
  assign n3572 = ~n3526 & ~n3571;
  assign n3573 = ~n3369 & n3572;
  assign n3574 = pi027 & n3221;
  assign n3575 = pi065 & ~n3221;
  assign n3576 = ~n3574 & ~n3575;
  assign n3577 = n3217 & ~n3576;
  assign n3578 = pi025 & n3221;
  assign n3579 = pi026 & ~n3221;
  assign n3580 = ~n3578 & ~n3579;
  assign n3581 = ~n3217 & ~n3580;
  assign n3582 = ~n3577 & ~n3581;
  assign n3583 = n3255 & ~n3582;
  assign n3584 = pi049 & n3221;
  assign n3585 = pi050 & ~n3221;
  assign n3586 = ~n3584 & ~n3585;
  assign n3587 = n3217 & ~n3586;
  assign n3588 = pi051 & n3221;
  assign n3589 = pi059 & ~n3221;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = ~n3217 & ~n3590;
  assign n3592 = ~n3587 & ~n3591;
  assign n3593 = n3254 & ~n3592;
  assign n3594 = pi055 & ~n3221;
  assign n3595 = pi054 & n3221;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = n3217 & ~n3596;
  assign n3598 = pi053 & n3221;
  assign n3599 = pi052 & ~n3221;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = ~n3217 & ~n3600;
  assign n3602 = ~n3597 & ~n3601;
  assign n3603 = ~n3254 & ~n3602;
  assign n3604 = ~n3593 & ~n3603;
  assign n3605 = ~n3246 & ~n3604;
  assign n3606 = pi030 & ~n3221;
  assign n3607 = pi067 & n3221;
  assign n3608 = ~n3606 & ~n3607;
  assign n3609 = n3217 & ~n3608;
  assign n3610 = pi066 & ~n3221;
  assign n3611 = pi029 & n3221;
  assign n3612 = ~n3610 & ~n3611;
  assign n3613 = ~n3217 & ~n3612;
  assign n3614 = ~n3609 & ~n3613;
  assign n3615 = n3266 & ~n3614;
  assign n3616 = ~n3605 & ~n3615;
  assign n3617 = ~n3583 & n3616;
  assign n3618 = ~n3306 & ~n3617;
  assign n3619 = pi056 & n3221;
  assign n3620 = pi063 & ~n3221;
  assign n3621 = ~n3619 & ~n3620;
  assign n3622 = n3217 & ~n3621;
  assign n3623 = pi022 & n3221;
  assign n3624 = pi064 & ~n3221;
  assign n3625 = ~n3623 & ~n3624;
  assign n3626 = ~n3217 & ~n3625;
  assign n3627 = ~n3622 & ~n3626;
  assign n3628 = n3254 & ~n3627;
  assign n3629 = pi024 & ~n3221;
  assign n3630 = pi023 & n3221;
  assign n3631 = ~n3629 & ~n3630;
  assign n3632 = n3217 & ~n3631;
  assign n3633 = pi062 & ~n3221;
  assign n3634 = pi061 & n3221;
  assign n3635 = ~n3633 & ~n3634;
  assign n3636 = ~n3217 & ~n3635;
  assign n3637 = ~n3632 & ~n3636;
  assign n3638 = ~n3254 & ~n3637;
  assign n3639 = ~n3628 & ~n3638;
  assign n3640 = ~n3246 & ~n3639;
  assign n3641 = pi060 & n3221;
  assign n3642 = pi021 & ~n3221;
  assign n3643 = ~n3641 & ~n3642;
  assign n3644 = n3217 & ~n3643;
  assign n3645 = pi020 & n3221;
  assign n3646 = pi058 & ~n3221;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~n3217 & ~n3647;
  assign n3649 = ~n3644 & ~n3648;
  assign n3650 = n3266 & ~n3649;
  assign n3651 = ~n3640 & ~n3650;
  assign n3652 = pi019 & n3221;
  assign n3653 = pi057 & ~n3221;
  assign n3654 = ~n3652 & ~n3653;
  assign n3655 = n3217 & ~n3654;
  assign n3656 = pi018 & n3221;
  assign n3657 = pi028 & ~n3221;
  assign n3658 = ~n3656 & ~n3657;
  assign n3659 = ~n3217 & ~n3658;
  assign n3660 = ~n3655 & ~n3659;
  assign n3661 = n3255 & ~n3660;
  assign n3662 = n3651 & ~n3661;
  assign n3663 = n3306 & ~n3662;
  assign n3664 = ~n3618 & ~n3663;
  assign n3665 = n3369 & n3664;
  assign n3666 = ~n3573 & ~n3665;
  assign n3667 = n3480 & ~n3666;
  assign n3668 = ~n3481 & ~n3667;
  assign n3669 = ~n3206 & n3668;
  assign po175 = n3207 | n3669;
  assign n3671 = pi136 & ~n594;
  assign n3672 = ~pi169 & ~pi191;
  assign n3673 = ~pi141 & ~pi159;
  assign n3674 = n3672 & n3673;
  assign n3675 = ~pi164 & ~pi186;
  assign n3676 = ~pi167 & ~pi168;
  assign n3677 = n3675 & n3676;
  assign n3678 = n3674 & n3677;
  assign n3679 = ~pi149 & ~pi154;
  assign n3680 = ~pi162 & ~pi166;
  assign n3681 = ~pi132 & ~pi147;
  assign n3682 = n3680 & n3681;
  assign n3683 = n3679 & n3682;
  assign n3684 = ~pi170 & n3683;
  assign n3685 = ~pi165 & n3684;
  assign n3686 = n3678 & n3685;
  assign n3687 = n3671 & n3686;
  assign n3688 = pi129 & ~n3687;
  assign n3689 = ~pi129 & n3687;
  assign po176 = n3688 | n3689;
  assign n3691 = ~pi133 & ~pi140;
  assign n3692 = n666 & n3691;
  assign n3693 = n678 & n3692;
  assign n3694 = pi130 & ~n3693;
  assign n3695 = ~pi130 & n3693;
  assign n3696 = ~n3694 & ~n3695;
  assign n3697 = pi145 & ~n3696;
  assign n3698 = pi130 & ~pi145;
  assign n3699 = ~n3697 & ~n3698;
  assign n3700 = pi136 & ~n3699;
  assign n3701 = ~pi176 & ~pi177;
  assign n3702 = ~pi178 & n3701;
  assign n3703 = ~pi161 & n3702;
  assign n3704 = ~pi150 & n3703;
  assign n3705 = ~pi156 & ~pi171;
  assign n3706 = n3704 & n3705;
  assign n3707 = ~pi136 & n3706;
  assign po177 = n3700 | n3707;
  assign n3709 = ~pi131 & ~pi136;
  assign n3710 = pi145 & n593;
  assign n3711 = ~pi131 & ~n3710;
  assign n3712 = ~n3709 & ~n3711;
  assign n3713 = ~pi236 & pi237;
  assign n3714 = ~pi136 & pi233;
  assign n3715 = n3713 & n3714;
  assign n3716 = n575 & n3715;
  assign n3717 = ~n3712 & ~n3716;
  assign n3718 = ~pi131 & ~pi271;
  assign n3719 = ~n1600 & ~n3718;
  assign n3720 = n3716 & ~n3719;
  assign po178 = n3717 | n3720;
  assign n3722 = pi136 & ~n3686;
  assign n3723 = pi157 & ~n3722;
  assign n3724 = ~pi165 & ~pi170;
  assign n3725 = ~pi166 & n3724;
  assign n3726 = ~pi162 & n3725;
  assign n3727 = n3675 & n3726;
  assign n3728 = ~pi168 & n3727;
  assign n3729 = ~pi167 & n3728;
  assign n3730 = n3672 & n3729;
  assign n3731 = ~pi159 & n3730;
  assign n3732 = ~pi141 & n3731;
  assign n3733 = ~pi154 & n3732;
  assign n3734 = ~pi147 & n3733;
  assign n3735 = ~pi149 & n3734;
  assign n3736 = pi132 & n3735;
  assign n3737 = ~pi132 & ~n3735;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = n3722 & n3738;
  assign po179 = n3723 | n3739;
  assign n3741 = ~pi136 & pi178;
  assign n3742 = ~n3706 & n3741;
  assign n3743 = ~pi133 & ~pi145;
  assign n3744 = pi145 & n946;
  assign n3745 = ~n3743 & ~n3744;
  assign n3746 = pi136 & n3745;
  assign po180 = n3742 | n3746;
  assign n3748 = ~pi151 & n3710;
  assign n3749 = pi136 & n3748;
  assign n3750 = pi134 & ~pi228;
  assign po181 = n3749 | n3750;
  assign n3752 = ~pi235 & ~pi237;
  assign n3753 = pi236 & n3752;
  assign n3754 = pi038 & n3753;
  assign n3755 = pi235 & ~pi237;
  assign n3756 = ~pi236 & n3755;
  assign n3757 = pi100 & n3756;
  assign n3758 = ~n3754 & ~n3757;
  assign n3759 = ~pi236 & n3752;
  assign n3760 = pi064 & n3759;
  assign n3761 = pi235 & pi237;
  assign n3762 = ~pi236 & n3761;
  assign n3763 = pi185 & n3762;
  assign n3764 = ~pi235 & pi237;
  assign n3765 = ~pi236 & n3764;
  assign n3766 = pi138 & n3765;
  assign n3767 = ~n3763 & ~n3766;
  assign n3768 = pi236 & n3755;
  assign n3769 = pi103 & n3768;
  assign n3770 = n3767 & ~n3769;
  assign n3771 = ~n3760 & n3770;
  assign po182 = ~n3758 | ~n3771;
  assign n3773 = pi136 & ~n3710;
  assign po183 = n3709 | n3773;
  assign n3775 = pi009 & n3753;
  assign n3776 = pi075 & n3756;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = pi063 & n3759;
  assign n3779 = pi153 & n3762;
  assign n3780 = pi143 & n3765;
  assign n3781 = ~n3779 & ~n3780;
  assign n3782 = pi124 & n3768;
  assign n3783 = n3781 & ~n3782;
  assign n3784 = ~n3778 & n3783;
  assign po184 = ~n3777 | ~n3784;
  assign n3786 = n1874 & n3716;
  assign n3787 = pi271 & n3716;
  assign n3788 = pi138 & ~n3787;
  assign po185 = n3786 | n3788;
  assign n3790 = pi177 & ~n3706;
  assign n3791 = ~pi136 & n3790;
  assign n3792 = ~pi139 & ~pi145;
  assign n3793 = pi145 & ~n682;
  assign n3794 = ~n3792 & ~n3793;
  assign n3795 = pi136 & n3794;
  assign po186 = n3791 | n3795;
  assign n3797 = ~pi136 & pi161;
  assign n3798 = ~n3706 & n3797;
  assign n3799 = ~pi140 & ~pi145;
  assign n3800 = pi145 & n672;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = pi136 & n3801;
  assign po187 = n3798 | n3802;
  assign n3804 = pi153 & ~n3722;
  assign n3805 = pi141 & ~n3731;
  assign n3806 = ~n3732 & ~n3805;
  assign n3807 = n3722 & ~n3806;
  assign po188 = n3804 | n3807;
  assign n3809 = pi176 & ~n3706;
  assign n3810 = ~pi136 & n3809;
  assign n3811 = pi145 & n702;
  assign n3812 = ~pi142 & ~pi145;
  assign n3813 = ~n3811 & ~n3812;
  assign n3814 = pi136 & n3813;
  assign po189 = n3810 | n3814;
  assign n3816 = n1349 & n3716;
  assign n3817 = pi143 & ~n3787;
  assign po190 = n3816 | n3817;
  assign n3819 = pi144 & ~n3787;
  assign n3820 = n1329 & n3716;
  assign po191 = n3819 | n3820;
  assign n3822 = ~pi153 & ~pi173;
  assign n3823 = ~pi160 & ~pi185;
  assign n3824 = ~pi163 & ~pi172;
  assign n3825 = ~pi157 & ~pi180;
  assign n3826 = n3824 & n3825;
  assign n3827 = n3823 & n3826;
  assign n3828 = n3822 & n3827;
  assign n3829 = ~pi174 & ~pi179;
  assign n3830 = ~pi175 & ~pi181;
  assign n3831 = ~pi155 & ~pi182;
  assign n3832 = ~pi183 & ~pi184;
  assign n3833 = n3831 & n3832;
  assign n3834 = n3830 & n3833;
  assign n3835 = n3829 & n3834;
  assign n3836 = n3828 & n3835;
  assign n3837 = n3709 & n3836;
  assign n3838 = ~pi129 & pi136;
  assign n3839 = pi165 & n3678;
  assign n3840 = ~pi170 & n3839;
  assign n3841 = n3683 & n3840;
  assign n3842 = n3838 & n3841;
  assign n3843 = pi129 & n3836;
  assign n3844 = ~n3842 & ~n3843;
  assign po192 = n3837 | ~n3844;
  assign n3846 = pi129 & n3841;
  assign n3847 = ~pi129 & n3836;
  assign n3848 = ~n3846 & ~n3847;
  assign po193 = pi136 & ~n3848;
  assign n3850 = pi180 & ~n3722;
  assign n3851 = n3675 & n3724;
  assign n3852 = n3680 & n3851;
  assign n3853 = n3676 & n3852;
  assign n3854 = n3672 & n3853;
  assign n3855 = n3673 & n3854;
  assign n3856 = n3679 & n3855;
  assign n3857 = pi147 & n3856;
  assign n3858 = ~pi147 & ~n3856;
  assign n3859 = ~n3857 & ~n3858;
  assign n3860 = n3722 & n3859;
  assign po194 = n3850 | n3860;
  assign n3862 = ~pi136 & pi156;
  assign n3863 = ~n3706 & n3862;
  assign n3864 = ~pi145 & ~pi148;
  assign n3865 = pi145 & n721;
  assign n3866 = ~n3864 & ~n3865;
  assign n3867 = pi136 & n3866;
  assign po195 = n3863 | n3867;
  assign n3869 = pi163 & ~n3722;
  assign n3870 = ~pi154 & ~pi169;
  assign n3871 = ~pi165 & ~pi186;
  assign n3872 = n3680 & n3871;
  assign n3873 = ~pi170 & n3872;
  assign n3874 = n3676 & n3873;
  assign n3875 = ~pi191 & n3874;
  assign n3876 = ~pi164 & n3875;
  assign n3877 = n3870 & n3876;
  assign n3878 = n3673 & n3877;
  assign n3879 = pi149 & n3878;
  assign n3880 = ~pi149 & ~n3878;
  assign n3881 = ~n3879 & ~n3880;
  assign n3882 = n3722 & n3881;
  assign po196 = n3869 | n3882;
  assign n3884 = pi270 & n3716;
  assign n3885 = pi150 & ~n3884;
  assign n3886 = pi150 & pi270;
  assign n3887 = ~n1233 & ~n3886;
  assign n3888 = n3716 & ~n3887;
  assign po197 = n3885 | n3888;
  assign n3890 = n1367 & n3716;
  assign n3891 = ~pi151 & ~n3787;
  assign po198 = n3890 | n3891;
  assign n3893 = n1892 & n3716;
  assign n3894 = ~pi152 & ~n3787;
  assign po199 = n3893 | n3894;
  assign n3896 = n581 & n3713;
  assign n3897 = pi231 & n3896;
  assign n3898 = n3714 & n3897;
  assign n3899 = pi271 & n3898;
  assign n3900 = pi153 & ~n3899;
  assign n3901 = n1349 & n3898;
  assign po200 = n3900 | n3901;
  assign n3903 = n3677 & n3726;
  assign n3904 = n3674 & n3903;
  assign n3905 = pi154 & ~n3904;
  assign n3906 = ~pi154 & n3904;
  assign n3907 = ~n3905 & ~n3906;
  assign n3908 = n3722 & ~n3907;
  assign n3909 = pi172 & ~n3722;
  assign po201 = n3908 | n3909;
  assign n3911 = pi270 & n3898;
  assign n3912 = pi155 & ~n3911;
  assign n3913 = n1293 & n3898;
  assign po202 = n3912 | n3913;
  assign n3915 = n1274 & n3716;
  assign n3916 = pi156 & ~n3884;
  assign po203 = n3915 | n3916;
  assign n3918 = pi157 & ~n3899;
  assign n3919 = n1635 & n3898;
  assign po204 = n3918 | n3919;
  assign n3921 = n571 & n3716;
  assign n3922 = ~pi158 & ~n3884;
  assign po205 = n3921 | n3922;
  assign n3924 = ~pi159 & n3854;
  assign n3925 = pi159 & ~n3854;
  assign n3926 = ~n3924 & ~n3925;
  assign n3927 = n3722 & ~n3926;
  assign n3928 = pi173 & ~n3722;
  assign po206 = n3927 | n3928;
  assign n3930 = pi160 & ~n3899;
  assign n3931 = n1600 & n3898;
  assign po207 = n3930 | n3931;
  assign n3933 = n1819 & n3716;
  assign n3934 = pi161 & ~n3884;
  assign po208 = n3933 | n3934;
  assign n3936 = pi181 & ~n3722;
  assign n3937 = pi162 & ~n3725;
  assign n3938 = ~n3726 & ~n3937;
  assign n3939 = n3722 & ~n3938;
  assign po209 = n3936 | n3939;
  assign n3941 = pi163 & ~n3899;
  assign n3942 = n1892 & n3898;
  assign po210 = n3941 | n3942;
  assign n3944 = pi182 & ~n3722;
  assign n3945 = pi164 & n3873;
  assign n3946 = ~pi164 & ~n3873;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = n3722 & n3947;
  assign po211 = n3944 | n3948;
  assign n3950 = pi179 & ~n3722;
  assign n3951 = ~pi165 & n3722;
  assign po212 = n3950 | n3951;
  assign n3953 = pi175 & ~n3722;
  assign n3954 = pi166 & ~n3724;
  assign n3955 = ~n3725 & ~n3954;
  assign n3956 = n3722 & ~n3955;
  assign po213 = n3953 | n3956;
  assign n3958 = pi184 & ~n3722;
  assign n3959 = pi167 & ~n3728;
  assign n3960 = ~n3729 & ~n3959;
  assign n3961 = n3722 & ~n3960;
  assign po214 = n3958 | n3961;
  assign n3963 = pi183 & ~n3722;
  assign n3964 = pi168 & n3852;
  assign n3965 = ~pi168 & ~n3852;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = n3722 & n3966;
  assign po215 = n3963 | n3967;
  assign n3969 = pi185 & ~n3722;
  assign n3970 = pi169 & n3876;
  assign n3971 = ~pi169 & ~n3876;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = n3722 & n3972;
  assign po216 = n3969 | n3973;
  assign n3975 = pi174 & ~n3722;
  assign n3976 = pi165 & pi170;
  assign n3977 = ~n3724 & ~n3976;
  assign n3978 = n3722 & ~n3977;
  assign po217 = n3975 | n3978;
  assign n3980 = n1252 & n3716;
  assign n3981 = pi171 & ~n3884;
  assign po218 = n3980 | n3981;
  assign n3983 = pi172 & ~n3899;
  assign n3984 = n1367 & n3898;
  assign po219 = n3983 | n3984;
  assign n3986 = pi173 & ~n3899;
  assign n3987 = n1329 & n3898;
  assign po220 = n3986 | n3987;
  assign n3989 = pi174 & ~n3911;
  assign n3990 = n1252 & n3898;
  assign po221 = n3989 | n3990;
  assign n3992 = pi175 & ~n3911;
  assign n3993 = n1274 & n3898;
  assign po222 = n3992 | n3993;
  assign n3995 = n1800 & n3716;
  assign n3996 = pi176 & ~n3884;
  assign po223 = n3995 | n3996;
  assign n3998 = n1293 & n3716;
  assign n3999 = pi177 & ~n3884;
  assign po224 = n3998 | n3999;
  assign n4001 = n1838 & n3716;
  assign n4002 = pi178 & ~n3884;
  assign po225 = n4001 | n4002;
  assign n4004 = pi179 & ~n3911;
  assign n4005 = n1233 & n3898;
  assign po226 = n4004 | n4005;
  assign n4007 = pi180 & ~n3899;
  assign n4008 = n1605 & n3898;
  assign po227 = n4007 | n4008;
  assign n4010 = pi181 & ~n3911;
  assign n4011 = n1800 & n3898;
  assign po228 = n4010 | n4011;
  assign n4013 = pi182 & ~n3911;
  assign n4014 = n1819 & n3898;
  assign po229 = n4013 | n4014;
  assign n4016 = pi183 & ~n3911;
  assign n4017 = n1838 & n3898;
  assign po230 = n4016 | n4017;
  assign n4019 = pi184 & ~n3911;
  assign n4020 = n571 & n3898;
  assign po231 = n4019 | n4020;
  assign n4022 = pi185 & ~n3899;
  assign n4023 = n1874 & n3898;
  assign po232 = n4022 | n4023;
  assign n4025 = pi186 & ~n3726;
  assign n4026 = ~pi186 & n3726;
  assign n4027 = ~n4025 & ~n4026;
  assign n4028 = n3722 & ~n4027;
  assign n4029 = pi155 & ~n3722;
  assign po233 = n4028 | n4029;
  assign n4031 = ~pi136 & pi171;
  assign n4032 = ~n3706 & n4031;
  assign n4033 = ~pi145 & ~pi187;
  assign n4034 = pi145 & n732;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = pi136 & n4035;
  assign po234 = n4032 | n4036;
  assign n4038 = pi184 & n3762;
  assign n4039 = pi236 & n3764;
  assign n4040 = ~pi195 & n4039;
  assign n4041 = ~n4038 & ~n4040;
  assign n4042 = ~pi158 & n3765;
  assign n4043 = pi115 & n3768;
  assign n4044 = ~n4042 & ~n4043;
  assign n4045 = pi007 & n3753;
  assign n4046 = pi000 & n3756;
  assign n4047 = ~n4045 & ~n4046;
  assign n4048 = pi021 & n3759;
  assign n4049 = n4047 & ~n4048;
  assign n4050 = n4044 & n4049;
  assign po235 = ~n4041 | ~n4050;
  assign n4052 = pi181 & n3762;
  assign n4053 = ~pi193 & n4039;
  assign n4054 = ~n4052 & ~n4053;
  assign n4055 = pi176 & n3765;
  assign n4056 = pi119 & n3768;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = pi034 & n3753;
  assign n4059 = pi073 & n3756;
  assign n4060 = ~n4058 & ~n4059;
  assign n4061 = pi057 & n3759;
  assign n4062 = n4060 & ~n4061;
  assign n4063 = n4057 & n4062;
  assign po236 = ~n4054 | ~n4063;
  assign n4065 = ~pi145 & pi190;
  assign n4066 = pi145 & ~pi190;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = pi136 & ~n4067;
  assign n4069 = pi150 & ~n3706;
  assign n4070 = ~pi136 & n4069;
  assign po237 = n4068 | n4070;
  assign n4072 = pi191 & ~n3903;
  assign n4073 = ~pi191 & n3903;
  assign n4074 = ~n4072 & ~n4073;
  assign n4075 = n3722 & ~n4074;
  assign n4076 = pi160 & ~n3722;
  assign po238 = n4075 | n4076;
  assign n4078 = n574 & n3714;
  assign n4079 = pi231 & n4078;
  assign n4080 = pi237 & n4079;
  assign n4081 = pi236 & n4080;
  assign n4082 = n1819 & n4081;
  assign n4083 = pi270 & n4081;
  assign n4084 = ~pi192 & ~n4083;
  assign po239 = n4082 | n4084;
  assign n4086 = n1800 & n4081;
  assign n4087 = ~pi193 & ~n4083;
  assign po240 = n4086 | n4087;
  assign n4089 = n1252 & n4081;
  assign n4090 = ~pi194 & ~n4083;
  assign po241 = n4089 | n4090;
  assign n4092 = n571 & n4081;
  assign n4093 = ~pi195 & ~n4083;
  assign po242 = n4092 | n4093;
  assign n4095 = n1233 & n4081;
  assign n4096 = ~pi196 & ~n4083;
  assign po243 = n4095 | n4096;
  assign n4098 = n1274 & n4081;
  assign n4099 = ~pi197 & ~n4083;
  assign po244 = n4098 | n4099;
  assign n4101 = n1293 & n4081;
  assign n4102 = ~pi198 & ~n4083;
  assign po245 = n4101 | n4102;
  assign n4104 = n1838 & n4081;
  assign n4105 = ~pi199 & ~n4083;
  assign po246 = n4104 | n4105;
  assign n4107 = pi006 & n3753;
  assign n4108 = pi074 & n3756;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = pi020 & n3759;
  assign n4111 = pi155 & n3762;
  assign n4112 = ~pi198 & n4039;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = pi177 & n3765;
  assign n4115 = pi116 & n3768;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = n4113 & n4116;
  assign n4118 = ~n4110 & n4117;
  assign po247 = ~n4109 | ~n4118;
  assign n4120 = pi035 & n3753;
  assign n4121 = pi106 & n3756;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = pi058 & n3759;
  assign n4124 = pi182 & n3762;
  assign n4125 = ~pi192 & n4039;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = pi161 & n3765;
  assign n4128 = pi122 & n3768;
  assign n4129 = ~n4127 & ~n4128;
  assign n4130 = n4126 & n4129;
  assign n4131 = ~n4123 & n4130;
  assign po248 = ~n4122 | ~n4131;
  assign n4133 = pi033 & n3753;
  assign n4134 = pi003 & n3756;
  assign n4135 = ~n4133 & ~n4134;
  assign n4136 = pi018 & n3759;
  assign n4137 = pi179 & n3762;
  assign n4138 = ~pi196 & n4039;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = pi150 & n3765;
  assign n4141 = pi118 & n3768;
  assign n4142 = ~n4140 & ~n4141;
  assign n4143 = n4139 & n4142;
  assign n4144 = ~n4136 & n4143;
  assign po249 = ~n4135 | ~n4144;
  assign n4146 = pi004 & n3753;
  assign n4147 = pi071 & n3756;
  assign n4148 = ~n4146 & ~n4147;
  assign n4149 = pi028 & n3759;
  assign n4150 = pi174 & n3762;
  assign n4151 = ~pi194 & n4039;
  assign n4152 = ~n4150 & ~n4151;
  assign n4153 = pi171 & n3765;
  assign n4154 = pi089 & n3768;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = n4152 & n4155;
  assign n4157 = ~n4149 & n4156;
  assign po250 = ~n4148 | ~n4157;
  assign n4159 = pi036 & n3753;
  assign n4160 = pi107 & n3756;
  assign n4161 = ~n4159 & ~n4160;
  assign n4162 = pi060 & n3759;
  assign n4163 = pi183 & n3762;
  assign n4164 = ~pi199 & n4039;
  assign n4165 = ~n4163 & ~n4164;
  assign n4166 = pi178 & n3765;
  assign n4167 = pi123 & n3768;
  assign n4168 = ~n4166 & ~n4167;
  assign n4169 = n4165 & n4168;
  assign n4170 = ~n4162 & n4169;
  assign po251 = ~n4161 | ~n4170;
  assign n4172 = pi005 & n3753;
  assign n4173 = pi072 & n3756;
  assign n4174 = ~n4172 & ~n4173;
  assign n4175 = pi019 & n3759;
  assign n4176 = pi175 & n3762;
  assign n4177 = ~pi197 & n4039;
  assign n4178 = ~n4176 & ~n4177;
  assign n4179 = pi156 & n3765;
  assign n4180 = pi096 & n3768;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = n4178 & n4181;
  assign n4183 = ~n4175 & n4182;
  assign po252 = ~n4174 | ~n4183;
  assign n4185 = pi008 & n3753;
  assign n4186 = pi109 & n3756;
  assign n4187 = ~n4185 & ~n4186;
  assign n4188 = pi056 & n3759;
  assign n4189 = pi173 & n3762;
  assign n4190 = pi144 & n3765;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = pi117 & n3768;
  assign n4193 = n4191 & ~n4192;
  assign n4194 = ~n4188 & n4193;
  assign po253 = ~n4187 | ~n4194;
  assign n4196 = pi039 & n3753;
  assign n4197 = pi076 & n3756;
  assign n4198 = ~n4196 & ~n4197;
  assign n4199 = pi062 & n3759;
  assign n4200 = pi163 & n3762;
  assign n4201 = ~pi152 & n3765;
  assign n4202 = ~n4200 & ~n4201;
  assign n4203 = pi125 & n3768;
  assign n4204 = n4202 & ~n4203;
  assign n4205 = ~n4199 & n4204;
  assign po254 = ~n4198 | ~n4205;
  assign n4207 = pi180 & n3762;
  assign n4208 = pi023 & n3759;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = pi126 & n3768;
  assign n4211 = pi048 & n3753;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = pi077 & n3756;
  assign n4214 = n4212 & ~n4213;
  assign po255 = ~n4209 | ~n4214;
  assign n4216 = pi010 & n3753;
  assign n4217 = pi112 & n3756;
  assign n4218 = ~n4216 & ~n4217;
  assign n4219 = pi061 & n3759;
  assign n4220 = pi172 & n3762;
  assign n4221 = ~pi151 & n3765;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = pi105 & n3768;
  assign n4224 = n4222 & ~n4223;
  assign n4225 = ~n4219 & n4224;
  assign po256 = ~n4218 | ~n4225;
  assign n4227 = pi037 & n3753;
  assign n4228 = pi101 & n3756;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = pi022 & n3759;
  assign n4231 = pi160 & n3762;
  assign n4232 = ~pi131 & n3765;
  assign n4233 = ~n4231 & ~n4232;
  assign n4234 = pi084 & n3768;
  assign n4235 = n4233 & ~n4234;
  assign n4236 = ~n4230 & n4235;
  assign po257 = ~n4229 | ~n4236;
  assign n4238 = pi157 & n3762;
  assign n4239 = pi024 & n3759;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = pi085 & n3768;
  assign n4242 = pi047 & n3753;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = pi078 & n3756;
  assign n4245 = n4243 & ~n4244;
  assign po258 = ~n4240 | ~n4245;
  assign n4247 = pi080 & n3756;
  assign n4248 = pi046 & n3753;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = pi093 & n3768;
  assign n4251 = pi049 & n3759;
  assign n4252 = ~n4250 & ~n4251;
  assign po259 = ~n4249 | ~n4252;
  assign n4254 = pi086 & n3768;
  assign n4255 = pi040 & n3753;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = pi025 & n3759;
  assign n4258 = pi099 & n3756;
  assign n4259 = ~n4257 & ~n4258;
  assign po260 = ~n4256 | ~n4259;
  assign n4261 = pi027 & n3759;
  assign n4262 = pi111 & n3756;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = pi097 & n3768;
  assign n4265 = pi045 & n3753;
  assign n4266 = ~n4264 & ~n4265;
  assign po261 = ~n4263 | ~n4266;
  assign n4268 = pi104 & n3768;
  assign n4269 = pi043 & n3753;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = pi026 & n3759;
  assign n4272 = pi110 & n3756;
  assign n4273 = ~n4271 & ~n4272;
  assign po262 = ~n4270 | ~n4273;
  assign n4275 = pi121 & n3768;
  assign n4276 = pi041 & n3753;
  assign n4277 = ~n4275 & ~n4276;
  assign n4278 = pi065 & n3759;
  assign n4279 = pi070 & n3756;
  assign n4280 = ~n4278 & ~n4279;
  assign po263 = ~n4277 | ~n4280;
  assign n4282 = pi120 & n3768;
  assign n4283 = pi012 & n3753;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = pi067 & n3759;
  assign n4286 = pi069 & n3756;
  assign n4287 = ~n4285 & ~n4286;
  assign po264 = ~n4284 | ~n4287;
  assign n4289 = pi050 & n3759;
  assign n4290 = pi081 & n3756;
  assign n4291 = ~n4289 & ~n4290;
  assign n4292 = pi090 & n3768;
  assign n4293 = pi014 & n3753;
  assign n4294 = ~n4292 & ~n4293;
  assign po265 = ~n4291 | ~n4294;
  assign n4296 = pi066 & n3759;
  assign n4297 = pi068 & n3756;
  assign n4298 = ~n4296 & ~n4297;
  assign n4299 = pi127 & n3768;
  assign n4300 = pi011 & n3753;
  assign n4301 = ~n4299 & ~n4300;
  assign po266 = ~n4298 | ~n4301;
  assign n4303 = pi055 & n3759;
  assign n4304 = pi002 & n3756;
  assign n4305 = ~n4303 & ~n4304;
  assign n4306 = pi094 & n3768;
  assign n4307 = pi017 & n3753;
  assign n4308 = ~n4306 & ~n4307;
  assign po267 = ~n4305 | ~n4308;
  assign n4310 = pi053 & n3759;
  assign n4311 = pi098 & n3756;
  assign n4312 = ~n4310 & ~n4311;
  assign n4313 = pi095 & n3768;
  assign n4314 = pi031 & n3753;
  assign n4315 = ~n4313 & ~n4314;
  assign po268 = ~n4312 | ~n4315;
  assign n4317 = pi051 & n3759;
  assign n4318 = pi001 & n3756;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = pi102 & n3768;
  assign n4321 = pi044 & n3753;
  assign n4322 = ~n4320 & ~n4321;
  assign po269 = ~n4319 | ~n4322;
  assign n4324 = pi030 & n3759;
  assign n4325 = pi114 & n3756;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = pi087 & n3768;
  assign n4328 = pi013 & n3753;
  assign n4329 = ~n4327 & ~n4328;
  assign po270 = ~n4326 | ~n4329;
  assign n4331 = pi054 & n3759;
  assign n4332 = pi083 & n3756;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = pi092 & n3768;
  assign n4335 = pi016 & n3753;
  assign n4336 = ~n4334 & ~n4335;
  assign po271 = ~n4333 | ~n4336;
  assign n4338 = pi029 & n3759;
  assign n4339 = pi113 & n3756;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = pi108 & n3768;
  assign n4342 = pi042 & n3753;
  assign n4343 = ~n4341 & ~n4342;
  assign po272 = ~n4340 | ~n4343;
  assign n4345 = pi052 & n3759;
  assign n4346 = pi082 & n3756;
  assign n4347 = ~n4345 & ~n4346;
  assign n4348 = pi091 & n3768;
  assign n4349 = pi015 & n3753;
  assign n4350 = ~n4348 & ~n4349;
  assign po273 = ~n4347 | ~n4350;
  assign n4352 = pi059 & n3759;
  assign n4353 = pi079 & n3756;
  assign n4354 = ~n4352 & ~n4353;
  assign n4355 = pi088 & n3768;
  assign n4356 = pi032 & n3753;
  assign n4357 = ~n4355 & ~n4356;
  assign po274 = ~n4354 | ~n4357;
  assign po275 = ~pi228 & n561;
  assign po045 = 1'b1;
  assign po044 = ~pi230;
  assign po000 = pi202;
  assign po001 = pi203;
  assign po002 = pi205;
  assign po003 = pi189;
  assign po004 = pi200;
  assign po005 = pi201;
  assign po006 = pi204;
  assign po007 = pi188;
  assign po008 = pi210;
  assign po009 = pi135;
  assign po010 = pi206;
  assign po011 = pi137;
  assign po012 = pi209;
  assign po013 = pi207;
  assign po014 = pi208;
  assign po015 = pi211;
  assign po016 = pi213;
  assign po017 = pi215;
  assign po018 = pi214;
  assign po019 = pi216;
  assign po020 = pi225;
  assign po021 = pi219;
  assign po022 = pi217;
  assign po023 = pi223;
  assign po024 = pi222;
  assign po025 = pi227;
  assign po026 = pi212;
  assign po027 = pi218;
  assign po028 = pi221;
  assign po029 = pi226;
  assign po030 = pi224;
  assign po031 = pi220;
  assign po032 = pi228;
  assign po033 = pi134;
  assign po034 = pi129;
  assign po035 = pi128;
  assign po046 = pi229;
endmodule


